* SPICE3 file created from nand4_x.ext - technology: sky130B

.subckt nand4 A B C D VSS VDD Y
X0 Y.t4 D.t0 VDD.t2 w_n37_916.t3 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1 Y.t5 D.t1 a_284_88.t0 VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2 a_284_88.t1 C.t0 a_188_88.t0 VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3 a_92_88.t0 A.t0 VSS.t0 VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X4 a_188_88.t1 B.t0 a_92_88.t1 VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X5 a_572_88.t1 C.t1 a_476_88.t1 VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X6 a_476_88.t0 D.t2 Y.t2 VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X7 Y.t1 B.t1 VDD.t1 w_n37_916.t1 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X8 VDD.t5 C.t2 Y.t7 w_n37_916.t5 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X9 VSS.t1 A.t1 a_668_88.t0 VSUBS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X10 a_668_88.t1 B.t2 a_572_88.t0 VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X11 VDD.t0 A.t2 Y.t0 w_n37_916.t0 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X12 Y.t6 C.t3 VDD.t4 w_n37_916.t4 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X13 Y.t9 A.t3 VDD.t7 w_n37_916.t7 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X14 VDD.t3 D.t3 Y.t3 w_n37_916.t2 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X15 VDD.t6 B.t3 Y.t8 w_n37_916.t6 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
R0 D.n1 D.t2 396.372
R1 D.n1 D.t1 395.014
R2 D.n0 D.t3 378.589
R3 D.n0 D.t0 308.481
R4 D.n2 D.n0 162.359
R5 D.n2 D.n1 161.3
R6 D D.n2 0.813906
R7 VDD.n3 VDD.t7 205.349
R8 VDD.n0 VDD.t3 205.349
R9 VDD.n5 VDD.n4 185.16
R10 VDD VDD.n6 185.16
R11 VDD.n2 VDD.n1 185.16
R12 VDD.n4 VDD.t1 20.1899
R13 VDD.n4 VDD.t0 20.1899
R14 VDD.n6 VDD.t4 20.1899
R15 VDD.n6 VDD.t6 20.1899
R16 VDD.n1 VDD.t2 20.1899
R17 VDD.n1 VDD.t5 20.1899
R18 VDD.n0 VDD 0.813226
R19 VDD.n2 VDD.n0 0.122949
R20 VDD VDD.n2 0.122949
R21 VDD VDD.n5 0.122949
R22 VDD.n5 VDD.n3 0.122949
R23 VDD.n3 VDD 0.0189949
R24 Y.n2 Y.n0 187.373
R25 Y.n2 Y.n1 187.192
R26 Y.n4 Y.n3 187.192
R27 Y.n6 Y.n5 187.192
R28 Y Y.n8 32.908
R29 Y.n0 Y.t0 20.1899
R30 Y.n0 Y.t9 20.1899
R31 Y.n1 Y.t8 20.1899
R32 Y.n1 Y.t1 20.1899
R33 Y.n3 Y.t7 20.1899
R34 Y.n3 Y.t6 20.1899
R35 Y.n5 Y.t3 20.1899
R36 Y.n5 Y.t4 20.1899
R37 Y.n8 Y.t2 9.9005
R38 Y.n8 Y.t5 9.9005
R39 Y.n6 Y.n4 0.179604
R40 Y.n4 Y.n2 0.179604
R41 Y.n7 Y.n6 0.169597
R42 Y.n7 Y 0.00298344
R43 Y Y.n7 0.00202439
R44 w_n37_916.n0 w_n37_916.t7 219.835
R45 w_n37_916.t3 w_n37_916.t2 188.43
R46 w_n37_916.t5 w_n37_916.t3 188.43
R47 w_n37_916.t4 w_n37_916.t5 188.43
R48 w_n37_916.t6 w_n37_916.t4 188.43
R49 w_n37_916.t1 w_n37_916.t6 188.43
R50 w_n37_916.t0 w_n37_916.t1 188.43
R51 w_n37_916.t7 w_n37_916.t0 188.43
R52 a_284_88.t0 a_284_88.t1 19.8005
R53 C.n1 C.t1 659.222
R54 C.n1 C.t0 631.28
R55 C.n0 C.t2 378.589
R56 C.n0 C.t3 308.481
R57 C.n2 C.n0 161.922
R58 C.n2 C.n1 161.3
R59 C C.n2 0.779486
R60 a_188_88.t0 a_188_88.t1 19.8005
R61 A.t0 A.n0 676.337
R62 A.n1 A.t1 596.697
R63 A.n1 A.t0 495.663
R64 A.n0 A.t2 361.062
R65 A.n0 A.t3 331.533
R66 A.n2 A.n1 158.75
R67 A.n2 A.n0 152
R68 A A.n2 9.38979
R69 VSS VSS.t1 43.6442
R70 VSS.n0 VSS.t0 42.5938
R71 VSS.n1 VSS 0.393978
R72 VSS.n1 VSS.n0 0.0720206
R73 VSS.n1 VSS 0.0559348
R74 VSS VSS.n1 0.0114536
R75 VSS.n0 VSS 0.00672852
R76 a_92_88.t0 a_92_88.t1 19.8005
R77 B.t0 B.n1 633.284
R78 B.n2 B.t2 530.331
R79 B.n2 B.t0 514.096
R80 B.n0 B.t3 353.029
R81 B.n0 B.t1 330.974
R82 B.n4 B.n0 161.76
R83 B.n3 B.n1 152
R84 B.n1 B.n0 94.0247
R85 B.n3 B.n2 68.0971
R86 B.n4 B.n3 9.3005
R87 B B.n4 0.413543
R88 a_476_88.t0 a_476_88.t1 19.8005
R89 a_572_88.t0 a_572_88.t1 19.8005
R90 a_668_88.t0 a_668_88.t1 19.8005
C0 D A 0.120842f
C1 D Y 1.1806f
C2 A Y 0.368563f
C3 D B 0.234677f
C4 B A 3.01059f
C5 VDD C 0.023317f
C6 D VSS 0.413731f
C7 A VSS 1.12039f
C8 B Y 0.637694f
C9 Y VSS 1.27567f
C10 B VSS 0.400149f
C11 D VDD 0.024765f
C12 VDD A 0.056468f
C13 VDD Y 1.98533f
C14 VDD B 0.025356f
C15 VDD VSS 0.003468f
C16 D C 1.44042f
C17 C A 0.133449f
C18 C Y 0.142092f
C19 C B 1.14663f
C20 C VSS 0.004517f
C21 VSS VSUBS 0.622116f
C22 Y VSUBS 0.348866f
C23 VDD VSUBS 0.471795f
C24 D VSUBS 0.31561f
C25 C VSUBS 0.476083f
C26 B VSUBS 0.838493f
C27 A VSUBS 1.833005f
C28 B.t3 VSUBS 0.062553f
C29 B.t1 VSUBS 0.058765f
C30 B.n0 VSUBS 0.155388f
C31 B.n1 VSUBS 0.235096f
C32 B.t2 VSUBS 0.120805f
C33 B.t0 VSUBS 0.130739f
C34 B.n2 VSUBS 0.773955f
C35 B.n3 VSUBS 1.15399f
C36 B.n4 VSUBS 0.244581f
C37 A.t2 VSUBS 0.070188f
C38 A.t3 VSUBS 0.064546f
C39 A.n0 VSUBS 0.336828f
C40 A.t1 VSUBS 0.197923f
C41 A.t0 VSUBS 0.227883f
C42 A.n1 VSUBS 1.20419f
C43 A.n2 VSUBS 0.686187f
.ends

