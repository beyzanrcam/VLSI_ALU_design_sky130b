magic
tech sky130B
magscale 1 2
timestamp 1734792667
<< error_s >>
rect 892 683 6297 684
rect 126 266 6297 683
rect 6298 266 7237 684
rect 126 265 5531 266
rect 226 139 426 197
rect 616 139 816 197
rect 1117 139 1317 197
rect 1507 139 1707 197
rect 2029 139 2229 197
rect 2419 139 2619 197
rect 2921 140 3121 198
rect 3311 140 3511 198
rect 3813 140 4013 198
rect 4203 140 4403 198
rect 4712 140 4912 198
rect 5102 140 5302 198
rect 5631 140 5831 198
rect 6021 140 6221 198
rect 6571 140 6771 198
rect 6961 140 7161 198
rect 226 51 426 109
rect 616 51 816 109
rect 1117 51 1317 109
rect 1507 51 1707 109
rect 2029 51 2229 109
rect 2419 51 2619 109
rect 2921 52 3121 110
rect 3311 52 3511 110
rect 3813 52 4013 110
rect 4203 52 4403 110
rect 4712 52 4912 110
rect 5102 52 5302 110
rect 5631 52 5831 110
rect 6021 52 6221 110
rect 6571 52 6771 110
rect 6961 52 7161 110
<< nwell >>
rect 892 265 5531 684
rect 6298 266 6551 684
<< metal1 >>
rect 112 603 179 816
rect 1003 603 1070 816
rect 1915 603 1982 816
rect 2807 604 2874 817
rect 3699 604 3766 817
rect 4598 604 4665 817
rect 5517 604 5584 817
rect 6457 604 6524 817
rect 892 16 975 603
rect 1783 16 1866 603
rect 2695 16 2778 603
rect 3587 16 3670 604
rect 4479 16 4562 604
rect 5378 16 5461 604
rect 6297 16 6380 604
rect 7237 16 7320 604
use buffer  buffer_0 ~/Documents/Dersler/VLSI/vlsi_sky130b/design/mag/inv
timestamp 1734791363
transform 1 0 -1346 0 1 312
box 1458 -297 2238 371
use buffer  buffer_1
timestamp 1734791363
transform 1 0 -455 0 1 312
box 1458 -297 2238 371
use buffer  buffer_2
timestamp 1734791363
transform 1 0 2241 0 1 313
box 1458 -297 2238 371
use buffer  buffer_3
timestamp 1734791363
transform 1 0 457 0 1 312
box 1458 -297 2238 371
use buffer  buffer_4
timestamp 1734791363
transform 1 0 1349 0 1 313
box 1458 -297 2238 371
use buffer  buffer_5
timestamp 1734791363
transform 1 0 4059 0 1 313
box 1458 -297 2238 371
use buffer  buffer_6
timestamp 1734791363
transform 1 0 3140 0 1 313
box 1458 -297 2238 371
use buffer  buffer_7
timestamp 1734791363
transform 1 0 4999 0 1 313
box 1458 -297 2238 371
<< end >>
