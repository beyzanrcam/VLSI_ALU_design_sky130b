magic
tech sky130B
magscale 1 2
timestamp 1735226356
<< error_s >>
rect 1472 -47 2227 371
rect 1572 -173 1772 -115
rect 1951 -173 2151 -115
rect 1572 -261 1772 -203
rect 1951 -261 2151 -203
rect 1697 -294 2017 -270
rect 1697 -566 1721 -294
rect 1697 -590 2017 -566
<< nwell >>
rect 1848 -47 1851 371
<< metal1 >>
rect 1572 527 2165 547
rect 1572 405 1801 527
rect 1923 405 2165 527
rect 1572 371 2165 405
rect 1786 319 1951 371
rect 1848 -222 1851 291
rect 1772 -297 1951 -250
rect 1833 -398 1880 -297
rect 1831 -404 1883 -398
rect 1831 -462 1883 -456
<< via1 >>
rect 1801 405 1923 527
rect 1831 -456 1883 -404
<< metal2 >>
rect 1790 527 1934 533
rect 1790 405 1801 527
rect 1923 405 1934 527
rect 1790 399 1934 405
rect 1820 -402 1894 -401
rect 1820 -458 1829 -402
rect 1885 -458 1894 -402
<< via2 >>
rect 1801 405 1923 527
rect 1829 -404 1885 -402
rect 1829 -456 1831 -404
rect 1831 -456 1883 -404
rect 1883 -456 1885 -404
rect 1829 -458 1885 -456
<< metal3 >>
rect 1790 532 1934 533
rect 1790 400 1796 532
rect 1928 400 1934 532
rect 1790 399 1934 400
rect 1787 -397 1927 -396
rect 1787 -463 1824 -397
rect 1890 -463 1927 -397
rect 1787 -465 1927 -463
<< via3 >>
rect 1796 527 1928 532
rect 1796 405 1801 527
rect 1801 405 1923 527
rect 1923 405 1928 527
rect 1796 400 1928 405
rect 1824 -402 1890 -397
rect 1824 -458 1829 -402
rect 1829 -458 1885 -402
rect 1885 -458 1890 -402
rect 1824 -463 1890 -458
<< metal4 >>
rect 1795 532 1929 533
rect 1795 400 1796 532
rect 1928 400 1929 532
rect 1795 399 1929 400
<< via4 >>
rect 1721 -397 1993 -294
rect 1721 -463 1824 -397
rect 1824 -463 1890 -397
rect 1890 -463 1993 -397
rect 1721 -566 1993 -463
<< metal5 >>
rect 1697 -294 2017 -270
rect 1697 -566 1721 -294
rect 1993 -566 2017 -294
rect 1697 -590 2017 -566
use inv  inv_0
timestamp 1735171245
transform 1 0 1472 0 1 -47
box 0 -250 376 418
use inv  inv_1
timestamp 1735171245
transform 1 0 1851 0 1 -47
box 0 -250 376 418
<< end >>
