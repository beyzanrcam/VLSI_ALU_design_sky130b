magic
tech sky130B
magscale 1 2
timestamp 1732965435
<< error_p >>
rect -77 472 -19 478
rect 115 472 173 478
rect -77 438 -65 472
rect 115 438 127 472
rect -77 432 -19 438
rect 115 432 173 438
rect -173 -438 -115 -432
rect 19 -438 77 -432
rect -173 -472 -161 -438
rect 19 -472 31 -438
rect -173 -478 -115 -472
rect 19 -478 77 -472
<< nmos >>
rect -159 -400 -129 400
rect -63 -400 -33 400
rect 33 -400 63 400
rect 129 -400 159 400
<< ndiff >>
rect -221 388 -159 400
rect -221 -388 -209 388
rect -175 -388 -159 388
rect -221 -400 -159 -388
rect -129 388 -63 400
rect -129 -388 -113 388
rect -79 -388 -63 388
rect -129 -400 -63 -388
rect -33 388 33 400
rect -33 -388 -17 388
rect 17 -388 33 388
rect -33 -400 33 -388
rect 63 388 129 400
rect 63 -388 79 388
rect 113 -388 129 388
rect 63 -400 129 -388
rect 159 388 221 400
rect 159 -388 175 388
rect 209 -388 221 388
rect 159 -400 221 -388
<< ndiffc >>
rect -209 -388 -175 388
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
rect 175 -388 209 388
<< poly >>
rect -81 472 -15 488
rect -81 438 -65 472
rect -31 438 -15 472
rect -159 400 -129 426
rect -81 422 -15 438
rect 111 472 177 488
rect 111 438 127 472
rect 161 438 177 472
rect -63 400 -33 422
rect 33 400 63 426
rect 111 422 177 438
rect 129 400 159 422
rect -159 -422 -129 -400
rect -177 -438 -111 -422
rect -63 -426 -33 -400
rect 33 -422 63 -400
rect -177 -472 -161 -438
rect -127 -472 -111 -438
rect -177 -488 -111 -472
rect 15 -438 81 -422
rect 129 -426 159 -400
rect 15 -472 31 -438
rect 65 -472 81 -438
rect 15 -488 81 -472
<< polycont >>
rect -65 438 -31 472
rect 127 438 161 472
rect -161 -472 -127 -438
rect 31 -472 65 -438
<< locali >>
rect -81 438 -65 472
rect -31 438 -15 472
rect 111 438 127 472
rect 161 438 177 472
rect -209 388 -175 404
rect -209 -404 -175 -388
rect -113 388 -79 404
rect -113 -404 -79 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 79 388 113 404
rect 79 -404 113 -388
rect 175 388 209 404
rect 175 -404 209 -388
rect -177 -472 -161 -438
rect -127 -472 -111 -438
rect 15 -472 31 -438
rect 65 -472 81 -438
<< viali >>
rect -65 438 -31 472
rect 127 438 161 472
rect -209 -388 -175 388
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
rect 175 -388 209 388
rect -161 -472 -127 -438
rect 31 -472 65 -438
<< metal1 >>
rect -77 472 -19 478
rect -77 438 -65 472
rect -31 438 -19 472
rect -77 432 -19 438
rect 115 472 173 478
rect 115 438 127 472
rect 161 438 173 472
rect 115 432 173 438
rect -215 388 -169 400
rect -215 -388 -209 388
rect -175 -388 -169 388
rect -215 -400 -169 -388
rect -119 388 -73 400
rect -119 -388 -113 388
rect -79 -388 -73 388
rect -119 -400 -73 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 73 388 119 400
rect 73 -388 79 388
rect 113 -388 119 388
rect 73 -400 119 -388
rect 169 388 215 400
rect 169 -388 175 388
rect 209 -388 215 388
rect 169 -400 215 -388
rect -173 -438 -115 -432
rect -173 -472 -161 -438
rect -127 -472 -115 -438
rect -173 -478 -115 -472
rect 19 -438 77 -432
rect 19 -472 31 -438
rect 65 -472 77 -438
rect 19 -478 77 -472
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 0.150 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
