magic
tech sky130B
magscale 1 2
timestamp 1734801607
<< error_s >>
rect 1472 -47 2238 371
rect 1572 -173 1772 -115
rect 1962 -173 2162 -115
rect 1572 -261 1772 -203
rect 1962 -261 2162 -203
rect 1709 -286 2029 -262
rect 1709 -558 1733 -286
rect 1709 -582 2029 -558
<< nwell >>
rect 1790 319 1958 371
rect 1813 -47 1936 319
<< metal1 >>
rect 1568 496 2180 516
rect 1568 374 1807 496
rect 1929 374 2180 496
rect 1568 340 2180 374
rect 1689 -297 2065 -262
rect 1568 -334 2166 -297
rect 1568 -473 1781 -334
rect 1774 -510 1781 -473
rect 1957 -473 2166 -334
rect 1957 -510 1964 -473
<< via1 >>
rect 1807 374 1929 496
rect 1781 -510 1957 -334
<< metal2 >>
rect 1796 496 1940 502
rect 1796 374 1807 496
rect 1929 374 1940 496
rect 1796 368 1940 374
rect 1770 -334 1968 -329
rect 1770 -510 1781 -334
rect 1957 -510 1968 -334
rect 1770 -515 1968 -510
<< via2 >>
rect 1807 374 1929 496
rect 1781 -510 1957 -334
<< metal3 >>
rect 1796 501 1940 502
rect 1796 369 1802 501
rect 1934 369 1940 501
rect 1796 368 1940 369
rect 1770 -515 1776 -329
rect 1962 -515 1968 -329
<< via3 >>
rect 1802 496 1934 501
rect 1802 374 1807 496
rect 1807 374 1929 496
rect 1929 374 1934 496
rect 1802 369 1934 374
rect 1776 -334 1962 -329
rect 1776 -510 1781 -334
rect 1781 -510 1957 -334
rect 1957 -510 1962 -334
rect 1776 -515 1962 -510
<< metal4 >>
rect 1801 501 1935 502
rect 1801 369 1802 501
rect 1934 369 1935 501
rect 1801 368 1935 369
rect 1684 -286 2055 -285
rect 1684 -558 1733 -286
rect 2005 -558 2055 -286
<< via4 >>
rect 1733 -329 2005 -286
rect 1733 -515 1776 -329
rect 1776 -515 1962 -329
rect 1962 -515 2005 -329
rect 1733 -558 2005 -515
<< metal5 >>
rect 1709 -286 2029 -262
rect 1709 -558 1733 -286
rect 2005 -558 2029 -286
rect 1709 -582 2029 -558
use inv  inv_0
timestamp 1734798227
transform 1 0 1472 0 1 -47
box -14 -250 376 418
use inv  inv_1
timestamp 1734798227
transform 1 0 1862 0 1 -47
box -14 -250 376 418
<< end >>
