magic
tech sky130B
magscale 1 2
timestamp 1734801607
<< error_s >>
rect 781 683 782 828
rect 809 683 810 856
rect 1672 684 1673 828
rect 1700 684 1701 856
rect 2584 684 2585 828
rect 2612 684 2613 856
rect 3476 684 3477 829
rect 3504 684 3505 857
rect 4368 684 4369 829
rect 4396 684 4397 857
rect 5267 684 5268 829
rect 5295 684 5296 857
rect 6186 684 6187 829
rect 6214 684 6215 857
rect 7126 684 7127 829
rect 7154 684 7155 857
rect 878 683 7223 684
rect 112 266 7223 683
rect 112 265 6457 266
rect 188 139 388 197
rect 578 139 778 197
rect 1079 139 1279 197
rect 1469 139 1669 197
rect 1991 139 2191 197
rect 2381 139 2581 197
rect 2883 140 3083 198
rect 3273 140 3473 198
rect 3775 140 3975 198
rect 4165 140 4365 198
rect 4674 140 4874 198
rect 5064 140 5264 198
rect 5593 140 5793 198
rect 5983 140 6183 198
rect 6533 140 6733 198
rect 6923 140 7123 198
rect 188 51 388 109
rect 578 51 778 109
rect 1079 51 1279 109
rect 1469 51 1669 109
rect 1991 51 2191 109
rect 2381 51 2581 109
rect 2883 52 3083 110
rect 3273 52 3473 110
rect 3775 52 3975 110
rect 4165 52 4365 110
rect 4674 52 4874 110
rect 5064 52 5264 110
rect 5593 52 5793 110
rect 5983 52 6183 110
rect 6533 52 6733 110
rect 6923 52 7123 110
rect 321 26 641 50
rect 1212 26 1532 50
rect 2124 26 2444 50
rect 3016 27 3336 51
rect 3908 27 4228 51
rect 4807 27 5127 51
rect 5726 27 6046 51
rect 6666 27 6986 51
rect 321 -246 345 26
rect 1212 -246 1236 26
rect 2124 -246 2148 26
rect 3016 -245 3040 27
rect 3908 -245 3932 27
rect 4807 -245 4831 27
rect 5726 -245 5750 27
rect 6666 -245 6690 27
rect 321 -270 641 -246
rect 1212 -270 1532 -246
rect 2124 -270 2444 -246
rect 3016 -269 3336 -245
rect 3908 -269 4228 -245
rect 4807 -269 5127 -245
rect 5726 -269 6046 -245
rect 6666 -269 6986 -245
<< nwell >>
rect 878 265 6457 684
<< metal1 >>
rect 809 603 892 923
rect 1700 603 1783 923
rect 2612 603 2695 923
rect 3504 604 3587 924
rect 4396 604 4479 924
rect 5295 604 5378 924
rect 6214 604 6297 924
rect 7154 604 7237 924
rect 107 90 112 603
rect 948 528 1003 603
rect 107 62 155 90
rect 948 62 1031 528
rect 1860 90 1963 603
rect 2752 91 2855 604
rect 3644 91 3747 604
rect 4543 91 4646 604
rect 5462 91 5565 604
rect 6402 91 6505 604
rect 1860 62 1943 90
rect 2752 62 2835 91
rect 3644 63 3727 91
rect 4543 63 4626 91
rect 5462 63 5545 91
rect 6402 63 6485 91
rect 74 -161 155 62
rect 73 -376 155 -161
rect 810 2 1031 62
rect 1701 2 1943 62
rect 2613 3 2835 62
rect 810 -376 892 2
rect 1701 -376 1783 2
rect 2613 -376 2695 3
rect 3505 2 3727 63
rect 4397 3 4626 63
rect 5296 3 5545 63
rect 6215 3 6485 63
rect 3505 -375 3587 2
rect 4397 -375 4479 3
rect 5296 -377 5378 3
rect 6215 -376 6297 3
rect 7127 -160 7238 56
rect 7155 -376 7238 -160
use buffer  buffer_0 ~/Documents/Dersler/VLSI/vlsi_sky130b/design/mag/inv
timestamp 1734801607
transform -1 0 2350 0 1 312
box 1458 -582 2238 516
use buffer  buffer_1
timestamp 1734801607
transform -1 0 3241 0 1 312
box 1458 -582 2238 516
use buffer  buffer_2
timestamp 1734801607
transform -1 0 5937 0 1 313
box 1458 -582 2238 516
use buffer  buffer_3
timestamp 1734801607
transform -1 0 4153 0 1 312
box 1458 -582 2238 516
use buffer  buffer_4
timestamp 1734801607
transform -1 0 5045 0 1 313
box 1458 -582 2238 516
use buffer  buffer_5
timestamp 1734801607
transform -1 0 7755 0 1 313
box 1458 -582 2238 516
use buffer  buffer_6
timestamp 1734801607
transform -1 0 6836 0 1 313
box 1458 -582 2238 516
use buffer  buffer_7
timestamp 1734801607
transform -1 0 8695 0 1 313
box 1458 -582 2238 516
<< end >>
