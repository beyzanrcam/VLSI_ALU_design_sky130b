magic
tech sky130B
magscale 1 2
timestamp 1736620191
<< nwell >>
rect 356 684 1062 804
<< ndiff >>
rect 994 146 996 148
rect 626 54 1026 60
<< psubdiff >>
rect 626 28 1026 54
rect 626 -6 653 28
rect 988 -6 1026 28
rect 626 -17 1026 -6
<< nsubdiff >>
rect 396 761 1013 768
rect 396 714 420 761
rect 989 714 1013 761
rect 396 702 1013 714
<< psubdiffcont >>
rect 653 -6 988 28
<< nsubdiffcont >>
rect 420 714 989 761
<< poly >>
rect 453 387 520 408
rect 453 352 470 387
rect 504 352 520 387
rect 453 341 520 352
rect 742 387 809 408
rect 742 352 759 387
rect 793 352 809 387
rect 742 341 809 352
rect 453 146 496 341
rect 538 263 604 279
rect 538 228 554 263
rect 588 242 604 263
rect 588 228 714 242
rect 538 212 714 228
rect 453 130 604 146
rect 453 95 554 130
rect 588 95 604 130
rect 453 79 604 95
<< polycont >>
rect 470 352 504 387
rect 759 352 793 387
rect 554 228 588 263
rect 554 95 588 130
<< locali >>
rect 404 714 420 761
rect 989 714 1013 761
rect 453 352 470 387
rect 504 352 520 387
rect 742 381 759 387
rect 554 352 759 381
rect 793 352 809 387
rect 453 146 496 352
rect 554 347 809 352
rect 554 263 588 347
rect 554 212 588 228
rect 453 130 588 146
rect 453 95 554 130
rect 453 79 588 95
rect 626 -6 653 28
rect 988 -6 1026 28
<< viali >>
rect 420 714 989 761
rect 470 352 504 387
rect 759 352 793 387
rect 554 228 588 263
rect 653 -6 988 28
<< metal1 >>
rect 391 761 1025 768
rect 391 714 420 761
rect 989 714 1025 761
rect 391 555 1025 714
rect 485 434 1062 526
rect 356 387 520 405
rect 356 352 470 387
rect 504 352 520 387
rect 356 270 520 352
rect 548 387 808 406
rect 548 352 759 387
rect 793 352 808 387
rect 548 332 808 352
rect 548 263 598 332
rect 884 304 1062 434
rect 548 241 554 263
rect 356 228 554 241
rect 588 228 598 263
rect 626 252 1062 304
rect 356 105 598 228
rect 626 28 1026 105
rect 626 -6 653 28
rect 988 -6 1026 28
rect 626 -17 1026 -6
use nmos_2shared_W200-L015-F1  nmos_2shared_W200-L015-F1_0
timestamp 1736620191
transform 0 1 826 -1 0 179
box -125 -226 125 226
use pmos_p2-w321-L015-f3  pmos_p2-w321-L015-f3_0
timestamp 1736620191
transform 1 0 709 0 -1 541
box -353 -143 353 169
<< labels >>
rlabel metal1 356 341 356 341 7 A
port 1 w
rlabel metal1 356 173 356 173 7 B
port 2 w
rlabel metal1 826 54 826 54 5 VSS
port 3 s
rlabel metal1 709 684 709 684 1 VDD
port 4 n
rlabel metal1 1062 451 1062 451 3 Y
port 5 e
<< end >>
