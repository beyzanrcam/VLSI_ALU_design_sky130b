magic
tech sky130B
magscale 1 2
timestamp 1736181444
<< error_p >>
rect 0 0 376 418
rect 100 -126 300 -68
rect 100 -214 300 -156
<< nwell >>
rect 0 0 376 418
<< nmos >>
rect 100 -156 300 -126
<< pmos >>
rect 100 290 314 320
rect 100 194 314 224
rect 100 98 314 128
<< ndiff >>
rect 100 -80 300 -68
rect 100 -114 112 -80
rect 288 -114 300 -80
rect 100 -126 300 -114
rect 100 -168 300 -156
rect 100 -202 112 -168
rect 288 -202 300 -168
rect 100 -214 300 -202
<< pdiff >>
rect 100 370 314 382
rect 100 336 112 370
rect 302 336 314 370
rect 100 320 314 336
rect 100 274 314 290
rect 100 240 112 274
rect 306 240 314 274
rect 100 224 314 240
rect 100 178 314 194
rect 100 144 112 178
rect 302 144 314 178
rect 100 128 314 144
rect 100 82 314 98
rect 100 48 112 82
rect 306 48 314 82
rect 100 36 314 48
<< ndiffc >>
rect 112 -114 288 -80
rect 112 -202 288 -168
<< pdiffc >>
rect 112 336 302 370
rect 112 240 306 274
rect 112 144 302 178
rect 112 48 306 82
<< poly >>
rect 3 322 69 338
rect 3 96 19 322
rect 53 320 69 322
rect 53 290 100 320
rect 314 290 340 320
rect 53 224 69 290
rect 53 194 100 224
rect 314 194 340 224
rect 53 128 69 194
rect 53 98 100 128
rect 314 98 340 128
rect 53 96 69 98
rect 3 80 69 96
rect 3 -124 70 -108
rect 3 -158 19 -124
rect 53 -126 70 -124
rect 53 -156 100 -126
rect 300 -156 326 -126
rect 53 -158 70 -156
rect 3 -174 70 -158
<< polycont >>
rect 19 96 53 322
rect 19 -158 53 -124
<< locali >>
rect 3 322 53 339
rect 96 336 106 370
rect 302 336 318 370
rect 3 96 19 322
rect 96 240 112 274
rect 306 240 324 274
rect 96 144 106 178
rect 302 144 318 178
rect 3 -124 53 96
rect 96 48 112 82
rect 306 48 324 82
rect 96 -114 112 -80
rect 288 -114 304 -80
rect 3 -158 19 -124
rect 3 -174 53 -158
rect 96 -202 112 -168
rect 288 -202 304 -168
<< viali >>
rect 106 336 112 370
rect 112 336 185 370
rect 19 96 53 322
rect 229 240 306 274
rect 106 144 112 178
rect 112 144 185 178
rect 229 48 306 82
rect 112 -114 288 -80
rect 19 -158 53 -124
rect 112 -202 288 -168
<< metal1 >>
rect 96 370 318 418
rect 96 366 106 370
rect -14 322 69 338
rect -14 96 19 322
rect 53 96 69 322
rect 100 336 106 366
rect 185 366 318 370
rect 185 336 191 366
rect 100 178 191 336
rect 100 144 106 178
rect 185 144 191 178
rect 100 128 191 144
rect 223 274 376 338
rect 223 240 229 274
rect 306 240 376 274
rect -14 -124 69 96
rect 223 82 376 240
rect 100 48 229 82
rect 306 48 376 82
rect 100 -80 376 48
rect 100 -114 112 -80
rect 288 -114 376 -80
rect 100 -120 300 -114
rect -14 -158 19 -124
rect 53 -158 69 -124
rect -14 -175 69 -158
rect 100 -168 300 -161
rect 100 -202 112 -168
rect 288 -202 300 -168
rect 328 -175 376 -114
rect 100 -203 300 -202
rect 96 -250 304 -203
<< labels >>
rlabel metal1 376 -31 376 -31 3 Y
port 3 e
rlabel metal1 0 -31 0 -31 7 A
port 2 e
rlabel metal1 144 418 144 418 1 VDD
port 1 n
rlabel metal1 201 -250 201 -250 5 VSS
port 4 s
<< end >>
