magic
tech sky130B
magscale 1 2
timestamp 1735388107
<< error_s >>
rect -40 250 3696 668
rect 60 124 260 182
rect 540 124 740 182
rect 1000 124 1200 182
rect 1460 124 1660 182
rect 1940 124 2140 182
rect 2440 124 2640 182
rect 2920 124 3120 182
rect 3420 124 3620 182
rect 60 36 260 94
rect 540 36 740 94
rect 1000 36 1200 94
rect 1460 36 1660 94
rect 1940 36 2140 94
rect 2440 36 2640 94
rect 2920 36 3120 94
rect 3420 36 3620 94
<< nwell >>
rect -40 250 3696 668
<< metal1 >>
rect -40 588 29 883
rect 113 814 165 820
rect 113 616 165 762
rect 440 588 509 883
rect 594 818 646 824
rect 594 616 646 766
rect 900 588 969 883
rect 1059 820 1111 826
rect 1059 616 1111 768
rect 1360 588 1429 883
rect 1516 822 1568 828
rect 1516 616 1568 770
rect 1840 588 1909 883
rect 1985 825 2037 831
rect 1985 616 2037 773
rect 2340 588 2409 883
rect 2507 825 2559 831
rect 2507 616 2559 773
rect 2820 588 2889 883
rect 2990 825 3042 831
rect 2990 616 3042 773
rect 3320 588 3389 883
rect 3499 819 3551 825
rect 3499 616 3551 767
rect 122 -195 211 89
rect 122 -290 211 -284
rect 288 -501 336 87
rect 603 -201 692 89
rect 603 -296 692 -290
rect 768 -501 816 75
rect 1045 -201 1134 89
rect 1045 -296 1134 -290
rect 1228 -501 1276 75
rect 1497 -196 1586 89
rect 1497 -291 1586 -285
rect 1688 -501 1736 75
rect 1972 -195 2061 89
rect 1972 -290 2061 -284
rect 2168 -501 2216 75
rect 2479 -199 2568 89
rect 2479 -294 2568 -288
rect 2668 -501 2716 75
rect 2965 -200 3054 89
rect 2965 -295 3054 -289
rect 3148 -501 3196 75
rect 3458 -207 3547 89
rect 3458 -302 3547 -296
rect 3648 -501 3696 75
<< via1 >>
rect 113 762 165 814
rect 594 766 646 818
rect 1059 768 1111 820
rect 1516 770 1568 822
rect 1985 773 2037 825
rect 2507 773 2559 825
rect 2990 773 3042 825
rect 3499 767 3551 819
rect 122 -284 211 -195
rect 603 -290 692 -201
rect 1045 -290 1134 -201
rect 1497 -285 1586 -196
rect 1972 -284 2061 -195
rect 2479 -288 2568 -199
rect 2965 -289 3054 -200
rect 3458 -296 3547 -207
<< metal2 >>
rect 98 818 180 829
rect 98 758 109 818
rect 169 758 180 818
rect 98 747 180 758
rect 579 822 661 833
rect 579 762 590 822
rect 650 762 661 822
rect 579 751 661 762
rect 1044 824 1126 835
rect 1044 764 1055 824
rect 1115 764 1126 824
rect 1044 753 1126 764
rect 1501 826 1583 837
rect 1501 766 1512 826
rect 1572 766 1583 826
rect 1501 755 1583 766
rect 1970 829 2052 840
rect 1970 769 1981 829
rect 2041 769 2052 829
rect 1970 758 2052 769
rect 2492 829 2574 840
rect 2492 769 2503 829
rect 2563 769 2574 829
rect 2492 758 2574 769
rect 2975 829 3057 840
rect 2975 769 2986 829
rect 3046 769 3057 829
rect 2975 758 3057 769
rect 3484 823 3566 834
rect 3484 763 3495 823
rect 3555 763 3566 823
rect 3484 752 3566 763
rect 113 -284 122 -195
rect 211 -284 220 -195
rect 598 -201 697 -190
rect 1040 -201 1139 -190
rect 1492 -196 1591 -185
rect 1967 -195 2066 -184
rect 597 -290 603 -201
rect 692 -290 698 -201
rect 1039 -290 1045 -201
rect 1134 -290 1140 -201
rect 1491 -285 1497 -196
rect 1586 -285 1592 -196
rect 1966 -284 1972 -195
rect 2061 -284 2067 -195
rect 2474 -199 2573 -188
rect 598 -301 697 -290
rect 1040 -301 1139 -290
rect 1492 -296 1591 -285
rect 1967 -295 2066 -284
rect 2473 -288 2479 -199
rect 2568 -288 2574 -199
rect 2960 -200 3059 -189
rect 2474 -299 2573 -288
rect 2959 -289 2965 -200
rect 3054 -289 3060 -200
rect 3453 -207 3552 -196
rect 2960 -300 3059 -289
rect 3452 -296 3458 -207
rect 3547 -296 3553 -207
rect 3453 -307 3552 -296
<< via2 >>
rect 109 814 169 818
rect 109 762 113 814
rect 113 762 165 814
rect 165 762 169 814
rect 109 758 169 762
rect 590 818 650 822
rect 590 766 594 818
rect 594 766 646 818
rect 646 766 650 818
rect 590 762 650 766
rect 1055 820 1115 824
rect 1055 768 1059 820
rect 1059 768 1111 820
rect 1111 768 1115 820
rect 1055 764 1115 768
rect 1512 822 1572 826
rect 1512 770 1516 822
rect 1516 770 1568 822
rect 1568 770 1572 822
rect 1512 766 1572 770
rect 1981 825 2041 829
rect 1981 773 1985 825
rect 1985 773 2037 825
rect 2037 773 2041 825
rect 1981 769 2041 773
rect 2503 825 2563 829
rect 2503 773 2507 825
rect 2507 773 2559 825
rect 2559 773 2563 825
rect 2503 769 2563 773
rect 2986 825 3046 829
rect 2986 773 2990 825
rect 2990 773 3042 825
rect 3042 773 3046 825
rect 2986 769 3046 773
rect 3495 819 3555 823
rect 3495 767 3499 819
rect 3499 767 3551 819
rect 3551 767 3555 819
rect 3495 763 3555 767
rect 122 -284 211 -195
rect 603 -290 692 -201
rect 1045 -290 1134 -201
rect 1497 -285 1586 -196
rect 1972 -284 2061 -195
rect 2479 -288 2568 -199
rect 2965 -289 3054 -200
rect 3458 -296 3547 -207
<< metal3 >>
rect 63 823 227 859
rect 63 753 104 823
rect 174 753 227 823
rect 63 720 227 753
rect 563 827 674 842
rect 563 757 585 827
rect 655 757 674 827
rect 563 742 674 757
rect 1027 829 1142 849
rect 1027 759 1050 829
rect 1120 759 1142 829
rect 1027 738 1142 759
rect 1469 831 1624 854
rect 1469 761 1507 831
rect 1577 761 1624 831
rect 1469 737 1624 761
rect 1939 834 2090 864
rect 1939 764 1976 834
rect 2046 764 2090 834
rect 1939 737 2090 764
rect 2455 834 2624 864
rect 2455 764 2498 834
rect 2568 764 2624 834
rect 2455 737 2624 764
rect 2943 834 3098 864
rect 2943 764 2981 834
rect 3051 764 3098 834
rect 2943 737 3098 764
rect 3440 828 3606 862
rect 3440 758 3490 828
rect 3560 758 3606 828
rect 3440 737 3606 758
rect 92 -190 242 -168
rect 92 -289 117 -190
rect 216 -289 242 -190
rect 92 -315 242 -289
rect 592 -295 598 -196
rect 697 -295 703 -196
rect 1034 -295 1040 -196
rect 1139 -295 1145 -196
rect 1486 -290 1492 -191
rect 1591 -290 1597 -191
rect 1961 -289 1967 -190
rect 2066 -289 2072 -190
rect 2468 -293 2474 -194
rect 2573 -293 2579 -194
rect 2954 -294 2960 -195
rect 3059 -294 3065 -195
rect 3447 -301 3453 -202
rect 3552 -301 3558 -202
<< via3 >>
rect 104 818 174 823
rect 104 758 109 818
rect 109 758 169 818
rect 169 758 174 818
rect 104 753 174 758
rect 585 822 655 827
rect 585 762 590 822
rect 590 762 650 822
rect 650 762 655 822
rect 585 757 655 762
rect 1050 824 1120 829
rect 1050 764 1055 824
rect 1055 764 1115 824
rect 1115 764 1120 824
rect 1050 759 1120 764
rect 1507 826 1577 831
rect 1507 766 1512 826
rect 1512 766 1572 826
rect 1572 766 1577 826
rect 1507 761 1577 766
rect 1976 829 2046 834
rect 1976 769 1981 829
rect 1981 769 2041 829
rect 2041 769 2046 829
rect 1976 764 2046 769
rect 2498 829 2568 834
rect 2498 769 2503 829
rect 2503 769 2563 829
rect 2563 769 2568 829
rect 2498 764 2568 769
rect 2981 829 3051 834
rect 2981 769 2986 829
rect 2986 769 3046 829
rect 3046 769 3051 829
rect 2981 764 3051 769
rect 3490 823 3560 828
rect 3490 763 3495 823
rect 3495 763 3555 823
rect 3555 763 3560 823
rect 3490 758 3560 763
rect 117 -195 216 -190
rect 117 -284 122 -195
rect 122 -284 211 -195
rect 211 -284 216 -195
rect 117 -289 216 -284
rect 598 -201 697 -196
rect 598 -290 603 -201
rect 603 -290 692 -201
rect 692 -290 697 -201
rect 598 -295 697 -290
rect 1040 -201 1139 -196
rect 1040 -290 1045 -201
rect 1045 -290 1134 -201
rect 1134 -290 1139 -201
rect 1040 -295 1139 -290
rect 1492 -196 1591 -191
rect 1492 -285 1497 -196
rect 1497 -285 1586 -196
rect 1586 -285 1591 -196
rect 1492 -290 1591 -285
rect 1967 -195 2066 -190
rect 1967 -284 1972 -195
rect 1972 -284 2061 -195
rect 2061 -284 2066 -195
rect 1967 -289 2066 -284
rect 2474 -199 2573 -194
rect 2474 -288 2479 -199
rect 2479 -288 2568 -199
rect 2568 -288 2573 -199
rect 2474 -293 2573 -288
rect 2960 -200 3059 -195
rect 2960 -289 2965 -200
rect 2965 -289 3054 -200
rect 3054 -289 3059 -200
rect 2960 -294 3059 -289
rect 3453 -207 3552 -202
rect 3453 -296 3458 -207
rect 3458 -296 3547 -207
rect 3547 -296 3552 -207
rect 3453 -301 3552 -296
<< metal4 >>
rect 63 834 3606 883
rect 63 831 1976 834
rect 63 829 1507 831
rect 63 827 1050 829
rect 63 823 585 827
rect 63 753 104 823
rect 174 757 585 823
rect 655 759 1050 827
rect 1120 761 1507 829
rect 1577 764 1976 831
rect 2046 764 2498 834
rect 2568 764 2981 834
rect 3051 828 3606 834
rect 3051 764 3490 828
rect 1577 761 3490 764
rect 1120 759 3490 761
rect 655 758 3490 759
rect 3560 758 3606 828
rect 655 757 3606 758
rect 174 753 3606 757
rect 63 737 3606 753
rect 63 720 3604 737
<< via4 >>
rect 7 -190 327 -79
rect 7 -289 117 -190
rect 117 -289 216 -190
rect 216 -289 327 -190
rect 7 -399 327 -289
rect 488 -196 808 -85
rect 488 -295 598 -196
rect 598 -295 697 -196
rect 697 -295 808 -196
rect 488 -405 808 -295
rect 930 -196 1250 -85
rect 930 -295 1040 -196
rect 1040 -295 1139 -196
rect 1139 -295 1250 -196
rect 930 -405 1250 -295
rect 1382 -191 1702 -80
rect 1382 -290 1492 -191
rect 1492 -290 1591 -191
rect 1591 -290 1702 -191
rect 1382 -400 1702 -290
rect 1857 -190 2177 -79
rect 1857 -289 1967 -190
rect 1967 -289 2066 -190
rect 2066 -289 2177 -190
rect 1857 -399 2177 -289
rect 2364 -194 2684 -83
rect 2364 -293 2474 -194
rect 2474 -293 2573 -194
rect 2573 -293 2684 -194
rect 2364 -403 2684 -293
rect 2850 -195 3170 -84
rect 2850 -294 2960 -195
rect 2960 -294 3059 -195
rect 3059 -294 3170 -195
rect 2850 -404 3170 -294
rect 3343 -202 3663 -91
rect 3343 -301 3453 -202
rect 3453 -301 3552 -202
rect 3552 -301 3663 -202
rect 3343 -411 3663 -301
<< metal5 >>
rect -110 -24 435 -22
rect -110 -79 3853 -24
rect -110 -399 7 -79
rect 327 -80 1857 -79
rect 327 -85 1382 -80
rect 327 -399 488 -85
rect -110 -405 488 -399
rect 808 -405 930 -85
rect 1250 -400 1382 -85
rect 1702 -399 1857 -80
rect 2177 -83 3853 -79
rect 2177 -399 2364 -83
rect 1702 -400 2364 -399
rect 1250 -403 2364 -400
rect 2684 -84 3853 -83
rect 2684 -403 2850 -84
rect 1250 -404 2850 -403
rect 3170 -91 3853 -84
rect 3170 -404 3343 -91
rect 1250 -405 3343 -404
rect -110 -411 3343 -405
rect 3663 -411 3853 -91
rect -110 -501 3853 -411
use inv  inv_0 ~/Desktop/vlsi_sky130b/design/mag/inv
timestamp 1735380995
transform 1 0 3320 0 1 250
box 0 -250 376 418
use inv  inv_1
timestamp 1735380995
transform 1 0 -40 0 1 250
box 0 -250 376 418
use inv  inv_2
timestamp 1735380995
transform 1 0 440 0 1 250
box 0 -250 376 418
use inv  inv_3
timestamp 1735380995
transform 1 0 900 0 1 250
box 0 -250 376 418
use inv  inv_4
timestamp 1735380995
transform 1 0 1360 0 1 250
box 0 -250 376 418
use inv  inv_5
timestamp 1735380995
transform 1 0 1840 0 1 250
box 0 -250 376 418
use inv  inv_6
timestamp 1735380995
transform 1 0 2340 0 1 250
box 0 -250 376 418
use inv  inv_7
timestamp 1735380995
transform 1 0 2820 0 1 250
box 0 -250 376 418
<< labels >>
rlabel metal1 -32 831 19 878 5 A7
port 1 s
rlabel metal1 449 831 500 878 5 A6
port 2 s
rlabel metal1 908 828 959 875 5 A5
port 3 s
rlabel metal1 1368 829 1419 876 5 A4
port 4 s
rlabel metal1 1849 830 1900 877 5 A3
port 5 s
rlabel metal1 2348 831 2399 878 5 A2
port 6 s
rlabel metal1 2829 830 2880 877 5 A1
port 7 s
rlabel metal1 3329 828 3380 875 5 A0
port 8 s
rlabel metal1 3652 -495 3687 -462 1 S0
port 9 n
rlabel metal1 3153 -488 3188 -455 1 S1
port 10 n
rlabel metal1 2674 -495 2709 -462 1 S2
port 11 n
rlabel metal1 2174 -496 2209 -463 1 S3
port 12 n
rlabel metal1 1694 -496 1729 -463 1 S4
port 13 n
rlabel metal1 1235 -496 1270 -463 1 S5
port 14 n
rlabel metal1 774 -496 809 -463 1 S6
port 15 n
rlabel metal1 294 -495 329 -462 1 S7
port 16 n
<< end >>
