** sch_path: /home/ubuntu/Desktop/examples/xschem/five_T_OTA_noise_TB.sch
**.subckt five_T_OTA_noise_TB
x1 OUT net2 net1 IBIAS GND VDD five_T_OTA
V1 VDD GND 1.8
I0 VDD IBIAS 50u
V2 net1 net2 0 AC 1
V3 net1 GND 0.9
C1 OUT GND 1p m=1
.save  v(out)
**** begin user architecture code



.control

save all

op
write five_T_OTA_noise_TB.raw

noise v(out) v2 dec 10 1e3 1e9
set appendwrite
write five_T_OTA_noise_TB.raw

plot noise1.v(onoise_spectrum)
print noise2.v(onoise_total)

.endc



** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  five_T_OTA.sym # of pins=6
** sym_path: /home/ubuntu/Desktop/examples/xschem/five_T_OTA.sym
** sch_path: /home/ubuntu/Desktop/examples/xschem/five_T_OTA.sch
.subckt five_T_OTA  OUT MINUS PLUS IBIAS VSS VDD
*.iopin VDD
*.iopin VSS
*.iopin MINUS
*.iopin PLUS
*.iopin OUT
*.iopin IBIAS
XM2 IBIAS IBIAS VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 IBIAS VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
.save  v(ibias)
.save  v(out)
.save  v(net2)
.save  v(net1)
XM4 net2 PLUS net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.3 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM5 OUT MINUS net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.3 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM3 net2 net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.7 W=2.3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM6 OUT net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.7 W=2.3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
.ends

.GLOBAL GND
.end
