** sch_path: /home/efeler_gibi/Documents/vlsi/vlsi_sky130b/design/xschem/From Layout/NAND/nand_TB.sch
**.subckt nand_TB OUTPUT VDD VSS OUTPUT2
*.opin OUTPUT
*.iopin VDD
*.iopin VSS
*.opin OUTPUT2
V1 VDD GND 1.2
V2 VSS GND 0
V4 INPUT GND pulse(0,1.2,0.01u,0 ,0,0.01u,0.02u)
x1 INPUT INPUT INPUT INPUT VSS VDD OUTPUT nand4
x2 OUTPUT VSS VDD net1 inv
x3 OUTPUT VSS VDD net2 inv
x4 OUTPUT VSS VDD net3 inv
x5 OUTPUT VSS VDD net4 inv
x6 OUTPUT2 VSS VDD net5 inv
x7 OUTPUT2 VSS VDD net6 inv
x8 OUTPUT2 VSS VDD net7 inv
x9 OUTPUT2 VSS VDD net8 inv
x10 INPUT VSS VDD INPUT2 inv
x11 INPUT2 GND GND GND VSS VDD OUTPUT2 nand4
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice tt_mm




.include '../mag/NAND/NAND4/nand4_x.spice'v
.incluce '../mag/inv/inv_x.spice'
.control
set color0 = white

save all
tran 0.001n 0.03u
plot INPUT OUTPUT title 'a'
plot INPUT2 OUTPUT2 title 'a'


meas tran t_input when V(INPUT)=0.6 RISE=1
meas tran t_output when V(OUTPUT)=0.6 FALL=1
let tpdr = (t_output - t_input) * 1e9
echo tpdr (ns) is:
print tpdr
meas tran t_input when V(INPUT)=0.6 FALL=1
meas tran t_output when V(OUTPUT)=0.6 RISE=1
let tpdf = (t_output - t_input) * 1e9
echo tpdf (ns) is:
print tpdf
let tpd = (tpdf + tpdr)/2
echo tpd (ns) is:
print tpd



meas tran t_input when V(INPUT2)=0.6 RISE=1
meas tran t_output when V(OUTPUT2)=0.6 FALL=1
let tpdr = (t_output - t_input) * 1e9
echo tpdr (ns) is:
print tpdr
meas tran t_input when V(INPUT2)=0.6 FALL=1
meas tran t_output when V(OUTPUT2)=0.6 RISE=1
let tpdf = (t_output - t_input) * 1e9
echo tpdf (ns) is:
print tpdf
let tpd = (tpdf + tpdr)/2
echo tpd (ns) is:
print tpd
.endc


**** end user architecture code
**.ends

* expanding   symbol:  INV/inv.sym # of pins=2
** sym_path: /home/efeler_gibi/Documents/vlsi/vlsi_sky130b/design/xschem/INV/inv.sym
** sch_path: /home/efeler_gibi/Documents/vlsi/vlsi_sky130b/design/xschem/INV/inv.sch
.subckt inv A VSS VDD Y
*.ipin A
*.opin Y
XM1 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.21 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
