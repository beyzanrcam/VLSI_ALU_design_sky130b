magic
tech sky130B
magscale 1 2
timestamp 1736450894
<< nwell >>
rect -1843 2757 -550 3243
rect 493 2013 3416 2590
<< metal1 >>
rect -1841 2505 -1772 2751
rect -1842 2446 -1772 2505
rect -1499 2530 -1430 2751
rect -1499 2440 -1430 2461
rect -1402 1988 -1333 2751
rect -1059 2528 -990 2590
rect -1059 2446 -990 2459
rect -962 2446 -893 2587
rect -619 2537 -550 2597
rect -620 2527 -550 2537
rect -551 2506 -550 2527
rect -620 2446 -551 2458
rect -294 2077 -242 2083
rect -294 2019 -242 2025
rect -1402 1922 -232 1988
rect -1402 1829 -1333 1922
<< via1 >>
rect -1499 2461 -1430 2530
rect -1059 2459 -990 2528
rect -620 2458 -551 2527
rect -294 2025 -242 2077
rect 669 2024 722 2076
rect 1602 2025 1655 2077
rect 2533 2025 2586 2077
rect 1600 1927 1652 1979
rect 2535 1927 2587 1979
<< metal2 >>
rect -1499 2641 -287 2710
rect -1499 2530 -1430 2641
rect -1499 2455 -1430 2461
rect -1065 2459 -1059 2528
rect -990 2459 -984 2528
rect -1059 2363 -990 2459
rect -626 2458 -620 2527
rect -551 2458 -545 2527
rect -620 2315 -551 2458
rect -1059 2295 -990 2304
rect -356 2086 -287 2641
rect -356 2077 2740 2086
rect -356 2025 -294 2077
rect -242 2076 1602 2077
rect -242 2025 669 2076
rect -356 2024 669 2025
rect 722 2025 1602 2076
rect 1655 2025 2533 2077
rect 2586 2025 2740 2077
rect 722 2024 2740 2025
rect -356 2017 2740 2024
rect 2529 1983 2600 1985
rect 1589 1925 1598 1981
rect 1654 1925 1663 1981
rect 2523 1927 2535 1983
rect 2591 1927 2600 1983
rect 2529 1921 2593 1927
<< via2 >>
rect -1059 2304 -990 2363
rect 1598 1979 1654 1981
rect 1598 1927 1600 1979
rect 1600 1927 1652 1979
rect 1652 1927 1654 1979
rect 1598 1925 1654 1927
rect 2535 1979 2591 1983
rect 2535 1927 2587 1979
rect 2587 1927 2591 1979
<< metal3 >>
rect -1064 2363 -985 2368
rect -1064 2304 -1059 2363
rect -990 2304 -985 2363
rect -1064 2299 -985 2304
rect -1058 1990 -989 2299
rect -1058 1983 2602 1990
rect -1058 1981 2535 1983
rect -1058 1925 1598 1981
rect 1654 1927 2535 1981
rect 2591 1927 2602 1983
rect 1654 1925 2602 1927
rect -1058 1920 2602 1925
use inv  inv_1 ~/Documents/vlsi/vlsi_sky130b/design/mag/inv
timestamp 1735843251
transform 1 0 -1402 0 1 2757
box 0 -311 412 486
use inv  inv_2
timestamp 1735843251
transform 1 0 -962 0 1 2757
box 0 -311 412 486
use inv  inv_3
timestamp 1735843251
transform 1 0 -1842 0 1 2757
box 0 -311 412 486
use NAND4F  NAND4F_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NAND/NAND4
timestamp 1736096163
transform 1 0 2507 0 1 2017
box 10 -1175 909 571
use NAND4F  NAND4F_1
timestamp 1736096163
transform 1 0 -308 0 1 2017
box 10 -1175 909 571
use NAND4F  NAND4F_2
timestamp 1736096163
transform 1 0 640 0 1 2017
box 10 -1175 909 571
use NAND4F  NAND4F_3
timestamp 1736096163
transform 1 0 1576 0 1 2017
box 10 -1175 909 571
<< end >>
