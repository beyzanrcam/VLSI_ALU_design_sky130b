magic
tech sky130A
magscale 1 2
timestamp 1733250542
<< nwell >>
rect 2 6 1284 922
<< nmos >>
rect 100 -657 130 -527
rect 196 -657 226 -527
rect 292 -657 322 -527
rect 388 -657 418 -527
rect 484 -657 514 -527
rect 580 -657 610 -527
rect 676 -657 706 -527
rect 772 -657 802 -527
rect 868 -657 898 -527
rect 964 -657 994 -527
rect 1060 -657 1090 -527
rect 1156 -657 1186 -527
<< pmos >>
rect 100 129 130 679
rect 196 129 226 679
rect 292 129 322 679
rect 388 129 418 679
rect 484 129 514 679
rect 580 129 610 679
rect 676 129 706 679
rect 772 129 802 679
rect 868 129 898 679
rect 964 129 994 679
rect 1060 129 1090 679
rect 1156 129 1186 679
<< ndiff >>
rect 38 -539 100 -527
rect 38 -645 50 -539
rect 84 -645 100 -539
rect 38 -657 100 -645
rect 130 -539 196 -527
rect 130 -645 146 -539
rect 180 -645 196 -539
rect 130 -657 196 -645
rect 226 -539 292 -527
rect 226 -645 242 -539
rect 276 -645 292 -539
rect 226 -657 292 -645
rect 322 -539 388 -527
rect 322 -645 338 -539
rect 372 -645 388 -539
rect 322 -657 388 -645
rect 418 -539 484 -527
rect 418 -645 434 -539
rect 468 -645 484 -539
rect 418 -657 484 -645
rect 514 -539 580 -527
rect 514 -645 530 -539
rect 564 -645 580 -539
rect 514 -657 580 -645
rect 610 -539 676 -527
rect 610 -645 626 -539
rect 660 -645 676 -539
rect 610 -657 676 -645
rect 706 -539 772 -527
rect 706 -645 722 -539
rect 756 -645 772 -539
rect 706 -657 772 -645
rect 802 -539 868 -527
rect 802 -645 818 -539
rect 852 -645 868 -539
rect 802 -657 868 -645
rect 898 -539 964 -527
rect 898 -645 914 -539
rect 948 -645 964 -539
rect 898 -657 964 -645
rect 994 -539 1060 -527
rect 994 -645 1010 -539
rect 1044 -645 1060 -539
rect 994 -657 1060 -645
rect 1090 -539 1156 -527
rect 1090 -645 1106 -539
rect 1140 -645 1156 -539
rect 1090 -657 1156 -645
rect 1186 -539 1248 -527
rect 1186 -645 1202 -539
rect 1236 -645 1248 -539
rect 1186 -657 1248 -645
<< pdiff >>
rect 38 667 100 679
rect 38 141 50 667
rect 84 141 100 667
rect 38 129 100 141
rect 130 667 196 679
rect 130 141 146 667
rect 180 141 196 667
rect 130 129 196 141
rect 226 667 292 679
rect 226 141 242 667
rect 276 141 292 667
rect 226 129 292 141
rect 322 667 388 679
rect 322 141 338 667
rect 372 141 388 667
rect 322 129 388 141
rect 418 667 484 679
rect 418 141 434 667
rect 468 141 484 667
rect 418 129 484 141
rect 514 667 580 679
rect 514 141 530 667
rect 564 141 580 667
rect 514 129 580 141
rect 610 667 676 679
rect 610 141 626 667
rect 660 141 676 667
rect 610 129 676 141
rect 706 667 772 679
rect 706 141 722 667
rect 756 141 772 667
rect 706 129 772 141
rect 802 667 868 679
rect 802 141 818 667
rect 852 141 868 667
rect 802 129 868 141
rect 898 667 964 679
rect 898 141 914 667
rect 948 141 964 667
rect 898 129 964 141
rect 994 667 1060 679
rect 994 141 1010 667
rect 1044 141 1060 667
rect 994 129 1060 141
rect 1090 667 1156 679
rect 1090 141 1106 667
rect 1140 141 1156 667
rect 1090 129 1156 141
rect 1186 667 1248 679
rect 1186 141 1202 667
rect 1236 141 1248 667
rect 1186 129 1248 141
<< ndiffc >>
rect 50 -645 84 -539
rect 146 -645 180 -539
rect 242 -645 276 -539
rect 338 -645 372 -539
rect 434 -645 468 -539
rect 530 -645 564 -539
rect 626 -645 660 -539
rect 722 -645 756 -539
rect 818 -645 852 -539
rect 914 -645 948 -539
rect 1010 -645 1044 -539
rect 1106 -645 1140 -539
rect 1202 -645 1236 -539
<< pdiffc >>
rect 50 141 84 667
rect 146 141 180 667
rect 242 141 276 667
rect 338 141 372 667
rect 434 141 468 667
rect 530 141 564 667
rect 626 141 660 667
rect 722 141 756 667
rect 818 141 852 667
rect 914 141 948 667
rect 1010 141 1044 667
rect 1106 141 1140 667
rect 1202 141 1236 667
<< psubdiff >>
rect 38 -777 1248 -761
rect 38 -843 100 -777
rect 1186 -843 1248 -777
rect 38 -858 1248 -843
<< nsubdiff >>
rect 38 869 1248 886
rect 38 803 100 869
rect 1186 803 1248 869
rect 38 787 1248 803
<< psubdiffcont >>
rect 100 -843 1186 -777
<< nsubdiffcont >>
rect 100 803 1186 869
<< poly >>
rect 100 679 130 710
rect 196 679 226 710
rect 292 679 322 710
rect 388 679 418 710
rect 484 679 514 710
rect 580 679 610 710
rect 676 679 706 710
rect 772 679 802 710
rect 868 679 898 710
rect 964 679 994 710
rect 1060 679 1090 710
rect 1156 679 1186 710
rect 100 98 130 129
rect 196 98 226 129
rect 292 98 322 129
rect 100 74 322 98
rect 100 40 130 74
rect 292 40 322 74
rect 100 16 322 40
rect 388 98 418 129
rect 484 98 514 129
rect 580 98 610 129
rect 388 74 610 98
rect 388 40 418 74
rect 580 40 610 74
rect 388 16 610 40
rect 676 98 706 129
rect 772 98 802 129
rect 868 98 898 129
rect 676 74 898 98
rect 676 40 706 74
rect 868 40 898 74
rect 676 16 898 40
rect 964 98 994 129
rect 1060 98 1090 129
rect 1156 98 1186 129
rect 964 74 1186 98
rect 964 40 994 74
rect 1156 40 1186 74
rect 964 16 1186 40
rect 100 -440 322 -422
rect 100 -474 130 -440
rect 292 -474 322 -440
rect 100 -505 322 -474
rect 100 -527 130 -505
rect 196 -527 226 -505
rect 292 -527 322 -505
rect 388 -440 610 -422
rect 388 -474 418 -440
rect 580 -474 610 -440
rect 388 -505 610 -474
rect 388 -527 418 -505
rect 484 -527 514 -505
rect 580 -527 610 -505
rect 676 -440 898 -422
rect 676 -474 706 -440
rect 868 -474 898 -440
rect 676 -505 898 -474
rect 676 -527 706 -505
rect 772 -527 802 -505
rect 868 -527 898 -505
rect 964 -440 1186 -422
rect 964 -474 994 -440
rect 1156 -474 1186 -440
rect 964 -505 1186 -474
rect 964 -527 994 -505
rect 1060 -527 1090 -505
rect 1156 -527 1186 -505
rect 100 -683 130 -657
rect 196 -683 226 -657
rect 292 -683 322 -657
rect 388 -683 418 -657
rect 484 -683 514 -657
rect 580 -683 610 -657
rect 676 -683 706 -657
rect 772 -683 802 -657
rect 868 -683 898 -657
rect 964 -683 994 -657
rect 1060 -683 1090 -657
rect 1156 -683 1186 -657
<< polycont >>
rect 130 40 292 74
rect 418 40 580 74
rect 706 40 868 74
rect 994 40 1156 74
rect 130 -474 292 -440
rect 418 -474 580 -440
rect 706 -474 868 -440
rect 994 -474 1156 -440
<< locali >>
rect 38 869 1248 886
rect 38 803 100 869
rect 1186 803 1248 869
rect 38 787 1248 803
rect 50 667 84 683
rect 50 125 84 141
rect 146 667 180 683
rect 146 125 180 141
rect 242 667 276 683
rect 242 125 276 141
rect 338 667 372 683
rect 338 125 372 141
rect 434 667 468 683
rect 434 125 468 141
rect 530 667 564 683
rect 530 125 564 141
rect 626 667 660 683
rect 626 125 660 141
rect 722 667 756 683
rect 722 125 756 141
rect 818 667 852 683
rect 818 125 852 141
rect 914 667 948 683
rect 914 125 948 141
rect 1010 667 1044 683
rect 1010 125 1044 141
rect 1106 667 1140 683
rect 1106 125 1140 141
rect 1202 667 1236 683
rect 1202 125 1236 141
rect 114 74 308 90
rect 114 55 130 74
rect 1 40 130 55
rect 292 40 308 74
rect 1 21 308 40
rect 402 74 596 90
rect 402 40 418 74
rect 580 40 596 74
rect 402 -13 596 40
rect 1 -47 596 -13
rect 690 74 884 90
rect 690 40 706 74
rect 868 40 884 74
rect 690 -81 884 40
rect 1 -115 884 -81
rect 978 74 1172 90
rect 978 40 994 74
rect 1156 40 1172 74
rect 978 -149 1172 40
rect 1 -183 1172 -149
rect 1 -251 1172 -217
rect 1 -319 884 -285
rect 1 -387 596 -353
rect 1 -440 308 -421
rect 1 -455 130 -440
rect 114 -474 130 -455
rect 292 -474 308 -440
rect 114 -488 308 -474
rect 402 -440 596 -387
rect 402 -474 418 -440
rect 580 -474 596 -440
rect 402 -488 596 -474
rect 690 -440 884 -319
rect 690 -474 706 -440
rect 868 -474 884 -440
rect 690 -488 884 -474
rect 978 -440 1172 -251
rect 978 -474 994 -440
rect 1156 -474 1172 -440
rect 978 -488 1172 -474
rect 50 -661 84 -645
rect 146 -539 180 -523
rect 242 -661 276 -645
rect 338 -539 372 -523
rect 434 -661 468 -645
rect 530 -539 564 -523
rect 626 -661 660 -645
rect 722 -539 756 -523
rect 818 -661 852 -645
rect 914 -539 948 -523
rect 1010 -661 1044 -645
rect 1106 -539 1140 -523
rect 1202 -661 1236 -645
rect 38 -777 1248 -761
rect 38 -843 100 -777
rect 1186 -843 1248 -777
rect 38 -858 1248 -843
<< viali >>
rect 100 803 1186 869
rect 50 559 84 661
rect 50 164 84 266
rect 146 351 180 475
rect 242 559 276 661
rect 242 164 276 266
rect 338 351 372 475
rect 434 557 468 659
rect 434 158 468 260
rect 530 351 564 475
rect 626 556 660 658
rect 626 141 660 243
rect 722 351 756 475
rect 818 556 852 658
rect 818 158 852 260
rect 914 351 948 475
rect 1010 556 1044 658
rect 1010 165 1044 267
rect 1106 350 1140 474
rect 1202 556 1236 658
rect 1202 165 1236 267
rect 50 -539 84 -523
rect 50 -557 84 -539
rect 146 -645 180 -627
rect 146 -661 180 -645
rect 242 -539 276 -523
rect 242 -557 276 -539
rect 338 -645 372 -627
rect 338 -661 372 -645
rect 434 -539 468 -523
rect 434 -557 468 -539
rect 530 -645 564 -628
rect 530 -662 564 -645
rect 626 -539 660 -523
rect 626 -557 660 -539
rect 722 -645 756 -627
rect 722 -661 756 -645
rect 818 -539 852 -523
rect 818 -557 852 -539
rect 914 -645 948 -627
rect 914 -661 948 -645
rect 1010 -539 1044 -523
rect 1010 -557 1044 -539
rect 1106 -645 1140 -627
rect 1106 -661 1140 -645
rect 1202 -539 1236 -523
rect 1202 -557 1236 -539
rect 100 -843 1186 -777
<< metal1 >>
rect 2 869 1284 886
rect 2 803 100 869
rect 1186 803 1284 869
rect 2 787 1284 803
rect 38 661 292 787
rect 38 559 50 661
rect 84 559 242 661
rect 276 559 292 661
rect 38 538 292 559
rect 418 659 868 685
rect 418 557 434 659
rect 468 658 868 659
rect 468 557 626 658
rect 418 556 626 557
rect 660 556 818 658
rect 852 556 868 658
rect 418 538 868 556
rect 994 658 1248 787
rect 994 556 1010 658
rect 1044 556 1202 658
rect 1236 556 1248 658
rect 994 538 1248 556
rect 130 475 1156 500
rect 130 351 146 475
rect 180 351 338 475
rect 372 351 530 475
rect 564 351 722 475
rect 756 351 914 475
rect 948 474 1156 475
rect 948 351 1106 474
rect 130 350 1106 351
rect 1140 350 1156 474
rect 130 321 1156 350
rect 38 266 292 288
rect 38 164 50 266
rect 84 164 242 266
rect 276 164 292 266
rect 38 141 292 164
rect 418 260 867 277
rect 418 158 434 260
rect 468 243 818 260
rect 468 158 626 243
rect 418 141 626 158
rect 660 158 818 243
rect 852 158 867 260
rect 660 141 867 158
rect 994 267 1249 288
rect 994 165 1010 267
rect 1044 165 1202 267
rect 1236 165 1249 267
rect 994 141 1249 165
rect 610 -148 676 141
rect 610 -251 1284 -148
rect 610 -505 676 -251
rect 38 -523 292 -505
rect 38 -557 50 -523
rect 84 -557 242 -523
rect 276 -557 292 -523
rect 38 -573 292 -557
rect 418 -523 868 -505
rect 418 -557 434 -523
rect 468 -557 626 -523
rect 660 -557 818 -523
rect 852 -557 868 -523
rect 418 -573 868 -557
rect 994 -523 1248 -505
rect 994 -557 1010 -523
rect 1044 -557 1202 -523
rect 1236 -557 1248 -523
rect 994 -573 1248 -557
rect 38 -761 100 -573
rect 130 -627 580 -615
rect 130 -661 146 -627
rect 180 -661 338 -627
rect 372 -628 580 -627
rect 372 -661 530 -628
rect 130 -662 530 -661
rect 564 -662 580 -628
rect 130 -683 580 -662
rect 706 -627 1156 -615
rect 706 -661 722 -627
rect 756 -661 914 -627
rect 948 -661 1106 -627
rect 1140 -661 1156 -627
rect 706 -683 1156 -661
rect 1186 -761 1248 -573
rect 2 -777 1284 -761
rect 2 -843 100 -777
rect 1186 -843 1284 -777
rect 2 -858 1284 -843
<< labels >>
flabel metal1 602 818 756 870 1 FreeSerif 80 0 0 0 VDD
port 1 n
flabel metal1 592 -835 746 -783 1 FreeSerif 80 0 0 0 VSS
port 2 n
flabel locali 13 -243 34 -223 1 FreeSerif 80 0 0 0 N1
port 3 n
flabel locali 12 -311 33 -291 1 FreeSerif 80 0 0 0 N2
port 4 n
flabel locali 12 -380 33 -360 1 FreeSerif 80 0 0 0 N3
port 5 n
flabel locali 12 -448 33 -428 1 FreeSerif 80 0 0 0 N4
port 6 n
flabel locali 13 -177 34 -157 1 FreeSerif 80 0 0 0 P1
port 7 n
flabel locali 13 -108 34 -88 1 FreeSerif 80 0 0 0 P2
port 8 n
flabel locali 13 -39 34 -19 1 FreeSerif 80 0 0 0 P3
port 9 n
flabel locali 13 28 34 48 1 FreeSerif 80 0 0 0 P4
port 10 n
flabel metal1 1183 -228 1257 -164 1 FreeSerif 80 0 0 0 OUT
port 11 n
<< end >>
