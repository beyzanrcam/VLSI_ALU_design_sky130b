magic
tech sky130B
magscale 1 2
timestamp 1736019943
<< nwell >>
rect -602 1489 -492 1966
rect -602 1467 -482 1489
rect -602 1047 -456 1467
rect -602 1023 -461 1047
rect -602 991 -492 1023
<< psubdiff >>
rect -72 307 370 375
rect -72 194 -8 307
rect 322 194 370 307
rect -72 118 370 194
<< nsubdiff >>
rect -566 1413 -456 1903
rect -566 1059 -516 1413
rect -482 1059 -456 1413
rect -566 1047 -456 1059
<< psubdiffcont >>
rect -8 194 322 307
<< nsubdiffcont >>
rect -516 1059 -482 1413
<< poly >>
rect -238 1000 -172 1016
rect -238 966 -222 1000
rect -188 966 -172 1000
rect -238 950 -172 966
rect 50 1000 116 1016
rect 50 966 66 1000
rect 100 966 116 1000
rect 50 950 116 966
rect -202 674 -172 950
rect -202 644 20 674
rect 86 650 116 950
rect 182 1000 248 1016
rect 182 966 198 1000
rect 232 966 248 1000
rect 182 950 248 966
rect 182 650 212 950
rect 470 734 500 991
rect 434 718 500 734
rect 434 697 450 718
rect 278 684 450 697
rect 484 684 500 718
rect 278 667 500 684
rect 278 655 308 667
<< polycont >>
rect -222 966 -188 1000
rect 66 966 100 1000
rect 198 966 232 1000
rect 450 684 484 718
<< locali >>
rect -516 1413 -482 1429
rect -516 1043 -482 1059
rect -238 966 -222 1000
rect -188 966 -172 1000
rect 50 966 66 1000
rect 100 966 116 1000
rect 182 966 198 1000
rect 232 966 248 1000
rect 434 684 450 718
rect 484 684 500 718
rect -60 375 -26 425
rect 132 375 166 425
rect 324 375 358 425
rect -60 307 358 375
rect -60 194 -8 307
rect 322 194 358 307
rect -60 146 358 194
<< viali >>
rect -516 1059 -482 1413
rect -222 966 -188 1000
rect 66 966 100 1000
rect 198 966 232 1000
rect 450 684 484 718
rect -8 194 322 307
<< metal1 >>
rect -308 1523 -162 1903
rect -116 1523 30 1903
rect 268 1523 606 1903
rect -531 1413 -450 1425
rect -531 1059 -516 1413
rect -482 1059 -450 1413
rect -531 1047 -450 1059
rect -404 1047 -258 1425
rect -20 1047 318 1425
rect 556 1047 702 1425
rect 611 1016 748 1047
rect -602 1000 -172 1016
rect -602 966 -222 1000
rect -188 966 -172 1000
rect -602 950 -172 966
rect -141 1000 116 1016
rect -141 966 66 1000
rect 100 966 116 1000
rect -141 950 116 966
rect 182 1000 248 1016
rect 182 966 198 1000
rect 232 966 248 1000
rect -141 922 -75 950
rect 182 922 248 966
rect -602 856 -75 922
rect -42 856 248 922
rect 611 950 790 1016
rect -42 828 25 856
rect -602 762 25 828
rect -602 718 500 734
rect -602 684 450 718
rect 484 684 500 718
rect -602 668 500 684
rect 611 629 748 950
rect 76 429 748 629
rect -20 307 334 317
rect -20 194 -8 307
rect 322 194 334 307
rect -20 187 334 194
use sky130_fd_pr__nfet_01v8_S9NJ5Q  sky130_fd_pr__nfet_01v8_S9NJ5Q_0
timestamp 1736016530
transform 1 0 149 0 1 529
box -221 -126 221 126
use sky130_fd_pr__pfet_01v8_64A2S3  sky130_fd_pr__pfet_01v8_64A2S3_0
timestamp 1736019897
transform 1 0 149 0 1 1475
box -641 -484 641 491
<< labels >>
rlabel metal1 -602 981 -602 981 3 A
port 6 e
rlabel metal1 -602 889 -602 889 3 B
port 7 e
rlabel metal1 -602 793 -602 793 3 C
port 8 e
rlabel metal1 -602 698 -602 698 3 D
port 9 e
rlabel metal1 158 187 158 187 5 VSS
port 10 s
rlabel metal1 -531 1235 -531 1235 5 VDD
port 11 s
rlabel metal1 790 982 790 982 3 Y
port 12 e
<< end >>
