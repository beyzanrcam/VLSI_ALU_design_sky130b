magic
tech sky130B
magscale 1 2
timestamp 1736515926
<< nwell >>
rect -1843 2757 -550 3243
rect 493 2013 3416 2590
rect -298 -904 3416 -328
<< metal1 >>
rect -1841 2505 -1772 2751
rect -1842 2446 -1772 2505
rect -1841 -332 -1772 2446
rect -1499 2530 -1430 2751
rect -1499 2440 -1430 2461
rect -1402 1997 -1333 2751
rect -1059 2528 -990 2590
rect -1059 2446 -990 2459
rect -1408 1991 -1327 1997
rect -1408 1922 -1402 1991
rect -1333 1988 -1327 1991
rect -1333 1922 -1315 1988
rect -1408 1916 -1327 1922
rect -1402 -238 -1333 1916
rect -962 1856 -893 2587
rect -619 2537 -550 2597
rect -962 1781 -893 1787
rect -620 2506 -550 2537
rect -620 1894 -551 2506
rect -294 2077 -242 2083
rect -294 2019 -242 2025
rect -303 1983 -232 1988
rect 705 1984 715 1986
rect -303 1931 -287 1983
rect -235 1931 -232 1983
rect 709 1932 715 1984
rect -303 1922 -232 1931
rect 705 1927 715 1932
rect 1018 1901 1099 1918
rect -620 1828 -231 1894
rect -79 1828 -73 1894
rect -7 1828 -1 1894
rect 1018 1849 1024 1901
rect 1093 1849 1099 1901
rect 1589 1888 1642 1894
rect 1589 1829 1642 1835
rect -620 -135 -551 1828
rect -626 -204 -620 -135
rect -551 -144 -545 -135
rect -551 -204 -232 -144
rect -620 -210 -232 -204
rect -1402 -302 -1334 -238
rect -1401 -304 -1334 -302
rect -1268 -304 -232 -238
rect -1841 -398 -459 -332
rect -393 -398 -229 -332
<< via1 >>
rect -1499 2461 -1430 2530
rect -1059 2459 -990 2528
rect -1402 1922 -1333 1991
rect -962 1787 -893 1856
rect -294 2025 -242 2077
rect 669 2024 722 2076
rect 1602 2025 1655 2077
rect 2533 2025 2586 2077
rect -287 1931 -235 1983
rect 657 1932 709 1984
rect 1600 1927 1652 1979
rect 2535 1927 2587 1979
rect -73 1828 -7 1894
rect 1024 1849 1093 1901
rect 1589 1835 1642 1888
rect 2862 1863 2931 1932
rect -620 -204 -551 -135
rect 1001 -215 1065 -151
rect 1593 -210 1659 -144
rect 2864 -211 2924 -151
rect -1334 -304 -1268 -238
rect 679 -299 731 -247
rect 1601 -304 1667 -238
rect 2537 -303 2603 -237
rect -459 -398 -393 -332
rect 663 -393 728 -341
rect 1592 -393 1657 -341
rect 2551 -393 2616 -341
<< metal2 >>
rect -1499 2641 -287 2710
rect -1499 2530 -1430 2641
rect -1499 2455 -1430 2461
rect -1065 2459 -1059 2528
rect -990 2459 -984 2528
rect -1059 2363 -990 2459
rect -1059 2295 -990 2304
rect -356 2086 -287 2641
rect -356 2077 2740 2086
rect -356 2025 -294 2077
rect -242 2076 1602 2077
rect -242 2025 669 2076
rect -356 2024 669 2025
rect 722 2025 1602 2076
rect 1655 2025 2533 2077
rect 2586 2025 2740 2077
rect 722 2024 2740 2025
rect -356 2017 2740 2024
rect -1408 1991 -1327 1997
rect -1408 1922 -1402 1991
rect -1333 1986 -1327 1991
rect -1333 1984 715 1986
rect -1333 1983 657 1984
rect -1333 1931 -287 1983
rect -235 1932 657 1983
rect 709 1932 715 1984
rect -235 1931 715 1932
rect -1333 1927 715 1931
rect 782 1936 1514 1989
rect 2529 1983 2600 1985
rect -1333 1922 -1327 1927
rect -1408 1916 -1327 1922
rect -79 1894 -7 1899
rect 782 1894 848 1936
rect -971 1856 -884 1865
rect -971 1787 -962 1856
rect -893 1787 -884 1856
rect -79 1828 -73 1894
rect -7 1828 848 1894
rect 1024 1901 1093 1907
rect 1461 1888 1514 1936
rect 1589 1925 1598 1981
rect 1654 1925 1663 1981
rect 2523 1927 2535 1983
rect 2591 1927 2600 1983
rect 2856 1932 2936 1938
rect 2529 1921 2593 1927
rect 1141 1856 1200 1860
rect 1093 1851 1205 1856
rect 1093 1849 1141 1851
rect -79 1822 -7 1828
rect 1024 1792 1141 1849
rect 1200 1792 1205 1851
rect 1461 1835 1589 1888
rect 1642 1835 1648 1888
rect 2856 1863 2862 1932
rect 2931 1863 2936 1932
rect 2856 1856 2936 1863
rect 1024 1787 1205 1792
rect -971 1778 -884 1787
rect 1141 1783 1200 1787
rect 996 -116 1070 -110
rect -620 -135 -551 -129
rect -551 -188 806 -149
rect 996 -151 1005 -116
rect 1061 -151 1070 -116
rect 996 -180 1001 -151
rect -620 -210 -551 -204
rect -1334 -238 -1268 -232
rect -1268 -247 739 -238
rect -1268 -299 679 -247
rect 731 -299 739 -247
rect 767 -257 806 -188
rect 1065 -180 1070 -151
rect 1215 -210 1593 -144
rect 1659 -210 1665 -144
rect 2864 -151 2924 -145
rect 2857 -209 2864 -153
rect 2924 -209 2931 -153
rect 1001 -221 1065 -215
rect 1216 -257 1255 -210
rect 2864 -217 2924 -211
rect 767 -296 1255 -257
rect -1268 -304 739 -299
rect 1592 -304 1601 -238
rect 1667 -304 1676 -238
rect 2531 -303 2537 -237
rect 2603 -303 2612 -237
rect -1334 -310 -1268 -304
rect -466 -398 -459 -332
rect -393 -341 2662 -332
rect -393 -393 663 -341
rect 728 -393 1592 -341
rect 1657 -393 2551 -341
rect 2616 -393 2662 -341
rect -393 -398 2662 -393
rect -459 -404 -393 -398
<< via2 >>
rect -1059 2304 -990 2363
rect -962 1787 -893 1856
rect 1598 1979 1654 1981
rect 1598 1927 1600 1979
rect 1600 1927 1652 1979
rect 1652 1927 1654 1979
rect 1598 1925 1654 1927
rect 2535 1979 2591 1983
rect 2535 1927 2587 1979
rect 2587 1927 2591 1979
rect 1141 1792 1200 1851
rect 2867 1868 2926 1927
rect 1005 -151 1061 -116
rect 1005 -172 1061 -151
rect 2866 -209 2922 -153
rect 1601 -304 1667 -242
rect 2547 -303 2603 -242
<< metal3 >>
rect -1064 2363 -985 2368
rect -1064 2304 -1059 2363
rect -990 2304 -985 2363
rect -1064 2299 -985 2304
rect -1058 2040 -989 2299
rect -1109 1990 -988 2040
rect -1109 1983 2602 1990
rect -1109 1981 2535 1983
rect -1109 1971 1598 1981
rect -1101 1925 1598 1971
rect 1654 1927 2535 1981
rect 2591 1927 2602 1983
rect 1654 1925 2602 1927
rect -1101 1922 2602 1925
rect -1101 -237 -1035 1922
rect -827 1920 2602 1922
rect 2862 1927 2931 1932
rect 2862 1868 2867 1927
rect 2926 1868 2931 1927
rect -967 1856 -888 1861
rect 2862 1856 2931 1868
rect -967 1787 -962 1856
rect -893 1851 2931 1856
rect -893 1792 1141 1851
rect 1200 1792 2931 1851
rect -893 1787 2931 1792
rect -967 1782 -888 1787
rect -967 1709 -893 1782
rect -960 -117 -900 1709
rect 998 -116 1071 -111
rect 998 -117 1005 -116
rect -960 -172 1005 -117
rect 1061 -117 1071 -116
rect 1061 -148 2924 -117
rect 1061 -153 2927 -148
rect 1061 -172 2866 -153
rect -960 -177 2866 -172
rect 2861 -209 2866 -177
rect 2922 -209 2927 -153
rect 2861 -214 2927 -209
rect -1101 -242 2621 -237
rect -1101 -303 1601 -242
rect 1596 -304 1601 -303
rect 1667 -303 2547 -242
rect 2603 -303 2621 -242
rect 1667 -304 1672 -303
rect 1596 -309 1672 -304
rect 2542 -308 2621 -303
use inv  inv_1 ~/Documents/vlsi/vlsi_sky130b/design/mag/inv
timestamp 1735843251
transform 1 0 -1402 0 1 2757
box 0 -311 412 486
use inv  inv_2
timestamp 1735843251
transform 1 0 -962 0 1 2757
box 0 -311 412 486
use inv  inv_3
timestamp 1735843251
transform 1 0 -1842 0 1 2757
box 0 -311 412 486
use NAND4F  NAND4F_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NAND/NAND4
timestamp 1736096163
transform 1 0 2507 0 1 2017
box 10 -1175 909 571
use NAND4F  NAND4F_1
timestamp 1736096163
transform 1 0 1576 0 -1 -333
box 10 -1175 909 571
use NAND4F  NAND4F_2
timestamp 1736096163
transform 1 0 640 0 1 2017
box 10 -1175 909 571
use NAND4F  NAND4F_3
timestamp 1736096163
transform 1 0 1576 0 1 2017
box 10 -1175 909 571
use NAND4F  NAND4F_4
timestamp 1736096163
transform 1 0 -308 0 1 2017
box 10 -1175 909 571
use NAND4F  NAND4F_5
timestamp 1736096163
transform 1 0 -308 0 -1 -333
box 10 -1175 909 571
use NAND4F  NAND4F_6
timestamp 1736096163
transform 1 0 640 0 -1 -333
box 10 -1175 909 571
use NAND4F  NAND4F_7
timestamp 1736096163
transform 1 0 2507 0 -1 -332
box 10 -1175 909 571
<< end >>
