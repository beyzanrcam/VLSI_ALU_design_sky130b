magic
tech sky130B
magscale 1 2
timestamp 1645019219
<< nwell >>
rect 276 354 698 1122
<< pwell >>
rect 276 -204 698 354
<< nmos >>
rect 472 -56 502 144
<< pmos >>
rect 472 574 502 974
<< ndiff >>
rect 414 132 472 144
rect 414 -44 426 132
rect 460 -44 472 132
rect 414 -56 472 -44
rect 502 132 560 144
rect 502 -44 514 132
rect 548 -44 560 132
rect 502 -56 560 -44
<< pdiff >>
rect 414 962 472 974
rect 414 586 426 962
rect 460 586 472 962
rect 414 574 472 586
rect 502 962 560 974
rect 502 586 514 962
rect 548 586 560 962
rect 502 574 560 586
<< ndiffc >>
rect 426 -44 460 132
rect 514 -44 548 132
<< pdiffc >>
rect 426 586 460 962
rect 514 586 548 962
<< psubdiff >>
rect 312 284 662 318
rect 312 -134 346 284
rect 628 -134 662 284
rect 312 -168 408 -134
rect 566 -168 662 -134
<< nsubdiff >>
rect 312 1052 408 1086
rect 566 1052 662 1086
rect 312 424 346 1052
rect 628 424 662 1052
rect 312 390 662 424
<< psubdiffcont >>
rect 408 -168 566 -134
<< nsubdiffcont >>
rect 408 1052 566 1086
<< poly >>
rect 472 974 502 1000
rect 472 543 502 574
rect 454 527 520 543
rect 454 493 470 527
rect 504 493 520 527
rect 454 477 520 493
rect 454 216 520 232
rect 454 182 470 216
rect 504 182 520 216
rect 454 166 520 182
rect 472 144 502 166
rect 472 -82 502 -56
<< polycont >>
rect 470 493 504 527
rect 470 182 504 216
<< locali >>
rect 392 1052 408 1086
rect 566 1052 582 1086
rect 426 962 460 1052
rect 426 570 460 586
rect 514 962 548 978
rect 514 570 548 586
rect 454 493 470 527
rect 504 493 520 527
rect 454 182 470 216
rect 504 182 520 216
rect 426 132 460 148
rect 426 -134 460 -44
rect 514 132 548 148
rect 514 -60 548 -44
rect 392 -168 408 -134
rect 566 -168 582 -134
<< viali >>
rect 426 586 460 962
rect 514 586 548 962
rect 470 493 504 527
rect 470 182 504 216
rect 426 -44 460 132
rect 514 -44 548 132
<< metal1 >>
rect 420 962 466 974
rect -22 804 178 852
rect 420 804 426 962
rect -22 758 426 804
rect -22 652 178 758
rect 420 586 426 758
rect 460 586 466 962
rect 420 574 466 586
rect 508 962 554 974
rect 508 586 514 962
rect 548 828 554 962
rect 548 772 648 828
rect 548 586 554 772
rect 508 574 554 586
rect 458 527 516 533
rect 458 493 470 527
rect 504 493 516 527
rect -12 340 188 420
rect 458 340 516 493
rect -12 294 516 340
rect -12 220 188 294
rect 458 216 516 294
rect 458 182 470 216
rect 504 182 516 216
rect 458 176 516 182
rect 614 410 648 772
rect 784 410 984 478
rect 614 364 984 410
rect 420 132 466 144
rect -8 60 192 108
rect -8 58 254 60
rect 420 58 426 132
rect -8 12 426 58
rect -8 -92 192 12
rect 420 -44 426 12
rect 460 -44 466 132
rect 420 -56 466 -44
rect 508 132 554 144
rect 508 -44 514 132
rect 548 74 554 132
rect 614 74 648 364
rect 784 278 984 364
rect 548 18 656 74
rect 548 -44 554 18
rect 508 -56 554 -44
<< labels >>
flabel metal1 -22 652 178 852 0 FreeSans 256 0 0 0 VDD
port 2 nsew
flabel metal1 -12 220 188 420 0 FreeSans 256 0 0 0 A
port 1 nsew
flabel metal1 784 278 984 478 0 FreeSans 256 0 0 0 Y
port 3 nsew
flabel metal1 -8 -92 192 108 0 FreeSans 256 0 0 0 VSS
port 4 nsew
<< end >>
