magic
tech sky130A
magscale 1 2
timestamp 1736616668
<< nwell >>
rect -3439 3542 3242 4070
rect -3388 1730 -2206 2288
rect -1652 1730 -524 2272
rect -3388 438 -2260 980
rect -1652 438 -524 980
rect -3388 -1535 -2260 -993
rect -1651 -1535 -523 -993
rect -3388 -2827 -2260 -2285
rect -1652 -2827 -524 -2285
rect -3388 -4799 -2260 -4257
rect -1651 -4799 -523 -4257
rect -3388 -6091 -2260 -5549
rect -1651 -6091 -523 -5549
<< locali >>
rect 154 1006 264 1634
rect 154 942 596 1006
<< metal1 >>
rect -2781 3422 -2683 3696
rect -1749 3574 -1335 3576
rect -1749 3557 -1330 3574
rect -2305 3484 -2010 3524
rect -3544 3291 -3388 3372
rect -2305 3365 -2209 3484
rect -2077 3365 -2010 3484
rect -1749 3464 -1687 3557
rect -1369 3470 -1330 3557
rect -1369 3464 -1335 3470
rect -1749 3440 -1335 3464
rect -712 3422 -664 3696
rect 92 3556 400 3579
rect 92 3459 155 3556
rect 362 3459 400 3556
rect 92 3439 400 3459
rect 1030 3422 1078 3696
rect 1933 3558 2137 3578
rect 1933 3451 2001 3558
rect 1933 3439 2137 3451
rect 2792 3422 2856 3696
rect 3218 3535 3508 3553
rect -2305 3320 -2010 3365
rect -1583 3379 -1356 3412
rect -3559 3244 -3350 3291
rect -3559 3066 -3506 3244
rect -3384 3066 -3350 3244
rect -1583 3151 -1550 3379
rect -1387 3151 -1356 3379
rect 100 3265 328 3411
rect -1583 3118 -1356 3151
rect 99 3189 328 3265
rect 1752 3297 2088 3411
rect 3218 3379 3351 3535
rect 3465 3379 3508 3535
rect 3218 3366 3508 3379
rect -3559 3037 -3350 3066
rect 99 3066 127 3189
rect 303 3066 327 3189
rect 1752 3144 1803 3297
rect 2001 3144 2088 3297
rect 1752 3116 2088 3144
rect 99 3043 327 3066
rect -2260 2840 8008 2924
rect -3817 2215 -3534 2234
rect -3818 2167 -3534 2215
rect -3818 1894 -3763 2167
rect -3574 1894 -3534 2167
rect -3818 1852 -3534 1894
rect -3818 1763 -3652 1852
rect -3818 1628 -3388 1763
rect -3818 -1502 -3652 1628
rect -2687 1610 -2639 1884
rect -2260 1615 -2166 2840
rect -2044 2693 -3 2777
rect -3588 1580 -3377 1599
rect -3588 1478 -3551 1580
rect -3397 1478 -3377 1580
rect -3588 1449 -3377 1478
rect -2044 777 -1907 2693
rect -215 2545 -3 2629
rect -1844 1750 -1611 1762
rect -1844 1637 -1792 1750
rect -1646 1637 -1611 1750
rect -1844 1628 -1611 1637
rect -949 1610 -901 1884
rect -215 1702 -84 2545
rect -1867 1592 -1565 1599
rect -1867 1475 -1827 1592
rect -1591 1475 -1565 1592
rect -528 1555 -84 1702
rect -1867 1463 -1565 1475
rect -3588 451 -3274 471
rect -3588 351 -3559 451
rect -3305 351 -3274 451
rect -3588 336 -3274 351
rect -2689 318 -2641 592
rect -3593 182 -3388 307
rect -2308 265 -1907 777
rect -1861 457 -1595 471
rect -1861 348 -1828 457
rect -1624 348 -1595 457
rect -1861 336 -1595 348
rect -956 318 -908 592
rect -566 500 -260 526
rect -566 309 -516 500
rect -303 309 -260 500
rect -1868 295 -1580 307
rect -2308 263 -1968 265
rect -3593 -16 -3568 182
rect -3422 -16 -3388 182
rect -1868 185 -1840 295
rect -1608 185 -1580 295
rect -566 263 -260 309
rect -1868 172 -1580 185
rect -3593 -31 -3388 -16
rect -2260 -341 -2166 -340
rect -2260 -425 9761 -341
rect -3818 -1637 -3388 -1502
rect -3818 -4766 -3652 -1637
rect -2688 -1655 -2640 -1381
rect -2260 -1649 -2166 -425
rect -2044 -572 -3 -488
rect -3588 -1680 -3298 -1666
rect -3588 -1784 -3567 -1680
rect -3324 -1784 -3298 -1680
rect -3588 -1802 -3298 -1784
rect -3588 -2808 -3388 -2794
rect -3588 -2915 -3557 -2808
rect -3401 -2915 -3388 -2808
rect -3588 -2929 -3388 -2915
rect -2687 -2947 -2639 -2673
rect -2044 -2674 -1907 -572
rect -215 -720 -3 -636
rect -1798 -1518 -1623 -1502
rect -1798 -1625 -1764 -1518
rect -1644 -1625 -1623 -1518
rect -1798 -1637 -1623 -1625
rect -949 -1655 -901 -1381
rect -215 -1563 -84 -720
rect -1866 -1676 -1570 -1666
rect -1866 -1784 -1813 -1676
rect -1584 -1784 -1570 -1676
rect -531 -1710 -84 -1563
rect -1866 -1807 -1570 -1784
rect -3593 -3083 -3388 -2958
rect -2307 -3000 -1907 -2674
rect -1866 -2795 -1644 -2794
rect -1866 -2806 -1614 -2795
rect -1866 -2917 -1841 -2806
rect -1639 -2917 -1614 -2806
rect -1866 -2929 -1614 -2917
rect -950 -2947 -902 -2673
rect -566 -2788 -260 -2739
rect -1869 -2980 -1609 -2958
rect -2307 -3002 -1968 -3000
rect -3593 -3281 -3568 -3083
rect -3422 -3281 -3388 -3083
rect -1869 -3072 -1847 -2980
rect -1642 -3072 -1609 -2980
rect -566 -2962 -529 -2788
rect -307 -2962 -260 -2788
rect -566 -3002 -260 -2962
rect -1869 -3094 -1609 -3072
rect -3593 -3296 -3388 -3281
rect -2260 -3689 -3 -3605
rect -3818 -4901 -3388 -4766
rect -2687 -4919 -2639 -4645
rect -3588 -4956 -3225 -4930
rect -3588 -5047 -3519 -4956
rect -3291 -5047 -3225 -4956
rect -2260 -4974 -2167 -3689
rect -2044 -3836 -3 -3752
rect -3588 -5066 -3225 -5047
rect -2044 -5783 -1907 -3836
rect -215 -3984 -3 -3900
rect -951 -4919 -903 -4645
rect -215 -4827 -84 -3984
rect -528 -4974 -84 -4827
rect -3588 -6082 -3281 -6058
rect -3588 -6169 -3526 -6082
rect -3309 -6169 -3281 -6082
rect -3588 -6193 -3281 -6169
rect -2685 -6211 -2637 -5937
rect -3593 -6347 -3388 -6222
rect -2307 -6264 -1907 -5783
rect -1866 -6085 -1593 -6058
rect -1866 -6177 -1824 -6085
rect -1626 -6177 -1593 -6085
rect -1866 -6193 -1593 -6177
rect -958 -6211 -910 -5937
rect -566 -6045 -260 -6003
rect -1729 -6241 -1528 -6223
rect -2307 -6266 -1968 -6264
rect -3593 -6545 -3568 -6347
rect -3422 -6545 -3388 -6347
rect -1729 -6329 -1686 -6241
rect -1567 -6329 -1528 -6241
rect -566 -6231 -510 -6045
rect -311 -6231 -260 -6045
rect -566 -6266 -260 -6231
rect -1729 -6358 -1528 -6329
rect -3593 -6560 -3388 -6545
<< via1 >>
rect -2209 3365 -2077 3484
rect -1687 3464 -1369 3557
rect 155 3459 362 3556
rect 2001 3451 2150 3558
rect -3506 3066 -3384 3244
rect -1550 3151 -1387 3379
rect 3351 3379 3465 3535
rect 127 3066 303 3189
rect 1803 3144 2001 3297
rect -3763 1894 -3574 2167
rect -3551 1478 -3397 1580
rect -1792 1637 -1646 1750
rect -1827 1475 -1591 1592
rect -3559 351 -3305 451
rect -1828 348 -1624 457
rect -516 309 -303 500
rect -3568 -16 -3422 182
rect -1840 185 -1608 295
rect -3567 -1784 -3324 -1680
rect -3557 -2915 -3401 -2808
rect -1764 -1625 -1644 -1518
rect -1813 -1784 -1584 -1676
rect -1841 -2917 -1639 -2806
rect -3568 -3281 -3422 -3083
rect -1847 -3072 -1642 -2980
rect -529 -2962 -307 -2788
rect -3519 -5047 -3291 -4956
rect -3526 -6169 -3309 -6082
rect -1824 -6177 -1626 -6085
rect -3568 -6545 -3422 -6347
rect -1686 -6329 -1567 -6241
rect -510 -6231 -311 -6045
<< metal2 >>
rect -3591 4118 2084 4255
rect -3591 3625 -3448 4118
rect -1749 3576 -1606 4118
rect 92 3579 235 4118
rect -1749 3557 -1335 3576
rect -2251 3511 -2177 3515
rect -2251 3484 -2030 3511
rect -2251 3365 -2209 3484
rect -2077 3365 -2030 3484
rect -1749 3464 -1687 3557
rect -1369 3464 -1335 3557
rect 92 3556 400 3579
rect -1749 3440 -1335 3464
rect -364 3511 -244 3515
rect -2251 3324 -2030 3365
rect -3559 3244 -3350 3291
rect -3559 3066 -3506 3244
rect -3384 3066 -3350 3244
rect -3559 3037 -3350 3066
rect -2216 2727 -2030 3324
rect -1583 3379 -1356 3412
rect -1583 3151 -1550 3379
rect -1387 3151 -1356 3379
rect -364 3327 -135 3511
rect 92 3459 155 3556
rect 362 3459 400 3556
rect 1933 3578 2076 4118
rect 1933 3558 2238 3578
rect 92 3439 400 3459
rect 1477 3510 1516 3515
rect 1477 3327 1600 3510
rect 1933 3451 2001 3558
rect 2150 3451 2238 3558
rect 1933 3439 2238 3451
rect 3318 3535 3608 3554
rect 3318 3379 3351 3535
rect 3465 3379 3608 3535
rect 3318 3367 3608 3379
rect -1583 3118 -1356 3151
rect -275 2833 -135 3327
rect 100 3189 318 3210
rect 100 3066 127 3189
rect 303 3066 318 3189
rect 100 3045 318 3066
rect 1505 2985 1600 3327
rect 1752 3297 2032 3323
rect 1752 3144 1803 3297
rect 2001 3144 2032 3297
rect 1752 3116 2032 3144
rect 3453 3186 3608 3367
rect 3453 3064 13159 3186
rect 3458 3036 13159 3064
rect 1505 2984 10159 2985
rect 1505 2876 10170 2984
rect -1285 2727 -968 2736
rect -2216 2666 -968 2727
rect -285 2722 6879 2833
rect -2216 2614 3582 2666
rect -1285 2553 3582 2614
rect -1285 2544 -968 2553
rect -1869 2517 -1700 2527
rect -1869 2489 -1407 2517
rect -1869 2383 -1556 2489
rect -1432 2383 -1407 2489
rect 3458 2408 3581 2553
rect -1869 2354 -1407 2383
rect 6750 2376 6878 2722
rect 10028 2388 10170 2876
rect -3817 2167 -3534 2234
rect -3817 1894 -3763 2167
rect -3574 1894 -3534 2167
rect -3817 1852 -3534 1894
rect -1869 1763 -1700 2354
rect -2166 1762 -1692 1763
rect -2166 1751 -1611 1762
rect -2166 1637 -2151 1751
rect -2020 1750 -1611 1751
rect -2020 1637 -1792 1750
rect -1646 1637 -1611 1750
rect -2166 1628 -1611 1637
rect -3588 1580 -3377 1599
rect -3588 1478 -3551 1580
rect -3397 1478 -3377 1580
rect -3588 1449 -3377 1478
rect -1867 1592 -1565 1599
rect -1867 1475 -1827 1592
rect -1591 1475 -1565 1592
rect -1867 1463 -1565 1475
rect -312 1468 -3 1475
rect -3588 1204 -3412 1449
rect -1866 1204 -1692 1463
rect -3590 1069 -1692 1204
rect -3588 483 -3412 1069
rect -3588 471 -3410 483
rect -1866 471 -1692 1069
rect -351 1335 -3 1468
rect -518 526 -433 528
rect -351 526 -260 1335
rect -566 500 -260 526
rect -3588 451 -3274 471
rect -3588 351 -3559 451
rect -3305 351 -3274 451
rect -3588 336 -3274 351
rect -1866 457 -1595 471
rect -1866 348 -1828 457
rect -1624 348 -1595 457
rect -1866 336 -1595 348
rect -566 309 -516 500
rect -303 309 -260 500
rect -1868 295 -1580 307
rect -3593 182 -3395 211
rect -3593 -16 -3568 182
rect -3422 -16 -3395 182
rect -3593 -31 -3395 -16
rect -1868 185 -1840 295
rect -1608 185 -1580 295
rect -566 263 -260 309
rect -1868 -210 -1818 185
rect -1729 172 -1580 185
rect -1729 -108 -1692 172
rect -1729 -210 -1693 -108
rect -1868 -254 -1693 -210
rect 10 -200 287 -196
rect 10 -401 315 -200
rect 3275 -213 3407 -128
rect 6574 -187 6881 -83
rect 3275 -343 3638 -213
rect 3342 -344 3638 -343
rect -3604 -447 -299 -427
rect -3604 -453 -471 -447
rect -3604 -593 -3575 -453
rect -3446 -587 -471 -453
rect -342 -587 -299 -447
rect -3446 -593 -299 -587
rect -3604 -614 -299 -593
rect 171 -822 315 -401
rect 3452 -848 3636 -344
rect 6755 -863 6878 -187
rect 9870 -241 9997 -101
rect 13154 -136 13282 56
rect 10040 -241 10168 -240
rect 9865 -397 10168 -241
rect 9870 -398 9997 -397
rect 10040 -839 10168 -397
rect -2166 -1512 -1623 -1502
rect -2166 -1626 -2154 -1512
rect -2023 -1514 -1623 -1512
rect -2020 -1518 -1623 -1514
rect -2020 -1625 -1764 -1518
rect -1644 -1625 -1623 -1518
rect -2166 -1628 -2151 -1626
rect -2020 -1628 -1623 -1625
rect -2166 -1637 -1623 -1628
rect -3588 -1680 -3298 -1666
rect -3588 -1784 -3567 -1680
rect -3324 -1784 -3298 -1680
rect -3588 -1802 -3298 -1784
rect -1866 -1676 -1570 -1666
rect -1866 -1784 -1813 -1676
rect -1584 -1784 -1570 -1676
rect -3588 -2061 -3412 -1802
rect -1866 -1807 -1570 -1784
rect -312 -1797 -3 -1790
rect -1866 -2061 -1690 -1807
rect -3590 -2196 -1690 -2061
rect -3588 -2794 -3412 -2196
rect -1866 -2794 -1690 -2196
rect -351 -1930 -3 -1797
rect -518 -2739 -433 -2737
rect -351 -2739 -260 -1930
rect -566 -2788 -260 -2739
rect -3588 -2808 -3388 -2794
rect -3588 -2915 -3557 -2808
rect -3401 -2915 -3388 -2808
rect -3588 -2929 -3388 -2915
rect -1866 -2795 -1644 -2794
rect -1866 -2806 -1614 -2795
rect -1866 -2917 -1841 -2806
rect -1639 -2917 -1614 -2806
rect -1866 -2929 -1614 -2917
rect -1869 -2980 -1609 -2958
rect -3593 -3083 -3395 -3054
rect -3593 -3281 -3568 -3083
rect -3422 -3281 -3395 -3083
rect -1869 -3072 -1847 -2980
rect -1642 -3072 -1609 -2980
rect -566 -2962 -529 -2788
rect -307 -2962 -260 -2788
rect -566 -3002 -260 -2962
rect -1869 -3094 -1822 -3072
rect -3593 -3296 -3395 -3281
rect -1867 -3454 -1822 -3094
rect -1729 -3094 -1609 -3072
rect -1729 -3373 -1692 -3094
rect -1867 -3475 -1818 -3454
rect -1729 -3475 -1693 -3373
rect -1867 -3519 -1693 -3475
rect -11 -3621 314 -3495
rect 3281 -3497 3615 -3375
rect 169 -4142 299 -3621
rect 3456 -4161 3592 -3497
rect 6570 -3532 6886 -3387
rect 9874 -3505 10165 -3369
rect 13156 -3414 13288 -3296
rect 6744 -4189 6874 -3532
rect 10040 -4161 10164 -3505
rect -2166 -4776 -1533 -4766
rect -2166 -4890 -2154 -4776
rect -2017 -4890 -1533 -4776
rect -2166 -4892 -2151 -4890
rect -2020 -4892 -1533 -4890
rect -2166 -4901 -1533 -4892
rect -3588 -4956 -3225 -4930
rect -3588 -5047 -3519 -4956
rect -3291 -5047 -3225 -4956
rect -3588 -5066 -3225 -5047
rect -1866 -5066 -1547 -4930
rect -312 -5061 -3 -5054
rect -3588 -5325 -3412 -5066
rect -1866 -5325 -1690 -5066
rect -3590 -5460 -1690 -5325
rect -3588 -6058 -3412 -5460
rect -1866 -6058 -1690 -5460
rect -351 -5194 -3 -5061
rect -518 -6003 -433 -6001
rect -351 -6003 -260 -5194
rect -566 -6045 -260 -6003
rect -3588 -6082 -3281 -6058
rect -3588 -6169 -3526 -6082
rect -3309 -6169 -3281 -6082
rect -3588 -6193 -3281 -6169
rect -1866 -6085 -1593 -6058
rect -1866 -6177 -1824 -6085
rect -1626 -6177 -1593 -6085
rect -1866 -6193 -1593 -6177
rect -1867 -6229 -1528 -6223
rect -1868 -6241 -1528 -6229
rect -1868 -6272 -1686 -6241
rect -1868 -6287 -1822 -6272
rect -3593 -6347 -3395 -6318
rect -3593 -6545 -3568 -6347
rect -3422 -6545 -3395 -6347
rect -3593 -6560 -3395 -6545
rect -1868 -6733 -1825 -6287
rect -1733 -6293 -1686 -6272
rect -1729 -6329 -1686 -6293
rect -1567 -6329 -1528 -6241
rect -566 -6231 -510 -6045
rect -311 -6231 -260 -6045
rect -566 -6266 -260 -6231
rect -1729 -6358 -1528 -6329
rect -1729 -6637 -1692 -6358
rect -1868 -6739 -1818 -6733
rect -1729 -6739 -1693 -6637
rect -1868 -6783 -1693 -6739
rect 5 -6819 190 -6596
rect 3288 -6679 3396 -6550
rect 6579 -6679 6688 -6554
rect 9870 -6679 9978 -6550
rect 13156 -6678 13288 -6560
<< via2 >>
rect -3506 3066 -3384 3244
rect -1550 3151 -1387 3379
rect 127 3066 303 3189
rect 1803 3144 2001 3297
rect -1556 2383 -1432 2489
rect -3763 1894 -3574 2167
rect -2151 1637 -2020 1751
rect -3568 -16 -3422 182
rect -1818 185 -1729 236
rect -1818 -210 -1729 185
rect -3575 -593 -3446 -453
rect -471 -587 -342 -447
rect -2154 -1514 -2023 -1512
rect -2154 -1626 -2020 -1514
rect -2151 -1628 -2020 -1626
rect -3568 -3281 -3422 -3083
rect -1822 -3029 -1733 -3008
rect -1822 -3072 -1729 -3029
rect -1822 -3454 -1729 -3072
rect -1818 -3475 -1729 -3454
rect -2154 -4890 -2017 -4776
rect -2151 -4892 -2020 -4890
rect -1822 -6287 -1733 -6272
rect -3568 -6545 -3422 -6347
rect -1825 -6293 -1733 -6287
rect -1825 -6733 -1729 -6293
rect -1818 -6739 -1729 -6733
<< metal3 >>
rect -3817 4255 -3635 4259
rect -3817 4090 1969 4255
rect -3817 2234 -3635 4090
rect -1583 3379 -1356 3412
rect -3544 3291 -3354 3372
rect -3559 3244 -3350 3291
rect -3559 3066 -3506 3244
rect -3384 3066 -3350 3244
rect -3559 3037 -3350 3066
rect -1583 3151 -1550 3379
rect -1387 3151 -1356 3379
rect 1752 3323 1969 4090
rect 1752 3297 2032 3323
rect -1583 3118 -1356 3151
rect 100 3189 318 3210
rect -3542 2836 -3358 3037
rect -3542 2832 -1710 2836
rect -3542 2636 -1708 2832
rect -3817 2167 -3534 2234
rect -3817 1894 -3763 2167
rect -3574 1894 -3534 2167
rect -3817 1852 -3534 1894
rect -2166 1751 -2007 1796
rect -2166 1637 -2151 1751
rect -2020 1637 -2007 1751
rect -3607 211 -3416 332
rect -3607 182 -3395 211
rect -3607 -16 -3568 182
rect -3422 -16 -3395 182
rect -3607 -31 -3395 -16
rect -3607 -453 -3416 -31
rect -3607 -593 -3575 -453
rect -3446 -593 -3416 -453
rect -3607 -3054 -3416 -593
rect -2166 -1512 -2007 1637
rect -2166 -1626 -2154 -1512
rect -2023 -1514 -2007 -1512
rect -2166 -1628 -2151 -1626
rect -2020 -1628 -2007 -1514
rect -3607 -3083 -3395 -3054
rect -3607 -3281 -3568 -3083
rect -3422 -3281 -3395 -3083
rect -3607 -3296 -3395 -3281
rect -3607 -6318 -3416 -3296
rect -2166 -4776 -2007 -1628
rect -2166 -4890 -2154 -4776
rect -2017 -4890 -2007 -4776
rect -2166 -4892 -2151 -4890
rect -2020 -4892 -2007 -4890
rect -2166 -4901 -2007 -4892
rect -1893 236 -1708 2636
rect -1583 2489 -1415 3118
rect 100 3066 127 3189
rect 303 3066 318 3189
rect 1752 3144 1803 3297
rect 2001 3144 2032 3297
rect 1752 3116 2032 3144
rect 100 3052 318 3066
rect -480 3045 318 3052
rect -480 3033 271 3045
rect -1583 2383 -1556 2489
rect -1432 2383 -1415 2489
rect -1583 2362 -1415 2383
rect -481 2868 271 3033
rect -481 2858 265 2868
rect -1893 -210 -1818 236
rect -1729 -210 -1708 236
rect -1893 -3008 -1708 -210
rect -481 -447 -301 2858
rect -481 -587 -471 -447
rect -342 -587 -301 -447
rect -481 -623 -301 -587
rect -1893 -3454 -1822 -3008
rect -1733 -3029 -1708 -3008
rect -1893 -3475 -1818 -3454
rect -1729 -3475 -1708 -3029
rect -1893 -6272 -1708 -3475
rect -1893 -6287 -1822 -6272
rect -3607 -6347 -3395 -6318
rect -3607 -6545 -3568 -6347
rect -3422 -6545 -3395 -6347
rect -3607 -6560 -3395 -6545
rect -3607 -6772 -3416 -6560
rect -1893 -6733 -1825 -6287
rect -1733 -6293 -1708 -6272
rect -1893 -6739 -1818 -6733
rect -1729 -6739 -1708 -6293
rect -1893 -6782 -1708 -6739
<< metal5 >>
rect -3818 -7001 13360 4259
use 4bit_ADDER  4bit_ADDER_0
timestamp 1736616668
transform 1 0 171 0 1 -165
box -174 -307 13189 3089
use 4bit_ADDER  4bit_ADDER_1
timestamp 1736616668
transform 1 0 171 0 1 -3430
box -174 -307 13189 3089
use 4bit_ADDER  4bit_ADDER_2
timestamp 1736616668
transform 1 0 171 0 1 -6694
box -174 -307 13189 3089
use INV  INV_0
timestamp 1735843251
transform 1 0 -2684 0 1 3542
box 0 -311 412 486
use INV  INV_1
timestamp 1735843251
transform 1 0 -664 0 1 3542
box 0 -311 412 486
use INV  INV_2
timestamp 1735843251
transform 1 0 1077 0 1 3542
box 0 -311 412 486
use INV  INV_3
timestamp 1735843251
transform 1 0 2856 0 1 3542
box 0 -311 412 486
use INV  INV_4
timestamp 1735843251
transform 1 0 -2642 0 1 438
box 0 -311 412 486
use INV  INV_5
timestamp 1735843251
transform 1 0 -2640 0 1 1730
box 0 -311 412 486
use INV  INV_6
timestamp 1735843251
transform 1 0 -2640 0 1 -1535
box 0 -311 412 486
use INV  INV_7
timestamp 1735843251
transform 1 0 -2639 0 1 -2827
box 0 -311 412 486
use INV  INV_8
timestamp 1735843251
transform 1 0 -2639 0 1 -4799
box 0 -311 412 486
use INV  INV_9
timestamp 1735843251
transform 1 0 -2639 0 1 -6091
box 0 -311 412 486
use INV  INV_10
timestamp 1735843251
transform 1 0 -902 0 1 1730
box 0 -311 412 486
use INV  INV_11
timestamp 1735843251
transform 1 0 -908 0 1 438
box 0 -311 412 486
use INV  INV_12
timestamp 1735843251
transform 1 0 -906 0 1 -1535
box 0 -311 412 486
use INV  INV_13
timestamp 1735843251
transform 1 0 -902 0 1 -2827
box 0 -311 412 486
use INV  INV_14
timestamp 1735843251
transform 1 0 -906 0 1 -4799
box 0 -311 412 486
use INV  INV_15
timestamp 1735843251
transform 1 0 -910 0 1 -6091
box 0 -311 412 486
use NAND2  NAND2_0
timestamp 1736436273
transform 1 0 -3795 0 1 3170
box 356 -17 1062 804
use NAND2  NAND2_1
timestamp 1736436273
transform 1 0 -1758 0 1 3170
box 356 -17 1062 804
use NAND2  NAND2_2
timestamp 1736436273
transform 1 0 -28 0 1 3170
box 356 -17 1062 804
use NAND2  NAND2_3
timestamp 1736436273
transform 1 0 1732 0 1 3170
box 356 -17 1062 804
use NAND2  NAND2_4
timestamp 1736436273
transform 1 0 -3744 0 1 1358
box 356 -17 1062 804
use NAND2  NAND2_5
timestamp 1736436273
transform 1 0 -3744 0 1 66
box 356 -17 1062 804
use NAND2  NAND2_6
timestamp 1736436273
transform 1 0 -3744 0 1 -1907
box 356 -17 1062 804
use NAND2  NAND2_7
timestamp 1736436273
transform 1 0 -3744 0 1 -3199
box 356 -17 1062 804
use NAND2  NAND2_8
timestamp 1736436273
transform 1 0 -3744 0 1 -5171
box 356 -17 1062 804
use NAND2  NAND2_9
timestamp 1736436273
transform 1 0 -3744 0 1 -6463
box 356 -17 1062 804
use NAND2  NAND2_10
timestamp 1736436273
transform 1 0 -2008 0 1 1358
box 356 -17 1062 804
use NAND2  NAND2_11
timestamp 1736436273
transform 1 0 -2008 0 1 66
box 356 -17 1062 804
use NAND2  NAND2_12
timestamp 1736436273
transform 1 0 -2007 0 1 -1907
box 356 -17 1062 804
use NAND2  NAND2_13
timestamp 1736436273
transform 1 0 -2008 0 1 -3199
box 356 -17 1062 804
use NAND2  NAND2_14
timestamp 1736436273
transform 1 0 -2007 0 1 -5171
box 356 -17 1062 804
use NAND2  NAND2_15
timestamp 1736436273
transform 1 0 -2007 0 1 -6463
box 356 -17 1062 804
<< labels >>
flabel metal2 -3228 -2190 -3108 -2070 1 FreeSerif 160 0 0 0 B2
port 7 n
flabel metal2 -3220 -5452 -3100 -5332 1 FreeSerif 160 0 0 0 B3
port 9 n
flabel metal2 -2952 -576 -2832 -456 1 FreeSerif 160 0 0 0 A1
port 11 n
flabel metal2 12820 3054 12940 3174 1 FreeSerif 160 0 0 0 SO
port 13 n
flabel metal3 -2146 -202 -2026 -82 1 FreeSerif 160 0 0 0 A2
port 10 n
flabel metal1 -3794 1646 -3674 1766 1 FreeSerif 160 0 0 0 A0
port 6 n
flabel metal3 -3190 2678 -3070 2798 1 FreeSerif 160 0 0 0 A3
port 12 n
flabel metal2 -3584 3886 -3464 4006 1 FreeSerif 160 0 0 0 B0
port 8 n
rlabel metal2 -518 407 -518 407 3 Y
port 3 e
rlabel metal2 -518 -6122 -518 -6122 3 Y
port 3 e
flabel metal2 -3556 1080 -3436 1200 1 FreeSerif 160 0 0 0 B1
port 5 n
rlabel via1 -518 -2858 -518 -2858 3 Y
port 3 e
flabel metal2 54 -6728 150 -6642 1 FreeSerif 160 0 0 0 S7
port 19 n
flabel metal2 13182 -6664 13278 -6578 1 FreeSerif 160 0 0 0 S3
port 18 n
flabel metal2 9878 -6670 9974 -6584 1 FreeSerif 160 0 0 0 S4
port 17 n
flabel metal2 6586 -6668 6682 -6582 1 FreeSerif 160 0 0 0 S5
port 16 n
flabel metal2 13182 -3394 13278 -3308 1 FreeSerif 160 0 0 0 S2
port 15 n
flabel metal2 13166 -32 13262 54 1 FreeSerif 160 0 0 0 S1
port 14 n
flabel metal2 3294 -6664 3390 -6578 1 FreeSerif 160 0 0 0 S6
port 20 n
<< end >>
