* NGSPICE file created from nor4_pex.ext - technology: sky130B

.subckt nor4_pex A B C D VSS VDD Y
X0 Y.t3 D.t0 a_371_1047.t3 VDD.t5 sky130_fd_pr__pfet_01v8 ad=1.2412 pd=8.85 as=1.2412 ps=8.85 w=8.56 l=0.3
X1 VSS.t3 D.t1 Y.t4 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.3
X2 Y.t2 D.t2 a_371_1047.t1 VDD.t4 sky130_fd_pr__pfet_01v8 ad=2.4824 pd=17.7 as=1.2412 ps=8.85 w=8.56 l=0.3
X3 a_371_1047.t4 C.t0 a_17_1047.t2 VDD.t6 sky130_fd_pr__pfet_01v8 ad=1.2412 pd=8.85 as=1.2412 ps=8.85 w=8.56 l=0.3
X4 VSS.t5 B.t0 Y.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
X5 a_371_1047.t0 C.t1 a_17_1047.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.2412 pd=8.85 as=1.2412 ps=8.85 w=8.56 l=0.3
X6 a_n337_1047.t2 A.t0 VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=1.2412 pd=8.85 as=1.2412 ps=8.85 w=8.56 l=0.3
X7 Y.t6 A.t1 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.3
X8 Y.t0 C.t2 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
X9 a_n337_1047.t1 A.t2 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=1.2412 pd=8.85 as=2.4824 ps=17.7 w=8.56 l=0.3
X10 a_17_1047.t5 B.t1 a_n337_1047.t5 VDD.t11 sky130_fd_pr__pfet_01v8 ad=1.2412 pd=8.85 as=1.2412 ps=8.85 w=8.56 l=0.3
X11 a_17_1047.t0 C.t3 a_371_1047.t5 VDD.t14 sky130_fd_pr__pfet_01v8 ad=1.2412 pd=8.85 as=1.2412 ps=8.85 w=8.56 l=0.3
X12 a_371_1047.t2 D.t3 Y.t1 VDD.t3 sky130_fd_pr__pfet_01v8 ad=1.2412 pd=8.85 as=1.2412 ps=8.85 w=8.56 l=0.3
X13 VDD.t10 A.t3 a_n337_1047.t0 VDD.t9 sky130_fd_pr__pfet_01v8 ad=1.2412 pd=8.85 as=1.2412 ps=8.85 w=8.56 l=0.3
X14 a_n337_1047.t4 B.t2 a_17_1047.t4 VDD.t8 sky130_fd_pr__pfet_01v8 ad=1.2412 pd=8.85 as=1.2412 ps=8.85 w=8.56 l=0.3
X15 a_17_1047.t3 B.t3 a_n337_1047.t3 VDD.t7 sky130_fd_pr__pfet_01v8 ad=1.2412 pd=8.85 as=1.2412 ps=8.85 w=8.56 l=0.3
R0 D.n0 D.t0 920.658
R1 D.n0 D.t2 920.658
R2 D.n0 D.t3 888.658
R3 D.n1 D.t1 488.247
R4 D.n1 D.n0 18.6187
R5 D D.n1 11.3874
R6 a_371_1047.n2 a_371_1047.n1 198.589
R7 a_371_1047.n2 a_371_1047.n0 198.589
R8 a_371_1047.n3 a_371_1047.n2 198.552
R9 a_371_1047.n1 a_371_1047.t5 3.33753
R10 a_371_1047.n1 a_371_1047.t4 3.33753
R11 a_371_1047.n0 a_371_1047.t1 3.33753
R12 a_371_1047.n0 a_371_1047.t2 3.33753
R13 a_371_1047.n3 a_371_1047.t3 3.33753
R14 a_371_1047.t0 a_371_1047.n3 3.33753
R15 Y.n1 Y.t2 186.383
R16 Y.n1 Y.n0 183.047
R17 Y.n4 Y.n2 67.5725
R18 Y.n4 Y.n3 67.4397
R19 Y.n3 Y.t4 8.7005
R20 Y.n3 Y.t0 8.7005
R21 Y.n2 Y.t5 8.7005
R22 Y.n2 Y.t6 8.7005
R23 Y.n0 Y.t1 3.33753
R24 Y.n0 Y.t3 3.33753
R25 Y Y.n1 2.23104
R26 Y Y.n4 0.263392
R27 VDD.n1 VDD.t13 186.383
R28 VDD.n1 VDD.n0 183.047
R29 VDD VDD.n1 126.691
R30 VDD.t3 VDD.t4 50.8165
R31 VDD.t5 VDD.t3 50.8165
R32 VDD.t0 VDD.t5 50.8165
R33 VDD.t14 VDD.t0 50.8165
R34 VDD.t6 VDD.t14 50.8165
R35 VDD.t7 VDD.t6 50.8165
R36 VDD.t8 VDD.t7 50.8165
R37 VDD.t11 VDD.t8 50.8165
R38 VDD.t1 VDD.t11 50.8165
R39 VDD.t9 VDD.t1 50.8165
R40 VDD VDD.t12 26.2698
R41 VDD VDD.t9 24.5472
R42 VDD.n0 VDD.t2 3.33753
R43 VDD.n0 VDD.t10 3.33753
R44 VDD.t12 VDD 0.861787
R45 VSS.t0 VSS.t2 445.666
R46 VSS.t4 VSS.t6 445.666
R47 VSS.n3 VSS.t0 253.048
R48 VSS.n3 VSS.t4 192.619
R49 VSS.n1 VSS.t3 148.349
R50 VSS VSS.t7 144.772
R51 VSS.n1 VSS.n0 126.457
R52 VSS.n5 VSS.n4 48.7505
R53 VSS.n4 VSS.n3 48.7505
R54 VSS.n4 VSS.n2 42.9266
R55 VSS.n0 VSS.t1 8.7005
R56 VSS.n0 VSS.t5 8.7005
R57 VSS.n5 VSS 3.13063
R58 VSS VSS.n5 0.391766
R59 VSS VSS.n1 0.0563952
R60 C.n0 C.t0 920.658
R61 C.n0 C.t1 920.658
R62 C.n0 C.t3 888.658
R63 C.n1 C.t2 403.702
R64 C.n1 C.n0 54.5383
R65 C C.n1 10.5749
R66 a_17_1047.n2 a_17_1047.n1 183.081
R67 a_17_1047.n2 a_17_1047.n0 183.081
R68 a_17_1047.n3 a_17_1047.n2 183.047
R69 a_17_1047.n1 a_17_1047.t4 3.33753
R70 a_17_1047.n1 a_17_1047.t5 3.33753
R71 a_17_1047.n0 a_17_1047.t1 3.33753
R72 a_17_1047.n0 a_17_1047.t0 3.33753
R73 a_17_1047.t2 a_17_1047.n3 3.33753
R74 a_17_1047.n3 a_17_1047.t3 3.33753
R75 B.n0 B.t1 920.658
R76 B.n0 B.t3 920.658
R77 B.n0 B.t2 888.658
R78 B.n1 B.t0 380.817
R79 B.n1 B.n0 77.4231
R80 B B.n1 10.4056
R81 A.n0 A.t2 920.658
R82 A.n0 A.t0 920.658
R83 A.n0 A.t3 888.658
R84 A.n1 A.t1 417.846
R85 A.n1 A.n0 89.0187
R86 A A.n1 9.73589
R87 a_n337_1047.n2 a_n337_1047.n1 198.589
R88 a_n337_1047.n2 a_n337_1047.n0 198.589
R89 a_n337_1047.n3 a_n337_1047.n2 198.552
R90 a_n337_1047.n1 a_n337_1047.t0 3.33753
R91 a_n337_1047.n1 a_n337_1047.t1 3.33753
R92 a_n337_1047.n0 a_n337_1047.t3 3.33753
R93 a_n337_1047.n0 a_n337_1047.t4 3.33753
R94 a_n337_1047.n3 a_n337_1047.t5 3.33753
R95 a_n337_1047.t2 a_n337_1047.n3 3.33753
C0 C VDD 0.028417f
C1 VDD B 0.052775f
C2 VDD Y 0.103029f
C3 C B 1.43522f
C4 VDD D 0.091693f
C5 C Y 0.096376f
C6 Y B 0.078972f
C7 C D 1.13157f
C8 B D 0.112523f
C9 Y D 0.512491f
C10 VDD A 0.266201f
C11 C A 0.063981f
C12 B A 0.804134f
C13 Y A 0.015958f
C14 A D 0.094438f
C15 Y VSS 2.648274f
C16 D VSS 0.819834f
C17 C VSS 0.51477f
C18 B VSS 0.558936f
C19 A VSS 0.822639f
C20 VDD VSS 11.712298f
C21 a_n337_1047.t5 VSS 0.121162f
C22 a_n337_1047.t3 VSS 0.121162f
C23 a_n337_1047.t4 VSS 0.121162f
C24 a_n337_1047.n0 VSS 0.40268f
C25 a_n337_1047.t0 VSS 0.121162f
C26 a_n337_1047.t1 VSS 0.121162f
C27 a_n337_1047.n1 VSS 0.40268f
C28 a_n337_1047.n2 VSS 2.36511f
C29 a_n337_1047.n3 VSS 0.402555f
C30 a_n337_1047.t2 VSS 0.121162f
C31 a_17_1047.t3 VSS 0.113028f
C32 a_17_1047.t1 VSS 0.113028f
C33 a_17_1047.t0 VSS 0.113028f
C34 a_17_1047.n0 VSS 0.371211f
C35 a_17_1047.t4 VSS 0.113028f
C36 a_17_1047.t5 VSS 0.113028f
C37 a_17_1047.n1 VSS 0.371211f
C38 a_17_1047.n2 VSS 2.40833f
C39 a_17_1047.n3 VSS 0.371085f
C40 a_17_1047.t2 VSS 0.113028f
C41 VDD.t4 VSS 0.263427f
C42 VDD.t3 VSS 0.136936f
C43 VDD.t5 VSS 0.136936f
C44 VDD.t0 VSS 0.136936f
C45 VDD.t14 VSS 0.136936f
C46 VDD.t6 VSS 0.136936f
C47 VDD.t7 VSS 0.136936f
C48 VDD.t8 VSS 0.136936f
C49 VDD.t11 VSS 0.136936f
C50 VDD.t1 VSS 0.136936f
C51 VDD.t9 VSS 0.101541f
C52 VDD.t2 VSS 0.013059f
C53 VDD.t10 VSS 0.013059f
C54 VDD.n0 VSS 0.042874f
C55 VDD.t13 VSS 0.067989f
C56 VDD.n1 VSS 0.187678f
C57 VDD.t12 VSS 0.036555f
C58 Y.t2 VSS 0.418546f
C59 Y.t1 VSS 0.08039f
C60 Y.t3 VSS 0.08039f
C61 Y.n0 VSS 0.263931f
C62 Y.n1 VSS 1.14787f
C63 Y.t5 VSS 0.018783f
C64 Y.t6 VSS 0.018783f
C65 Y.n2 VSS 0.053481f
C66 Y.t4 VSS 0.018783f
C67 Y.t0 VSS 0.018783f
C68 Y.n3 VSS 0.053224f
C69 Y.n4 VSS 0.413916f
C70 a_371_1047.t3 VSS 0.146522f
C71 a_371_1047.t1 VSS 0.146522f
C72 a_371_1047.t2 VSS 0.146522f
C73 a_371_1047.n0 VSS 0.486962f
C74 a_371_1047.t5 VSS 0.146522f
C75 a_371_1047.t4 VSS 0.146522f
C76 a_371_1047.n1 VSS 0.486962f
C77 a_371_1047.n2 VSS 2.86013f
C78 a_371_1047.n3 VSS 0.48681f
C79 a_371_1047.t0 VSS 0.146522f
.ends

