** sch_path: /home/erhangok/Documents/Dersler/VLSI/vlsi_sky130b/design/xschem/inv_TB.sch
**.subckt inv_TB OUTPUT
*.opin OUTPUT
V1 VDD GND 1.2
V2 VSS GND 0
V4 INPUT GND pulse(0,1.2,0.01u,1p,1p,0.01u,0.02u)
x1 VSS OUTPUT INPUT VDD inv
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice tt_mm




.control
set color0 = white

save all
tran 0.01n 0.03u
plot INPUT OUTPUT title 'a'

meas tran t_input when V(INPUT)=0.6 RISE=1
meas tran t_output when V(OUTPUT)=0.6 FALL=1
let tpdr = (t_output - t_input) * 1e9
echo (a) tpdr (ns) is:
print tpdr
meas tran t_input when V(INPUT)=0.6 FALL=1
meas tran t_output when V(OUTPUT)=0.6 RISE=1
let tpdf = (t_output - t_input) * 1e9
echo (a) tpdf (ns) is:
print tpdf
let tpd = (tpdf + tpdr)/2
echo (a) tpd (ns) is:
print tpd

.endc


**** end user architecture code
**.ends

* expanding   symbol:  inv.sym # of pins=4
** sym_path: /home/erhangok/Documents/Dersler/VLSI/vlsi_sky130b/design/xschem/inv.sym
** sch_path: /home/erhangok/Documents/Dersler/VLSI/vlsi_sky130b/design/xschem/inv.sch
.subckt inv VSS OUT IN VDD
*.iopin VDD
*.iopin VSS
*.iopin IN
*.iopin OUT
XM1 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT IN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
