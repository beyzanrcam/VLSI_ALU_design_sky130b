* NGSPICE file created from nor2_pex.ext - technology: sky130B

.subckt nor2 A B VSS VDD Y
X0 a_154_100.t1 B.t0 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.3103 pd=2.43 as=0.6206 ps=4.86 w=2.14 l=0.3
X1 a_1098_100.t1 A.t0 Y.t3 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.3103 pd=2.43 as=0.3103 ps=2.43 w=2.14 l=0.3
X2 Y.t1 A.t1 a_862_100.t1 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.3103 pd=2.43 as=0.3103 ps=2.43 w=2.14 l=0.3
X3 a_272_100.t1 B.t1 a_626_100.t1 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.3103 pd=2.43 as=0.3103 ps=2.43 w=2.14 l=0.3
X4 a_862_100.t0 A.t2 a_272_100.t5 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.3103 pd=2.43 as=0.3103 ps=2.43 w=2.14 l=0.3
X5 a_626_100.t0 B.t2 VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.3103 pd=2.43 as=0.3103 ps=2.43 w=2.14 l=0.3
X6 VDD.t4 B.t3 a_390_100.t0 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.3103 pd=2.43 as=0.3103 ps=2.43 w=2.14 l=0.3
X7 Y.t4 A.t3 a_1334_100.t1 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.6206 pd=4.86 as=0.3103 ps=2.43 w=2.14 l=0.3
X8 VSS.t3 A.t4 Y.t2 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.3
X9 a_390_100.t1 B.t4 a_272_100.t2 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.3103 pd=2.43 as=0.3103 ps=2.43 w=2.14 l=0.3
X10 Y.t0 B.t5 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.3
X11 a_1334_100.t0 A.t5 a_272_100.t4 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.3103 pd=2.43 as=0.3103 ps=2.43 w=2.14 l=0.3
X12 a_272_100.t0 B.t6 a_154_100.t0 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.3103 pd=2.43 as=0.3103 ps=2.43 w=2.14 l=0.3
X13 a_272_100.t3 A.t6 a_1098_100.t0 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.3103 pd=2.43 as=0.3103 ps=2.43 w=2.14 l=0.3
R0 B.n5 B.t5 535.899
R1 B.n2 B.t1 417.341
R2 B.n0 B.t0 417.341
R3 B.n3 B.t3 372.918
R4 B.n2 B.t2 372.918
R5 B.n0 B.t6 372.918
R6 B.n1 B.t4 372.918
R7 B B.n4 113.737
R8 B.n1 B.n0 44.424
R9 B.n3 B.n2 44.424
R10 B.n4 B.n3 16.1887
R11 B.n4 B.n1 15.0593
R12 B.n5 B 6.02403
R13 B B.n5 5.48621
R14 B.n5 B 4.75479
R15 VDD.n2 VDD.t9 158.858
R16 VDD.n2 VDD.n1 145.48
R17 VDD.t0 VDD.t11 110.01
R18 VDD.t10 VDD.t0 110.01
R19 VDD.t13 VDD.t10 110.01
R20 VDD.t14 VDD.t13 110.01
R21 VDD.t12 VDD.t14 110.01
R22 VDD.t7 VDD.t12 110.01
R23 VDD.t5 VDD.t7 110.01
R24 VDD.t3 VDD.t5 110.01
R25 VDD.t2 VDD.t3 110.01
R26 VDD.t1 VDD.t8 110.01
R27 VDD.n0 VDD.t1 78.3126
R28 VDD VDD.n0 47.4658
R29 VDD.n0 VDD.t2 31.6982
R30 VDD.n1 VDD.t6 13.3486
R31 VDD.n1 VDD.t4 13.3486
R32 VDD VDD.n2 0.0655794
R33 a_154_100.t0 a_154_100.t1 26.6968
R34 A.n0 A.t3 417.341
R35 A A.t4 384.558
R36 A.n4 A.t2 372.918
R37 A.n3 A.t1 372.918
R38 A.n2 A.t0 372.918
R39 A.n1 A.t6 372.918
R40 A.n0 A.t5 372.918
R41 A.n5 A.n4 65.5064
R42 A.n1 A.n0 44.424
R43 A.n2 A.n1 44.424
R44 A.n3 A.n2 44.424
R45 A.n4 A.n3 44.424
R46 A.n5 A 4.89462
R47 A A.n5 1.88285
R48 Y.n1 Y.t4 158.811
R49 Y.n1 Y.n0 145.726
R50 Y Y.n2 83.3758
R51 Y.n0 Y.t3 13.3486
R52 Y.n0 Y.t1 13.3486
R53 Y.n2 Y.t2 8.7005
R54 Y.n2 Y.t0 8.7005
R55 Y Y.n1 0.43199
R56 a_1098_100.t0 a_1098_100.t1 26.6968
R57 a_862_100.t0 a_862_100.t1 26.6968
R58 a_626_100.t0 a_626_100.t1 26.6968
R59 a_272_100.n3 a_272_100.n2 146.124
R60 a_272_100.n2 a_272_100.n0 146.123
R61 a_272_100.n2 a_272_100.n1 145.821
R62 a_272_100.n1 a_272_100.t5 13.3486
R63 a_272_100.n1 a_272_100.t1 13.3486
R64 a_272_100.n0 a_272_100.t4 13.3486
R65 a_272_100.n0 a_272_100.t3 13.3486
R66 a_272_100.n3 a_272_100.t2 13.3486
R67 a_272_100.t0 a_272_100.n3 13.3486
R68 a_390_100.t0 a_390_100.t1 26.6968
R69 a_1334_100.t0 a_1334_100.t1 26.6968
R70 VSS VSS.t0 974.856
R71 VSS.t0 VSS.t2 323.49
R72 VSS.n0 VSS.t3 41.6266
R73 VSS.n0 VSS.t1 41.3938
R74 VSS VSS.n0 0.023
C0 Y A 0.204858f
C1 B A 0.159179f
C2 VDD A 0.049461f
C3 Y B 0.019228f
C4 Y VDD 0.113724f
C5 B VDD 0.249656f
C6 Y VSS 1.05355f
C7 A VSS 0.788605f
C8 B VSS 0.907937f
C9 VDD VSS 5.18777f
.ends

