magic
tech sky130B
magscale 1 2
timestamp 1736620191
<< nwell >>
rect 22 787 20462 1687
<< poly >>
rect 18 709 131 729
rect -64 692 131 709
rect -64 658 -48 692
rect -14 658 131 692
rect -64 642 131 658
rect 18 620 131 642
rect 2509 708 2647 727
rect 2509 698 2732 708
rect 2509 647 2531 698
rect 2582 647 2732 698
rect 2509 637 2732 647
rect 5054 706 5259 719
rect 7687 708 7890 720
rect 5054 696 5339 706
rect 5054 648 5076 696
rect 5124 648 5339 696
rect 5054 638 5339 648
rect 7687 698 7974 708
rect 7687 646 7709 698
rect 7761 646 7974 698
rect 2509 618 2647 637
rect 5054 626 5259 638
rect 7687 636 7974 646
rect 10484 707 10669 719
rect 10484 697 10741 707
rect 10484 648 10500 697
rect 10549 648 10741 697
rect 10484 638 10741 648
rect 13072 703 13242 715
rect 16036 709 16194 721
rect 18845 711 19005 723
rect 13072 693 13316 703
rect 13072 651 13088 693
rect 13130 651 13316 693
rect 13072 641 13316 651
rect 16036 699 16279 709
rect 16036 645 16052 699
rect 16106 645 16279 699
rect 7687 624 7890 636
rect 10484 626 10669 638
rect 13072 629 13242 641
rect 16036 635 16279 645
rect 18845 701 19095 711
rect 18845 647 18861 701
rect 18915 647 19095 701
rect 18845 637 19095 647
rect 16036 623 16194 635
rect 18845 625 19005 637
<< polycont >>
rect -48 658 -14 692
rect 2531 647 2582 698
rect 5076 648 5124 696
rect 7709 646 7761 698
rect 10500 648 10549 697
rect 13088 651 13130 693
rect 16052 645 16106 699
rect 18861 647 18915 701
<< locali >>
rect 2531 708 2582 714
rect -48 697 -14 708
rect 5076 706 5124 712
rect 7709 708 7761 714
rect -48 642 -14 654
rect 10500 707 10549 713
rect 16052 709 16106 715
rect 18861 711 18915 717
rect 2531 631 2582 637
rect 5076 632 5124 638
rect 13088 703 13130 709
rect 7709 630 7761 636
rect 10500 632 10549 638
rect 13088 635 13130 641
rect 16052 629 16106 635
rect 18861 631 18915 637
<< viali >>
rect 2521 698 2592 708
rect -52 692 -9 697
rect -52 658 -48 692
rect -48 658 -14 692
rect -14 658 -9 692
rect -52 654 -9 658
rect 2521 647 2531 698
rect 2531 647 2582 698
rect 2582 647 2592 698
rect 2521 637 2592 647
rect 5066 696 5134 706
rect 5066 648 5076 696
rect 5076 648 5124 696
rect 5124 648 5134 696
rect 5066 638 5134 648
rect 7699 698 7771 708
rect 7699 646 7709 698
rect 7709 646 7761 698
rect 7761 646 7771 698
rect 7699 636 7771 646
rect 10490 697 10559 707
rect 10490 648 10500 697
rect 10500 648 10549 697
rect 10549 648 10559 697
rect 10490 638 10559 648
rect 13078 693 13140 703
rect 13078 651 13088 693
rect 13088 651 13130 693
rect 13130 651 13140 693
rect 13078 641 13140 651
rect 16042 699 16116 709
rect 16042 645 16052 699
rect 16052 645 16106 699
rect 16106 645 16116 699
rect 16042 635 16116 645
rect 18851 701 18925 711
rect 18851 647 18861 701
rect 18861 647 18915 701
rect 18915 647 18925 701
rect 18851 637 18925 647
<< metal1 >>
rect -239 608 -147 1756
rect -64 697 21 1756
rect 2386 720 2472 1756
rect 2521 720 2592 1756
rect -64 654 -52 697
rect -9 654 21 697
rect -64 642 21 654
rect -239 465 143 608
rect 1343 504 1603 641
rect 1510 -77 1603 504
rect 2387 576 2471 720
rect 2509 708 2604 720
rect 2509 637 2521 708
rect 2592 637 2604 708
rect 2509 631 2604 637
rect 2387 492 2733 576
rect 3979 492 4286 596
rect 4182 -77 4286 492
rect 4905 581 4999 1756
rect 5054 706 5146 1756
rect 5054 638 5066 706
rect 5134 638 5146 706
rect 5054 632 5146 638
rect 4905 487 5347 581
rect 6597 512 6845 598
rect 6759 -77 6845 512
rect 7510 580 7602 1756
rect 7687 708 7783 1756
rect 7687 636 7699 708
rect 7771 636 7783 708
rect 7687 624 7783 636
rect 7510 488 7979 580
rect 9232 518 9532 601
rect 9449 -77 9532 518
rect 10354 579 10443 1756
rect 10484 707 10570 1756
rect 10484 638 10490 707
rect 10559 638 10570 707
rect 10484 626 10570 638
rect 10354 490 10746 579
rect 11997 514 12274 603
rect 12185 -77 12274 514
rect 12943 578 13030 1756
rect 13072 703 13152 1756
rect 13072 641 13078 703
rect 13140 641 13152 703
rect 13072 629 13152 641
rect 12943 491 13324 578
rect 14573 505 14897 600
rect 14802 -77 14897 505
rect 15869 580 15960 1756
rect 16036 709 16128 1756
rect 16036 635 16042 709
rect 16116 635 16128 709
rect 16036 623 16128 635
rect 15869 489 16283 580
rect 17533 508 17838 597
rect 17749 -77 17838 508
rect 18682 586 18781 1756
rect 18845 711 18937 1756
rect 18845 637 18851 711
rect 18925 637 18937 711
rect 18845 625 18937 637
rect 18682 487 19103 586
rect 20355 509 20622 585
rect 20546 -77 20622 509
<< metal4 >>
rect 146 1519 20338 1645
<< metal5 >>
rect 505 1 19917 394
use XOR2  XOR2_0
timestamp 1736620191
transform 1 0 19091 0 1 -77
box -109 77 1371 1764
use XOR2  XOR2_1
timestamp 1736620191
transform 1 0 109 0 1 -77
box -109 77 1371 1764
use XOR2  XOR2_2
timestamp 1736620191
transform 1 0 2729 0 1 -79
box -109 77 1371 1764
use XOR2  XOR2_3
timestamp 1736620191
transform 1 0 5338 0 1 -79
box -109 77 1371 1764
use XOR2  XOR2_4
timestamp 1736620191
transform 1 0 7971 0 1 -79
box -109 77 1371 1764
use XOR2  XOR2_5
timestamp 1736620191
transform 1 0 10739 0 1 -79
box -109 77 1371 1764
use XOR2  XOR2_6
timestamp 1736620191
transform 1 0 13318 0 1 -79
box -109 77 1371 1764
use XOR2  XOR2_7
timestamp 1736620191
transform 1 0 16275 0 1 -79
box -109 77 1371 1764
<< labels >>
flabel metal1 -235 1689 -156 1751 0 FreeSans 160 0 0 0 B7
port 1 nsew
flabel metal1 -53 1696 4 1742 0 FreeSans 160 0 0 0 A7
port 3 nsew
flabel metal1 2529 1704 2586 1750 0 FreeSans 160 0 0 0 A6
port 4 nsew
flabel metal1 5070 1698 5127 1744 0 FreeSans 160 0 0 0 A5
port 5 nsew
flabel metal1 7702 1696 7759 1742 0 FreeSans 160 0 0 0 A4
port 6 nsew
flabel metal1 10495 1702 10552 1748 0 FreeSans 160 0 0 0 A3
port 7 nsew
flabel metal1 13081 1701 13138 1747 0 FreeSans 160 0 0 0 A2
port 8 nsew
flabel metal1 16051 1700 16108 1746 0 FreeSans 160 0 0 0 A1
port 9 nsew
flabel metal1 18859 1699 18916 1745 0 FreeSans 160 0 0 0 A0
port 10 nsew
flabel metal1 18703 1698 18760 1744 0 FreeSans 160 0 0 0 B0
port 11 nsew
flabel metal1 15884 1702 15941 1748 0 FreeSans 160 0 0 0 B1
port 12 nsew
flabel metal1 12956 1699 13013 1745 0 FreeSans 160 0 0 0 B2
port 13 nsew
flabel metal1 10370 1704 10427 1750 0 FreeSans 160 0 0 0 B3
port 14 nsew
flabel metal1 7525 1698 7582 1744 0 FreeSans 160 0 0 0 B4
port 15 nsew
flabel metal1 4921 1699 4978 1745 0 FreeSans 160 0 0 0 B5
port 16 nsew
flabel metal1 2399 1702 2456 1748 0 FreeSans 160 0 0 0 B6
port 17 nsew
flabel metal1 1525 -65 1582 -19 0 FreeSans 160 0 0 0 S7
port 18 nsew
flabel metal1 4206 -63 4263 -17 0 FreeSans 160 0 0 0 S6
port 19 nsew
flabel metal1 6774 -70 6831 -24 0 FreeSans 160 0 0 0 S5
port 20 nsew
flabel metal1 9464 -67 9521 -21 0 FreeSans 160 0 0 0 S4
port 21 nsew
flabel metal1 12200 -70 12257 -24 0 FreeSans 160 0 0 0 S3
port 22 nsew
flabel metal1 14824 -63 14881 -17 0 FreeSans 160 0 0 0 S2
port 23 nsew
flabel metal1 17763 -68 17820 -22 0 FreeSans 160 0 0 0 S1
port 24 nsew
flabel metal1 20558 -66 20615 -20 0 FreeSans 160 0 0 0 S0
port 25 nsew
<< end >>
