** sch_path: /home/ubuntu/Desktop/examples/xschem/inv_TB.sch
**.subckt inv_TB
V2 VDD GND 1.8
V1 A GND pulse 0 1.8 2n 1n 1n 10n 20n
x2 A VDD Y GND inv
**** begin user architecture code



.include ../mag/inv_pex.spice

.options KEEPOPINFO

.control

save all

tran 0.1n 200n
write inv_TB.raw

.endc



** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends
.GLOBAL GND
.end
