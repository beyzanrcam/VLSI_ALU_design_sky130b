magic
tech sky130B
magscale 1 2
timestamp 1736026236
<< nwell >>
rect 1387 1327 1465 1856
rect 1380 1223 1465 1327
rect 1380 1034 1488 1223
rect 1380 1019 1465 1034
rect 1387 906 1465 1019
rect 1387 881 1469 906
<< metal1 >>
rect 65 1090 71 1142
rect 123 1090 129 1142
rect -5 866 -2 875
rect 1312 840 1321 906
rect 1387 840 1393 906
rect 3943 870 3947 885
rect -5 773 -2 782
rect -5 681 -2 690
rect -5 586 -2 595
rect -5 450 1 516
rect 67 450 73 516
rect 3377 503 3429 509
rect 3377 445 3429 451
rect -5 349 1 415
rect 67 349 73 415
rect -5 248 1 314
rect 67 248 73 314
rect -5 154 1 220
rect 67 154 73 220
rect 725 107 777 113
rect 725 49 777 55
rect 2193 107 2258 114
rect 2193 55 2199 107
rect 2251 55 2258 107
rect 2193 49 2258 55
<< via1 >>
rect 3084 1399 3136 1451
rect 71 1090 123 1142
rect 1541 1087 1593 1139
rect 2877 945 2943 1011
rect 1321 840 1387 906
rect 1471 840 1537 906
rect 1567 746 1633 812
rect 1673 652 1739 718
rect 1773 558 1839 624
rect 1 450 67 516
rect 3377 451 3429 503
rect 1 349 67 415
rect 1 248 67 314
rect 1 154 67 220
rect 725 55 777 107
rect 2199 55 2251 107
<< metal2 >>
rect 3062 1453 3160 1475
rect 3062 1397 3082 1453
rect 3138 1397 3160 1453
rect 3062 1378 3160 1397
rect 53 1144 142 1157
rect 53 1088 69 1144
rect 125 1088 142 1144
rect 53 1074 142 1088
rect 1525 1141 1609 1152
rect 1525 1085 1539 1141
rect 1595 1085 1609 1141
rect 1525 1071 1609 1085
rect 2871 945 2877 1011
rect 2943 945 2949 1011
rect 1312 840 1321 906
rect 1387 840 1396 906
rect 1465 840 1471 906
rect 1537 840 1543 906
rect 1467 516 1533 840
rect 1561 746 1567 812
rect 1633 746 1639 812
rect -5 450 1 516
rect 67 450 1533 516
rect 1567 415 1633 746
rect 1667 652 1673 718
rect 1739 652 1745 718
rect -5 349 1 415
rect 67 349 1633 415
rect 1673 314 1739 652
rect 1767 558 1773 624
rect 1839 558 1845 624
rect -5 248 1 314
rect 67 248 1739 314
rect 1769 220 1835 558
rect 3355 505 3452 522
rect 3355 449 3375 505
rect 3431 449 3452 505
rect 3355 428 3452 449
rect -5 154 1 220
rect 67 154 1835 220
rect 702 109 798 123
rect 702 53 723 109
rect 779 53 798 109
rect 702 27 798 53
rect 2176 109 2273 128
rect 2176 53 2197 109
rect 2253 53 2273 109
rect 2176 33 2273 53
<< via2 >>
rect 3082 1451 3138 1453
rect 3082 1399 3084 1451
rect 3084 1399 3136 1451
rect 3136 1399 3138 1451
rect 3082 1397 3138 1399
rect 69 1142 125 1144
rect 69 1090 71 1142
rect 71 1090 123 1142
rect 123 1090 125 1142
rect 69 1088 125 1090
rect 1539 1139 1595 1141
rect 1539 1087 1541 1139
rect 1541 1087 1593 1139
rect 1593 1087 1595 1139
rect 1539 1085 1595 1087
rect 2882 950 2938 1006
rect 1321 840 1387 906
rect 3375 503 3431 505
rect 3375 451 3377 503
rect 3377 451 3429 503
rect 3429 451 3431 503
rect 3375 449 3431 451
rect 723 107 779 109
rect 723 55 725 107
rect 725 55 777 107
rect 777 55 779 107
rect 723 53 779 55
rect 2197 107 2253 109
rect 2197 55 2199 107
rect 2199 55 2251 107
rect 2251 55 2253 107
rect 2197 53 2253 55
<< metal3 >>
rect 3051 1458 3176 1482
rect 3051 1392 3077 1458
rect 3143 1392 3176 1458
rect 3051 1370 3176 1392
rect 35 1149 160 1167
rect 35 1083 64 1149
rect 130 1083 160 1149
rect 35 1055 160 1083
rect 1503 1146 1628 1168
rect 1503 1080 1534 1146
rect 1600 1080 1628 1146
rect 1503 1056 1628 1080
rect 2877 1006 2943 1011
rect 2877 950 2882 1006
rect 2938 950 2943 1006
rect 1316 906 1392 911
rect 2877 906 2943 950
rect 1316 840 1321 906
rect 1387 840 2943 906
rect 1316 835 1392 840
rect 3347 510 3452 522
rect 3347 444 3370 510
rect 3436 444 3452 510
rect 3347 428 3452 444
rect 696 114 814 132
rect 696 48 718 114
rect 784 48 814 114
rect 696 17 814 48
rect 2170 114 2273 128
rect 2170 48 2192 114
rect 2258 48 2273 114
rect 2170 33 2273 48
<< via3 >>
rect 3077 1453 3143 1458
rect 3077 1397 3082 1453
rect 3082 1397 3138 1453
rect 3138 1397 3143 1453
rect 3077 1392 3143 1397
rect 64 1144 130 1149
rect 64 1088 69 1144
rect 69 1088 125 1144
rect 125 1088 130 1144
rect 64 1083 130 1088
rect 1534 1141 1600 1146
rect 1534 1085 1539 1141
rect 1539 1085 1595 1141
rect 1595 1085 1600 1141
rect 1534 1080 1600 1085
rect 3370 505 3436 510
rect 3370 449 3375 505
rect 3375 449 3431 505
rect 3431 449 3436 505
rect 3370 444 3436 449
rect 718 109 784 114
rect 718 53 723 109
rect 723 53 779 109
rect 779 53 784 109
rect 718 48 784 53
rect 2192 109 2258 114
rect 2192 53 2197 109
rect 2197 53 2253 109
rect 2253 53 2258 109
rect 2192 48 2258 53
<< metal4 >>
rect 2597 1458 3192 1515
rect 2597 1392 3077 1458
rect 3143 1392 3192 1458
rect 2597 1342 3192 1392
rect 2597 1203 2770 1342
rect 31 1149 2770 1203
rect 31 1083 64 1149
rect 130 1146 2770 1149
rect 130 1083 1534 1146
rect 31 1080 1534 1083
rect 1600 1080 2770 1146
rect 31 1030 2770 1080
<< via4 >>
rect 3267 510 3539 613
rect 3267 444 3370 510
rect 3370 444 3436 510
rect 3436 444 3539 510
rect 3267 341 3539 444
rect 615 114 887 217
rect 615 48 718 114
rect 718 48 784 114
rect 784 48 887 114
rect 615 -55 887 48
rect 2089 114 2361 217
rect 2089 48 2192 114
rect 2192 48 2258 114
rect 2258 48 2361 114
rect 2089 -55 2361 48
<< metal5 >>
rect 3243 613 3563 637
rect 3243 341 3267 613
rect 3539 341 3563 613
rect 3243 241 3563 341
rect 591 217 3563 241
rect 591 -55 615 217
rect 887 -55 2089 217
rect 2361 -55 3563 217
rect 591 -79 3563 -55
use nor2  nor2_0 ~/Documents/Dersler/VLSI/vlsi_sky130b/design/mag/NOR/NOR2
timestamp 1736020690
transform 1 0 2857 0 1 942
box 0 -480 1090 580
use nor4  nor4_0 ~/Documents/Dersler/VLSI/vlsi_sky130b/design/mag/NOR/NOR4
timestamp 1736019943
transform 1 0 2067 0 1 -110
box -602 118 790 1966
use nor4  nor4_1
timestamp 1736019943
transform 1 0 597 0 1 -110
box -602 118 790 1966
<< labels >>
rlabel metal1 -5 872 -5 872 3 A0
port 1 e
rlabel metal1 -5 780 -5 780 3 A1
port 2 e
rlabel metal1 -5 687 -5 687 3 A2
port 3 e
rlabel metal1 -5 591 -5 591 3 A3
port 4 e
rlabel metal1 -5 479 -5 479 3 A4
port 5 e
rlabel metal1 -5 380 -5 380 3 A5
port 6 e
rlabel metal1 -5 279 -5 279 3 A6
port 7 e
rlabel metal1 -5 182 -5 182 3 A7
port 8 e
rlabel metal5 2271 -79 2271 -79 5 VSS
rlabel metal4 1424 1203 1424 1203 5 VDD
rlabel metal1 3947 879 3947 879 3 Y
port 11 e
<< end >>
