magic
tech sky130B
magscale 1 2
timestamp 1733168276
<< nwell >>
rect -37 954 861 1400
rect -37 916 765 954
<< nmos >>
rect 62 88 92 488
rect 158 88 188 488
rect 254 88 284 488
rect 350 88 380 488
rect 446 88 476 488
rect 542 88 572 488
rect 638 88 668 488
rect 734 88 764 488
<< pmos >>
rect 61 1016 91 1338
rect 157 1016 187 1338
rect 253 1016 283 1338
rect 349 1016 379 1338
rect 445 1016 475 1338
rect 541 1016 571 1338
rect 637 1016 667 1338
rect 733 1016 763 1338
<< ndiff >>
rect 0 476 62 488
rect 0 100 12 476
rect 46 100 62 476
rect 0 88 62 100
rect 92 88 158 488
rect 188 88 254 488
rect 284 88 350 488
rect 380 476 446 488
rect 380 100 396 476
rect 430 100 446 476
rect 380 88 446 100
rect 476 88 542 488
rect 572 88 638 488
rect 668 88 734 488
rect 764 476 826 488
rect 764 100 780 476
rect 814 100 826 476
rect 764 88 826 100
<< pdiff >>
rect -1 1326 61 1338
rect -1 1028 11 1326
rect 45 1028 61 1326
rect -1 1016 61 1028
rect 91 1326 157 1338
rect 91 1028 107 1326
rect 141 1028 157 1326
rect 91 1016 157 1028
rect 187 1326 253 1338
rect 187 1028 203 1326
rect 237 1028 253 1326
rect 187 1016 253 1028
rect 283 1326 349 1338
rect 283 1028 299 1326
rect 333 1028 349 1326
rect 283 1016 349 1028
rect 379 1326 445 1338
rect 379 1028 395 1326
rect 429 1028 445 1326
rect 379 1016 445 1028
rect 475 1326 541 1338
rect 475 1028 491 1326
rect 525 1028 541 1326
rect 475 1016 541 1028
rect 571 1326 637 1338
rect 571 1028 587 1326
rect 621 1028 637 1326
rect 571 1016 637 1028
rect 667 1326 733 1338
rect 667 1028 683 1326
rect 717 1028 733 1326
rect 667 1016 733 1028
rect 763 1326 825 1338
rect 763 1028 779 1326
rect 813 1028 825 1326
rect 763 1016 825 1028
<< ndiffc >>
rect 12 100 46 476
rect 396 100 430 476
rect 780 100 814 476
<< pdiffc >>
rect 11 1028 45 1326
rect 107 1028 141 1326
rect 203 1028 237 1326
rect 299 1028 333 1326
rect 395 1028 429 1326
rect 491 1028 525 1326
rect 587 1028 621 1326
rect 683 1028 717 1326
rect 779 1028 813 1326
<< poly >>
rect 61 1338 91 1364
rect 157 1338 187 1364
rect 253 1338 283 1364
rect 349 1338 379 1364
rect 445 1338 475 1364
rect 541 1338 571 1364
rect 637 1338 667 1364
rect 733 1338 763 1364
rect 61 985 91 1016
rect 157 985 187 1016
rect 253 986 283 1016
rect 31 969 187 985
rect 31 935 59 969
rect 93 935 187 969
rect 31 919 187 935
rect 235 985 303 986
rect 349 985 379 1016
rect 445 985 475 1016
rect 541 985 571 1016
rect 637 985 667 1016
rect 733 985 763 1016
rect 235 969 379 985
rect 235 935 251 969
rect 285 935 379 969
rect 235 919 379 935
rect 427 969 571 985
rect 427 935 443 969
rect 477 935 571 969
rect 427 919 571 935
rect 619 969 763 985
rect 619 935 635 969
rect 669 935 763 969
rect 619 919 763 935
rect 31 522 100 919
rect 235 870 303 919
rect 158 779 303 870
rect 158 745 174 779
rect 208 745 303 779
rect 158 738 303 745
rect 158 732 216 738
rect 157 730 216 732
rect 62 488 92 522
rect 157 508 212 730
rect 254 674 572 696
rect 254 638 344 674
rect 442 638 572 674
rect 254 627 572 638
rect 158 488 188 508
rect 254 488 284 627
rect 350 569 476 585
rect 350 530 385 569
rect 439 530 476 569
rect 350 514 476 530
rect 350 488 380 514
rect 446 488 476 514
rect 542 488 572 627
rect 638 488 668 514
rect 734 488 764 514
rect 62 62 92 88
rect 0 44 106 62
rect 158 48 188 88
rect 254 62 284 88
rect 350 61 380 88
rect 446 61 476 88
rect 542 62 572 88
rect 638 48 668 88
rect 734 62 764 88
rect 720 48 826 62
rect 0 -76 20 44
rect 87 -53 106 44
rect 148 36 214 48
rect 148 2 164 36
rect 198 19 214 36
rect 612 36 678 48
rect 612 19 628 36
rect 198 2 628 19
rect 662 2 678 36
rect 148 -11 678 2
rect 720 44 827 48
rect 720 -53 741 44
rect 87 -76 741 -53
rect 808 -76 827 44
rect 0 -94 827 -76
<< polycont >>
rect 59 935 93 969
rect 251 935 285 969
rect 443 935 477 969
rect 635 935 669 969
rect 174 745 208 779
rect 344 638 442 674
rect 385 530 439 569
rect 20 -76 87 44
rect 164 2 198 36
rect 628 2 662 36
rect 741 -76 808 44
<< locali >>
rect 11 1326 45 1342
rect 107 1326 141 1342
rect 11 1012 45 1028
rect 107 1012 141 1023
rect 203 1326 237 1342
rect 203 1012 237 1028
rect 299 1326 333 1342
rect 395 1326 429 1342
rect 299 1012 333 1023
rect 395 1012 429 1028
rect 491 1326 525 1342
rect 587 1326 621 1342
rect 491 1012 525 1023
rect 587 1012 621 1028
rect 683 1326 717 1342
rect 779 1326 813 1342
rect 683 1012 717 1023
rect 779 1012 813 1028
rect 235 969 300 974
rect 43 935 59 969
rect 93 935 110 969
rect 235 935 251 969
rect 285 935 301 969
rect 427 935 443 969
rect 477 935 493 969
rect 619 935 635 969
rect 669 935 685 969
rect 43 884 110 935
rect 42 813 746 884
rect 63 526 114 813
rect 12 476 46 492
rect 12 84 46 100
rect 80 50 114 526
rect 0 44 114 50
rect 0 -76 20 44
rect 87 -53 114 44
rect 148 745 174 779
rect 208 745 678 779
rect 148 725 678 745
rect 148 48 300 725
rect 334 674 458 691
rect 334 638 344 674
rect 442 638 458 674
rect 334 621 458 638
rect 350 530 385 569
rect 439 530 476 569
rect 396 476 430 492
rect 396 84 430 100
rect 594 48 678 725
rect 148 36 678 48
rect 148 2 164 36
rect 198 2 628 36
rect 662 2 678 36
rect 148 -11 678 2
rect 712 48 746 813
rect 780 476 814 492
rect 780 84 814 100
rect 712 44 827 48
rect 712 -53 741 44
rect 87 -76 741 -53
rect 808 -76 827 44
rect 0 -94 827 -76
<< viali >>
rect 11 1213 45 1323
rect 106 1028 107 1135
rect 107 1028 141 1135
rect 106 1023 141 1028
rect 203 1213 237 1323
rect 395 1213 429 1323
rect 299 1028 333 1135
rect 333 1028 334 1135
rect 299 1023 334 1028
rect 587 1213 621 1323
rect 491 1028 525 1135
rect 525 1028 526 1135
rect 491 1023 526 1028
rect 779 1213 813 1323
rect 683 1028 717 1135
rect 717 1028 718 1135
rect 683 1023 718 1028
rect 59 935 93 969
rect 251 935 285 969
rect 443 935 477 969
rect 635 935 669 969
rect 12 100 46 476
rect 174 745 208 779
rect 344 638 442 674
rect 385 530 439 569
rect 396 100 430 476
rect 780 100 814 476
<< metal1 >>
rect -1 1335 826 1400
rect -1 1323 825 1335
rect -1 1213 11 1323
rect 45 1213 203 1323
rect 237 1213 395 1323
rect 429 1213 587 1323
rect 621 1213 779 1323
rect 813 1213 825 1323
rect -1 1204 825 1213
rect -1 1135 861 1150
rect -1 1023 106 1135
rect 141 1023 299 1135
rect 334 1023 491 1135
rect 526 1023 683 1135
rect 718 1023 861 1135
rect -1 1016 861 1023
rect -37 969 110 975
rect -37 935 59 969
rect 93 935 110 969
rect -37 813 110 935
rect 235 974 298 975
rect 235 969 300 974
rect 235 935 251 969
rect 285 935 300 969
rect 235 785 300 935
rect 427 969 493 985
rect 427 935 443 969
rect 477 935 493 969
rect -37 779 301 785
rect -37 745 174 779
rect 208 745 301 779
rect -37 716 301 745
rect 427 688 493 935
rect -37 674 493 688
rect -37 638 344 674
rect 442 638 493 674
rect -37 619 493 638
rect 521 969 681 985
rect 521 935 635 969
rect 669 935 681 969
rect 521 918 681 935
rect 521 591 587 918
rect 710 890 861 1016
rect -37 569 587 591
rect -37 530 385 569
rect 439 530 587 569
rect -37 522 587 530
rect 615 625 861 890
rect 615 488 746 625
rect 0 476 362 488
rect 0 100 12 476
rect 46 100 362 476
rect 0 21 362 100
rect 390 476 746 488
rect 390 100 396 476
rect 430 100 746 476
rect 390 88 746 100
rect 774 476 827 488
rect 774 100 780 476
rect 814 100 827 476
rect 774 21 827 100
rect 0 -94 827 21
<< labels >>
rlabel metal1 -37 813 -4 882 7 A
port 1 w
rlabel metal1 -37 716 -5 785 7 B
port 2 w
rlabel metal1 -37 619 -4 688 7 C
port 3 w
rlabel metal1 -37 522 -5 591 7 D
port 4 w
rlabel metal1 0 -94 827 21 5 VSS
port 5 s
rlabel metal1 -1 1366 826 1400 5 VDD
port 6 n
rlabel metal1 815 625 861 1150 5 Y
port 7 e
<< end >>
