* NGSPICE file created from nor3_pex.ext - technology: sky130B

.subckt nor3 A B C VSS VDD Y
X0 a_n77_875.t2 A.t0 VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.52965 pd=3.54 as=0.52965 ps=3.54 w=3.21 l=0.15
X1 Y.t2 A.t1 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X2 VDD.t4 A.t2 a_n77_875.t1 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.52965 pd=3.54 as=0.52965 ps=3.54 w=3.21 l=0.15
X3 VSS.t5 B.t0 Y.t4 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X4 Y.t0 C.t0 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X5 a_n77_875.t0 A.t3 VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.52965 pd=3.54 as=0.9951 ps=7.04 w=3.21 l=0.15
X6 a_211_875.t2 B.t1 a_n77_875.t4 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.52965 pd=3.54 as=0.52965 ps=3.54 w=3.21 l=0.15
X7 a_n77_875.t3 B.t2 a_211_875.t1 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.52965 pd=3.54 as=0.52965 ps=3.54 w=3.21 l=0.15
X8 a_211_875.t0 B.t3 a_n77_875.t5 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.52965 pd=3.54 as=0.52965 ps=3.54 w=3.21 l=0.15
X9 a_211_875.t5 C.t1 Y.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.52965 pd=3.54 as=0.52965 ps=3.54 w=3.21 l=0.15
X10 Y.t5 C.t2 a_211_875.t4 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.9951 pd=7.04 as=0.52965 ps=3.54 w=3.21 l=0.15
X11 Y.t3 C.t3 a_211_875.t3 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.52965 pd=3.54 as=0.52965 ps=3.54 w=3.21 l=0.15
R0 A.n0 A.t3 719.788
R1 A.n2 A.t1 696.418
R2 A.n1 A.t0 576.501
R3 A.n0 A.t2 565.548
R4 A A.n2 162.031
R5 A.n1 A.n0 72.3005
R6 A.n2 A.n1 34.3247
R7 VDD.n1 VDD.t2 138.853
R8 VDD.n1 VDD.n0 128.728
R9 VDD.n4 VDD.n3 123.334
R10 VDD.t0 VDD.t11 94.0211
R11 VDD.t9 VDD.t0 94.0211
R12 VDD.t10 VDD.t9 94.0211
R13 VDD.t7 VDD.t10 94.0211
R14 VDD.t8 VDD.t7 94.0211
R15 VDD.t5 VDD.t8 94.0211
R16 VDD.t3 VDD.t5 94.0211
R17 VDD.n3 VDD.t1 61.7015
R18 VDD.n3 VDD.t3 32.3201
R19 VDD.n0 VDD.t6 10.1267
R20 VDD.n0 VDD.t4 10.1267
R21 VDD.n5 VDD.n4 3.1005
R22 VDD.n5 VDD.n1 0.0801569
R23 VDD.n4 VDD.n2 0.0144891
R24 VDD VDD.n5 0.00111275
R25 a_n77_875.n2 a_n77_875.n1 132.536
R26 a_n77_875.n2 a_n77_875.n0 132.536
R27 a_n77_875.n3 a_n77_875.n2 132.454
R28 a_n77_875.n1 a_n77_875.t1 10.1267
R29 a_n77_875.n1 a_n77_875.t0 10.1267
R30 a_n77_875.n0 a_n77_875.t5 10.1267
R31 a_n77_875.n0 a_n77_875.t3 10.1267
R32 a_n77_875.n3 a_n77_875.t4 10.1267
R33 a_n77_875.t2 a_n77_875.n3 10.1267
R34 VSS.t4 VSS.t0 606.898
R35 VSS.n2 VSS.t2 543.678
R36 VSS VSS.t3 153.87
R37 VSS.n4 VSS.n0 130.333
R38 VSS.n4 VSS.n3 73.1255
R39 VSS.n3 VSS.n2 73.1255
R40 VSS.n2 VSS.t4 63.2189
R41 VSS.n3 VSS.n1 44.0502
R42 VSS.n0 VSS.t1 19.8005
R43 VSS.n0 VSS.t5 19.8005
R44 VSS VSS.n4 3.364
R45 Y.n1 Y.t5 142.603
R46 Y.n1 Y.n0 132.513
R47 Y.n3 Y.t0 86.1172
R48 Y.n3 Y.n2 66.4372
R49 Y.n2 Y.t4 19.8005
R50 Y.n2 Y.t2 19.8005
R51 Y.n0 Y.t1 10.1267
R52 Y.n0 Y.t3 10.1267
R53 Y Y.n3 0.264151
R54 Y Y.n1 0.195401
R55 B.n0 B.t3 719.788
R56 B.n0 B.t1 719.788
R57 B.n0 B.t2 565.548
R58 B.n1 B.t0 435.408
R59 B.n1 B.n0 178.34
R60 B B.n1 162.44
R61 C.n0 C.t2 719.788
R62 C.n1 C.t3 565.548
R63 C.n0 C.t1 565.548
R64 C.n2 C.n1 456.293
R65 C.n2 C.t0 218.799
R66 C C.n2 162.656
R67 C.n1 C.n0 154.24
R68 a_211_875.n2 a_211_875.n0 128.767
R69 a_211_875.n3 a_211_875.n2 128.767
R70 a_211_875.n2 a_211_875.n1 128.69
R71 a_211_875.n1 a_211_875.t3 10.1267
R72 a_211_875.n1 a_211_875.t0 10.1267
R73 a_211_875.n0 a_211_875.t4 10.1267
R74 a_211_875.n0 a_211_875.t5 10.1267
R75 a_211_875.n3 a_211_875.t1 10.1267
R76 a_211_875.t2 a_211_875.n3 10.1267
C0 B C 0.471635f
C1 B A 0.652088f
C2 Y C 0.416086f
C3 A Y 0.012402f
C4 B VDD 0.033186f
C5 A C 0.017562f
C6 VDD Y 0.070002f
C7 VDD C 0.024197f
C8 A VDD 0.121157f
C9 B Y 0.030731f
C10 Y VSS 1.06787f
C11 C VSS 0.561586f
C12 B VSS 0.345794f
C13 A VSS 0.43138f
C14 VDD VSS 3.30718f
.ends

