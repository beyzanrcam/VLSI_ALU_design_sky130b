magic
tech sky130B
magscale 1 2
timestamp 1734016331
<< nwell >>
rect -37 -16 1286 559
<< nmos >>
rect 578 -339 608 -139
rect 674 -339 704 -139
<< pmos >>
rect 98 100 128 314
rect 194 100 224 314
rect 290 100 320 314
rect 386 100 416 314
rect 482 100 512 314
rect 578 100 608 314
rect 674 100 704 314
rect 770 100 800 314
rect 866 100 896 314
rect 962 100 992 314
rect 1058 100 1088 314
rect 1154 100 1184 314
<< ndiff >>
rect 516 -151 578 -139
rect 516 -327 528 -151
rect 562 -327 578 -151
rect 516 -339 578 -327
rect 608 -151 674 -139
rect 608 -327 624 -151
rect 658 -327 674 -151
rect 608 -339 674 -327
rect 704 -151 766 -139
rect 704 -327 720 -151
rect 754 -327 766 -151
rect 704 -339 766 -327
<< pdiff >>
rect 36 302 98 314
rect 36 112 48 302
rect 82 112 98 302
rect 36 100 98 112
rect 128 100 194 314
rect 224 302 290 314
rect 224 112 240 302
rect 274 112 290 302
rect 224 100 290 112
rect 320 100 386 314
rect 416 302 482 314
rect 416 112 432 302
rect 466 112 482 302
rect 416 100 482 112
rect 512 100 578 314
rect 608 302 674 314
rect 608 112 624 302
rect 658 112 674 302
rect 608 100 674 112
rect 704 100 770 314
rect 800 302 866 314
rect 800 112 816 302
rect 850 112 866 302
rect 800 100 866 112
rect 896 100 962 314
rect 992 302 1058 314
rect 992 112 1008 302
rect 1042 112 1058 302
rect 992 100 1058 112
rect 1088 100 1154 314
rect 1184 302 1246 314
rect 1184 112 1200 302
rect 1234 112 1246 302
rect 1184 100 1246 112
<< ndiffc >>
rect 528 -327 562 -151
rect 624 -327 658 -151
rect 720 -327 754 -151
<< pdiffc >>
rect 48 112 82 302
rect 240 112 274 302
rect 432 112 466 302
rect 624 112 658 302
rect 816 112 850 302
rect 1008 112 1042 302
rect 1200 112 1234 302
<< psubdiff >>
rect 516 -430 766 -394
rect 516 -494 563 -430
rect 725 -494 766 -430
rect 516 -527 766 -494
<< nsubdiff >>
rect 46 481 466 523
rect 46 430 89 481
rect 257 430 466 481
rect 46 392 466 430
<< psubdiffcont >>
rect 563 -494 725 -430
<< nsubdiffcont >>
rect 89 430 257 481
<< poly >>
rect 98 314 128 340
rect 194 314 224 340
rect 290 314 320 340
rect 386 314 416 340
rect 482 314 512 340
rect 578 314 608 340
rect 674 314 704 340
rect 770 314 800 340
rect 866 314 896 340
rect 962 314 992 340
rect 1058 314 1088 340
rect 1154 314 1184 340
rect 98 69 128 100
rect 194 69 224 100
rect 290 69 320 100
rect 386 69 416 100
rect 482 69 512 100
rect 578 69 608 100
rect 98 53 608 69
rect 98 19 480 53
rect 514 19 608 53
rect 98 3 608 19
rect 578 -139 608 3
rect 674 69 704 100
rect 770 69 800 100
rect 866 69 896 100
rect 962 69 992 100
rect 1058 69 1088 100
rect 1154 69 1184 100
rect 674 3 1184 69
rect 674 -39 704 3
rect 656 -55 722 -39
rect 656 -89 672 -55
rect 706 -89 722 -55
rect 656 -105 722 -89
rect 674 -139 704 -105
rect 578 -365 608 -339
rect 674 -365 704 -339
<< polycont >>
rect 480 19 514 53
rect 672 -89 706 -55
<< locali >>
rect 46 481 466 501
rect 46 430 89 481
rect 257 430 466 481
rect 46 411 466 430
rect 48 302 82 411
rect 48 96 82 112
rect 240 302 274 318
rect 240 96 274 112
rect 432 302 466 411
rect 432 96 466 112
rect 624 302 658 318
rect 624 96 658 112
rect 816 302 850 318
rect 816 96 850 112
rect 1008 302 1042 318
rect 1008 96 1042 112
rect 1200 302 1234 318
rect 1200 96 1234 112
rect 464 19 480 53
rect 514 19 530 53
rect 656 -89 672 -55
rect 706 -89 722 -55
rect 528 -151 562 -135
rect 528 -410 562 -327
rect 624 -151 658 -135
rect 624 -343 658 -327
rect 720 -151 754 -135
rect 720 -410 754 -327
rect 516 -430 766 -410
rect 516 -494 563 -430
rect 725 -494 766 -430
rect 516 -512 766 -494
<< viali >>
rect 48 112 82 302
rect 240 112 274 302
rect 432 112 466 302
rect 624 112 658 302
rect 816 112 850 302
rect 1008 112 1042 302
rect 1200 112 1234 302
rect 480 19 514 53
rect 672 -89 706 -55
rect 624 -327 658 -151
<< metal1 >>
rect 234 362 1048 421
rect 42 302 88 314
rect 42 112 48 302
rect 82 112 88 302
rect 42 100 88 112
rect 234 302 280 362
rect 234 112 240 302
rect 274 112 280 302
rect 234 100 280 112
rect 426 302 472 314
rect 426 112 432 302
rect 466 112 472 302
rect 426 100 472 112
rect 618 302 664 362
rect 618 112 624 302
rect 658 112 664 302
rect 618 100 664 112
rect 810 302 856 314
rect 810 112 816 302
rect 850 112 856 302
rect 810 69 856 112
rect 1002 302 1048 362
rect 1002 112 1008 302
rect 1042 112 1048 302
rect 1002 100 1048 112
rect 1194 302 1240 314
rect 1194 112 1200 302
rect 1234 112 1240 302
rect 1194 69 1240 112
rect -68 53 526 69
rect -68 19 480 53
rect 514 19 526 53
rect -68 3 526 19
rect 810 8 1240 69
rect -68 -55 722 -39
rect -68 -89 672 -55
rect 706 -89 722 -55
rect -68 -105 722 -89
rect 810 -139 856 8
rect 618 -151 856 -139
rect 618 -327 624 -151
rect 658 -327 856 -151
rect 618 -339 856 -327
<< labels >>
flabel metal1 -61 10 16 62 1 FreeSerif 320 0 0 0 A
port 1 w
flabel metal1 -60 -99 17 -47 1 FreeSerif 320 0 0 0 B
port 2 w
flabel metal1 777 -236 854 -184 1 FreeSerif 320 0 0 0 Y
port 5 s
rlabel locali 562 -494 732 -426 5 VSS
port 3 s
rlabel locali 82 424 262 486 1 VDD
port 4 n
<< end >>
