magic
tech sky130B
magscale 1 2
timestamp 1736595726
<< nwell >>
rect 3025 865 4210 866
rect 1812 860 4210 865
rect 693 845 4210 860
rect -501 843 4210 845
rect -5019 812 -3004 813
rect -1701 812 4210 843
rect -5019 434 4210 812
rect -5019 433 3706 434
rect -5019 428 2521 433
rect -5019 413 1308 428
rect -5019 411 189 413
rect -5019 381 -1005 411
rect -2982 380 -1005 381
rect -2982 379 -2205 380
<< metal1 >>
rect -5260 250 -5171 1197
rect -5090 279 -5018 1197
rect -4732 1086 -4620 1094
rect -4732 990 -4724 1086
rect -4628 990 -4620 1086
rect -4732 982 -4620 990
rect -4724 712 -4628 982
rect -4380 313 -4172 395
rect -5260 114 -4997 250
rect -4615 -367 -4514 26
rect -4615 -474 -4514 -468
rect -4250 -734 -4172 313
rect -3950 250 -3861 1197
rect -3780 279 -3708 1197
rect -3426 1066 -3314 1074
rect -3426 970 -3418 1066
rect -3322 970 -3314 1066
rect -3426 962 -3314 970
rect -3419 717 -3322 962
rect -3008 305 -2867 387
rect -3950 114 -3708 250
rect -3299 -407 -3198 42
rect -3299 -514 -3198 -508
rect -2945 -734 -2867 305
rect -2649 249 -2560 1197
rect -2479 278 -2407 1197
rect -2118 1076 -2006 1084
rect -2118 980 -2110 1076
rect -2014 980 -2006 1076
rect -2118 972 -2006 980
rect -2110 751 -2014 972
rect -1701 307 -1565 389
rect -2649 113 -2407 249
rect -2005 -410 -1904 69
rect -2005 -517 -1904 -511
rect -1643 -734 -1565 307
rect -1443 280 -1354 1197
rect -1273 309 -1201 1197
rect -922 1076 -810 1084
rect -922 980 -914 1076
rect -818 980 -810 1076
rect -922 972 -810 980
rect -914 771 -818 972
rect -512 323 -365 405
rect -1443 144 -1201 280
rect -807 -401 -706 77
rect -807 -508 -706 -502
rect -443 -734 -365 323
rect -255 282 -166 1197
rect -85 311 -13 1197
rect 272 1076 384 1084
rect 272 980 280 1076
rect 376 980 384 1076
rect 272 972 384 980
rect 280 776 376 972
rect 691 376 824 458
rect -255 146 -13 282
rect 365 -378 466 87
rect 365 -485 466 -479
rect 746 -734 824 376
rect 873 297 962 1197
rect 1036 427 1106 1197
rect 1386 1090 1498 1098
rect 1386 994 1394 1090
rect 1490 994 1498 1090
rect 1386 986 1498 994
rect 1394 759 1490 986
rect 1114 427 1115 461
rect 1036 326 1115 427
rect 1802 360 1926 442
rect 873 161 1115 297
rect 1506 -370 1607 96
rect 1506 -477 1607 -471
rect 1848 -734 1926 360
rect 2078 302 2167 1197
rect 2248 331 2320 1197
rect 2618 1096 2730 1104
rect 2618 1000 2626 1096
rect 2722 1000 2730 1096
rect 2618 992 2730 1000
rect 2626 792 2722 992
rect 3022 368 3131 450
rect 2078 166 2320 302
rect 2718 -361 2819 108
rect 2718 -468 2819 -462
rect 3053 -734 3131 368
rect 3262 303 3351 1197
rect 3432 332 3504 1197
rect 3792 1100 3904 1108
rect 3792 1004 3800 1100
rect 3896 1004 3904 1100
rect 3792 996 3904 1004
rect 3800 785 3896 996
rect 4204 376 4324 458
rect 3262 167 3504 303
rect 3914 -318 4015 103
rect 3914 -425 4015 -419
rect 4246 -734 4324 376
<< via1 >>
rect -4724 990 -4628 1086
rect -4615 -468 -4514 -367
rect -3418 970 -3322 1066
rect -3299 -508 -3198 -407
rect -2110 980 -2014 1076
rect -2005 -511 -1904 -410
rect -914 980 -818 1076
rect -807 -502 -706 -401
rect 280 980 376 1076
rect 365 -479 466 -378
rect 1394 994 1490 1090
rect 1506 -471 1607 -370
rect 2626 1000 2722 1096
rect 2718 -462 2819 -361
rect 3800 1004 3896 1100
rect 3914 -419 4015 -318
<< metal2 >>
rect -4734 1086 -4618 1096
rect 1384 1090 1500 1100
rect -4734 990 -4724 1086
rect -4628 990 -4618 1086
rect -2120 1076 -2004 1086
rect -4734 980 -4618 990
rect -3428 1066 -3312 1076
rect -3428 970 -3418 1066
rect -3322 970 -3312 1066
rect -2120 980 -2110 1076
rect -2014 980 -2004 1076
rect -2120 970 -2004 980
rect -924 1076 -808 1086
rect -924 980 -914 1076
rect -818 980 -808 1076
rect -924 970 -808 980
rect 270 1076 386 1086
rect 270 980 280 1076
rect 376 980 386 1076
rect 1384 994 1394 1090
rect 1490 994 1500 1090
rect 1384 984 1500 994
rect 2616 1096 2732 1106
rect 2616 1000 2626 1096
rect 2722 1000 2732 1096
rect 2616 990 2732 1000
rect 3790 1100 3906 1110
rect 3790 1004 3800 1100
rect 3896 1004 3906 1100
rect 3790 994 3906 1004
rect 270 970 386 980
rect -3428 960 -3312 970
rect 3899 -318 4027 -306
rect -4630 -367 -4502 -355
rect -4630 -468 -4615 -367
rect -4514 -468 -4502 -367
rect 350 -378 478 -366
rect -4630 -478 -4502 -468
rect -3314 -407 -3186 -395
rect -3314 -508 -3299 -407
rect -3198 -508 -3186 -407
rect -3314 -518 -3186 -508
rect -2020 -410 -1892 -398
rect -2020 -511 -2005 -410
rect -1904 -511 -1892 -410
rect -2020 -521 -1892 -511
rect -822 -401 -694 -389
rect -822 -502 -807 -401
rect -706 -502 -694 -401
rect 350 -479 365 -378
rect 466 -479 478 -378
rect 350 -489 478 -479
rect 1491 -370 1619 -358
rect 1491 -471 1506 -370
rect 1607 -471 1619 -370
rect 1491 -481 1619 -471
rect 2703 -361 2831 -349
rect 2703 -462 2718 -361
rect 2819 -462 2831 -361
rect 3899 -419 3914 -318
rect 4015 -419 4027 -318
rect 3899 -429 4027 -419
rect 2703 -472 2831 -462
rect -822 -512 -694 -502
<< via2 >>
rect -4724 990 -4628 1086
rect -3418 970 -3322 1066
rect -2110 980 -2014 1076
rect -914 980 -818 1076
rect 280 980 376 1076
rect 1394 994 1490 1090
rect 2626 1000 2722 1096
rect 3800 1004 3896 1100
rect -4615 -468 -4514 -367
rect -3299 -508 -3198 -407
rect -2005 -511 -1904 -410
rect -807 -502 -706 -401
rect 365 -479 466 -378
rect 1506 -471 1607 -370
rect 2718 -462 2819 -361
rect 3914 -419 4015 -318
<< metal3 >>
rect -4736 1091 -4616 1098
rect -4736 985 -4729 1091
rect -4623 985 -4616 1091
rect 1382 1095 1502 1102
rect -2122 1081 -2002 1088
rect -4736 978 -4616 985
rect -3430 1071 -3310 1078
rect -3430 965 -3423 1071
rect -3317 965 -3310 1071
rect -2122 975 -2115 1081
rect -2009 975 -2002 1081
rect -2122 968 -2002 975
rect -926 1081 -806 1088
rect -926 975 -919 1081
rect -813 975 -806 1081
rect -926 968 -806 975
rect 268 1081 388 1088
rect 268 975 275 1081
rect 381 975 388 1081
rect 1382 989 1389 1095
rect 1495 989 1502 1095
rect 1382 982 1502 989
rect 2614 1101 2734 1108
rect 2614 995 2621 1101
rect 2727 995 2734 1101
rect 2614 988 2734 995
rect 3788 1105 3908 1112
rect 3788 999 3795 1105
rect 3901 999 3908 1105
rect 3788 992 3908 999
rect 268 968 388 975
rect -3430 958 -3310 965
rect 3883 -313 4039 -289
rect -4646 -362 -4490 -338
rect -4646 -473 -4620 -362
rect -4509 -473 -4490 -362
rect -4646 -501 -4490 -473
rect -3330 -402 -3174 -378
rect -3330 -513 -3304 -402
rect -3193 -513 -3174 -402
rect -3330 -541 -3174 -513
rect -2036 -405 -1880 -381
rect -2036 -516 -2010 -405
rect -1899 -516 -1880 -405
rect -2036 -544 -1880 -516
rect -838 -396 -682 -372
rect -838 -507 -812 -396
rect -701 -507 -682 -396
rect -838 -535 -682 -507
rect 334 -373 490 -349
rect 334 -484 360 -373
rect 471 -484 490 -373
rect 334 -512 490 -484
rect 1475 -365 1631 -341
rect 1475 -476 1501 -365
rect 1612 -476 1631 -365
rect 1475 -504 1631 -476
rect 2687 -356 2843 -332
rect 2687 -467 2713 -356
rect 2824 -467 2843 -356
rect 3883 -424 3909 -313
rect 4020 -424 4039 -313
rect 3883 -452 4039 -424
rect 2687 -495 2843 -467
<< via3 >>
rect -4729 1086 -4623 1091
rect -4729 990 -4724 1086
rect -4724 990 -4628 1086
rect -4628 990 -4623 1086
rect -4729 985 -4623 990
rect -3423 1066 -3317 1071
rect -3423 970 -3418 1066
rect -3418 970 -3322 1066
rect -3322 970 -3317 1066
rect -3423 965 -3317 970
rect -2115 1076 -2009 1081
rect -2115 980 -2110 1076
rect -2110 980 -2014 1076
rect -2014 980 -2009 1076
rect -2115 975 -2009 980
rect -919 1076 -813 1081
rect -919 980 -914 1076
rect -914 980 -818 1076
rect -818 980 -813 1076
rect -919 975 -813 980
rect 275 1076 381 1081
rect 275 980 280 1076
rect 280 980 376 1076
rect 376 980 381 1076
rect 275 975 381 980
rect 1389 1090 1495 1095
rect 1389 994 1394 1090
rect 1394 994 1490 1090
rect 1490 994 1495 1090
rect 1389 989 1495 994
rect 2621 1096 2727 1101
rect 2621 1000 2626 1096
rect 2626 1000 2722 1096
rect 2722 1000 2727 1096
rect 2621 995 2727 1000
rect 3795 1100 3901 1105
rect 3795 1004 3800 1100
rect 3800 1004 3896 1100
rect 3896 1004 3901 1100
rect 3795 999 3901 1004
rect -4620 -367 -4509 -362
rect -4620 -468 -4615 -367
rect -4615 -468 -4514 -367
rect -4514 -468 -4509 -367
rect -4620 -473 -4509 -468
rect -3304 -407 -3193 -402
rect -3304 -508 -3299 -407
rect -3299 -508 -3198 -407
rect -3198 -508 -3193 -407
rect -3304 -513 -3193 -508
rect -2010 -410 -1899 -405
rect -2010 -511 -2005 -410
rect -2005 -511 -1904 -410
rect -1904 -511 -1899 -410
rect -2010 -516 -1899 -511
rect -812 -401 -701 -396
rect -812 -502 -807 -401
rect -807 -502 -706 -401
rect -706 -502 -701 -401
rect -812 -507 -701 -502
rect 360 -378 471 -373
rect 360 -479 365 -378
rect 365 -479 466 -378
rect 466 -479 471 -378
rect 360 -484 471 -479
rect 1501 -370 1612 -365
rect 1501 -471 1506 -370
rect 1506 -471 1607 -370
rect 1607 -471 1612 -370
rect 1501 -476 1612 -471
rect 2713 -361 2824 -356
rect 2713 -462 2718 -361
rect 2718 -462 2819 -361
rect 2819 -462 2824 -361
rect 2713 -467 2824 -462
rect 3909 -318 4020 -313
rect 3909 -419 3914 -318
rect 3914 -419 4015 -318
rect 4015 -419 4020 -318
rect 3909 -424 4020 -419
<< metal4 >>
rect -4970 1105 4122 1197
rect -4970 1101 3795 1105
rect -4970 1095 2621 1101
rect -4970 1091 1389 1095
rect -4970 985 -4729 1091
rect -4623 1081 1389 1091
rect -4623 1071 -2115 1081
rect -4623 985 -3423 1071
rect -4970 965 -3423 985
rect -3317 975 -2115 1071
rect -2009 975 -919 1081
rect -813 975 275 1081
rect 381 989 1389 1081
rect 1495 995 2621 1095
rect 2727 999 3795 1101
rect 3901 999 4122 1105
rect 2727 995 4122 999
rect 1495 989 4122 995
rect 381 975 4122 989
rect -3317 965 4122 975
rect -4970 927 4122 965
<< via4 >>
rect -4724 -362 -4404 -257
rect -4724 -473 -4620 -362
rect -4620 -473 -4509 -362
rect -4509 -473 -4404 -362
rect -4724 -577 -4404 -473
rect -3408 -402 -3088 -297
rect -3408 -513 -3304 -402
rect -3304 -513 -3193 -402
rect -3193 -513 -3088 -402
rect -3408 -617 -3088 -513
rect -2114 -405 -1794 -300
rect -2114 -516 -2010 -405
rect -2010 -516 -1899 -405
rect -1899 -516 -1794 -405
rect -2114 -620 -1794 -516
rect -916 -396 -596 -291
rect -916 -507 -812 -396
rect -812 -507 -701 -396
rect -701 -507 -596 -396
rect -916 -611 -596 -507
rect 256 -373 576 -268
rect 256 -484 360 -373
rect 360 -484 471 -373
rect 471 -484 576 -373
rect 256 -588 576 -484
rect 1397 -365 1717 -260
rect 1397 -476 1501 -365
rect 1501 -476 1612 -365
rect 1612 -476 1717 -365
rect 1397 -580 1717 -476
rect 2609 -356 2929 -251
rect 2609 -467 2713 -356
rect 2713 -467 2824 -356
rect 2824 -467 2929 -356
rect 2609 -571 2929 -467
rect 3805 -313 4125 -208
rect 3805 -424 3909 -313
rect 3909 -424 4020 -313
rect 4020 -424 4125 -313
rect 3805 -528 4125 -424
<< metal5 >>
rect -4930 -208 4221 -92
rect -4930 -251 3805 -208
rect -4930 -257 2609 -251
rect -4930 -577 -4724 -257
rect -4404 -260 2609 -257
rect -4404 -268 1397 -260
rect -4404 -291 256 -268
rect -4404 -297 -916 -291
rect -4404 -577 -3408 -297
rect -4930 -617 -3408 -577
rect -3088 -300 -916 -297
rect -3088 -617 -2114 -300
rect -4930 -620 -2114 -617
rect -1794 -611 -916 -300
rect -596 -588 256 -291
rect 576 -580 1397 -268
rect 1717 -571 2609 -260
rect 2929 -528 3805 -251
rect 4125 -528 4221 -208
rect 2929 -571 4221 -528
rect 1717 -580 4221 -571
rect 576 -588 4221 -580
rect -596 -611 4221 -588
rect -1794 -620 4221 -611
rect -4930 -734 4221 -620
use NAND2  NAND2_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NAND/NAND2
timestamp 1736436273
transform 1 0 3148 0 1 62
box 356 -17 1062 804
use NAND2  NAND2_1
timestamp 1736436273
transform 1 0 -369 0 1 41
box 356 -17 1062 804
use NAND2  NAND2_2
timestamp 1736436273
transform 1 0 -1563 0 1 39
box 356 -17 1062 804
use NAND2  NAND2_4
timestamp 1736436273
transform 1 0 -5375 0 1 9
box 356 -17 1062 804
use NAND2  NAND2_6
timestamp 1736436273
transform 1 0 750 0 1 56
box 356 -17 1062 804
use NAND2  NAND2_7
timestamp 1736436273
transform 1 0 1963 0 1 61
box 356 -17 1062 804
use NAND2  NAND2_8
timestamp 1736436273
transform 1 0 -4066 0 1 9
box 356 -17 1062 804
use NAND2  NAND2_9
timestamp 1736436273
transform 1 0 -2763 0 1 8
box 356 -17 1062 804
<< labels >>
rlabel metal1 -5251 1132 -5184 1189 1 A0
port 3 n
rlabel metal1 -5082 1132 -5026 1189 1 B0
port 4 n
rlabel metal1 -3945 1127 -3870 1191 1 A1
port 5 n
rlabel metal1 -3770 1127 -3716 1190 1 B1
port 6 n
rlabel metal1 -2641 1133 -2572 1189 1 A2
port 7 n
rlabel metal1 -2469 1133 -2413 1188 1 B2
port 8 n
rlabel metal1 -1435 1120 -1362 1188 1 A3
port 9 n
rlabel metal1 -1265 1121 -1209 1188 1 B3
port 10 n
rlabel metal1 -247 1121 -175 1190 1 A4
port 11 n
rlabel metal1 -80 1121 -18 1190 1 B4
port 12 n
rlabel metal1 879 1110 953 1191 1 A5
port 13 n
rlabel metal1 1045 1113 1099 1191 1 B5
port 14 n
rlabel metal1 2082 1109 2161 1192 1 A6
port 15 n
rlabel metal1 2256 1109 2316 1191 1 B6
port 16 n
rlabel metal1 3268 1107 3342 1189 1 A7
port 17 n
rlabel metal1 3439 1107 3498 1188 1 B7
port 18 n
rlabel metal1 -4244 -729 -4179 -660 5 P0
port 19 s
rlabel metal1 -2938 -728 -2873 -659 5 P1
port 20 s
rlabel metal1 -1637 -729 -1572 -660 5 P2
port 21 s
rlabel metal1 -438 -730 -373 -661 5 P3
port 22 s
rlabel metal1 752 -729 817 -660 5 P4
port 23 s
rlabel metal1 1854 -730 1919 -661 5 P5
port 24 s
rlabel metal1 3057 -729 3122 -660 5 P6
port 25 s
rlabel metal1 4253 -729 4318 -660 5 P7
port 26 s
<< end >>
