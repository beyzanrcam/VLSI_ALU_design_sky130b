magic
tech sky130B
magscale 1 2
timestamp 1733246765
<< error_p >>
rect -678 937 -620 943
rect -560 937 -502 943
rect -442 937 -384 943
rect -324 937 -266 943
rect -206 937 -148 943
rect -88 937 -30 943
rect 30 937 88 943
rect 148 937 206 943
rect 266 937 324 943
rect 384 937 442 943
rect 502 937 560 943
rect 620 937 678 943
rect -678 903 -666 937
rect -560 903 -548 937
rect -442 903 -430 937
rect -324 903 -312 937
rect -206 903 -194 937
rect -88 903 -76 937
rect 30 903 42 937
rect 148 903 160 937
rect 266 903 278 937
rect 384 903 396 937
rect 502 903 514 937
rect 620 903 632 937
rect -678 897 -620 903
rect -560 897 -502 903
rect -442 897 -384 903
rect -324 897 -266 903
rect -206 897 -148 903
rect -88 897 -30 903
rect 30 897 88 903
rect 148 897 206 903
rect 266 897 324 903
rect 384 897 442 903
rect 502 897 560 903
rect 620 897 678 903
rect -678 -903 -620 -897
rect -560 -903 -502 -897
rect -442 -903 -384 -897
rect -324 -903 -266 -897
rect -206 -903 -148 -897
rect -88 -903 -30 -897
rect 30 -903 88 -897
rect 148 -903 206 -897
rect 266 -903 324 -897
rect 384 -903 442 -897
rect 502 -903 560 -897
rect 620 -903 678 -897
rect -678 -937 -666 -903
rect -560 -937 -548 -903
rect -442 -937 -430 -903
rect -324 -937 -312 -903
rect -206 -937 -194 -903
rect -88 -937 -76 -903
rect 30 -937 42 -903
rect 148 -937 160 -903
rect 266 -937 278 -903
rect 384 -937 396 -903
rect 502 -937 514 -903
rect 620 -937 632 -903
rect -678 -943 -620 -937
rect -560 -943 -502 -937
rect -442 -943 -384 -937
rect -324 -943 -266 -937
rect -206 -943 -148 -937
rect -88 -943 -30 -937
rect 30 -943 88 -937
rect 148 -943 206 -937
rect 266 -943 324 -937
rect 384 -943 442 -937
rect 502 -943 560 -937
rect 620 -943 678 -937
<< nwell >>
rect -875 -1075 875 1075
<< pmos >>
rect -679 -856 -619 856
rect -561 -856 -501 856
rect -443 -856 -383 856
rect -325 -856 -265 856
rect -207 -856 -147 856
rect -89 -856 -29 856
rect 29 -856 89 856
rect 147 -856 207 856
rect 265 -856 325 856
rect 383 -856 443 856
rect 501 -856 561 856
rect 619 -856 679 856
<< pdiff >>
rect -737 844 -679 856
rect -737 -844 -725 844
rect -691 -844 -679 844
rect -737 -856 -679 -844
rect -619 844 -561 856
rect -619 -844 -607 844
rect -573 -844 -561 844
rect -619 -856 -561 -844
rect -501 844 -443 856
rect -501 -844 -489 844
rect -455 -844 -443 844
rect -501 -856 -443 -844
rect -383 844 -325 856
rect -383 -844 -371 844
rect -337 -844 -325 844
rect -383 -856 -325 -844
rect -265 844 -207 856
rect -265 -844 -253 844
rect -219 -844 -207 844
rect -265 -856 -207 -844
rect -147 844 -89 856
rect -147 -844 -135 844
rect -101 -844 -89 844
rect -147 -856 -89 -844
rect -29 844 29 856
rect -29 -844 -17 844
rect 17 -844 29 844
rect -29 -856 29 -844
rect 89 844 147 856
rect 89 -844 101 844
rect 135 -844 147 844
rect 89 -856 147 -844
rect 207 844 265 856
rect 207 -844 219 844
rect 253 -844 265 844
rect 207 -856 265 -844
rect 325 844 383 856
rect 325 -844 337 844
rect 371 -844 383 844
rect 325 -856 383 -844
rect 443 844 501 856
rect 443 -844 455 844
rect 489 -844 501 844
rect 443 -856 501 -844
rect 561 844 619 856
rect 561 -844 573 844
rect 607 -844 619 844
rect 561 -856 619 -844
rect 679 844 737 856
rect 679 -844 691 844
rect 725 -844 737 844
rect 679 -856 737 -844
<< pdiffc >>
rect -725 -844 -691 844
rect -607 -844 -573 844
rect -489 -844 -455 844
rect -371 -844 -337 844
rect -253 -844 -219 844
rect -135 -844 -101 844
rect -17 -844 17 844
rect 101 -844 135 844
rect 219 -844 253 844
rect 337 -844 371 844
rect 455 -844 489 844
rect 573 -844 607 844
rect 691 -844 725 844
<< nsubdiff >>
rect -839 1005 -743 1039
rect 743 1005 839 1039
rect -839 943 -805 1005
rect 805 943 839 1005
rect -839 -1005 -805 -943
rect 805 -1005 839 -943
rect -839 -1039 -743 -1005
rect 743 -1039 839 -1005
<< nsubdiffcont >>
rect -743 1005 743 1039
rect -839 -943 -805 943
rect 805 -943 839 943
rect -743 -1039 743 -1005
<< poly >>
rect -682 937 -616 953
rect -682 903 -666 937
rect -632 903 -616 937
rect -682 887 -616 903
rect -564 937 -498 953
rect -564 903 -548 937
rect -514 903 -498 937
rect -564 887 -498 903
rect -446 937 -380 953
rect -446 903 -430 937
rect -396 903 -380 937
rect -446 887 -380 903
rect -328 937 -262 953
rect -328 903 -312 937
rect -278 903 -262 937
rect -328 887 -262 903
rect -210 937 -144 953
rect -210 903 -194 937
rect -160 903 -144 937
rect -210 887 -144 903
rect -92 937 -26 953
rect -92 903 -76 937
rect -42 903 -26 937
rect -92 887 -26 903
rect 26 937 92 953
rect 26 903 42 937
rect 76 903 92 937
rect 26 887 92 903
rect 144 937 210 953
rect 144 903 160 937
rect 194 903 210 937
rect 144 887 210 903
rect 262 937 328 953
rect 262 903 278 937
rect 312 903 328 937
rect 262 887 328 903
rect 380 937 446 953
rect 380 903 396 937
rect 430 903 446 937
rect 380 887 446 903
rect 498 937 564 953
rect 498 903 514 937
rect 548 903 564 937
rect 498 887 564 903
rect 616 937 682 953
rect 616 903 632 937
rect 666 903 682 937
rect 616 887 682 903
rect -679 856 -619 887
rect -561 856 -501 887
rect -443 856 -383 887
rect -325 856 -265 887
rect -207 856 -147 887
rect -89 856 -29 887
rect 29 856 89 887
rect 147 856 207 887
rect 265 856 325 887
rect 383 856 443 887
rect 501 856 561 887
rect 619 856 679 887
rect -679 -887 -619 -856
rect -561 -887 -501 -856
rect -443 -887 -383 -856
rect -325 -887 -265 -856
rect -207 -887 -147 -856
rect -89 -887 -29 -856
rect 29 -887 89 -856
rect 147 -887 207 -856
rect 265 -887 325 -856
rect 383 -887 443 -856
rect 501 -887 561 -856
rect 619 -887 679 -856
rect -682 -903 -616 -887
rect -682 -937 -666 -903
rect -632 -937 -616 -903
rect -682 -953 -616 -937
rect -564 -903 -498 -887
rect -564 -937 -548 -903
rect -514 -937 -498 -903
rect -564 -953 -498 -937
rect -446 -903 -380 -887
rect -446 -937 -430 -903
rect -396 -937 -380 -903
rect -446 -953 -380 -937
rect -328 -903 -262 -887
rect -328 -937 -312 -903
rect -278 -937 -262 -903
rect -328 -953 -262 -937
rect -210 -903 -144 -887
rect -210 -937 -194 -903
rect -160 -937 -144 -903
rect -210 -953 -144 -937
rect -92 -903 -26 -887
rect -92 -937 -76 -903
rect -42 -937 -26 -903
rect -92 -953 -26 -937
rect 26 -903 92 -887
rect 26 -937 42 -903
rect 76 -937 92 -903
rect 26 -953 92 -937
rect 144 -903 210 -887
rect 144 -937 160 -903
rect 194 -937 210 -903
rect 144 -953 210 -937
rect 262 -903 328 -887
rect 262 -937 278 -903
rect 312 -937 328 -903
rect 262 -953 328 -937
rect 380 -903 446 -887
rect 380 -937 396 -903
rect 430 -937 446 -903
rect 380 -953 446 -937
rect 498 -903 564 -887
rect 498 -937 514 -903
rect 548 -937 564 -903
rect 498 -953 564 -937
rect 616 -903 682 -887
rect 616 -937 632 -903
rect 666 -937 682 -903
rect 616 -953 682 -937
<< polycont >>
rect -666 903 -632 937
rect -548 903 -514 937
rect -430 903 -396 937
rect -312 903 -278 937
rect -194 903 -160 937
rect -76 903 -42 937
rect 42 903 76 937
rect 160 903 194 937
rect 278 903 312 937
rect 396 903 430 937
rect 514 903 548 937
rect 632 903 666 937
rect -666 -937 -632 -903
rect -548 -937 -514 -903
rect -430 -937 -396 -903
rect -312 -937 -278 -903
rect -194 -937 -160 -903
rect -76 -937 -42 -903
rect 42 -937 76 -903
rect 160 -937 194 -903
rect 278 -937 312 -903
rect 396 -937 430 -903
rect 514 -937 548 -903
rect 632 -937 666 -903
<< locali >>
rect -839 1005 -743 1039
rect 743 1005 839 1039
rect -839 943 -805 1005
rect 805 943 839 1005
rect -682 903 -666 937
rect -632 903 -616 937
rect -564 903 -548 937
rect -514 903 -498 937
rect -446 903 -430 937
rect -396 903 -380 937
rect -328 903 -312 937
rect -278 903 -262 937
rect -210 903 -194 937
rect -160 903 -144 937
rect -92 903 -76 937
rect -42 903 -26 937
rect 26 903 42 937
rect 76 903 92 937
rect 144 903 160 937
rect 194 903 210 937
rect 262 903 278 937
rect 312 903 328 937
rect 380 903 396 937
rect 430 903 446 937
rect 498 903 514 937
rect 548 903 564 937
rect 616 903 632 937
rect 666 903 682 937
rect -725 844 -691 860
rect -725 -860 -691 -844
rect -607 844 -573 860
rect -607 -860 -573 -844
rect -489 844 -455 860
rect -489 -860 -455 -844
rect -371 844 -337 860
rect -371 -860 -337 -844
rect -253 844 -219 860
rect -253 -860 -219 -844
rect -135 844 -101 860
rect -135 -860 -101 -844
rect -17 844 17 860
rect -17 -860 17 -844
rect 101 844 135 860
rect 101 -860 135 -844
rect 219 844 253 860
rect 219 -860 253 -844
rect 337 844 371 860
rect 337 -860 371 -844
rect 455 844 489 860
rect 455 -860 489 -844
rect 573 844 607 860
rect 573 -860 607 -844
rect 691 844 725 860
rect 691 -860 725 -844
rect -682 -937 -666 -903
rect -632 -937 -616 -903
rect -564 -937 -548 -903
rect -514 -937 -498 -903
rect -446 -937 -430 -903
rect -396 -937 -380 -903
rect -328 -937 -312 -903
rect -278 -937 -262 -903
rect -210 -937 -194 -903
rect -160 -937 -144 -903
rect -92 -937 -76 -903
rect -42 -937 -26 -903
rect 26 -937 42 -903
rect 76 -937 92 -903
rect 144 -937 160 -903
rect 194 -937 210 -903
rect 262 -937 278 -903
rect 312 -937 328 -903
rect 380 -937 396 -903
rect 430 -937 446 -903
rect 498 -937 514 -903
rect 548 -937 564 -903
rect 616 -937 632 -903
rect 666 -937 682 -903
rect -839 -1005 -805 -943
rect 805 -1005 839 -943
rect -839 -1039 -743 -1005
rect 743 -1039 839 -1005
<< viali >>
rect -666 903 -632 937
rect -548 903 -514 937
rect -430 903 -396 937
rect -312 903 -278 937
rect -194 903 -160 937
rect -76 903 -42 937
rect 42 903 76 937
rect 160 903 194 937
rect 278 903 312 937
rect 396 903 430 937
rect 514 903 548 937
rect 632 903 666 937
rect -725 -844 -691 844
rect -607 -844 -573 844
rect -489 -844 -455 844
rect -371 -844 -337 844
rect -253 -844 -219 844
rect -135 -844 -101 844
rect -17 -844 17 844
rect 101 -844 135 844
rect 219 -844 253 844
rect 337 -844 371 844
rect 455 -844 489 844
rect 573 -844 607 844
rect 691 -844 725 844
rect -666 -937 -632 -903
rect -548 -937 -514 -903
rect -430 -937 -396 -903
rect -312 -937 -278 -903
rect -194 -937 -160 -903
rect -76 -937 -42 -903
rect 42 -937 76 -903
rect 160 -937 194 -903
rect 278 -937 312 -903
rect 396 -937 430 -903
rect 514 -937 548 -903
rect 632 -937 666 -903
<< metal1 >>
rect -678 937 -620 943
rect -678 903 -666 937
rect -632 903 -620 937
rect -678 897 -620 903
rect -560 937 -502 943
rect -560 903 -548 937
rect -514 903 -502 937
rect -560 897 -502 903
rect -442 937 -384 943
rect -442 903 -430 937
rect -396 903 -384 937
rect -442 897 -384 903
rect -324 937 -266 943
rect -324 903 -312 937
rect -278 903 -266 937
rect -324 897 -266 903
rect -206 937 -148 943
rect -206 903 -194 937
rect -160 903 -148 937
rect -206 897 -148 903
rect -88 937 -30 943
rect -88 903 -76 937
rect -42 903 -30 937
rect -88 897 -30 903
rect 30 937 88 943
rect 30 903 42 937
rect 76 903 88 937
rect 30 897 88 903
rect 148 937 206 943
rect 148 903 160 937
rect 194 903 206 937
rect 148 897 206 903
rect 266 937 324 943
rect 266 903 278 937
rect 312 903 324 937
rect 266 897 324 903
rect 384 937 442 943
rect 384 903 396 937
rect 430 903 442 937
rect 384 897 442 903
rect 502 937 560 943
rect 502 903 514 937
rect 548 903 560 937
rect 502 897 560 903
rect 620 937 678 943
rect 620 903 632 937
rect 666 903 678 937
rect 620 897 678 903
rect -731 844 -685 856
rect -731 -844 -725 844
rect -691 -844 -685 844
rect -731 -856 -685 -844
rect -613 844 -567 856
rect -613 -844 -607 844
rect -573 -844 -567 844
rect -613 -856 -567 -844
rect -495 844 -449 856
rect -495 -844 -489 844
rect -455 -844 -449 844
rect -495 -856 -449 -844
rect -377 844 -331 856
rect -377 -844 -371 844
rect -337 -844 -331 844
rect -377 -856 -331 -844
rect -259 844 -213 856
rect -259 -844 -253 844
rect -219 -844 -213 844
rect -259 -856 -213 -844
rect -141 844 -95 856
rect -141 -844 -135 844
rect -101 -844 -95 844
rect -141 -856 -95 -844
rect -23 844 23 856
rect -23 -844 -17 844
rect 17 -844 23 844
rect -23 -856 23 -844
rect 95 844 141 856
rect 95 -844 101 844
rect 135 -844 141 844
rect 95 -856 141 -844
rect 213 844 259 856
rect 213 -844 219 844
rect 253 -844 259 844
rect 213 -856 259 -844
rect 331 844 377 856
rect 331 -844 337 844
rect 371 -844 377 844
rect 331 -856 377 -844
rect 449 844 495 856
rect 449 -844 455 844
rect 489 -844 495 844
rect 449 -856 495 -844
rect 567 844 613 856
rect 567 -844 573 844
rect 607 -844 613 844
rect 567 -856 613 -844
rect 685 844 731 856
rect 685 -844 691 844
rect 725 -844 731 844
rect 685 -856 731 -844
rect -678 -903 -620 -897
rect -678 -937 -666 -903
rect -632 -937 -620 -903
rect -678 -943 -620 -937
rect -560 -903 -502 -897
rect -560 -937 -548 -903
rect -514 -937 -502 -903
rect -560 -943 -502 -937
rect -442 -903 -384 -897
rect -442 -937 -430 -903
rect -396 -937 -384 -903
rect -442 -943 -384 -937
rect -324 -903 -266 -897
rect -324 -937 -312 -903
rect -278 -937 -266 -903
rect -324 -943 -266 -937
rect -206 -903 -148 -897
rect -206 -937 -194 -903
rect -160 -937 -148 -903
rect -206 -943 -148 -937
rect -88 -903 -30 -897
rect -88 -937 -76 -903
rect -42 -937 -30 -903
rect -88 -943 -30 -937
rect 30 -903 88 -897
rect 30 -937 42 -903
rect 76 -937 88 -903
rect 30 -943 88 -937
rect 148 -903 206 -897
rect 148 -937 160 -903
rect 194 -937 206 -903
rect 148 -943 206 -937
rect 266 -903 324 -897
rect 266 -937 278 -903
rect 312 -937 324 -903
rect 266 -943 324 -937
rect 384 -903 442 -897
rect 384 -937 396 -903
rect 430 -937 442 -903
rect 384 -943 442 -937
rect 502 -903 560 -897
rect 502 -937 514 -903
rect 548 -937 560 -903
rect 502 -943 560 -937
rect 620 -903 678 -897
rect 620 -937 632 -903
rect 666 -937 678 -903
rect 620 -943 678 -937
<< properties >>
string FIXED_BBOX -822 -1022 822 1022
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.56 l 0.30 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
