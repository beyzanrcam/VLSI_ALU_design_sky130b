magic
tech sky130B
magscale 1 2
timestamp 1736012282
<< nwell >>
rect 1 459 1090 580
rect 0 3 1090 459
<< nmos >>
rect 482 -330 512 -130
rect 578 -330 608 -130
<< pmos >>
rect 98 103 128 359
rect 194 103 224 359
rect 290 103 320 359
rect 386 103 416 359
rect 482 103 512 359
rect 578 103 608 359
rect 674 103 704 359
rect 770 103 800 359
rect 866 103 896 359
rect 962 103 992 359
<< ndiff >>
rect 420 -142 482 -130
rect 420 -318 432 -142
rect 466 -318 482 -142
rect 420 -330 482 -318
rect 512 -142 578 -130
rect 512 -318 528 -142
rect 562 -318 578 -142
rect 512 -330 578 -318
rect 608 -142 670 -130
rect 608 -318 624 -142
rect 658 -318 670 -142
rect 608 -330 670 -318
<< pdiff >>
rect 36 347 98 359
rect 36 115 48 347
rect 82 115 98 347
rect 36 103 98 115
rect 128 347 194 359
rect 128 115 144 347
rect 178 115 194 347
rect 128 103 194 115
rect 224 347 290 359
rect 224 115 240 347
rect 274 115 290 347
rect 224 103 290 115
rect 320 347 386 359
rect 320 115 336 347
rect 370 115 386 347
rect 320 103 386 115
rect 416 347 482 359
rect 416 115 432 347
rect 466 115 482 347
rect 416 103 482 115
rect 512 347 578 359
rect 512 115 528 347
rect 562 115 578 347
rect 512 103 578 115
rect 608 347 674 359
rect 608 115 624 347
rect 658 115 674 347
rect 608 103 674 115
rect 704 347 770 359
rect 704 115 720 347
rect 754 115 770 347
rect 704 103 770 115
rect 800 347 866 359
rect 800 115 816 347
rect 850 115 866 347
rect 800 103 866 115
rect 896 347 962 359
rect 896 115 912 347
rect 946 115 962 347
rect 896 103 962 115
rect 992 347 1054 359
rect 992 115 1008 347
rect 1042 115 1054 347
rect 992 103 1054 115
<< ndiffc >>
rect 432 -318 466 -142
rect 528 -318 562 -142
rect 624 -318 658 -142
<< pdiffc >>
rect 48 115 82 347
rect 144 115 178 347
rect 240 115 274 347
rect 336 115 370 347
rect 432 115 466 347
rect 528 115 562 347
rect 624 115 658 347
rect 720 115 754 347
rect 816 115 850 347
rect 912 115 946 347
rect 1008 115 1042 347
<< psubdiff >>
rect 420 -401 670 -384
rect 420 -462 446 -401
rect 645 -462 670 -401
rect 420 -480 670 -462
<< nsubdiff >>
rect 46 502 466 544
rect 46 451 74 502
rect 431 451 466 502
rect 46 413 466 451
<< psubdiffcont >>
rect 446 -462 645 -401
<< nsubdiffcont >>
rect 74 451 431 502
<< poly >>
rect 98 359 128 385
rect 194 359 224 385
rect 290 359 320 385
rect 386 359 416 385
rect 482 359 512 385
rect 578 359 608 385
rect 674 359 704 385
rect 770 359 800 385
rect 866 359 896 385
rect 962 359 992 385
rect 98 77 128 103
rect 194 77 224 103
rect 290 77 320 103
rect 386 77 416 103
rect 482 77 512 103
rect 98 53 512 77
rect 98 19 433 53
rect 467 19 512 53
rect 98 6 512 19
rect 482 -130 512 6
rect 578 77 608 103
rect 674 77 704 103
rect 770 77 800 103
rect 866 77 896 103
rect 962 77 992 103
rect 578 6 992 77
rect 578 -36 608 6
rect 560 -52 626 -36
rect 560 -86 576 -52
rect 610 -86 626 -52
rect 560 -102 626 -86
rect 578 -130 608 -102
rect 482 -356 512 -330
rect 578 -356 608 -330
<< polycont >>
rect 433 19 467 53
rect 576 -86 610 -52
<< locali >>
rect 46 502 466 522
rect 46 451 74 502
rect 431 451 466 502
rect 46 432 466 451
rect 48 347 82 432
rect 48 99 82 115
rect 144 347 178 363
rect 144 99 178 115
rect 240 347 274 432
rect 240 99 274 115
rect 336 347 370 363
rect 336 99 370 115
rect 432 347 466 432
rect 432 99 466 115
rect 528 347 562 363
rect 528 99 562 115
rect 624 347 658 363
rect 624 99 658 115
rect 720 347 754 363
rect 720 99 754 115
rect 816 347 850 363
rect 816 99 850 115
rect 912 347 946 363
rect 912 99 946 115
rect 1008 347 1042 363
rect 1008 99 1042 115
rect 417 19 433 53
rect 467 19 483 53
rect 560 -86 576 -52
rect 610 -86 626 -52
rect 432 -142 466 -126
rect 432 -390 466 -318
rect 528 -142 562 -126
rect 528 -334 562 -318
rect 624 -142 658 -126
rect 624 -390 658 -318
rect 420 -401 670 -390
rect 420 -462 446 -401
rect 645 -462 670 -401
rect 420 -474 670 -462
<< viali >>
rect 74 451 431 502
rect 48 115 82 205
rect 144 257 178 347
rect 240 115 274 205
rect 336 257 370 347
rect 432 115 466 205
rect 528 257 562 347
rect 624 115 658 205
rect 720 257 754 347
rect 816 115 850 205
rect 912 257 946 347
rect 1008 115 1042 205
rect 433 19 467 53
rect 576 -86 610 -52
rect 528 -318 562 -142
rect 446 -462 645 -401
<< metal1 >>
rect 62 502 443 510
rect 62 451 74 502
rect 431 451 443 502
rect 62 444 443 451
rect 138 347 952 359
rect 138 257 144 347
rect 178 257 336 347
rect 370 257 528 347
rect 562 257 720 347
rect 754 257 912 347
rect 946 257 952 347
rect 138 245 952 257
rect 42 205 472 217
rect 42 115 48 205
rect 82 115 240 205
rect 274 115 432 205
rect 466 115 472 205
rect 42 103 472 115
rect 618 205 1090 217
rect 618 115 624 205
rect 658 115 816 205
rect 850 115 1008 205
rect 1042 115 1090 205
rect 618 103 1090 115
rect 0 53 526 69
rect 0 19 433 53
rect 467 19 526 53
rect 0 3 526 19
rect 0 -52 626 -36
rect 0 -86 576 -52
rect 610 -86 626 -52
rect 0 -102 626 -86
rect 522 -136 568 -130
rect 965 -136 1090 103
rect 522 -142 1090 -136
rect 522 -318 528 -142
rect 562 -318 1090 -142
rect 522 -330 1090 -318
rect 568 -334 1090 -330
rect 568 -335 1088 -334
rect 568 -336 1037 -335
rect 434 -401 657 -394
rect 434 -462 446 -401
rect 645 -462 657 -401
rect 434 -468 657 -462
<< labels >>
flabel metal1 7 10 84 62 1 FreeSerif 320 0 0 0 A
port 1 e
rlabel metal1 253 510 253 510 5 VDD
port 4 s
flabel metal1 8 -96 85 -44 1 FreeSerif 320 0 0 0 B
port 2 e
flabel metal1 1012 -102 1089 -50 1 FreeSerif 320 0 0 0 Y
port 5 e
rlabel metal1 549 -468 549 -468 5 VSS
port 3 s
<< end >>
