magic
tech sky130B
magscale 1 2
timestamp 1733166153
<< error_p >>
rect -596 -706 596 740
<< nwell >>
rect -596 -706 596 740
<< pmos >>
rect -502 -606 -442 678
rect -384 -606 -324 678
rect -266 -606 -206 678
rect -148 -606 -88 678
rect -30 -606 30 678
rect 88 -606 148 678
rect 206 -606 266 678
rect 324 -606 384 678
rect 442 -606 502 678
<< pdiff >>
rect -560 666 -502 678
rect -560 -594 -548 666
rect -514 -594 -502 666
rect -560 -606 -502 -594
rect -442 666 -384 678
rect -442 -594 -430 666
rect -396 -594 -384 666
rect -442 -606 -384 -594
rect -324 666 -266 678
rect -324 -594 -312 666
rect -278 -594 -266 666
rect -324 -606 -266 -594
rect -206 666 -148 678
rect -206 -594 -194 666
rect -160 -594 -148 666
rect -206 -606 -148 -594
rect -88 666 -30 678
rect -88 -594 -76 666
rect -42 -594 -30 666
rect -88 -606 -30 -594
rect 30 666 88 678
rect 30 -594 42 666
rect 76 -594 88 666
rect 30 -606 88 -594
rect 148 666 206 678
rect 148 -594 160 666
rect 194 -594 206 666
rect 148 -606 206 -594
rect 266 666 324 678
rect 266 -594 278 666
rect 312 -594 324 666
rect 266 -606 324 -594
rect 384 666 442 678
rect 384 -594 396 666
rect 430 -594 442 666
rect 384 -606 442 -594
rect 502 666 560 678
rect 502 -594 514 666
rect 548 -594 560 666
rect 502 -606 560 -594
<< pdiffc >>
rect -548 -594 -514 666
rect -430 -594 -396 666
rect -312 -594 -278 666
rect -194 -594 -160 666
rect -76 -594 -42 666
rect 42 -594 76 666
rect 160 -594 194 666
rect 278 -594 312 666
rect 396 -594 430 666
rect 514 -594 548 666
<< poly >>
rect -502 678 -442 704
rect -384 678 -324 704
rect -266 678 -206 704
rect -148 678 -88 704
rect -30 678 30 704
rect 88 678 148 704
rect 206 678 266 704
rect 324 678 384 704
rect 442 678 502 704
rect -502 -637 -442 -606
rect -384 -637 -324 -606
rect -266 -637 -206 -606
rect -148 -637 -88 -606
rect -30 -637 30 -606
rect 88 -637 148 -606
rect 206 -637 266 -606
rect 324 -637 384 -606
rect 442 -637 502 -606
rect -505 -653 -439 -637
rect -505 -687 -489 -653
rect -455 -687 -439 -653
rect -505 -703 -439 -687
rect -387 -653 -321 -637
rect -387 -687 -371 -653
rect -337 -687 -321 -653
rect -387 -703 -321 -687
rect -269 -653 -203 -637
rect -269 -687 -253 -653
rect -219 -687 -203 -653
rect -269 -703 -203 -687
rect -151 -653 -85 -637
rect -151 -687 -135 -653
rect -101 -687 -85 -653
rect -151 -703 -85 -687
rect -33 -653 33 -637
rect -33 -687 -17 -653
rect 17 -687 33 -653
rect -33 -703 33 -687
rect 85 -653 151 -637
rect 85 -687 101 -653
rect 135 -687 151 -653
rect 85 -703 151 -687
rect 203 -653 269 -637
rect 203 -687 219 -653
rect 253 -687 269 -653
rect 203 -703 269 -687
rect 321 -653 387 -637
rect 321 -687 337 -653
rect 371 -687 387 -653
rect 321 -703 387 -687
rect 439 -653 505 -637
rect 439 -687 455 -653
rect 489 -687 505 -653
rect 439 -703 505 -687
<< polycont >>
rect -489 -687 -455 -653
rect -371 -687 -337 -653
rect -253 -687 -219 -653
rect -135 -687 -101 -653
rect -17 -687 17 -653
rect 101 -687 135 -653
rect 219 -687 253 -653
rect 337 -687 371 -653
rect 455 -687 489 -653
<< locali >>
rect -548 666 -514 682
rect -548 -610 -514 -594
rect -430 666 -396 682
rect -430 -610 -396 -594
rect -312 666 -278 682
rect -312 -610 -278 -594
rect -194 666 -160 682
rect -194 -610 -160 -594
rect -76 666 -42 682
rect -76 -610 -42 -594
rect 42 666 76 682
rect 42 -610 76 -594
rect 160 666 194 682
rect 160 -610 194 -594
rect 278 666 312 682
rect 278 -610 312 -594
rect 396 666 430 682
rect 396 -610 430 -594
rect 514 666 548 682
rect 514 -610 548 -594
rect -505 -687 -489 -653
rect -455 -687 -439 -653
rect -387 -687 -371 -653
rect -337 -687 -321 -653
rect -269 -687 -253 -653
rect -219 -687 -203 -653
rect -151 -687 -135 -653
rect -101 -687 -85 -653
rect -33 -687 -17 -653
rect 17 -687 33 -653
rect 85 -687 101 -653
rect 135 -687 151 -653
rect 203 -687 219 -653
rect 253 -687 269 -653
rect 321 -687 337 -653
rect 371 -687 387 -653
rect 439 -687 455 -653
rect 489 -687 505 -653
<< viali >>
rect -548 -594 -514 666
rect -430 -594 -396 666
rect -312 -594 -278 666
rect -194 -594 -160 666
rect -76 -594 -42 666
rect 42 -594 76 666
rect 160 -594 194 666
rect 278 -594 312 666
rect 396 -594 430 666
rect 514 -594 548 666
<< metal1 >>
rect -554 666 -508 678
rect -554 -594 -548 666
rect -514 -594 -508 666
rect -554 -606 -508 -594
rect -436 666 -390 678
rect -436 -594 -430 666
rect -396 -594 -390 666
rect -436 -606 -390 -594
rect -318 666 -272 678
rect -318 -594 -312 666
rect -278 -594 -272 666
rect -318 -606 -272 -594
rect -200 666 -154 678
rect -200 -594 -194 666
rect -160 -594 -154 666
rect -200 -606 -154 -594
rect -82 666 -36 678
rect -82 -594 -76 666
rect -42 -594 -36 666
rect -82 -606 -36 -594
rect 36 666 82 678
rect 36 -594 42 666
rect 76 -594 82 666
rect 36 -606 82 -594
rect 154 666 200 678
rect 154 -594 160 666
rect 194 -594 200 666
rect 154 -606 200 -594
rect 272 666 318 678
rect 272 -594 278 666
rect 312 -594 318 666
rect 272 -606 318 -594
rect 390 666 436 678
rect 390 -594 396 666
rect 430 -594 436 666
rect 390 -606 436 -594
rect 508 666 554 678
rect 508 -594 514 666
rect 548 -594 554 666
rect 508 -606 554 -594
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.42 l 0.30 m 1 nf 9 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
