magic
tech sky130A
magscale 1 2
timestamp 1736606925
<< nwell >>
rect -3447 3502 -2268 4023
rect -1606 3502 -427 4023
rect 235 3502 1414 4023
rect 2076 3502 3255 4023
rect -3423 1730 -2244 2251
rect -1697 1730 -518 2251
rect -3423 438 -2244 959
rect -1697 438 -518 959
rect -3423 -1535 -2244 -1014
rect -1697 -1535 -518 -1014
rect -3423 -2827 -2244 -2306
rect -1697 -2827 -518 -2306
rect -3423 -4799 -2244 -4278
rect -1697 -4799 -518 -4278
rect -3423 -6091 -2244 -5570
rect -1697 -6091 -518 -5570
<< nmos >>
rect -3177 3342 -2777 3372
rect -2544 3346 -2344 3376
rect -1336 3342 -936 3372
rect -703 3346 -503 3376
rect 505 3342 905 3372
rect 1138 3346 1338 3376
rect 2346 3342 2746 3372
rect 2979 3346 3179 3376
rect -3177 3246 -2777 3276
rect -1336 3246 -936 3276
rect 505 3246 905 3276
rect 2346 3246 2746 3276
rect -3153 1570 -2753 1600
rect -2520 1574 -2320 1604
rect -1427 1570 -1027 1600
rect -794 1574 -594 1604
rect -3153 1474 -2753 1504
rect -1427 1474 -1027 1504
rect -3153 278 -2753 308
rect -2520 282 -2320 312
rect -1427 278 -1027 308
rect -794 282 -594 312
rect -3153 182 -2753 212
rect -1427 182 -1027 212
rect -3153 -1695 -2753 -1665
rect -2520 -1691 -2320 -1661
rect -1427 -1695 -1027 -1665
rect -794 -1691 -594 -1661
rect -3153 -1791 -2753 -1761
rect -1427 -1791 -1027 -1761
rect -3153 -2987 -2753 -2957
rect -2520 -2983 -2320 -2953
rect -1427 -2987 -1027 -2957
rect -794 -2983 -594 -2953
rect -3153 -3083 -2753 -3053
rect -1427 -3083 -1027 -3053
rect -3153 -4959 -2753 -4929
rect -2520 -4955 -2320 -4925
rect -1427 -4959 -1027 -4929
rect -794 -4955 -594 -4925
rect -3153 -5055 -2753 -5025
rect -1427 -5055 -1027 -5025
rect -3153 -6251 -2753 -6221
rect -2520 -6247 -2320 -6217
rect -1427 -6251 -1027 -6221
rect -794 -6247 -594 -6217
rect -3153 -6347 -2753 -6317
rect -1427 -6347 -1027 -6317
<< pmos >>
rect -3349 3564 -3319 3778
rect -3253 3564 -3223 3778
rect -3157 3564 -3127 3778
rect -3061 3564 -3031 3778
rect -2965 3564 -2935 3778
rect -2869 3564 -2839 3778
rect -2544 3792 -2330 3822
rect -2544 3696 -2330 3726
rect -2544 3600 -2330 3630
rect -1508 3564 -1478 3778
rect -1412 3564 -1382 3778
rect -1316 3564 -1286 3778
rect -1220 3564 -1190 3778
rect -1124 3564 -1094 3778
rect -1028 3564 -998 3778
rect -703 3792 -489 3822
rect -703 3696 -489 3726
rect -703 3600 -489 3630
rect 333 3564 363 3778
rect 429 3564 459 3778
rect 525 3564 555 3778
rect 621 3564 651 3778
rect 717 3564 747 3778
rect 813 3564 843 3778
rect 1138 3792 1352 3822
rect 1138 3696 1352 3726
rect 1138 3600 1352 3630
rect 2174 3564 2204 3778
rect 2270 3564 2300 3778
rect 2366 3564 2396 3778
rect 2462 3564 2492 3778
rect 2558 3564 2588 3778
rect 2654 3564 2684 3778
rect 2979 3792 3193 3822
rect 2979 3696 3193 3726
rect 2979 3600 3193 3630
rect -3325 1792 -3295 2006
rect -3229 1792 -3199 2006
rect -3133 1792 -3103 2006
rect -3037 1792 -3007 2006
rect -2941 1792 -2911 2006
rect -2845 1792 -2815 2006
rect -2520 2020 -2306 2050
rect -2520 1924 -2306 1954
rect -2520 1828 -2306 1858
rect -1599 1792 -1569 2006
rect -1503 1792 -1473 2006
rect -1407 1792 -1377 2006
rect -1311 1792 -1281 2006
rect -1215 1792 -1185 2006
rect -1119 1792 -1089 2006
rect -794 2020 -580 2050
rect -794 1924 -580 1954
rect -794 1828 -580 1858
rect -3325 500 -3295 714
rect -3229 500 -3199 714
rect -3133 500 -3103 714
rect -3037 500 -3007 714
rect -2941 500 -2911 714
rect -2845 500 -2815 714
rect -2520 728 -2306 758
rect -2520 632 -2306 662
rect -2520 536 -2306 566
rect -1599 500 -1569 714
rect -1503 500 -1473 714
rect -1407 500 -1377 714
rect -1311 500 -1281 714
rect -1215 500 -1185 714
rect -1119 500 -1089 714
rect -794 728 -580 758
rect -794 632 -580 662
rect -794 536 -580 566
rect -3325 -1473 -3295 -1259
rect -3229 -1473 -3199 -1259
rect -3133 -1473 -3103 -1259
rect -3037 -1473 -3007 -1259
rect -2941 -1473 -2911 -1259
rect -2845 -1473 -2815 -1259
rect -2520 -1245 -2306 -1215
rect -2520 -1341 -2306 -1311
rect -2520 -1437 -2306 -1407
rect -1599 -1473 -1569 -1259
rect -1503 -1473 -1473 -1259
rect -1407 -1473 -1377 -1259
rect -1311 -1473 -1281 -1259
rect -1215 -1473 -1185 -1259
rect -1119 -1473 -1089 -1259
rect -794 -1245 -580 -1215
rect -794 -1341 -580 -1311
rect -794 -1437 -580 -1407
rect -3325 -2765 -3295 -2551
rect -3229 -2765 -3199 -2551
rect -3133 -2765 -3103 -2551
rect -3037 -2765 -3007 -2551
rect -2941 -2765 -2911 -2551
rect -2845 -2765 -2815 -2551
rect -2520 -2537 -2306 -2507
rect -2520 -2633 -2306 -2603
rect -2520 -2729 -2306 -2699
rect -1599 -2765 -1569 -2551
rect -1503 -2765 -1473 -2551
rect -1407 -2765 -1377 -2551
rect -1311 -2765 -1281 -2551
rect -1215 -2765 -1185 -2551
rect -1119 -2765 -1089 -2551
rect -794 -2537 -580 -2507
rect -794 -2633 -580 -2603
rect -794 -2729 -580 -2699
rect -3325 -4737 -3295 -4523
rect -3229 -4737 -3199 -4523
rect -3133 -4737 -3103 -4523
rect -3037 -4737 -3007 -4523
rect -2941 -4737 -2911 -4523
rect -2845 -4737 -2815 -4523
rect -2520 -4509 -2306 -4479
rect -2520 -4605 -2306 -4575
rect -2520 -4701 -2306 -4671
rect -1599 -4737 -1569 -4523
rect -1503 -4737 -1473 -4523
rect -1407 -4737 -1377 -4523
rect -1311 -4737 -1281 -4523
rect -1215 -4737 -1185 -4523
rect -1119 -4737 -1089 -4523
rect -794 -4509 -580 -4479
rect -794 -4605 -580 -4575
rect -794 -4701 -580 -4671
rect -3325 -6029 -3295 -5815
rect -3229 -6029 -3199 -5815
rect -3133 -6029 -3103 -5815
rect -3037 -6029 -3007 -5815
rect -2941 -6029 -2911 -5815
rect -2845 -6029 -2815 -5815
rect -2520 -5801 -2306 -5771
rect -2520 -5897 -2306 -5867
rect -2520 -5993 -2306 -5963
rect -1599 -6029 -1569 -5815
rect -1503 -6029 -1473 -5815
rect -1407 -6029 -1377 -5815
rect -1311 -6029 -1281 -5815
rect -1215 -6029 -1185 -5815
rect -1119 -6029 -1089 -5815
rect -794 -5801 -580 -5771
rect -794 -5897 -580 -5867
rect -794 -5993 -580 -5963
<< ndiff >>
rect -3177 3422 -2777 3434
rect -3177 3388 -3165 3422
rect -2789 3388 -2777 3422
rect -2544 3422 -2344 3434
rect -3177 3372 -2777 3388
rect -2544 3388 -2532 3422
rect -2356 3388 -2344 3422
rect -2544 3376 -2344 3388
rect -3177 3276 -2777 3342
rect -2544 3334 -2344 3346
rect -2544 3300 -2532 3334
rect -2356 3300 -2344 3334
rect -2544 3288 -2344 3300
rect -1336 3422 -936 3434
rect -1336 3388 -1324 3422
rect -948 3388 -936 3422
rect -703 3422 -503 3434
rect -1336 3372 -936 3388
rect -703 3388 -691 3422
rect -515 3388 -503 3422
rect -703 3376 -503 3388
rect -1336 3276 -936 3342
rect -703 3334 -503 3346
rect -703 3300 -691 3334
rect -515 3300 -503 3334
rect -703 3288 -503 3300
rect 505 3422 905 3434
rect 505 3388 517 3422
rect 893 3388 905 3422
rect 1138 3422 1338 3434
rect 505 3372 905 3388
rect 1138 3388 1150 3422
rect 1326 3388 1338 3422
rect 1138 3376 1338 3388
rect 505 3276 905 3342
rect 1138 3334 1338 3346
rect 1138 3300 1150 3334
rect 1326 3300 1338 3334
rect 1138 3288 1338 3300
rect 2346 3422 2746 3434
rect 2346 3388 2358 3422
rect 2734 3388 2746 3422
rect 2979 3422 3179 3434
rect 2346 3372 2746 3388
rect 2979 3388 2991 3422
rect 3167 3388 3179 3422
rect 2979 3376 3179 3388
rect 2346 3276 2746 3342
rect 2979 3334 3179 3346
rect 2979 3300 2991 3334
rect 3167 3300 3179 3334
rect 2979 3288 3179 3300
rect -3177 3230 -2777 3246
rect -3177 3196 -3165 3230
rect -2789 3196 -2777 3230
rect -1336 3230 -936 3246
rect -3177 3184 -2777 3196
rect -1336 3196 -1324 3230
rect -948 3196 -936 3230
rect 505 3230 905 3246
rect -1336 3184 -936 3196
rect 505 3196 517 3230
rect 893 3196 905 3230
rect 2346 3230 2746 3246
rect 505 3184 905 3196
rect 2346 3196 2358 3230
rect 2734 3196 2746 3230
rect 2346 3184 2746 3196
rect -3153 1650 -2753 1662
rect -3153 1616 -3141 1650
rect -2765 1616 -2753 1650
rect -2520 1650 -2320 1662
rect -3153 1600 -2753 1616
rect -2520 1616 -2508 1650
rect -2332 1616 -2320 1650
rect -2520 1604 -2320 1616
rect -3153 1504 -2753 1570
rect -2520 1562 -2320 1574
rect -2520 1528 -2508 1562
rect -2332 1528 -2320 1562
rect -2520 1516 -2320 1528
rect -1427 1650 -1027 1662
rect -1427 1616 -1415 1650
rect -1039 1616 -1027 1650
rect -794 1650 -594 1662
rect -1427 1600 -1027 1616
rect -794 1616 -782 1650
rect -606 1616 -594 1650
rect -794 1604 -594 1616
rect -1427 1504 -1027 1570
rect -794 1562 -594 1574
rect -794 1528 -782 1562
rect -606 1528 -594 1562
rect -794 1516 -594 1528
rect -3153 1458 -2753 1474
rect -3153 1424 -3141 1458
rect -2765 1424 -2753 1458
rect -1427 1458 -1027 1474
rect -3153 1412 -2753 1424
rect -1427 1424 -1415 1458
rect -1039 1424 -1027 1458
rect -1427 1412 -1027 1424
rect -3153 358 -2753 370
rect -3153 324 -3141 358
rect -2765 324 -2753 358
rect -2520 358 -2320 370
rect -3153 308 -2753 324
rect -2520 324 -2508 358
rect -2332 324 -2320 358
rect -2520 312 -2320 324
rect -3153 212 -2753 278
rect -2520 270 -2320 282
rect -2520 236 -2508 270
rect -2332 236 -2320 270
rect -2520 224 -2320 236
rect -1427 358 -1027 370
rect -1427 324 -1415 358
rect -1039 324 -1027 358
rect -794 358 -594 370
rect -1427 308 -1027 324
rect -794 324 -782 358
rect -606 324 -594 358
rect -794 312 -594 324
rect -1427 212 -1027 278
rect -794 270 -594 282
rect -794 236 -782 270
rect -606 236 -594 270
rect -794 224 -594 236
rect -3153 166 -2753 182
rect -3153 132 -3141 166
rect -2765 132 -2753 166
rect -1427 166 -1027 182
rect -3153 120 -2753 132
rect -1427 132 -1415 166
rect -1039 132 -1027 166
rect -1427 120 -1027 132
rect -3153 -1615 -2753 -1603
rect -3153 -1649 -3141 -1615
rect -2765 -1649 -2753 -1615
rect -2520 -1615 -2320 -1603
rect -3153 -1665 -2753 -1649
rect -2520 -1649 -2508 -1615
rect -2332 -1649 -2320 -1615
rect -2520 -1661 -2320 -1649
rect -3153 -1761 -2753 -1695
rect -2520 -1703 -2320 -1691
rect -2520 -1737 -2508 -1703
rect -2332 -1737 -2320 -1703
rect -2520 -1749 -2320 -1737
rect -1427 -1615 -1027 -1603
rect -1427 -1649 -1415 -1615
rect -1039 -1649 -1027 -1615
rect -794 -1615 -594 -1603
rect -1427 -1665 -1027 -1649
rect -794 -1649 -782 -1615
rect -606 -1649 -594 -1615
rect -794 -1661 -594 -1649
rect -1427 -1761 -1027 -1695
rect -794 -1703 -594 -1691
rect -794 -1737 -782 -1703
rect -606 -1737 -594 -1703
rect -794 -1749 -594 -1737
rect -3153 -1807 -2753 -1791
rect -3153 -1841 -3141 -1807
rect -2765 -1841 -2753 -1807
rect -1427 -1807 -1027 -1791
rect -3153 -1853 -2753 -1841
rect -1427 -1841 -1415 -1807
rect -1039 -1841 -1027 -1807
rect -1427 -1853 -1027 -1841
rect -3153 -2907 -2753 -2895
rect -3153 -2941 -3141 -2907
rect -2765 -2941 -2753 -2907
rect -2520 -2907 -2320 -2895
rect -3153 -2957 -2753 -2941
rect -2520 -2941 -2508 -2907
rect -2332 -2941 -2320 -2907
rect -2520 -2953 -2320 -2941
rect -3153 -3053 -2753 -2987
rect -2520 -2995 -2320 -2983
rect -2520 -3029 -2508 -2995
rect -2332 -3029 -2320 -2995
rect -2520 -3041 -2320 -3029
rect -1427 -2907 -1027 -2895
rect -1427 -2941 -1415 -2907
rect -1039 -2941 -1027 -2907
rect -794 -2907 -594 -2895
rect -1427 -2957 -1027 -2941
rect -794 -2941 -782 -2907
rect -606 -2941 -594 -2907
rect -794 -2953 -594 -2941
rect -1427 -3053 -1027 -2987
rect -794 -2995 -594 -2983
rect -794 -3029 -782 -2995
rect -606 -3029 -594 -2995
rect -794 -3041 -594 -3029
rect -3153 -3099 -2753 -3083
rect -3153 -3133 -3141 -3099
rect -2765 -3133 -2753 -3099
rect -1427 -3099 -1027 -3083
rect -3153 -3145 -2753 -3133
rect -1427 -3133 -1415 -3099
rect -1039 -3133 -1027 -3099
rect -1427 -3145 -1027 -3133
rect -3153 -4879 -2753 -4867
rect -3153 -4913 -3141 -4879
rect -2765 -4913 -2753 -4879
rect -2520 -4879 -2320 -4867
rect -3153 -4929 -2753 -4913
rect -2520 -4913 -2508 -4879
rect -2332 -4913 -2320 -4879
rect -2520 -4925 -2320 -4913
rect -3153 -5025 -2753 -4959
rect -2520 -4967 -2320 -4955
rect -2520 -5001 -2508 -4967
rect -2332 -5001 -2320 -4967
rect -2520 -5013 -2320 -5001
rect -1427 -4879 -1027 -4867
rect -1427 -4913 -1415 -4879
rect -1039 -4913 -1027 -4879
rect -794 -4879 -594 -4867
rect -1427 -4929 -1027 -4913
rect -794 -4913 -782 -4879
rect -606 -4913 -594 -4879
rect -794 -4925 -594 -4913
rect -1427 -5025 -1027 -4959
rect -794 -4967 -594 -4955
rect -794 -5001 -782 -4967
rect -606 -5001 -594 -4967
rect -794 -5013 -594 -5001
rect -3153 -5071 -2753 -5055
rect -3153 -5105 -3141 -5071
rect -2765 -5105 -2753 -5071
rect -1427 -5071 -1027 -5055
rect -3153 -5117 -2753 -5105
rect -1427 -5105 -1415 -5071
rect -1039 -5105 -1027 -5071
rect -1427 -5117 -1027 -5105
rect -3153 -6171 -2753 -6159
rect -3153 -6205 -3141 -6171
rect -2765 -6205 -2753 -6171
rect -2520 -6171 -2320 -6159
rect -3153 -6221 -2753 -6205
rect -2520 -6205 -2508 -6171
rect -2332 -6205 -2320 -6171
rect -2520 -6217 -2320 -6205
rect -3153 -6317 -2753 -6251
rect -2520 -6259 -2320 -6247
rect -2520 -6293 -2508 -6259
rect -2332 -6293 -2320 -6259
rect -2520 -6305 -2320 -6293
rect -1427 -6171 -1027 -6159
rect -1427 -6205 -1415 -6171
rect -1039 -6205 -1027 -6171
rect -794 -6171 -594 -6159
rect -1427 -6221 -1027 -6205
rect -794 -6205 -782 -6171
rect -606 -6205 -594 -6171
rect -794 -6217 -594 -6205
rect -1427 -6317 -1027 -6251
rect -794 -6259 -594 -6247
rect -794 -6293 -782 -6259
rect -606 -6293 -594 -6259
rect -794 -6305 -594 -6293
rect -3153 -6363 -2753 -6347
rect -3153 -6397 -3141 -6363
rect -2765 -6397 -2753 -6363
rect -1427 -6363 -1027 -6347
rect -3153 -6409 -2753 -6397
rect -1427 -6397 -1415 -6363
rect -1039 -6397 -1027 -6363
rect -1427 -6409 -1027 -6397
<< pdiff >>
rect -2544 3872 -2330 3884
rect -3411 3766 -3349 3778
rect -3411 3576 -3399 3766
rect -3365 3576 -3349 3766
rect -3411 3564 -3349 3576
rect -3319 3766 -3253 3778
rect -3319 3576 -3303 3766
rect -3269 3576 -3253 3766
rect -3319 3564 -3253 3576
rect -3223 3766 -3157 3778
rect -3223 3576 -3207 3766
rect -3173 3576 -3157 3766
rect -3223 3564 -3157 3576
rect -3127 3766 -3061 3778
rect -3127 3576 -3111 3766
rect -3077 3576 -3061 3766
rect -3127 3564 -3061 3576
rect -3031 3766 -2965 3778
rect -3031 3576 -3015 3766
rect -2981 3576 -2965 3766
rect -3031 3564 -2965 3576
rect -2935 3766 -2869 3778
rect -2935 3576 -2919 3766
rect -2885 3576 -2869 3766
rect -2935 3564 -2869 3576
rect -2839 3766 -2777 3778
rect -2839 3576 -2823 3766
rect -2789 3576 -2777 3766
rect -2544 3838 -2532 3872
rect -2342 3838 -2330 3872
rect -2544 3822 -2330 3838
rect -703 3872 -489 3884
rect -2544 3776 -2330 3792
rect -2544 3742 -2532 3776
rect -2338 3742 -2330 3776
rect -2544 3726 -2330 3742
rect -1570 3766 -1508 3778
rect -2544 3680 -2330 3696
rect -2544 3646 -2532 3680
rect -2342 3646 -2330 3680
rect -2544 3630 -2330 3646
rect -2544 3584 -2330 3600
rect -2839 3564 -2777 3576
rect -2544 3550 -2532 3584
rect -2338 3550 -2330 3584
rect -1570 3576 -1558 3766
rect -1524 3576 -1508 3766
rect -1570 3564 -1508 3576
rect -1478 3766 -1412 3778
rect -1478 3576 -1462 3766
rect -1428 3576 -1412 3766
rect -1478 3564 -1412 3576
rect -1382 3766 -1316 3778
rect -1382 3576 -1366 3766
rect -1332 3576 -1316 3766
rect -1382 3564 -1316 3576
rect -1286 3766 -1220 3778
rect -1286 3576 -1270 3766
rect -1236 3576 -1220 3766
rect -1286 3564 -1220 3576
rect -1190 3766 -1124 3778
rect -1190 3576 -1174 3766
rect -1140 3576 -1124 3766
rect -1190 3564 -1124 3576
rect -1094 3766 -1028 3778
rect -1094 3576 -1078 3766
rect -1044 3576 -1028 3766
rect -1094 3564 -1028 3576
rect -998 3766 -936 3778
rect -998 3576 -982 3766
rect -948 3576 -936 3766
rect -703 3838 -691 3872
rect -501 3838 -489 3872
rect -703 3822 -489 3838
rect 1138 3872 1352 3884
rect -703 3776 -489 3792
rect -703 3742 -691 3776
rect -497 3742 -489 3776
rect -703 3726 -489 3742
rect 271 3766 333 3778
rect -703 3680 -489 3696
rect -703 3646 -691 3680
rect -501 3646 -489 3680
rect -703 3630 -489 3646
rect -703 3584 -489 3600
rect -998 3564 -936 3576
rect -2544 3538 -2330 3550
rect -703 3550 -691 3584
rect -497 3550 -489 3584
rect 271 3576 283 3766
rect 317 3576 333 3766
rect 271 3564 333 3576
rect 363 3766 429 3778
rect 363 3576 379 3766
rect 413 3576 429 3766
rect 363 3564 429 3576
rect 459 3766 525 3778
rect 459 3576 475 3766
rect 509 3576 525 3766
rect 459 3564 525 3576
rect 555 3766 621 3778
rect 555 3576 571 3766
rect 605 3576 621 3766
rect 555 3564 621 3576
rect 651 3766 717 3778
rect 651 3576 667 3766
rect 701 3576 717 3766
rect 651 3564 717 3576
rect 747 3766 813 3778
rect 747 3576 763 3766
rect 797 3576 813 3766
rect 747 3564 813 3576
rect 843 3766 905 3778
rect 843 3576 859 3766
rect 893 3576 905 3766
rect 1138 3838 1150 3872
rect 1340 3838 1352 3872
rect 1138 3822 1352 3838
rect 2979 3872 3193 3884
rect 1138 3776 1352 3792
rect 1138 3742 1150 3776
rect 1344 3742 1352 3776
rect 1138 3726 1352 3742
rect 2112 3766 2174 3778
rect 1138 3680 1352 3696
rect 1138 3646 1150 3680
rect 1340 3646 1352 3680
rect 1138 3630 1352 3646
rect 1138 3584 1352 3600
rect 843 3564 905 3576
rect -703 3538 -489 3550
rect 1138 3550 1150 3584
rect 1344 3550 1352 3584
rect 2112 3576 2124 3766
rect 2158 3576 2174 3766
rect 2112 3564 2174 3576
rect 2204 3766 2270 3778
rect 2204 3576 2220 3766
rect 2254 3576 2270 3766
rect 2204 3564 2270 3576
rect 2300 3766 2366 3778
rect 2300 3576 2316 3766
rect 2350 3576 2366 3766
rect 2300 3564 2366 3576
rect 2396 3766 2462 3778
rect 2396 3576 2412 3766
rect 2446 3576 2462 3766
rect 2396 3564 2462 3576
rect 2492 3766 2558 3778
rect 2492 3576 2508 3766
rect 2542 3576 2558 3766
rect 2492 3564 2558 3576
rect 2588 3766 2654 3778
rect 2588 3576 2604 3766
rect 2638 3576 2654 3766
rect 2588 3564 2654 3576
rect 2684 3766 2746 3778
rect 2684 3576 2700 3766
rect 2734 3576 2746 3766
rect 2979 3838 2991 3872
rect 3181 3838 3193 3872
rect 2979 3822 3193 3838
rect 2979 3776 3193 3792
rect 2979 3742 2991 3776
rect 3185 3742 3193 3776
rect 2979 3726 3193 3742
rect 2979 3680 3193 3696
rect 2979 3646 2991 3680
rect 3181 3646 3193 3680
rect 2979 3630 3193 3646
rect 2979 3584 3193 3600
rect 2684 3564 2746 3576
rect 1138 3538 1352 3550
rect 2979 3550 2991 3584
rect 3185 3550 3193 3584
rect 2979 3538 3193 3550
rect -2520 2100 -2306 2112
rect -3387 1994 -3325 2006
rect -3387 1804 -3375 1994
rect -3341 1804 -3325 1994
rect -3387 1792 -3325 1804
rect -3295 1994 -3229 2006
rect -3295 1804 -3279 1994
rect -3245 1804 -3229 1994
rect -3295 1792 -3229 1804
rect -3199 1994 -3133 2006
rect -3199 1804 -3183 1994
rect -3149 1804 -3133 1994
rect -3199 1792 -3133 1804
rect -3103 1994 -3037 2006
rect -3103 1804 -3087 1994
rect -3053 1804 -3037 1994
rect -3103 1792 -3037 1804
rect -3007 1994 -2941 2006
rect -3007 1804 -2991 1994
rect -2957 1804 -2941 1994
rect -3007 1792 -2941 1804
rect -2911 1994 -2845 2006
rect -2911 1804 -2895 1994
rect -2861 1804 -2845 1994
rect -2911 1792 -2845 1804
rect -2815 1994 -2753 2006
rect -2815 1804 -2799 1994
rect -2765 1804 -2753 1994
rect -2520 2066 -2508 2100
rect -2318 2066 -2306 2100
rect -2520 2050 -2306 2066
rect -794 2100 -580 2112
rect -2520 2004 -2306 2020
rect -2520 1970 -2508 2004
rect -2314 1970 -2306 2004
rect -2520 1954 -2306 1970
rect -1661 1994 -1599 2006
rect -2520 1908 -2306 1924
rect -2520 1874 -2508 1908
rect -2318 1874 -2306 1908
rect -2520 1858 -2306 1874
rect -2520 1812 -2306 1828
rect -2815 1792 -2753 1804
rect -2520 1778 -2508 1812
rect -2314 1778 -2306 1812
rect -1661 1804 -1649 1994
rect -1615 1804 -1599 1994
rect -1661 1792 -1599 1804
rect -1569 1994 -1503 2006
rect -1569 1804 -1553 1994
rect -1519 1804 -1503 1994
rect -1569 1792 -1503 1804
rect -1473 1994 -1407 2006
rect -1473 1804 -1457 1994
rect -1423 1804 -1407 1994
rect -1473 1792 -1407 1804
rect -1377 1994 -1311 2006
rect -1377 1804 -1361 1994
rect -1327 1804 -1311 1994
rect -1377 1792 -1311 1804
rect -1281 1994 -1215 2006
rect -1281 1804 -1265 1994
rect -1231 1804 -1215 1994
rect -1281 1792 -1215 1804
rect -1185 1994 -1119 2006
rect -1185 1804 -1169 1994
rect -1135 1804 -1119 1994
rect -1185 1792 -1119 1804
rect -1089 1994 -1027 2006
rect -1089 1804 -1073 1994
rect -1039 1804 -1027 1994
rect -794 2066 -782 2100
rect -592 2066 -580 2100
rect -794 2050 -580 2066
rect -794 2004 -580 2020
rect -794 1970 -782 2004
rect -588 1970 -580 2004
rect -794 1954 -580 1970
rect -794 1908 -580 1924
rect -794 1874 -782 1908
rect -592 1874 -580 1908
rect -794 1858 -580 1874
rect -794 1812 -580 1828
rect -1089 1792 -1027 1804
rect -2520 1766 -2306 1778
rect -794 1778 -782 1812
rect -588 1778 -580 1812
rect -794 1766 -580 1778
rect -2520 808 -2306 820
rect -3387 702 -3325 714
rect -3387 512 -3375 702
rect -3341 512 -3325 702
rect -3387 500 -3325 512
rect -3295 702 -3229 714
rect -3295 512 -3279 702
rect -3245 512 -3229 702
rect -3295 500 -3229 512
rect -3199 702 -3133 714
rect -3199 512 -3183 702
rect -3149 512 -3133 702
rect -3199 500 -3133 512
rect -3103 702 -3037 714
rect -3103 512 -3087 702
rect -3053 512 -3037 702
rect -3103 500 -3037 512
rect -3007 702 -2941 714
rect -3007 512 -2991 702
rect -2957 512 -2941 702
rect -3007 500 -2941 512
rect -2911 702 -2845 714
rect -2911 512 -2895 702
rect -2861 512 -2845 702
rect -2911 500 -2845 512
rect -2815 702 -2753 714
rect -2815 512 -2799 702
rect -2765 512 -2753 702
rect -2520 774 -2508 808
rect -2318 774 -2306 808
rect -2520 758 -2306 774
rect -794 808 -580 820
rect -2520 712 -2306 728
rect -2520 678 -2508 712
rect -2314 678 -2306 712
rect -2520 662 -2306 678
rect -1661 702 -1599 714
rect -2520 616 -2306 632
rect -2520 582 -2508 616
rect -2318 582 -2306 616
rect -2520 566 -2306 582
rect -2520 520 -2306 536
rect -2815 500 -2753 512
rect -2520 486 -2508 520
rect -2314 486 -2306 520
rect -1661 512 -1649 702
rect -1615 512 -1599 702
rect -1661 500 -1599 512
rect -1569 702 -1503 714
rect -1569 512 -1553 702
rect -1519 512 -1503 702
rect -1569 500 -1503 512
rect -1473 702 -1407 714
rect -1473 512 -1457 702
rect -1423 512 -1407 702
rect -1473 500 -1407 512
rect -1377 702 -1311 714
rect -1377 512 -1361 702
rect -1327 512 -1311 702
rect -1377 500 -1311 512
rect -1281 702 -1215 714
rect -1281 512 -1265 702
rect -1231 512 -1215 702
rect -1281 500 -1215 512
rect -1185 702 -1119 714
rect -1185 512 -1169 702
rect -1135 512 -1119 702
rect -1185 500 -1119 512
rect -1089 702 -1027 714
rect -1089 512 -1073 702
rect -1039 512 -1027 702
rect -794 774 -782 808
rect -592 774 -580 808
rect -794 758 -580 774
rect -794 712 -580 728
rect -794 678 -782 712
rect -588 678 -580 712
rect -794 662 -580 678
rect -794 616 -580 632
rect -794 582 -782 616
rect -592 582 -580 616
rect -794 566 -580 582
rect -794 520 -580 536
rect -1089 500 -1027 512
rect -2520 474 -2306 486
rect -794 486 -782 520
rect -588 486 -580 520
rect -794 474 -580 486
rect -2520 -1165 -2306 -1153
rect -3387 -1271 -3325 -1259
rect -3387 -1461 -3375 -1271
rect -3341 -1461 -3325 -1271
rect -3387 -1473 -3325 -1461
rect -3295 -1271 -3229 -1259
rect -3295 -1461 -3279 -1271
rect -3245 -1461 -3229 -1271
rect -3295 -1473 -3229 -1461
rect -3199 -1271 -3133 -1259
rect -3199 -1461 -3183 -1271
rect -3149 -1461 -3133 -1271
rect -3199 -1473 -3133 -1461
rect -3103 -1271 -3037 -1259
rect -3103 -1461 -3087 -1271
rect -3053 -1461 -3037 -1271
rect -3103 -1473 -3037 -1461
rect -3007 -1271 -2941 -1259
rect -3007 -1461 -2991 -1271
rect -2957 -1461 -2941 -1271
rect -3007 -1473 -2941 -1461
rect -2911 -1271 -2845 -1259
rect -2911 -1461 -2895 -1271
rect -2861 -1461 -2845 -1271
rect -2911 -1473 -2845 -1461
rect -2815 -1271 -2753 -1259
rect -2815 -1461 -2799 -1271
rect -2765 -1461 -2753 -1271
rect -2520 -1199 -2508 -1165
rect -2318 -1199 -2306 -1165
rect -2520 -1215 -2306 -1199
rect -794 -1165 -580 -1153
rect -2520 -1261 -2306 -1245
rect -2520 -1295 -2508 -1261
rect -2314 -1295 -2306 -1261
rect -2520 -1311 -2306 -1295
rect -1661 -1271 -1599 -1259
rect -2520 -1357 -2306 -1341
rect -2520 -1391 -2508 -1357
rect -2318 -1391 -2306 -1357
rect -2520 -1407 -2306 -1391
rect -2520 -1453 -2306 -1437
rect -2815 -1473 -2753 -1461
rect -2520 -1487 -2508 -1453
rect -2314 -1487 -2306 -1453
rect -1661 -1461 -1649 -1271
rect -1615 -1461 -1599 -1271
rect -1661 -1473 -1599 -1461
rect -1569 -1271 -1503 -1259
rect -1569 -1461 -1553 -1271
rect -1519 -1461 -1503 -1271
rect -1569 -1473 -1503 -1461
rect -1473 -1271 -1407 -1259
rect -1473 -1461 -1457 -1271
rect -1423 -1461 -1407 -1271
rect -1473 -1473 -1407 -1461
rect -1377 -1271 -1311 -1259
rect -1377 -1461 -1361 -1271
rect -1327 -1461 -1311 -1271
rect -1377 -1473 -1311 -1461
rect -1281 -1271 -1215 -1259
rect -1281 -1461 -1265 -1271
rect -1231 -1461 -1215 -1271
rect -1281 -1473 -1215 -1461
rect -1185 -1271 -1119 -1259
rect -1185 -1461 -1169 -1271
rect -1135 -1461 -1119 -1271
rect -1185 -1473 -1119 -1461
rect -1089 -1271 -1027 -1259
rect -1089 -1461 -1073 -1271
rect -1039 -1461 -1027 -1271
rect -794 -1199 -782 -1165
rect -592 -1199 -580 -1165
rect -794 -1215 -580 -1199
rect -794 -1261 -580 -1245
rect -794 -1295 -782 -1261
rect -588 -1295 -580 -1261
rect -794 -1311 -580 -1295
rect -794 -1357 -580 -1341
rect -794 -1391 -782 -1357
rect -592 -1391 -580 -1357
rect -794 -1407 -580 -1391
rect -794 -1453 -580 -1437
rect -1089 -1473 -1027 -1461
rect -2520 -1499 -2306 -1487
rect -794 -1487 -782 -1453
rect -588 -1487 -580 -1453
rect -794 -1499 -580 -1487
rect -2520 -2457 -2306 -2445
rect -3387 -2563 -3325 -2551
rect -3387 -2753 -3375 -2563
rect -3341 -2753 -3325 -2563
rect -3387 -2765 -3325 -2753
rect -3295 -2563 -3229 -2551
rect -3295 -2753 -3279 -2563
rect -3245 -2753 -3229 -2563
rect -3295 -2765 -3229 -2753
rect -3199 -2563 -3133 -2551
rect -3199 -2753 -3183 -2563
rect -3149 -2753 -3133 -2563
rect -3199 -2765 -3133 -2753
rect -3103 -2563 -3037 -2551
rect -3103 -2753 -3087 -2563
rect -3053 -2753 -3037 -2563
rect -3103 -2765 -3037 -2753
rect -3007 -2563 -2941 -2551
rect -3007 -2753 -2991 -2563
rect -2957 -2753 -2941 -2563
rect -3007 -2765 -2941 -2753
rect -2911 -2563 -2845 -2551
rect -2911 -2753 -2895 -2563
rect -2861 -2753 -2845 -2563
rect -2911 -2765 -2845 -2753
rect -2815 -2563 -2753 -2551
rect -2815 -2753 -2799 -2563
rect -2765 -2753 -2753 -2563
rect -2520 -2491 -2508 -2457
rect -2318 -2491 -2306 -2457
rect -2520 -2507 -2306 -2491
rect -794 -2457 -580 -2445
rect -2520 -2553 -2306 -2537
rect -2520 -2587 -2508 -2553
rect -2314 -2587 -2306 -2553
rect -2520 -2603 -2306 -2587
rect -1661 -2563 -1599 -2551
rect -2520 -2649 -2306 -2633
rect -2520 -2683 -2508 -2649
rect -2318 -2683 -2306 -2649
rect -2520 -2699 -2306 -2683
rect -2520 -2745 -2306 -2729
rect -2815 -2765 -2753 -2753
rect -2520 -2779 -2508 -2745
rect -2314 -2779 -2306 -2745
rect -1661 -2753 -1649 -2563
rect -1615 -2753 -1599 -2563
rect -1661 -2765 -1599 -2753
rect -1569 -2563 -1503 -2551
rect -1569 -2753 -1553 -2563
rect -1519 -2753 -1503 -2563
rect -1569 -2765 -1503 -2753
rect -1473 -2563 -1407 -2551
rect -1473 -2753 -1457 -2563
rect -1423 -2753 -1407 -2563
rect -1473 -2765 -1407 -2753
rect -1377 -2563 -1311 -2551
rect -1377 -2753 -1361 -2563
rect -1327 -2753 -1311 -2563
rect -1377 -2765 -1311 -2753
rect -1281 -2563 -1215 -2551
rect -1281 -2753 -1265 -2563
rect -1231 -2753 -1215 -2563
rect -1281 -2765 -1215 -2753
rect -1185 -2563 -1119 -2551
rect -1185 -2753 -1169 -2563
rect -1135 -2753 -1119 -2563
rect -1185 -2765 -1119 -2753
rect -1089 -2563 -1027 -2551
rect -1089 -2753 -1073 -2563
rect -1039 -2753 -1027 -2563
rect -794 -2491 -782 -2457
rect -592 -2491 -580 -2457
rect -794 -2507 -580 -2491
rect -794 -2553 -580 -2537
rect -794 -2587 -782 -2553
rect -588 -2587 -580 -2553
rect -794 -2603 -580 -2587
rect -794 -2649 -580 -2633
rect -794 -2683 -782 -2649
rect -592 -2683 -580 -2649
rect -794 -2699 -580 -2683
rect -794 -2745 -580 -2729
rect -1089 -2765 -1027 -2753
rect -2520 -2791 -2306 -2779
rect -794 -2779 -782 -2745
rect -588 -2779 -580 -2745
rect -794 -2791 -580 -2779
rect -2520 -4429 -2306 -4417
rect -3387 -4535 -3325 -4523
rect -3387 -4725 -3375 -4535
rect -3341 -4725 -3325 -4535
rect -3387 -4737 -3325 -4725
rect -3295 -4535 -3229 -4523
rect -3295 -4725 -3279 -4535
rect -3245 -4725 -3229 -4535
rect -3295 -4737 -3229 -4725
rect -3199 -4535 -3133 -4523
rect -3199 -4725 -3183 -4535
rect -3149 -4725 -3133 -4535
rect -3199 -4737 -3133 -4725
rect -3103 -4535 -3037 -4523
rect -3103 -4725 -3087 -4535
rect -3053 -4725 -3037 -4535
rect -3103 -4737 -3037 -4725
rect -3007 -4535 -2941 -4523
rect -3007 -4725 -2991 -4535
rect -2957 -4725 -2941 -4535
rect -3007 -4737 -2941 -4725
rect -2911 -4535 -2845 -4523
rect -2911 -4725 -2895 -4535
rect -2861 -4725 -2845 -4535
rect -2911 -4737 -2845 -4725
rect -2815 -4535 -2753 -4523
rect -2815 -4725 -2799 -4535
rect -2765 -4725 -2753 -4535
rect -2520 -4463 -2508 -4429
rect -2318 -4463 -2306 -4429
rect -2520 -4479 -2306 -4463
rect -794 -4429 -580 -4417
rect -2520 -4525 -2306 -4509
rect -2520 -4559 -2508 -4525
rect -2314 -4559 -2306 -4525
rect -2520 -4575 -2306 -4559
rect -1661 -4535 -1599 -4523
rect -2520 -4621 -2306 -4605
rect -2520 -4655 -2508 -4621
rect -2318 -4655 -2306 -4621
rect -2520 -4671 -2306 -4655
rect -2520 -4717 -2306 -4701
rect -2815 -4737 -2753 -4725
rect -2520 -4751 -2508 -4717
rect -2314 -4751 -2306 -4717
rect -1661 -4725 -1649 -4535
rect -1615 -4725 -1599 -4535
rect -1661 -4737 -1599 -4725
rect -1569 -4535 -1503 -4523
rect -1569 -4725 -1553 -4535
rect -1519 -4725 -1503 -4535
rect -1569 -4737 -1503 -4725
rect -1473 -4535 -1407 -4523
rect -1473 -4725 -1457 -4535
rect -1423 -4725 -1407 -4535
rect -1473 -4737 -1407 -4725
rect -1377 -4535 -1311 -4523
rect -1377 -4725 -1361 -4535
rect -1327 -4725 -1311 -4535
rect -1377 -4737 -1311 -4725
rect -1281 -4535 -1215 -4523
rect -1281 -4725 -1265 -4535
rect -1231 -4725 -1215 -4535
rect -1281 -4737 -1215 -4725
rect -1185 -4535 -1119 -4523
rect -1185 -4725 -1169 -4535
rect -1135 -4725 -1119 -4535
rect -1185 -4737 -1119 -4725
rect -1089 -4535 -1027 -4523
rect -1089 -4725 -1073 -4535
rect -1039 -4725 -1027 -4535
rect -794 -4463 -782 -4429
rect -592 -4463 -580 -4429
rect -794 -4479 -580 -4463
rect -794 -4525 -580 -4509
rect -794 -4559 -782 -4525
rect -588 -4559 -580 -4525
rect -794 -4575 -580 -4559
rect -794 -4621 -580 -4605
rect -794 -4655 -782 -4621
rect -592 -4655 -580 -4621
rect -794 -4671 -580 -4655
rect -794 -4717 -580 -4701
rect -1089 -4737 -1027 -4725
rect -2520 -4763 -2306 -4751
rect -794 -4751 -782 -4717
rect -588 -4751 -580 -4717
rect -794 -4763 -580 -4751
rect -2520 -5721 -2306 -5709
rect -3387 -5827 -3325 -5815
rect -3387 -6017 -3375 -5827
rect -3341 -6017 -3325 -5827
rect -3387 -6029 -3325 -6017
rect -3295 -5827 -3229 -5815
rect -3295 -6017 -3279 -5827
rect -3245 -6017 -3229 -5827
rect -3295 -6029 -3229 -6017
rect -3199 -5827 -3133 -5815
rect -3199 -6017 -3183 -5827
rect -3149 -6017 -3133 -5827
rect -3199 -6029 -3133 -6017
rect -3103 -5827 -3037 -5815
rect -3103 -6017 -3087 -5827
rect -3053 -6017 -3037 -5827
rect -3103 -6029 -3037 -6017
rect -3007 -5827 -2941 -5815
rect -3007 -6017 -2991 -5827
rect -2957 -6017 -2941 -5827
rect -3007 -6029 -2941 -6017
rect -2911 -5827 -2845 -5815
rect -2911 -6017 -2895 -5827
rect -2861 -6017 -2845 -5827
rect -2911 -6029 -2845 -6017
rect -2815 -5827 -2753 -5815
rect -2815 -6017 -2799 -5827
rect -2765 -6017 -2753 -5827
rect -2520 -5755 -2508 -5721
rect -2318 -5755 -2306 -5721
rect -2520 -5771 -2306 -5755
rect -794 -5721 -580 -5709
rect -2520 -5817 -2306 -5801
rect -2520 -5851 -2508 -5817
rect -2314 -5851 -2306 -5817
rect -2520 -5867 -2306 -5851
rect -1661 -5827 -1599 -5815
rect -2520 -5913 -2306 -5897
rect -2520 -5947 -2508 -5913
rect -2318 -5947 -2306 -5913
rect -2520 -5963 -2306 -5947
rect -2520 -6009 -2306 -5993
rect -2815 -6029 -2753 -6017
rect -2520 -6043 -2508 -6009
rect -2314 -6043 -2306 -6009
rect -1661 -6017 -1649 -5827
rect -1615 -6017 -1599 -5827
rect -1661 -6029 -1599 -6017
rect -1569 -5827 -1503 -5815
rect -1569 -6017 -1553 -5827
rect -1519 -6017 -1503 -5827
rect -1569 -6029 -1503 -6017
rect -1473 -5827 -1407 -5815
rect -1473 -6017 -1457 -5827
rect -1423 -6017 -1407 -5827
rect -1473 -6029 -1407 -6017
rect -1377 -5827 -1311 -5815
rect -1377 -6017 -1361 -5827
rect -1327 -6017 -1311 -5827
rect -1377 -6029 -1311 -6017
rect -1281 -5827 -1215 -5815
rect -1281 -6017 -1265 -5827
rect -1231 -6017 -1215 -5827
rect -1281 -6029 -1215 -6017
rect -1185 -5827 -1119 -5815
rect -1185 -6017 -1169 -5827
rect -1135 -6017 -1119 -5827
rect -1185 -6029 -1119 -6017
rect -1089 -5827 -1027 -5815
rect -1089 -6017 -1073 -5827
rect -1039 -6017 -1027 -5827
rect -794 -5755 -782 -5721
rect -592 -5755 -580 -5721
rect -794 -5771 -580 -5755
rect -794 -5817 -580 -5801
rect -794 -5851 -782 -5817
rect -588 -5851 -580 -5817
rect -794 -5867 -580 -5851
rect -794 -5913 -580 -5897
rect -794 -5947 -782 -5913
rect -592 -5947 -580 -5913
rect -794 -5963 -580 -5947
rect -794 -6009 -580 -5993
rect -1089 -6029 -1027 -6017
rect -2520 -6055 -2306 -6043
rect -794 -6043 -782 -6009
rect -588 -6043 -580 -6009
rect -794 -6055 -580 -6043
<< ndiffc >>
rect -3165 3388 -2789 3422
rect -2532 3388 -2356 3422
rect -2532 3300 -2356 3334
rect -1324 3388 -948 3422
rect -691 3388 -515 3422
rect -691 3300 -515 3334
rect 517 3388 893 3422
rect 1150 3388 1326 3422
rect 1150 3300 1326 3334
rect 2358 3388 2734 3422
rect 2991 3388 3167 3422
rect 2991 3300 3167 3334
rect -3165 3196 -2789 3230
rect -1324 3196 -948 3230
rect 517 3196 893 3230
rect 2358 3196 2734 3230
rect -3141 1616 -2765 1650
rect -2508 1616 -2332 1650
rect -2508 1528 -2332 1562
rect -1415 1616 -1039 1650
rect -782 1616 -606 1650
rect -782 1528 -606 1562
rect -3141 1424 -2765 1458
rect -1415 1424 -1039 1458
rect -3141 324 -2765 358
rect -2508 324 -2332 358
rect -2508 236 -2332 270
rect -1415 324 -1039 358
rect -782 324 -606 358
rect -782 236 -606 270
rect -3141 132 -2765 166
rect -1415 132 -1039 166
rect -3141 -1649 -2765 -1615
rect -2508 -1649 -2332 -1615
rect -2508 -1737 -2332 -1703
rect -1415 -1649 -1039 -1615
rect -782 -1649 -606 -1615
rect -782 -1737 -606 -1703
rect -3141 -1841 -2765 -1807
rect -1415 -1841 -1039 -1807
rect -3141 -2941 -2765 -2907
rect -2508 -2941 -2332 -2907
rect -2508 -3029 -2332 -2995
rect -1415 -2941 -1039 -2907
rect -782 -2941 -606 -2907
rect -782 -3029 -606 -2995
rect -3141 -3133 -2765 -3099
rect -1415 -3133 -1039 -3099
rect -3141 -4913 -2765 -4879
rect -2508 -4913 -2332 -4879
rect -2508 -5001 -2332 -4967
rect -1415 -4913 -1039 -4879
rect -782 -4913 -606 -4879
rect -782 -5001 -606 -4967
rect -3141 -5105 -2765 -5071
rect -1415 -5105 -1039 -5071
rect -3141 -6205 -2765 -6171
rect -2508 -6205 -2332 -6171
rect -2508 -6293 -2332 -6259
rect -1415 -6205 -1039 -6171
rect -782 -6205 -606 -6171
rect -782 -6293 -606 -6259
rect -3141 -6397 -2765 -6363
rect -1415 -6397 -1039 -6363
<< pdiffc >>
rect -3399 3576 -3365 3766
rect -3303 3576 -3269 3766
rect -3207 3576 -3173 3766
rect -3111 3576 -3077 3766
rect -3015 3576 -2981 3766
rect -2919 3576 -2885 3766
rect -2823 3576 -2789 3766
rect -2532 3838 -2342 3872
rect -2532 3742 -2338 3776
rect -2532 3646 -2342 3680
rect -2532 3550 -2338 3584
rect -1558 3576 -1524 3766
rect -1462 3576 -1428 3766
rect -1366 3576 -1332 3766
rect -1270 3576 -1236 3766
rect -1174 3576 -1140 3766
rect -1078 3576 -1044 3766
rect -982 3576 -948 3766
rect -691 3838 -501 3872
rect -691 3742 -497 3776
rect -691 3646 -501 3680
rect -691 3550 -497 3584
rect 283 3576 317 3766
rect 379 3576 413 3766
rect 475 3576 509 3766
rect 571 3576 605 3766
rect 667 3576 701 3766
rect 763 3576 797 3766
rect 859 3576 893 3766
rect 1150 3838 1340 3872
rect 1150 3742 1344 3776
rect 1150 3646 1340 3680
rect 1150 3550 1344 3584
rect 2124 3576 2158 3766
rect 2220 3576 2254 3766
rect 2316 3576 2350 3766
rect 2412 3576 2446 3766
rect 2508 3576 2542 3766
rect 2604 3576 2638 3766
rect 2700 3576 2734 3766
rect 2991 3838 3181 3872
rect 2991 3742 3185 3776
rect 2991 3646 3181 3680
rect 2991 3550 3185 3584
rect -3375 1804 -3341 1994
rect -3279 1804 -3245 1994
rect -3183 1804 -3149 1994
rect -3087 1804 -3053 1994
rect -2991 1804 -2957 1994
rect -2895 1804 -2861 1994
rect -2799 1804 -2765 1994
rect -2508 2066 -2318 2100
rect -2508 1970 -2314 2004
rect -2508 1874 -2318 1908
rect -2508 1778 -2314 1812
rect -1649 1804 -1615 1994
rect -1553 1804 -1519 1994
rect -1457 1804 -1423 1994
rect -1361 1804 -1327 1994
rect -1265 1804 -1231 1994
rect -1169 1804 -1135 1994
rect -1073 1804 -1039 1994
rect -782 2066 -592 2100
rect -782 1970 -588 2004
rect -782 1874 -592 1908
rect -782 1778 -588 1812
rect -3375 512 -3341 702
rect -3279 512 -3245 702
rect -3183 512 -3149 702
rect -3087 512 -3053 702
rect -2991 512 -2957 702
rect -2895 512 -2861 702
rect -2799 512 -2765 702
rect -2508 774 -2318 808
rect -2508 678 -2314 712
rect -2508 582 -2318 616
rect -2508 486 -2314 520
rect -1649 512 -1615 702
rect -1553 512 -1519 702
rect -1457 512 -1423 702
rect -1361 512 -1327 702
rect -1265 512 -1231 702
rect -1169 512 -1135 702
rect -1073 512 -1039 702
rect -782 774 -592 808
rect -782 678 -588 712
rect -782 582 -592 616
rect -782 486 -588 520
rect -3375 -1461 -3341 -1271
rect -3279 -1461 -3245 -1271
rect -3183 -1461 -3149 -1271
rect -3087 -1461 -3053 -1271
rect -2991 -1461 -2957 -1271
rect -2895 -1461 -2861 -1271
rect -2799 -1461 -2765 -1271
rect -2508 -1199 -2318 -1165
rect -2508 -1295 -2314 -1261
rect -2508 -1391 -2318 -1357
rect -2508 -1487 -2314 -1453
rect -1649 -1461 -1615 -1271
rect -1553 -1461 -1519 -1271
rect -1457 -1461 -1423 -1271
rect -1361 -1461 -1327 -1271
rect -1265 -1461 -1231 -1271
rect -1169 -1461 -1135 -1271
rect -1073 -1461 -1039 -1271
rect -782 -1199 -592 -1165
rect -782 -1295 -588 -1261
rect -782 -1391 -592 -1357
rect -782 -1487 -588 -1453
rect -3375 -2753 -3341 -2563
rect -3279 -2753 -3245 -2563
rect -3183 -2753 -3149 -2563
rect -3087 -2753 -3053 -2563
rect -2991 -2753 -2957 -2563
rect -2895 -2753 -2861 -2563
rect -2799 -2753 -2765 -2563
rect -2508 -2491 -2318 -2457
rect -2508 -2587 -2314 -2553
rect -2508 -2683 -2318 -2649
rect -2508 -2779 -2314 -2745
rect -1649 -2753 -1615 -2563
rect -1553 -2753 -1519 -2563
rect -1457 -2753 -1423 -2563
rect -1361 -2753 -1327 -2563
rect -1265 -2753 -1231 -2563
rect -1169 -2753 -1135 -2563
rect -1073 -2753 -1039 -2563
rect -782 -2491 -592 -2457
rect -782 -2587 -588 -2553
rect -782 -2683 -592 -2649
rect -782 -2779 -588 -2745
rect -3375 -4725 -3341 -4535
rect -3279 -4725 -3245 -4535
rect -3183 -4725 -3149 -4535
rect -3087 -4725 -3053 -4535
rect -2991 -4725 -2957 -4535
rect -2895 -4725 -2861 -4535
rect -2799 -4725 -2765 -4535
rect -2508 -4463 -2318 -4429
rect -2508 -4559 -2314 -4525
rect -2508 -4655 -2318 -4621
rect -2508 -4751 -2314 -4717
rect -1649 -4725 -1615 -4535
rect -1553 -4725 -1519 -4535
rect -1457 -4725 -1423 -4535
rect -1361 -4725 -1327 -4535
rect -1265 -4725 -1231 -4535
rect -1169 -4725 -1135 -4535
rect -1073 -4725 -1039 -4535
rect -782 -4463 -592 -4429
rect -782 -4559 -588 -4525
rect -782 -4655 -592 -4621
rect -782 -4751 -588 -4717
rect -3375 -6017 -3341 -5827
rect -3279 -6017 -3245 -5827
rect -3183 -6017 -3149 -5827
rect -3087 -6017 -3053 -5827
rect -2991 -6017 -2957 -5827
rect -2895 -6017 -2861 -5827
rect -2799 -6017 -2765 -5827
rect -2508 -5755 -2318 -5721
rect -2508 -5851 -2314 -5817
rect -2508 -5947 -2318 -5913
rect -2508 -6043 -2314 -6009
rect -1649 -6017 -1615 -5827
rect -1553 -6017 -1519 -5827
rect -1457 -6017 -1423 -5827
rect -1361 -6017 -1327 -5827
rect -1265 -6017 -1231 -5827
rect -1169 -6017 -1135 -5827
rect -1073 -6017 -1039 -5827
rect -782 -5755 -592 -5721
rect -782 -5851 -588 -5817
rect -782 -5947 -592 -5913
rect -782 -6043 -588 -6009
<< psubdiff >>
rect -3177 3160 -2777 3184
rect -3177 3086 -3150 3160
rect -2815 3086 -2777 3160
rect -3177 3067 -2777 3086
rect -1336 3160 -936 3184
rect -1336 3086 -1309 3160
rect -974 3086 -936 3160
rect -1336 3067 -936 3086
rect 505 3160 905 3184
rect 505 3086 532 3160
rect 867 3086 905 3160
rect 505 3067 905 3086
rect 2346 3160 2746 3184
rect 2346 3086 2373 3160
rect 2708 3086 2746 3160
rect 2346 3067 2746 3086
rect -3153 1388 -2753 1412
rect -3153 1314 -3126 1388
rect -2791 1314 -2753 1388
rect -3153 1295 -2753 1314
rect -1427 1388 -1027 1412
rect -1427 1314 -1400 1388
rect -1065 1314 -1027 1388
rect -1427 1295 -1027 1314
rect -3153 96 -2753 120
rect -3153 22 -3126 96
rect -2791 22 -2753 96
rect -3153 3 -2753 22
rect -1427 96 -1027 120
rect -1427 22 -1400 96
rect -1065 22 -1027 96
rect -1427 3 -1027 22
rect -3153 -1877 -2753 -1853
rect -3153 -1951 -3126 -1877
rect -2791 -1951 -2753 -1877
rect -3153 -1970 -2753 -1951
rect -1427 -1877 -1027 -1853
rect -1427 -1951 -1400 -1877
rect -1065 -1951 -1027 -1877
rect -1427 -1970 -1027 -1951
rect -3153 -3169 -2753 -3145
rect -3153 -3243 -3126 -3169
rect -2791 -3243 -2753 -3169
rect -3153 -3262 -2753 -3243
rect -1427 -3169 -1027 -3145
rect -1427 -3243 -1400 -3169
rect -1065 -3243 -1027 -3169
rect -1427 -3262 -1027 -3243
rect -3153 -5141 -2753 -5117
rect -3153 -5215 -3126 -5141
rect -2791 -5215 -2753 -5141
rect -3153 -5234 -2753 -5215
rect -1427 -5141 -1027 -5117
rect -1427 -5215 -1400 -5141
rect -1065 -5215 -1027 -5141
rect -1427 -5234 -1027 -5215
rect -3153 -6433 -2753 -6409
rect -3153 -6507 -3126 -6433
rect -2791 -6507 -2753 -6433
rect -3153 -6526 -2753 -6507
rect -1427 -6433 -1027 -6409
rect -1427 -6507 -1400 -6433
rect -1065 -6507 -1027 -6433
rect -1427 -6526 -1027 -6507
<< nsubdiff >>
rect -3407 3921 -2790 3982
rect -3407 3874 -3197 3921
rect -2957 3874 -2790 3921
rect -1566 3921 -949 3982
rect -3407 3832 -2790 3874
rect -1566 3874 -1356 3921
rect -1116 3874 -949 3921
rect 275 3921 892 3982
rect -1566 3832 -949 3874
rect 275 3874 485 3921
rect 725 3874 892 3921
rect 2116 3921 2733 3982
rect 275 3832 892 3874
rect 2116 3874 2326 3921
rect 2566 3874 2733 3921
rect 2116 3832 2733 3874
rect -3383 2149 -2766 2210
rect -3383 2102 -3173 2149
rect -2933 2102 -2766 2149
rect -1657 2149 -1040 2210
rect -3383 2060 -2766 2102
rect -1657 2102 -1447 2149
rect -1207 2102 -1040 2149
rect -1657 2060 -1040 2102
rect -3383 857 -2766 918
rect -3383 810 -3173 857
rect -2933 810 -2766 857
rect -1657 857 -1040 918
rect -3383 768 -2766 810
rect -1657 810 -1447 857
rect -1207 810 -1040 857
rect -1657 768 -1040 810
rect -3383 -1116 -2766 -1055
rect -3383 -1163 -3173 -1116
rect -2933 -1163 -2766 -1116
rect -1657 -1116 -1040 -1055
rect -3383 -1205 -2766 -1163
rect -1657 -1163 -1447 -1116
rect -1207 -1163 -1040 -1116
rect -1657 -1205 -1040 -1163
rect -3383 -2408 -2766 -2347
rect -3383 -2455 -3173 -2408
rect -2933 -2455 -2766 -2408
rect -1657 -2408 -1040 -2347
rect -3383 -2497 -2766 -2455
rect -1657 -2455 -1447 -2408
rect -1207 -2455 -1040 -2408
rect -1657 -2497 -1040 -2455
rect -3383 -4380 -2766 -4319
rect -3383 -4427 -3173 -4380
rect -2933 -4427 -2766 -4380
rect -1657 -4380 -1040 -4319
rect -3383 -4469 -2766 -4427
rect -1657 -4427 -1447 -4380
rect -1207 -4427 -1040 -4380
rect -1657 -4469 -1040 -4427
rect -3383 -5672 -2766 -5611
rect -3383 -5719 -3173 -5672
rect -2933 -5719 -2766 -5672
rect -1657 -5672 -1040 -5611
rect -3383 -5761 -2766 -5719
rect -1657 -5719 -1447 -5672
rect -1207 -5719 -1040 -5672
rect -1657 -5761 -1040 -5719
<< psubdiffcont >>
rect -3150 3086 -2815 3160
rect -1309 3086 -974 3160
rect 532 3086 867 3160
rect 2373 3086 2708 3160
rect -3126 1314 -2791 1388
rect -1400 1314 -1065 1388
rect -3126 22 -2791 96
rect -1400 22 -1065 96
rect -3126 -1951 -2791 -1877
rect -1400 -1951 -1065 -1877
rect -3126 -3243 -2791 -3169
rect -1400 -3243 -1065 -3169
rect -3126 -5215 -2791 -5141
rect -1400 -5215 -1065 -5141
rect -3126 -6507 -2791 -6433
rect -1400 -6507 -1065 -6433
<< nsubdiffcont >>
rect -3197 3874 -2957 3921
rect -1356 3874 -1116 3921
rect 485 3874 725 3921
rect 2326 3874 2566 3921
rect -3173 2102 -2933 2149
rect -1447 2102 -1207 2149
rect -3173 810 -2933 857
rect -1447 810 -1207 857
rect -3173 -1163 -2933 -1116
rect -1447 -1163 -1207 -1116
rect -3173 -2455 -2933 -2408
rect -1447 -2455 -1207 -2408
rect -3173 -4427 -2933 -4380
rect -1447 -4427 -1207 -4380
rect -3173 -5719 -2933 -5672
rect -1447 -5719 -1207 -5672
<< poly >>
rect -2641 3824 -2575 3840
rect -3349 3778 -3319 3809
rect -3253 3778 -3223 3809
rect -3157 3778 -3127 3809
rect -3061 3778 -3031 3809
rect -2965 3778 -2935 3809
rect -2869 3778 -2839 3809
rect -2641 3598 -2625 3824
rect -2591 3822 -2575 3824
rect -800 3824 -734 3840
rect -2591 3792 -2544 3822
rect -2330 3792 -2304 3822
rect -2591 3726 -2575 3792
rect -1508 3778 -1478 3809
rect -1412 3778 -1382 3809
rect -1316 3778 -1286 3809
rect -1220 3778 -1190 3809
rect -1124 3778 -1094 3809
rect -1028 3778 -998 3809
rect -2591 3696 -2544 3726
rect -2330 3696 -2304 3726
rect -2591 3630 -2575 3696
rect -2591 3600 -2544 3630
rect -2330 3600 -2304 3630
rect -2591 3598 -2575 3600
rect -2641 3582 -2575 3598
rect -3349 3538 -3319 3564
rect -3253 3538 -3223 3564
rect -3157 3538 -3127 3564
rect -3350 3517 -3127 3538
rect -3350 3482 -3333 3517
rect -3299 3508 -3127 3517
rect -3061 3538 -3031 3564
rect -2965 3538 -2935 3564
rect -2869 3538 -2839 3564
rect -800 3598 -784 3824
rect -750 3822 -734 3824
rect 1041 3824 1107 3840
rect -750 3792 -703 3822
rect -489 3792 -463 3822
rect -750 3726 -734 3792
rect 333 3778 363 3809
rect 429 3778 459 3809
rect 525 3778 555 3809
rect 621 3778 651 3809
rect 717 3778 747 3809
rect 813 3778 843 3809
rect -750 3696 -703 3726
rect -489 3696 -463 3726
rect -750 3630 -734 3696
rect -750 3600 -703 3630
rect -489 3600 -463 3630
rect -750 3598 -734 3600
rect -800 3582 -734 3598
rect -1508 3538 -1478 3564
rect -1412 3538 -1382 3564
rect -1316 3538 -1286 3564
rect -3061 3517 -2839 3538
rect -3299 3482 -3283 3508
rect -3350 3471 -3283 3482
rect -3061 3482 -3044 3517
rect -3010 3508 -2839 3517
rect -1509 3517 -1286 3538
rect -3010 3482 -2994 3508
rect -3061 3471 -2994 3482
rect -1509 3482 -1492 3517
rect -1458 3508 -1286 3517
rect -1220 3538 -1190 3564
rect -1124 3538 -1094 3564
rect -1028 3538 -998 3564
rect 1041 3598 1057 3824
rect 1091 3822 1107 3824
rect 2882 3824 2948 3840
rect 1091 3792 1138 3822
rect 1352 3792 1378 3822
rect 1091 3726 1107 3792
rect 2174 3778 2204 3809
rect 2270 3778 2300 3809
rect 2366 3778 2396 3809
rect 2462 3778 2492 3809
rect 2558 3778 2588 3809
rect 2654 3778 2684 3809
rect 1091 3696 1138 3726
rect 1352 3696 1378 3726
rect 1091 3630 1107 3696
rect 1091 3600 1138 3630
rect 1352 3600 1378 3630
rect 1091 3598 1107 3600
rect 1041 3582 1107 3598
rect 333 3538 363 3564
rect 429 3538 459 3564
rect 525 3538 555 3564
rect -1220 3517 -998 3538
rect -1458 3482 -1442 3508
rect -1509 3471 -1442 3482
rect -1220 3482 -1203 3517
rect -1169 3508 -998 3517
rect 332 3517 555 3538
rect -1169 3482 -1153 3508
rect -1220 3471 -1153 3482
rect 332 3482 349 3517
rect 383 3508 555 3517
rect 621 3538 651 3564
rect 717 3538 747 3564
rect 813 3538 843 3564
rect 2882 3598 2898 3824
rect 2932 3822 2948 3824
rect 2932 3792 2979 3822
rect 3193 3792 3219 3822
rect 2932 3726 2948 3792
rect 2932 3696 2979 3726
rect 3193 3696 3219 3726
rect 2932 3630 2948 3696
rect 2932 3600 2979 3630
rect 3193 3600 3219 3630
rect 2932 3598 2948 3600
rect 2882 3582 2948 3598
rect 2174 3538 2204 3564
rect 2270 3538 2300 3564
rect 2366 3538 2396 3564
rect 621 3517 843 3538
rect 383 3482 399 3508
rect 332 3471 399 3482
rect 621 3482 638 3517
rect 672 3508 843 3517
rect 2173 3517 2396 3538
rect 672 3482 688 3508
rect 621 3471 688 3482
rect 2173 3482 2190 3517
rect 2224 3508 2396 3517
rect 2462 3538 2492 3564
rect 2558 3538 2588 3564
rect 2654 3538 2684 3564
rect 2462 3517 2684 3538
rect 2224 3482 2240 3508
rect 2173 3471 2240 3482
rect 2462 3482 2479 3517
rect 2513 3508 2684 3517
rect 2513 3482 2529 3508
rect 2462 3471 2529 3482
rect -3350 3276 -3307 3471
rect -3265 3393 -3199 3409
rect -3265 3358 -3249 3393
rect -3215 3372 -3199 3393
rect -2641 3378 -2574 3394
rect -3215 3358 -3177 3372
rect -3265 3342 -3177 3358
rect -2777 3342 -2751 3372
rect -2641 3344 -2625 3378
rect -2591 3376 -2574 3378
rect -2591 3346 -2544 3376
rect -2344 3346 -2318 3376
rect -2591 3344 -2574 3346
rect -2641 3328 -2574 3344
rect -1509 3276 -1466 3471
rect -1424 3393 -1358 3409
rect -1424 3358 -1408 3393
rect -1374 3372 -1358 3393
rect -800 3378 -733 3394
rect -1374 3358 -1336 3372
rect -1424 3342 -1336 3358
rect -936 3342 -910 3372
rect -800 3344 -784 3378
rect -750 3376 -733 3378
rect -750 3346 -703 3376
rect -503 3346 -477 3376
rect -750 3344 -733 3346
rect -800 3328 -733 3344
rect 332 3276 375 3471
rect 417 3393 483 3409
rect 417 3358 433 3393
rect 467 3372 483 3393
rect 1041 3378 1108 3394
rect 467 3358 505 3372
rect 417 3342 505 3358
rect 905 3342 931 3372
rect 1041 3344 1057 3378
rect 1091 3376 1108 3378
rect 1091 3346 1138 3376
rect 1338 3346 1364 3376
rect 1091 3344 1108 3346
rect 1041 3328 1108 3344
rect 2173 3276 2216 3471
rect 2258 3393 2324 3409
rect 2258 3358 2274 3393
rect 2308 3372 2324 3393
rect 2882 3378 2949 3394
rect 2308 3358 2346 3372
rect 2258 3342 2346 3358
rect 2746 3342 2772 3372
rect 2882 3344 2898 3378
rect 2932 3376 2949 3378
rect 2932 3346 2979 3376
rect 3179 3346 3205 3376
rect 2932 3344 2949 3346
rect 2882 3328 2949 3344
rect -3350 3260 -3177 3276
rect -3350 3225 -3249 3260
rect -3215 3246 -3177 3260
rect -2777 3246 -2751 3276
rect -1509 3260 -1336 3276
rect -3215 3225 -3199 3246
rect -3350 3209 -3199 3225
rect -1509 3225 -1408 3260
rect -1374 3246 -1336 3260
rect -936 3246 -910 3276
rect 332 3260 505 3276
rect -1374 3225 -1358 3246
rect -1509 3209 -1358 3225
rect 332 3225 433 3260
rect 467 3246 505 3260
rect 905 3246 931 3276
rect 2173 3260 2346 3276
rect 467 3225 483 3246
rect 332 3209 483 3225
rect 2173 3225 2274 3260
rect 2308 3246 2346 3260
rect 2746 3246 2772 3276
rect 2308 3225 2324 3246
rect 2173 3209 2324 3225
rect -2617 2052 -2551 2068
rect -3325 2006 -3295 2037
rect -3229 2006 -3199 2037
rect -3133 2006 -3103 2037
rect -3037 2006 -3007 2037
rect -2941 2006 -2911 2037
rect -2845 2006 -2815 2037
rect -2617 1826 -2601 2052
rect -2567 2050 -2551 2052
rect -891 2052 -825 2068
rect -2567 2020 -2520 2050
rect -2306 2020 -2280 2050
rect -2567 1954 -2551 2020
rect -1599 2006 -1569 2037
rect -1503 2006 -1473 2037
rect -1407 2006 -1377 2037
rect -1311 2006 -1281 2037
rect -1215 2006 -1185 2037
rect -1119 2006 -1089 2037
rect -2567 1924 -2520 1954
rect -2306 1924 -2280 1954
rect -2567 1858 -2551 1924
rect -2567 1828 -2520 1858
rect -2306 1828 -2280 1858
rect -2567 1826 -2551 1828
rect -2617 1810 -2551 1826
rect -3325 1766 -3295 1792
rect -3229 1766 -3199 1792
rect -3133 1766 -3103 1792
rect -3326 1745 -3103 1766
rect -3326 1710 -3309 1745
rect -3275 1736 -3103 1745
rect -3037 1766 -3007 1792
rect -2941 1766 -2911 1792
rect -2845 1766 -2815 1792
rect -891 1826 -875 2052
rect -841 2050 -825 2052
rect -841 2020 -794 2050
rect -580 2020 -554 2050
rect -841 1954 -825 2020
rect -841 1924 -794 1954
rect -580 1924 -554 1954
rect -841 1858 -825 1924
rect -841 1828 -794 1858
rect -580 1828 -554 1858
rect -841 1826 -825 1828
rect -891 1810 -825 1826
rect -1599 1766 -1569 1792
rect -1503 1766 -1473 1792
rect -1407 1766 -1377 1792
rect -3037 1745 -2815 1766
rect -3275 1710 -3259 1736
rect -3326 1699 -3259 1710
rect -3037 1710 -3020 1745
rect -2986 1736 -2815 1745
rect -1600 1745 -1377 1766
rect -2986 1710 -2970 1736
rect -3037 1699 -2970 1710
rect -1600 1710 -1583 1745
rect -1549 1736 -1377 1745
rect -1311 1766 -1281 1792
rect -1215 1766 -1185 1792
rect -1119 1766 -1089 1792
rect -1311 1745 -1089 1766
rect -1549 1710 -1533 1736
rect -1600 1699 -1533 1710
rect -1311 1710 -1294 1745
rect -1260 1736 -1089 1745
rect -1260 1710 -1244 1736
rect -1311 1699 -1244 1710
rect -3326 1504 -3283 1699
rect -3241 1621 -3175 1637
rect -3241 1586 -3225 1621
rect -3191 1600 -3175 1621
rect -2617 1606 -2550 1622
rect -3191 1586 -3153 1600
rect -3241 1570 -3153 1586
rect -2753 1570 -2727 1600
rect -2617 1572 -2601 1606
rect -2567 1604 -2550 1606
rect -2567 1574 -2520 1604
rect -2320 1574 -2294 1604
rect -2567 1572 -2550 1574
rect -2617 1556 -2550 1572
rect -1600 1504 -1557 1699
rect -1515 1621 -1449 1637
rect -1515 1586 -1499 1621
rect -1465 1600 -1449 1621
rect -891 1606 -824 1622
rect -1465 1586 -1427 1600
rect -1515 1570 -1427 1586
rect -1027 1570 -1001 1600
rect -891 1572 -875 1606
rect -841 1604 -824 1606
rect -841 1574 -794 1604
rect -594 1574 -568 1604
rect -841 1572 -824 1574
rect -891 1556 -824 1572
rect -3326 1488 -3153 1504
rect -3326 1453 -3225 1488
rect -3191 1474 -3153 1488
rect -2753 1474 -2727 1504
rect -1600 1488 -1427 1504
rect -3191 1453 -3175 1474
rect -3326 1437 -3175 1453
rect -1600 1453 -1499 1488
rect -1465 1474 -1427 1488
rect -1027 1474 -1001 1504
rect -1465 1453 -1449 1474
rect -1600 1437 -1449 1453
rect -2617 760 -2551 776
rect -3325 714 -3295 745
rect -3229 714 -3199 745
rect -3133 714 -3103 745
rect -3037 714 -3007 745
rect -2941 714 -2911 745
rect -2845 714 -2815 745
rect -2617 534 -2601 760
rect -2567 758 -2551 760
rect -891 760 -825 776
rect -2567 728 -2520 758
rect -2306 728 -2280 758
rect -2567 662 -2551 728
rect -1599 714 -1569 745
rect -1503 714 -1473 745
rect -1407 714 -1377 745
rect -1311 714 -1281 745
rect -1215 714 -1185 745
rect -1119 714 -1089 745
rect -2567 632 -2520 662
rect -2306 632 -2280 662
rect -2567 566 -2551 632
rect -2567 536 -2520 566
rect -2306 536 -2280 566
rect -2567 534 -2551 536
rect -2617 518 -2551 534
rect -3325 474 -3295 500
rect -3229 474 -3199 500
rect -3133 474 -3103 500
rect -3326 453 -3103 474
rect -3326 418 -3309 453
rect -3275 444 -3103 453
rect -3037 474 -3007 500
rect -2941 474 -2911 500
rect -2845 474 -2815 500
rect -891 534 -875 760
rect -841 758 -825 760
rect -841 728 -794 758
rect -580 728 -554 758
rect -841 662 -825 728
rect -841 632 -794 662
rect -580 632 -554 662
rect -841 566 -825 632
rect -841 536 -794 566
rect -580 536 -554 566
rect -841 534 -825 536
rect -891 518 -825 534
rect -1599 474 -1569 500
rect -1503 474 -1473 500
rect -1407 474 -1377 500
rect -3037 453 -2815 474
rect -3275 418 -3259 444
rect -3326 407 -3259 418
rect -3037 418 -3020 453
rect -2986 444 -2815 453
rect -1600 453 -1377 474
rect -2986 418 -2970 444
rect -3037 407 -2970 418
rect -1600 418 -1583 453
rect -1549 444 -1377 453
rect -1311 474 -1281 500
rect -1215 474 -1185 500
rect -1119 474 -1089 500
rect -1311 453 -1089 474
rect -1549 418 -1533 444
rect -1600 407 -1533 418
rect -1311 418 -1294 453
rect -1260 444 -1089 453
rect -1260 418 -1244 444
rect -1311 407 -1244 418
rect -3326 212 -3283 407
rect -3241 329 -3175 345
rect -3241 294 -3225 329
rect -3191 308 -3175 329
rect -2617 314 -2550 330
rect -3191 294 -3153 308
rect -3241 278 -3153 294
rect -2753 278 -2727 308
rect -2617 280 -2601 314
rect -2567 312 -2550 314
rect -2567 282 -2520 312
rect -2320 282 -2294 312
rect -2567 280 -2550 282
rect -2617 264 -2550 280
rect -1600 212 -1557 407
rect -1515 329 -1449 345
rect -1515 294 -1499 329
rect -1465 308 -1449 329
rect -891 314 -824 330
rect -1465 294 -1427 308
rect -1515 278 -1427 294
rect -1027 278 -1001 308
rect -891 280 -875 314
rect -841 312 -824 314
rect -841 282 -794 312
rect -594 282 -568 312
rect -841 280 -824 282
rect -891 264 -824 280
rect -3326 196 -3153 212
rect -3326 161 -3225 196
rect -3191 182 -3153 196
rect -2753 182 -2727 212
rect -1600 196 -1427 212
rect -3191 161 -3175 182
rect -3326 145 -3175 161
rect -1600 161 -1499 196
rect -1465 182 -1427 196
rect -1027 182 -1001 212
rect -1465 161 -1449 182
rect -1600 145 -1449 161
rect -2617 -1213 -2551 -1197
rect -3325 -1259 -3295 -1228
rect -3229 -1259 -3199 -1228
rect -3133 -1259 -3103 -1228
rect -3037 -1259 -3007 -1228
rect -2941 -1259 -2911 -1228
rect -2845 -1259 -2815 -1228
rect -2617 -1439 -2601 -1213
rect -2567 -1215 -2551 -1213
rect -891 -1213 -825 -1197
rect -2567 -1245 -2520 -1215
rect -2306 -1245 -2280 -1215
rect -2567 -1311 -2551 -1245
rect -1599 -1259 -1569 -1228
rect -1503 -1259 -1473 -1228
rect -1407 -1259 -1377 -1228
rect -1311 -1259 -1281 -1228
rect -1215 -1259 -1185 -1228
rect -1119 -1259 -1089 -1228
rect -2567 -1341 -2520 -1311
rect -2306 -1341 -2280 -1311
rect -2567 -1407 -2551 -1341
rect -2567 -1437 -2520 -1407
rect -2306 -1437 -2280 -1407
rect -2567 -1439 -2551 -1437
rect -2617 -1455 -2551 -1439
rect -3325 -1499 -3295 -1473
rect -3229 -1499 -3199 -1473
rect -3133 -1499 -3103 -1473
rect -3326 -1520 -3103 -1499
rect -3326 -1555 -3309 -1520
rect -3275 -1529 -3103 -1520
rect -3037 -1499 -3007 -1473
rect -2941 -1499 -2911 -1473
rect -2845 -1499 -2815 -1473
rect -891 -1439 -875 -1213
rect -841 -1215 -825 -1213
rect -841 -1245 -794 -1215
rect -580 -1245 -554 -1215
rect -841 -1311 -825 -1245
rect -841 -1341 -794 -1311
rect -580 -1341 -554 -1311
rect -841 -1407 -825 -1341
rect -841 -1437 -794 -1407
rect -580 -1437 -554 -1407
rect -841 -1439 -825 -1437
rect -891 -1455 -825 -1439
rect -1599 -1499 -1569 -1473
rect -1503 -1499 -1473 -1473
rect -1407 -1499 -1377 -1473
rect -3037 -1520 -2815 -1499
rect -3275 -1555 -3259 -1529
rect -3326 -1566 -3259 -1555
rect -3037 -1555 -3020 -1520
rect -2986 -1529 -2815 -1520
rect -1600 -1520 -1377 -1499
rect -2986 -1555 -2970 -1529
rect -3037 -1566 -2970 -1555
rect -1600 -1555 -1583 -1520
rect -1549 -1529 -1377 -1520
rect -1311 -1499 -1281 -1473
rect -1215 -1499 -1185 -1473
rect -1119 -1499 -1089 -1473
rect -1311 -1520 -1089 -1499
rect -1549 -1555 -1533 -1529
rect -1600 -1566 -1533 -1555
rect -1311 -1555 -1294 -1520
rect -1260 -1529 -1089 -1520
rect -1260 -1555 -1244 -1529
rect -1311 -1566 -1244 -1555
rect -3326 -1761 -3283 -1566
rect -3241 -1644 -3175 -1628
rect -3241 -1679 -3225 -1644
rect -3191 -1665 -3175 -1644
rect -2617 -1659 -2550 -1643
rect -3191 -1679 -3153 -1665
rect -3241 -1695 -3153 -1679
rect -2753 -1695 -2727 -1665
rect -2617 -1693 -2601 -1659
rect -2567 -1661 -2550 -1659
rect -2567 -1691 -2520 -1661
rect -2320 -1691 -2294 -1661
rect -2567 -1693 -2550 -1691
rect -2617 -1709 -2550 -1693
rect -1600 -1761 -1557 -1566
rect -1515 -1644 -1449 -1628
rect -1515 -1679 -1499 -1644
rect -1465 -1665 -1449 -1644
rect -891 -1659 -824 -1643
rect -1465 -1679 -1427 -1665
rect -1515 -1695 -1427 -1679
rect -1027 -1695 -1001 -1665
rect -891 -1693 -875 -1659
rect -841 -1661 -824 -1659
rect -841 -1691 -794 -1661
rect -594 -1691 -568 -1661
rect -841 -1693 -824 -1691
rect -891 -1709 -824 -1693
rect -3326 -1777 -3153 -1761
rect -3326 -1812 -3225 -1777
rect -3191 -1791 -3153 -1777
rect -2753 -1791 -2727 -1761
rect -1600 -1777 -1427 -1761
rect -3191 -1812 -3175 -1791
rect -3326 -1828 -3175 -1812
rect -1600 -1812 -1499 -1777
rect -1465 -1791 -1427 -1777
rect -1027 -1791 -1001 -1761
rect -1465 -1812 -1449 -1791
rect -1600 -1828 -1449 -1812
rect -2617 -2505 -2551 -2489
rect -3325 -2551 -3295 -2520
rect -3229 -2551 -3199 -2520
rect -3133 -2551 -3103 -2520
rect -3037 -2551 -3007 -2520
rect -2941 -2551 -2911 -2520
rect -2845 -2551 -2815 -2520
rect -2617 -2731 -2601 -2505
rect -2567 -2507 -2551 -2505
rect -891 -2505 -825 -2489
rect -2567 -2537 -2520 -2507
rect -2306 -2537 -2280 -2507
rect -2567 -2603 -2551 -2537
rect -1599 -2551 -1569 -2520
rect -1503 -2551 -1473 -2520
rect -1407 -2551 -1377 -2520
rect -1311 -2551 -1281 -2520
rect -1215 -2551 -1185 -2520
rect -1119 -2551 -1089 -2520
rect -2567 -2633 -2520 -2603
rect -2306 -2633 -2280 -2603
rect -2567 -2699 -2551 -2633
rect -2567 -2729 -2520 -2699
rect -2306 -2729 -2280 -2699
rect -2567 -2731 -2551 -2729
rect -2617 -2747 -2551 -2731
rect -3325 -2791 -3295 -2765
rect -3229 -2791 -3199 -2765
rect -3133 -2791 -3103 -2765
rect -3326 -2812 -3103 -2791
rect -3326 -2847 -3309 -2812
rect -3275 -2821 -3103 -2812
rect -3037 -2791 -3007 -2765
rect -2941 -2791 -2911 -2765
rect -2845 -2791 -2815 -2765
rect -891 -2731 -875 -2505
rect -841 -2507 -825 -2505
rect -841 -2537 -794 -2507
rect -580 -2537 -554 -2507
rect -841 -2603 -825 -2537
rect -841 -2633 -794 -2603
rect -580 -2633 -554 -2603
rect -841 -2699 -825 -2633
rect -841 -2729 -794 -2699
rect -580 -2729 -554 -2699
rect -841 -2731 -825 -2729
rect -891 -2747 -825 -2731
rect -1599 -2791 -1569 -2765
rect -1503 -2791 -1473 -2765
rect -1407 -2791 -1377 -2765
rect -3037 -2812 -2815 -2791
rect -3275 -2847 -3259 -2821
rect -3326 -2858 -3259 -2847
rect -3037 -2847 -3020 -2812
rect -2986 -2821 -2815 -2812
rect -1600 -2812 -1377 -2791
rect -2986 -2847 -2970 -2821
rect -3037 -2858 -2970 -2847
rect -1600 -2847 -1583 -2812
rect -1549 -2821 -1377 -2812
rect -1311 -2791 -1281 -2765
rect -1215 -2791 -1185 -2765
rect -1119 -2791 -1089 -2765
rect -1311 -2812 -1089 -2791
rect -1549 -2847 -1533 -2821
rect -1600 -2858 -1533 -2847
rect -1311 -2847 -1294 -2812
rect -1260 -2821 -1089 -2812
rect -1260 -2847 -1244 -2821
rect -1311 -2858 -1244 -2847
rect -3326 -3053 -3283 -2858
rect -3241 -2936 -3175 -2920
rect -3241 -2971 -3225 -2936
rect -3191 -2957 -3175 -2936
rect -2617 -2951 -2550 -2935
rect -3191 -2971 -3153 -2957
rect -3241 -2987 -3153 -2971
rect -2753 -2987 -2727 -2957
rect -2617 -2985 -2601 -2951
rect -2567 -2953 -2550 -2951
rect -2567 -2983 -2520 -2953
rect -2320 -2983 -2294 -2953
rect -2567 -2985 -2550 -2983
rect -2617 -3001 -2550 -2985
rect -1600 -3053 -1557 -2858
rect -1515 -2936 -1449 -2920
rect -1515 -2971 -1499 -2936
rect -1465 -2957 -1449 -2936
rect -891 -2951 -824 -2935
rect -1465 -2971 -1427 -2957
rect -1515 -2987 -1427 -2971
rect -1027 -2987 -1001 -2957
rect -891 -2985 -875 -2951
rect -841 -2953 -824 -2951
rect -841 -2983 -794 -2953
rect -594 -2983 -568 -2953
rect -841 -2985 -824 -2983
rect -891 -3001 -824 -2985
rect -3326 -3069 -3153 -3053
rect -3326 -3104 -3225 -3069
rect -3191 -3083 -3153 -3069
rect -2753 -3083 -2727 -3053
rect -1600 -3069 -1427 -3053
rect -3191 -3104 -3175 -3083
rect -3326 -3120 -3175 -3104
rect -1600 -3104 -1499 -3069
rect -1465 -3083 -1427 -3069
rect -1027 -3083 -1001 -3053
rect -1465 -3104 -1449 -3083
rect -1600 -3120 -1449 -3104
rect -2617 -4477 -2551 -4461
rect -3325 -4523 -3295 -4492
rect -3229 -4523 -3199 -4492
rect -3133 -4523 -3103 -4492
rect -3037 -4523 -3007 -4492
rect -2941 -4523 -2911 -4492
rect -2845 -4523 -2815 -4492
rect -2617 -4703 -2601 -4477
rect -2567 -4479 -2551 -4477
rect -891 -4477 -825 -4461
rect -2567 -4509 -2520 -4479
rect -2306 -4509 -2280 -4479
rect -2567 -4575 -2551 -4509
rect -1599 -4523 -1569 -4492
rect -1503 -4523 -1473 -4492
rect -1407 -4523 -1377 -4492
rect -1311 -4523 -1281 -4492
rect -1215 -4523 -1185 -4492
rect -1119 -4523 -1089 -4492
rect -2567 -4605 -2520 -4575
rect -2306 -4605 -2280 -4575
rect -2567 -4671 -2551 -4605
rect -2567 -4701 -2520 -4671
rect -2306 -4701 -2280 -4671
rect -2567 -4703 -2551 -4701
rect -2617 -4719 -2551 -4703
rect -3325 -4763 -3295 -4737
rect -3229 -4763 -3199 -4737
rect -3133 -4763 -3103 -4737
rect -3326 -4784 -3103 -4763
rect -3326 -4819 -3309 -4784
rect -3275 -4793 -3103 -4784
rect -3037 -4763 -3007 -4737
rect -2941 -4763 -2911 -4737
rect -2845 -4763 -2815 -4737
rect -891 -4703 -875 -4477
rect -841 -4479 -825 -4477
rect -841 -4509 -794 -4479
rect -580 -4509 -554 -4479
rect -841 -4575 -825 -4509
rect -841 -4605 -794 -4575
rect -580 -4605 -554 -4575
rect -841 -4671 -825 -4605
rect -841 -4701 -794 -4671
rect -580 -4701 -554 -4671
rect -841 -4703 -825 -4701
rect -891 -4719 -825 -4703
rect -1599 -4763 -1569 -4737
rect -1503 -4763 -1473 -4737
rect -1407 -4763 -1377 -4737
rect -3037 -4784 -2815 -4763
rect -3275 -4819 -3259 -4793
rect -3326 -4830 -3259 -4819
rect -3037 -4819 -3020 -4784
rect -2986 -4793 -2815 -4784
rect -1600 -4784 -1377 -4763
rect -2986 -4819 -2970 -4793
rect -3037 -4830 -2970 -4819
rect -1600 -4819 -1583 -4784
rect -1549 -4793 -1377 -4784
rect -1311 -4763 -1281 -4737
rect -1215 -4763 -1185 -4737
rect -1119 -4763 -1089 -4737
rect -1311 -4784 -1089 -4763
rect -1549 -4819 -1533 -4793
rect -1600 -4830 -1533 -4819
rect -1311 -4819 -1294 -4784
rect -1260 -4793 -1089 -4784
rect -1260 -4819 -1244 -4793
rect -1311 -4830 -1244 -4819
rect -3326 -5025 -3283 -4830
rect -3241 -4908 -3175 -4892
rect -3241 -4943 -3225 -4908
rect -3191 -4929 -3175 -4908
rect -2617 -4923 -2550 -4907
rect -3191 -4943 -3153 -4929
rect -3241 -4959 -3153 -4943
rect -2753 -4959 -2727 -4929
rect -2617 -4957 -2601 -4923
rect -2567 -4925 -2550 -4923
rect -2567 -4955 -2520 -4925
rect -2320 -4955 -2294 -4925
rect -2567 -4957 -2550 -4955
rect -2617 -4973 -2550 -4957
rect -1600 -5025 -1557 -4830
rect -1515 -4908 -1449 -4892
rect -1515 -4943 -1499 -4908
rect -1465 -4929 -1449 -4908
rect -891 -4923 -824 -4907
rect -1465 -4943 -1427 -4929
rect -1515 -4959 -1427 -4943
rect -1027 -4959 -1001 -4929
rect -891 -4957 -875 -4923
rect -841 -4925 -824 -4923
rect -841 -4955 -794 -4925
rect -594 -4955 -568 -4925
rect -841 -4957 -824 -4955
rect -891 -4973 -824 -4957
rect -3326 -5041 -3153 -5025
rect -3326 -5076 -3225 -5041
rect -3191 -5055 -3153 -5041
rect -2753 -5055 -2727 -5025
rect -1600 -5041 -1427 -5025
rect -3191 -5076 -3175 -5055
rect -3326 -5092 -3175 -5076
rect -1600 -5076 -1499 -5041
rect -1465 -5055 -1427 -5041
rect -1027 -5055 -1001 -5025
rect -1465 -5076 -1449 -5055
rect -1600 -5092 -1449 -5076
rect -2617 -5769 -2551 -5753
rect -3325 -5815 -3295 -5784
rect -3229 -5815 -3199 -5784
rect -3133 -5815 -3103 -5784
rect -3037 -5815 -3007 -5784
rect -2941 -5815 -2911 -5784
rect -2845 -5815 -2815 -5784
rect -2617 -5995 -2601 -5769
rect -2567 -5771 -2551 -5769
rect -891 -5769 -825 -5753
rect -2567 -5801 -2520 -5771
rect -2306 -5801 -2280 -5771
rect -2567 -5867 -2551 -5801
rect -1599 -5815 -1569 -5784
rect -1503 -5815 -1473 -5784
rect -1407 -5815 -1377 -5784
rect -1311 -5815 -1281 -5784
rect -1215 -5815 -1185 -5784
rect -1119 -5815 -1089 -5784
rect -2567 -5897 -2520 -5867
rect -2306 -5897 -2280 -5867
rect -2567 -5963 -2551 -5897
rect -2567 -5993 -2520 -5963
rect -2306 -5993 -2280 -5963
rect -2567 -5995 -2551 -5993
rect -2617 -6011 -2551 -5995
rect -3325 -6055 -3295 -6029
rect -3229 -6055 -3199 -6029
rect -3133 -6055 -3103 -6029
rect -3326 -6076 -3103 -6055
rect -3326 -6111 -3309 -6076
rect -3275 -6085 -3103 -6076
rect -3037 -6055 -3007 -6029
rect -2941 -6055 -2911 -6029
rect -2845 -6055 -2815 -6029
rect -891 -5995 -875 -5769
rect -841 -5771 -825 -5769
rect -841 -5801 -794 -5771
rect -580 -5801 -554 -5771
rect -841 -5867 -825 -5801
rect -841 -5897 -794 -5867
rect -580 -5897 -554 -5867
rect -841 -5963 -825 -5897
rect -841 -5993 -794 -5963
rect -580 -5993 -554 -5963
rect -841 -5995 -825 -5993
rect -891 -6011 -825 -5995
rect -1599 -6055 -1569 -6029
rect -1503 -6055 -1473 -6029
rect -1407 -6055 -1377 -6029
rect -3037 -6076 -2815 -6055
rect -3275 -6111 -3259 -6085
rect -3326 -6122 -3259 -6111
rect -3037 -6111 -3020 -6076
rect -2986 -6085 -2815 -6076
rect -1600 -6076 -1377 -6055
rect -2986 -6111 -2970 -6085
rect -3037 -6122 -2970 -6111
rect -1600 -6111 -1583 -6076
rect -1549 -6085 -1377 -6076
rect -1311 -6055 -1281 -6029
rect -1215 -6055 -1185 -6029
rect -1119 -6055 -1089 -6029
rect -1311 -6076 -1089 -6055
rect -1549 -6111 -1533 -6085
rect -1600 -6122 -1533 -6111
rect -1311 -6111 -1294 -6076
rect -1260 -6085 -1089 -6076
rect -1260 -6111 -1244 -6085
rect -1311 -6122 -1244 -6111
rect -3326 -6317 -3283 -6122
rect -3241 -6200 -3175 -6184
rect -3241 -6235 -3225 -6200
rect -3191 -6221 -3175 -6200
rect -2617 -6215 -2550 -6199
rect -3191 -6235 -3153 -6221
rect -3241 -6251 -3153 -6235
rect -2753 -6251 -2727 -6221
rect -2617 -6249 -2601 -6215
rect -2567 -6217 -2550 -6215
rect -2567 -6247 -2520 -6217
rect -2320 -6247 -2294 -6217
rect -2567 -6249 -2550 -6247
rect -2617 -6265 -2550 -6249
rect -1600 -6317 -1557 -6122
rect -1515 -6200 -1449 -6184
rect -1515 -6235 -1499 -6200
rect -1465 -6221 -1449 -6200
rect -891 -6215 -824 -6199
rect -1465 -6235 -1427 -6221
rect -1515 -6251 -1427 -6235
rect -1027 -6251 -1001 -6221
rect -891 -6249 -875 -6215
rect -841 -6217 -824 -6215
rect -841 -6247 -794 -6217
rect -594 -6247 -568 -6217
rect -841 -6249 -824 -6247
rect -891 -6265 -824 -6249
rect -3326 -6333 -3153 -6317
rect -3326 -6368 -3225 -6333
rect -3191 -6347 -3153 -6333
rect -2753 -6347 -2727 -6317
rect -1600 -6333 -1427 -6317
rect -3191 -6368 -3175 -6347
rect -3326 -6384 -3175 -6368
rect -1600 -6368 -1499 -6333
rect -1465 -6347 -1427 -6333
rect -1027 -6347 -1001 -6317
rect -1465 -6368 -1449 -6347
rect -1600 -6384 -1449 -6368
<< polycont >>
rect -2625 3598 -2591 3824
rect -3333 3482 -3299 3517
rect -784 3598 -750 3824
rect -3044 3482 -3010 3517
rect -1492 3482 -1458 3517
rect 1057 3598 1091 3824
rect -1203 3482 -1169 3517
rect 349 3482 383 3517
rect 2898 3598 2932 3824
rect 638 3482 672 3517
rect 2190 3482 2224 3517
rect 2479 3482 2513 3517
rect -3249 3358 -3215 3393
rect -2625 3344 -2591 3378
rect -1408 3358 -1374 3393
rect -784 3344 -750 3378
rect 433 3358 467 3393
rect 1057 3344 1091 3378
rect 2274 3358 2308 3393
rect 2898 3344 2932 3378
rect -3249 3225 -3215 3260
rect -1408 3225 -1374 3260
rect 433 3225 467 3260
rect 2274 3225 2308 3260
rect -2601 1826 -2567 2052
rect -3309 1710 -3275 1745
rect -875 1826 -841 2052
rect -3020 1710 -2986 1745
rect -1583 1710 -1549 1745
rect -1294 1710 -1260 1745
rect -3225 1586 -3191 1621
rect -2601 1572 -2567 1606
rect -1499 1586 -1465 1621
rect -875 1572 -841 1606
rect -3225 1453 -3191 1488
rect -1499 1453 -1465 1488
rect -2601 534 -2567 760
rect -3309 418 -3275 453
rect -875 534 -841 760
rect -3020 418 -2986 453
rect -1583 418 -1549 453
rect -1294 418 -1260 453
rect -3225 294 -3191 329
rect -2601 280 -2567 314
rect -1499 294 -1465 329
rect -875 280 -841 314
rect -3225 161 -3191 196
rect -1499 161 -1465 196
rect -2601 -1439 -2567 -1213
rect -3309 -1555 -3275 -1520
rect -875 -1439 -841 -1213
rect -3020 -1555 -2986 -1520
rect -1583 -1555 -1549 -1520
rect -1294 -1555 -1260 -1520
rect -3225 -1679 -3191 -1644
rect -2601 -1693 -2567 -1659
rect -1499 -1679 -1465 -1644
rect -875 -1693 -841 -1659
rect -3225 -1812 -3191 -1777
rect -1499 -1812 -1465 -1777
rect -2601 -2731 -2567 -2505
rect -3309 -2847 -3275 -2812
rect -875 -2731 -841 -2505
rect -3020 -2847 -2986 -2812
rect -1583 -2847 -1549 -2812
rect -1294 -2847 -1260 -2812
rect -3225 -2971 -3191 -2936
rect -2601 -2985 -2567 -2951
rect -1499 -2971 -1465 -2936
rect -875 -2985 -841 -2951
rect -3225 -3104 -3191 -3069
rect -1499 -3104 -1465 -3069
rect -2601 -4703 -2567 -4477
rect -3309 -4819 -3275 -4784
rect -875 -4703 -841 -4477
rect -3020 -4819 -2986 -4784
rect -1583 -4819 -1549 -4784
rect -1294 -4819 -1260 -4784
rect -3225 -4943 -3191 -4908
rect -2601 -4957 -2567 -4923
rect -1499 -4943 -1465 -4908
rect -875 -4957 -841 -4923
rect -3225 -5076 -3191 -5041
rect -1499 -5076 -1465 -5041
rect -2601 -5995 -2567 -5769
rect -3309 -6111 -3275 -6076
rect -875 -5995 -841 -5769
rect -3020 -6111 -2986 -6076
rect -1583 -6111 -1549 -6076
rect -1294 -6111 -1260 -6076
rect -3225 -6235 -3191 -6200
rect -2601 -6249 -2567 -6215
rect -1499 -6235 -1465 -6200
rect -875 -6249 -841 -6215
rect -3225 -6368 -3191 -6333
rect -1499 -6368 -1465 -6333
<< locali >>
rect -3271 3874 -3197 3921
rect -2957 3874 -2857 3921
rect -1430 3874 -1356 3921
rect -1116 3874 -1016 3921
rect 411 3874 485 3921
rect 725 3874 825 3921
rect 2252 3874 2326 3921
rect 2566 3874 2666 3921
rect -2641 3824 -2591 3841
rect -2548 3838 -2538 3872
rect -2342 3838 -2326 3872
rect -3399 3772 -3365 3782
rect -3399 3560 -3365 3576
rect -3303 3766 -3269 3782
rect -3303 3560 -3269 3570
rect -3207 3772 -3173 3782
rect -3207 3560 -3173 3576
rect -3111 3766 -3077 3782
rect -3111 3560 -3077 3570
rect -3015 3772 -2981 3782
rect -3015 3560 -2981 3576
rect -2919 3766 -2885 3782
rect -2919 3560 -2885 3570
rect -2823 3772 -2789 3782
rect -2823 3560 -2789 3576
rect -2641 3598 -2625 3824
rect -800 3824 -750 3841
rect -707 3838 -697 3872
rect -501 3838 -485 3872
rect -2548 3742 -2532 3776
rect -2338 3742 -2320 3776
rect -1558 3772 -1524 3782
rect -2548 3646 -2538 3680
rect -2342 3646 -2326 3680
rect -3350 3482 -3333 3517
rect -3299 3482 -3283 3517
rect -3061 3511 -3044 3517
rect -3249 3482 -3044 3511
rect -3010 3482 -2994 3517
rect -3350 3276 -3307 3482
rect -3249 3477 -2994 3482
rect -3249 3393 -3215 3477
rect -3181 3388 -3165 3422
rect -2789 3388 -2773 3422
rect -3249 3342 -3215 3358
rect -2641 3378 -2591 3598
rect -2548 3550 -2532 3584
rect -2338 3550 -2320 3584
rect -1558 3560 -1524 3576
rect -1462 3766 -1428 3782
rect -1462 3560 -1428 3570
rect -1366 3772 -1332 3782
rect -1366 3560 -1332 3576
rect -1270 3766 -1236 3782
rect -1270 3560 -1236 3570
rect -1174 3772 -1140 3782
rect -1174 3560 -1140 3576
rect -1078 3766 -1044 3782
rect -1078 3560 -1044 3570
rect -982 3772 -948 3782
rect -982 3560 -948 3576
rect -800 3598 -784 3824
rect 1041 3824 1091 3841
rect 1134 3838 1144 3872
rect 1340 3838 1356 3872
rect -707 3742 -691 3776
rect -497 3742 -479 3776
rect 283 3772 317 3782
rect -707 3646 -697 3680
rect -501 3646 -485 3680
rect -1509 3482 -1492 3517
rect -1458 3482 -1442 3517
rect -1220 3511 -1203 3517
rect -1408 3482 -1203 3511
rect -1169 3482 -1153 3517
rect -2548 3388 -2532 3422
rect -2356 3388 -2340 3422
rect -2641 3344 -2625 3378
rect -2641 3328 -2591 3344
rect -2548 3300 -2532 3334
rect -2356 3300 -2340 3334
rect -1509 3276 -1466 3482
rect -1408 3477 -1153 3482
rect -1408 3393 -1374 3477
rect -1340 3388 -1324 3422
rect -948 3388 -932 3422
rect -1408 3342 -1374 3358
rect -800 3378 -750 3598
rect -707 3550 -691 3584
rect -497 3550 -479 3584
rect 283 3560 317 3576
rect 379 3766 413 3782
rect 379 3560 413 3570
rect 475 3772 509 3782
rect 475 3560 509 3576
rect 571 3766 605 3782
rect 571 3560 605 3570
rect 667 3772 701 3782
rect 667 3560 701 3576
rect 763 3766 797 3782
rect 763 3560 797 3570
rect 859 3772 893 3782
rect 859 3560 893 3576
rect 1041 3598 1057 3824
rect 2882 3824 2932 3841
rect 2975 3838 2985 3872
rect 3181 3838 3197 3872
rect 1134 3742 1150 3776
rect 1344 3742 1362 3776
rect 2124 3772 2158 3782
rect 1134 3646 1144 3680
rect 1340 3646 1356 3680
rect 332 3482 349 3517
rect 383 3482 399 3517
rect 621 3511 638 3517
rect 433 3482 638 3511
rect 672 3482 688 3517
rect -707 3388 -691 3422
rect -515 3388 -499 3422
rect -800 3344 -784 3378
rect -800 3328 -750 3344
rect -707 3300 -691 3334
rect -515 3300 -499 3334
rect 332 3276 375 3482
rect 433 3477 688 3482
rect 433 3393 467 3477
rect 501 3388 517 3422
rect 893 3388 909 3422
rect 433 3342 467 3358
rect 1041 3378 1091 3598
rect 1134 3550 1150 3584
rect 1344 3550 1362 3584
rect 2124 3560 2158 3576
rect 2220 3766 2254 3782
rect 2220 3560 2254 3570
rect 2316 3772 2350 3782
rect 2316 3560 2350 3576
rect 2412 3766 2446 3782
rect 2412 3560 2446 3570
rect 2508 3772 2542 3782
rect 2508 3560 2542 3576
rect 2604 3766 2638 3782
rect 2604 3560 2638 3570
rect 2700 3772 2734 3782
rect 2700 3560 2734 3576
rect 2882 3598 2898 3824
rect 2975 3742 2991 3776
rect 3185 3742 3203 3776
rect 2975 3646 2985 3680
rect 3181 3646 3197 3680
rect 2173 3482 2190 3517
rect 2224 3482 2240 3517
rect 2462 3511 2479 3517
rect 2274 3482 2479 3511
rect 2513 3482 2529 3517
rect 1134 3388 1150 3422
rect 1326 3388 1342 3422
rect 1041 3344 1057 3378
rect 1041 3328 1091 3344
rect 1134 3300 1150 3334
rect 1326 3300 1342 3334
rect 2173 3276 2216 3482
rect 2274 3477 2529 3482
rect 2274 3393 2308 3477
rect 2342 3388 2358 3422
rect 2734 3388 2750 3422
rect 2274 3342 2308 3358
rect 2882 3378 2932 3598
rect 2975 3550 2991 3584
rect 3185 3550 3203 3584
rect 2975 3388 2991 3422
rect 3167 3388 3183 3422
rect 2882 3344 2898 3378
rect 2882 3328 2932 3344
rect 2975 3300 2991 3334
rect 3167 3300 3183 3334
rect -3350 3260 -3215 3276
rect -3350 3225 -3249 3260
rect -1509 3260 -1374 3276
rect -3350 3209 -3215 3225
rect -3181 3196 -3165 3230
rect -2789 3196 -2773 3230
rect -1509 3225 -1408 3260
rect 332 3260 467 3276
rect -1509 3209 -1374 3225
rect -1340 3196 -1324 3230
rect -948 3196 -932 3230
rect 332 3225 433 3260
rect 2173 3260 2308 3276
rect 332 3209 467 3225
rect 501 3196 517 3230
rect 893 3196 909 3230
rect 2173 3225 2274 3260
rect 2173 3209 2308 3225
rect 2342 3196 2358 3230
rect 2734 3196 2750 3230
rect -3177 3086 -3150 3160
rect -2815 3086 -2777 3160
rect -1336 3086 -1309 3160
rect -974 3086 -936 3160
rect 505 3086 532 3160
rect 867 3086 905 3160
rect 2346 3086 2373 3160
rect 2708 3086 2746 3160
rect -3247 2102 -3173 2149
rect -2933 2102 -2833 2149
rect -1521 2102 -1447 2149
rect -1207 2102 -1107 2149
rect -2617 2052 -2567 2069
rect -2524 2066 -2514 2100
rect -2318 2066 -2302 2100
rect -3375 2000 -3341 2010
rect -3375 1788 -3341 1804
rect -3279 1994 -3245 2010
rect -3279 1788 -3245 1798
rect -3183 2000 -3149 2010
rect -3183 1788 -3149 1804
rect -3087 1994 -3053 2010
rect -3087 1788 -3053 1798
rect -2991 2000 -2957 2010
rect -2991 1788 -2957 1804
rect -2895 1994 -2861 2010
rect -2895 1788 -2861 1798
rect -2799 2000 -2765 2010
rect -2799 1788 -2765 1804
rect -2617 1826 -2601 2052
rect -891 2052 -841 2069
rect -798 2066 -788 2100
rect -592 2066 -576 2100
rect -2524 1970 -2508 2004
rect -2314 1970 -2296 2004
rect -1649 2000 -1615 2010
rect -2524 1874 -2514 1908
rect -2318 1874 -2302 1908
rect -3326 1710 -3309 1745
rect -3275 1710 -3259 1745
rect -3037 1739 -3020 1745
rect -3225 1710 -3020 1739
rect -2986 1710 -2970 1745
rect -3326 1504 -3283 1710
rect -3225 1705 -2970 1710
rect -3225 1621 -3191 1705
rect -3157 1616 -3141 1650
rect -2765 1616 -2749 1650
rect -3225 1570 -3191 1586
rect -2617 1606 -2567 1826
rect -2524 1778 -2508 1812
rect -2314 1778 -2296 1812
rect -1649 1788 -1615 1804
rect -1553 1994 -1519 2010
rect -1553 1788 -1519 1798
rect -1457 2000 -1423 2010
rect -1457 1788 -1423 1804
rect -1361 1994 -1327 2010
rect -1361 1788 -1327 1798
rect -1265 2000 -1231 2010
rect -1265 1788 -1231 1804
rect -1169 1994 -1135 2010
rect -1169 1788 -1135 1798
rect -1073 2000 -1039 2010
rect -1073 1788 -1039 1804
rect -891 1826 -875 2052
rect -798 1970 -782 2004
rect -588 1970 -570 2004
rect -798 1874 -788 1908
rect -592 1874 -576 1908
rect -1600 1710 -1583 1745
rect -1549 1710 -1533 1745
rect -1311 1739 -1294 1745
rect -1499 1710 -1294 1739
rect -1260 1710 -1244 1745
rect -2524 1616 -2508 1650
rect -2332 1616 -2316 1650
rect -2617 1572 -2601 1606
rect -2617 1556 -2567 1572
rect -2524 1528 -2508 1562
rect -2332 1528 -2316 1562
rect -1600 1504 -1557 1710
rect -1499 1705 -1244 1710
rect -1499 1621 -1465 1705
rect -1431 1616 -1415 1650
rect -1039 1616 -1023 1650
rect -1499 1570 -1465 1586
rect -891 1606 -841 1826
rect -798 1778 -782 1812
rect -588 1778 -570 1812
rect -798 1616 -782 1650
rect -606 1616 -590 1650
rect -891 1572 -875 1606
rect -891 1556 -841 1572
rect -798 1528 -782 1562
rect -606 1528 -590 1562
rect -3326 1488 -3191 1504
rect -3326 1453 -3225 1488
rect -1600 1488 -1465 1504
rect -3326 1437 -3191 1453
rect -3157 1424 -3141 1458
rect -2765 1424 -2749 1458
rect -1600 1453 -1499 1488
rect -1600 1437 -1465 1453
rect -1431 1424 -1415 1458
rect -1039 1424 -1023 1458
rect -3153 1314 -3126 1388
rect -2791 1314 -2753 1388
rect -1427 1314 -1400 1388
rect -1065 1314 -1027 1388
rect 154 1006 264 1634
rect 154 942 596 1006
rect -3247 810 -3173 857
rect -2933 810 -2833 857
rect -1521 810 -1447 857
rect -1207 810 -1107 857
rect -2617 760 -2567 777
rect -2524 774 -2514 808
rect -2318 774 -2302 808
rect -3375 708 -3341 718
rect -3375 496 -3341 512
rect -3279 702 -3245 718
rect -3279 496 -3245 506
rect -3183 708 -3149 718
rect -3183 496 -3149 512
rect -3087 702 -3053 718
rect -3087 496 -3053 506
rect -2991 708 -2957 718
rect -2991 496 -2957 512
rect -2895 702 -2861 718
rect -2895 496 -2861 506
rect -2799 708 -2765 718
rect -2799 496 -2765 512
rect -2617 534 -2601 760
rect -891 760 -841 777
rect -798 774 -788 808
rect -592 774 -576 808
rect -2524 678 -2508 712
rect -2314 678 -2296 712
rect -1649 708 -1615 718
rect -2524 582 -2514 616
rect -2318 582 -2302 616
rect -3326 418 -3309 453
rect -3275 418 -3259 453
rect -3037 447 -3020 453
rect -3225 418 -3020 447
rect -2986 418 -2970 453
rect -3326 212 -3283 418
rect -3225 413 -2970 418
rect -3225 329 -3191 413
rect -3157 324 -3141 358
rect -2765 324 -2749 358
rect -3225 278 -3191 294
rect -2617 314 -2567 534
rect -2524 486 -2508 520
rect -2314 486 -2296 520
rect -1649 496 -1615 512
rect -1553 702 -1519 718
rect -1553 496 -1519 506
rect -1457 708 -1423 718
rect -1457 496 -1423 512
rect -1361 702 -1327 718
rect -1361 496 -1327 506
rect -1265 708 -1231 718
rect -1265 496 -1231 512
rect -1169 702 -1135 718
rect -1169 496 -1135 506
rect -1073 708 -1039 718
rect -1073 496 -1039 512
rect -891 534 -875 760
rect -798 678 -782 712
rect -588 678 -570 712
rect -798 582 -788 616
rect -592 582 -576 616
rect -1600 418 -1583 453
rect -1549 418 -1533 453
rect -1311 447 -1294 453
rect -1499 418 -1294 447
rect -1260 418 -1244 453
rect -2524 324 -2508 358
rect -2332 324 -2316 358
rect -2617 280 -2601 314
rect -2617 264 -2567 280
rect -2524 236 -2508 270
rect -2332 236 -2316 270
rect -1600 212 -1557 418
rect -1499 413 -1244 418
rect -1499 329 -1465 413
rect -1431 324 -1415 358
rect -1039 324 -1023 358
rect -1499 278 -1465 294
rect -891 314 -841 534
rect -798 486 -782 520
rect -588 486 -570 520
rect -798 324 -782 358
rect -606 324 -590 358
rect -891 280 -875 314
rect -891 264 -841 280
rect -798 236 -782 270
rect -606 236 -590 270
rect -3326 196 -3191 212
rect -3326 161 -3225 196
rect -1600 196 -1465 212
rect -3326 145 -3191 161
rect -3157 132 -3141 166
rect -2765 132 -2749 166
rect -1600 161 -1499 196
rect -1600 145 -1465 161
rect -1431 132 -1415 166
rect -1039 132 -1023 166
rect -3153 22 -3126 96
rect -2791 22 -2753 96
rect -1427 22 -1400 96
rect -1065 22 -1027 96
rect -3247 -1163 -3173 -1116
rect -2933 -1163 -2833 -1116
rect -1521 -1163 -1447 -1116
rect -1207 -1163 -1107 -1116
rect -2617 -1213 -2567 -1196
rect -2524 -1199 -2514 -1165
rect -2318 -1199 -2302 -1165
rect -3375 -1265 -3341 -1255
rect -3375 -1477 -3341 -1461
rect -3279 -1271 -3245 -1255
rect -3279 -1477 -3245 -1467
rect -3183 -1265 -3149 -1255
rect -3183 -1477 -3149 -1461
rect -3087 -1271 -3053 -1255
rect -3087 -1477 -3053 -1467
rect -2991 -1265 -2957 -1255
rect -2991 -1477 -2957 -1461
rect -2895 -1271 -2861 -1255
rect -2895 -1477 -2861 -1467
rect -2799 -1265 -2765 -1255
rect -2799 -1477 -2765 -1461
rect -2617 -1439 -2601 -1213
rect -891 -1213 -841 -1196
rect -798 -1199 -788 -1165
rect -592 -1199 -576 -1165
rect -2524 -1295 -2508 -1261
rect -2314 -1295 -2296 -1261
rect -1649 -1265 -1615 -1255
rect -2524 -1391 -2514 -1357
rect -2318 -1391 -2302 -1357
rect -3326 -1555 -3309 -1520
rect -3275 -1555 -3259 -1520
rect -3037 -1526 -3020 -1520
rect -3225 -1555 -3020 -1526
rect -2986 -1555 -2970 -1520
rect -3326 -1761 -3283 -1555
rect -3225 -1560 -2970 -1555
rect -3225 -1644 -3191 -1560
rect -3157 -1649 -3141 -1615
rect -2765 -1649 -2749 -1615
rect -3225 -1695 -3191 -1679
rect -2617 -1659 -2567 -1439
rect -2524 -1487 -2508 -1453
rect -2314 -1487 -2296 -1453
rect -1649 -1477 -1615 -1461
rect -1553 -1271 -1519 -1255
rect -1553 -1477 -1519 -1467
rect -1457 -1265 -1423 -1255
rect -1457 -1477 -1423 -1461
rect -1361 -1271 -1327 -1255
rect -1361 -1477 -1327 -1467
rect -1265 -1265 -1231 -1255
rect -1265 -1477 -1231 -1461
rect -1169 -1271 -1135 -1255
rect -1169 -1477 -1135 -1467
rect -1073 -1265 -1039 -1255
rect -1073 -1477 -1039 -1461
rect -891 -1439 -875 -1213
rect -798 -1295 -782 -1261
rect -588 -1295 -570 -1261
rect -798 -1391 -788 -1357
rect -592 -1391 -576 -1357
rect -1600 -1555 -1583 -1520
rect -1549 -1555 -1533 -1520
rect -1311 -1526 -1294 -1520
rect -1499 -1555 -1294 -1526
rect -1260 -1555 -1244 -1520
rect -2524 -1649 -2508 -1615
rect -2332 -1649 -2316 -1615
rect -2617 -1693 -2601 -1659
rect -2617 -1709 -2567 -1693
rect -2524 -1737 -2508 -1703
rect -2332 -1737 -2316 -1703
rect -1600 -1761 -1557 -1555
rect -1499 -1560 -1244 -1555
rect -1499 -1644 -1465 -1560
rect -1431 -1649 -1415 -1615
rect -1039 -1649 -1023 -1615
rect -1499 -1695 -1465 -1679
rect -891 -1659 -841 -1439
rect -798 -1487 -782 -1453
rect -588 -1487 -570 -1453
rect -798 -1649 -782 -1615
rect -606 -1649 -590 -1615
rect -891 -1693 -875 -1659
rect -891 -1709 -841 -1693
rect -798 -1737 -782 -1703
rect -606 -1737 -590 -1703
rect -3326 -1777 -3191 -1761
rect -3326 -1812 -3225 -1777
rect -1600 -1777 -1465 -1761
rect -3326 -1828 -3191 -1812
rect -3157 -1841 -3141 -1807
rect -2765 -1841 -2749 -1807
rect -1600 -1812 -1499 -1777
rect -1600 -1828 -1465 -1812
rect -1431 -1841 -1415 -1807
rect -1039 -1841 -1023 -1807
rect -3153 -1951 -3126 -1877
rect -2791 -1951 -2753 -1877
rect -1427 -1951 -1400 -1877
rect -1065 -1951 -1027 -1877
rect -3247 -2455 -3173 -2408
rect -2933 -2455 -2833 -2408
rect -1521 -2455 -1447 -2408
rect -1207 -2455 -1107 -2408
rect -2617 -2505 -2567 -2488
rect -2524 -2491 -2514 -2457
rect -2318 -2491 -2302 -2457
rect -3375 -2557 -3341 -2547
rect -3375 -2769 -3341 -2753
rect -3279 -2563 -3245 -2547
rect -3279 -2769 -3245 -2759
rect -3183 -2557 -3149 -2547
rect -3183 -2769 -3149 -2753
rect -3087 -2563 -3053 -2547
rect -3087 -2769 -3053 -2759
rect -2991 -2557 -2957 -2547
rect -2991 -2769 -2957 -2753
rect -2895 -2563 -2861 -2547
rect -2895 -2769 -2861 -2759
rect -2799 -2557 -2765 -2547
rect -2799 -2769 -2765 -2753
rect -2617 -2731 -2601 -2505
rect -891 -2505 -841 -2488
rect -798 -2491 -788 -2457
rect -592 -2491 -576 -2457
rect -2524 -2587 -2508 -2553
rect -2314 -2587 -2296 -2553
rect -1649 -2557 -1615 -2547
rect -2524 -2683 -2514 -2649
rect -2318 -2683 -2302 -2649
rect -3326 -2847 -3309 -2812
rect -3275 -2847 -3259 -2812
rect -3037 -2818 -3020 -2812
rect -3225 -2847 -3020 -2818
rect -2986 -2847 -2970 -2812
rect -3326 -3053 -3283 -2847
rect -3225 -2852 -2970 -2847
rect -3225 -2936 -3191 -2852
rect -3157 -2941 -3141 -2907
rect -2765 -2941 -2749 -2907
rect -3225 -2987 -3191 -2971
rect -2617 -2951 -2567 -2731
rect -2524 -2779 -2508 -2745
rect -2314 -2779 -2296 -2745
rect -1649 -2769 -1615 -2753
rect -1553 -2563 -1519 -2547
rect -1553 -2769 -1519 -2759
rect -1457 -2557 -1423 -2547
rect -1457 -2769 -1423 -2753
rect -1361 -2563 -1327 -2547
rect -1361 -2769 -1327 -2759
rect -1265 -2557 -1231 -2547
rect -1265 -2769 -1231 -2753
rect -1169 -2563 -1135 -2547
rect -1169 -2769 -1135 -2759
rect -1073 -2557 -1039 -2547
rect -1073 -2769 -1039 -2753
rect -891 -2731 -875 -2505
rect -798 -2587 -782 -2553
rect -588 -2587 -570 -2553
rect -798 -2683 -788 -2649
rect -592 -2683 -576 -2649
rect -1600 -2847 -1583 -2812
rect -1549 -2847 -1533 -2812
rect -1311 -2818 -1294 -2812
rect -1499 -2847 -1294 -2818
rect -1260 -2847 -1244 -2812
rect -2524 -2941 -2508 -2907
rect -2332 -2941 -2316 -2907
rect -2617 -2985 -2601 -2951
rect -2617 -3001 -2567 -2985
rect -2524 -3029 -2508 -2995
rect -2332 -3029 -2316 -2995
rect -1600 -3053 -1557 -2847
rect -1499 -2852 -1244 -2847
rect -1499 -2936 -1465 -2852
rect -1431 -2941 -1415 -2907
rect -1039 -2941 -1023 -2907
rect -1499 -2987 -1465 -2971
rect -891 -2951 -841 -2731
rect -798 -2779 -782 -2745
rect -588 -2779 -570 -2745
rect -798 -2941 -782 -2907
rect -606 -2941 -590 -2907
rect -891 -2985 -875 -2951
rect -891 -3001 -841 -2985
rect -798 -3029 -782 -2995
rect -606 -3029 -590 -2995
rect -3326 -3069 -3191 -3053
rect -3326 -3104 -3225 -3069
rect -1600 -3069 -1465 -3053
rect -3326 -3120 -3191 -3104
rect -3157 -3133 -3141 -3099
rect -2765 -3133 -2749 -3099
rect -1600 -3104 -1499 -3069
rect -1600 -3120 -1465 -3104
rect -1431 -3133 -1415 -3099
rect -1039 -3133 -1023 -3099
rect -3153 -3243 -3126 -3169
rect -2791 -3243 -2753 -3169
rect -1427 -3243 -1400 -3169
rect -1065 -3243 -1027 -3169
rect -3247 -4427 -3173 -4380
rect -2933 -4427 -2833 -4380
rect -1521 -4427 -1447 -4380
rect -1207 -4427 -1107 -4380
rect -2617 -4477 -2567 -4460
rect -2524 -4463 -2514 -4429
rect -2318 -4463 -2302 -4429
rect -3375 -4529 -3341 -4519
rect -3375 -4741 -3341 -4725
rect -3279 -4535 -3245 -4519
rect -3279 -4741 -3245 -4731
rect -3183 -4529 -3149 -4519
rect -3183 -4741 -3149 -4725
rect -3087 -4535 -3053 -4519
rect -3087 -4741 -3053 -4731
rect -2991 -4529 -2957 -4519
rect -2991 -4741 -2957 -4725
rect -2895 -4535 -2861 -4519
rect -2895 -4741 -2861 -4731
rect -2799 -4529 -2765 -4519
rect -2799 -4741 -2765 -4725
rect -2617 -4703 -2601 -4477
rect -891 -4477 -841 -4460
rect -798 -4463 -788 -4429
rect -592 -4463 -576 -4429
rect -2524 -4559 -2508 -4525
rect -2314 -4559 -2296 -4525
rect -1649 -4529 -1615 -4519
rect -2524 -4655 -2514 -4621
rect -2318 -4655 -2302 -4621
rect -3326 -4819 -3309 -4784
rect -3275 -4819 -3259 -4784
rect -3037 -4790 -3020 -4784
rect -3225 -4819 -3020 -4790
rect -2986 -4819 -2970 -4784
rect -3326 -5025 -3283 -4819
rect -3225 -4824 -2970 -4819
rect -3225 -4908 -3191 -4824
rect -3157 -4913 -3141 -4879
rect -2765 -4913 -2749 -4879
rect -3225 -4959 -3191 -4943
rect -2617 -4923 -2567 -4703
rect -2524 -4751 -2508 -4717
rect -2314 -4751 -2296 -4717
rect -1649 -4741 -1615 -4725
rect -1553 -4535 -1519 -4519
rect -1553 -4741 -1519 -4731
rect -1457 -4529 -1423 -4519
rect -1457 -4741 -1423 -4725
rect -1361 -4535 -1327 -4519
rect -1361 -4741 -1327 -4731
rect -1265 -4529 -1231 -4519
rect -1265 -4741 -1231 -4725
rect -1169 -4535 -1135 -4519
rect -1169 -4741 -1135 -4731
rect -1073 -4529 -1039 -4519
rect -1073 -4741 -1039 -4725
rect -891 -4703 -875 -4477
rect -798 -4559 -782 -4525
rect -588 -4559 -570 -4525
rect -798 -4655 -788 -4621
rect -592 -4655 -576 -4621
rect -1600 -4819 -1583 -4784
rect -1549 -4819 -1533 -4784
rect -1311 -4790 -1294 -4784
rect -1499 -4819 -1294 -4790
rect -1260 -4819 -1244 -4784
rect -2524 -4913 -2508 -4879
rect -2332 -4913 -2316 -4879
rect -2617 -4957 -2601 -4923
rect -2617 -4973 -2567 -4957
rect -2524 -5001 -2508 -4967
rect -2332 -5001 -2316 -4967
rect -1600 -5025 -1557 -4819
rect -1499 -4824 -1244 -4819
rect -1499 -4908 -1465 -4824
rect -1431 -4913 -1415 -4879
rect -1039 -4913 -1023 -4879
rect -1499 -4959 -1465 -4943
rect -891 -4923 -841 -4703
rect -798 -4751 -782 -4717
rect -588 -4751 -570 -4717
rect -798 -4913 -782 -4879
rect -606 -4913 -590 -4879
rect -891 -4957 -875 -4923
rect -891 -4973 -841 -4957
rect -798 -5001 -782 -4967
rect -606 -5001 -590 -4967
rect -3326 -5041 -3191 -5025
rect -3326 -5076 -3225 -5041
rect -1600 -5041 -1465 -5025
rect -3326 -5092 -3191 -5076
rect -3157 -5105 -3141 -5071
rect -2765 -5105 -2749 -5071
rect -1600 -5076 -1499 -5041
rect -1600 -5092 -1465 -5076
rect -1431 -5105 -1415 -5071
rect -1039 -5105 -1023 -5071
rect -3153 -5215 -3126 -5141
rect -2791 -5215 -2753 -5141
rect -1427 -5215 -1400 -5141
rect -1065 -5215 -1027 -5141
rect -3247 -5719 -3173 -5672
rect -2933 -5719 -2833 -5672
rect -1521 -5719 -1447 -5672
rect -1207 -5719 -1107 -5672
rect -2617 -5769 -2567 -5752
rect -2524 -5755 -2514 -5721
rect -2318 -5755 -2302 -5721
rect -3375 -5821 -3341 -5811
rect -3375 -6033 -3341 -6017
rect -3279 -5827 -3245 -5811
rect -3279 -6033 -3245 -6023
rect -3183 -5821 -3149 -5811
rect -3183 -6033 -3149 -6017
rect -3087 -5827 -3053 -5811
rect -3087 -6033 -3053 -6023
rect -2991 -5821 -2957 -5811
rect -2991 -6033 -2957 -6017
rect -2895 -5827 -2861 -5811
rect -2895 -6033 -2861 -6023
rect -2799 -5821 -2765 -5811
rect -2799 -6033 -2765 -6017
rect -2617 -5995 -2601 -5769
rect -891 -5769 -841 -5752
rect -798 -5755 -788 -5721
rect -592 -5755 -576 -5721
rect -2524 -5851 -2508 -5817
rect -2314 -5851 -2296 -5817
rect -1649 -5821 -1615 -5811
rect -2524 -5947 -2514 -5913
rect -2318 -5947 -2302 -5913
rect -3326 -6111 -3309 -6076
rect -3275 -6111 -3259 -6076
rect -3037 -6082 -3020 -6076
rect -3225 -6111 -3020 -6082
rect -2986 -6111 -2970 -6076
rect -3326 -6317 -3283 -6111
rect -3225 -6116 -2970 -6111
rect -3225 -6200 -3191 -6116
rect -3157 -6205 -3141 -6171
rect -2765 -6205 -2749 -6171
rect -3225 -6251 -3191 -6235
rect -2617 -6215 -2567 -5995
rect -2524 -6043 -2508 -6009
rect -2314 -6043 -2296 -6009
rect -1649 -6033 -1615 -6017
rect -1553 -5827 -1519 -5811
rect -1553 -6033 -1519 -6023
rect -1457 -5821 -1423 -5811
rect -1457 -6033 -1423 -6017
rect -1361 -5827 -1327 -5811
rect -1361 -6033 -1327 -6023
rect -1265 -5821 -1231 -5811
rect -1265 -6033 -1231 -6017
rect -1169 -5827 -1135 -5811
rect -1169 -6033 -1135 -6023
rect -1073 -5821 -1039 -5811
rect -1073 -6033 -1039 -6017
rect -891 -5995 -875 -5769
rect -798 -5851 -782 -5817
rect -588 -5851 -570 -5817
rect -798 -5947 -788 -5913
rect -592 -5947 -576 -5913
rect -1600 -6111 -1583 -6076
rect -1549 -6111 -1533 -6076
rect -1311 -6082 -1294 -6076
rect -1499 -6111 -1294 -6082
rect -1260 -6111 -1244 -6076
rect -2524 -6205 -2508 -6171
rect -2332 -6205 -2316 -6171
rect -2617 -6249 -2601 -6215
rect -2617 -6265 -2567 -6249
rect -2524 -6293 -2508 -6259
rect -2332 -6293 -2316 -6259
rect -1600 -6317 -1557 -6111
rect -1499 -6116 -1244 -6111
rect -1499 -6200 -1465 -6116
rect -1431 -6205 -1415 -6171
rect -1039 -6205 -1023 -6171
rect -1499 -6251 -1465 -6235
rect -891 -6215 -841 -5995
rect -798 -6043 -782 -6009
rect -588 -6043 -570 -6009
rect -798 -6205 -782 -6171
rect -606 -6205 -590 -6171
rect -891 -6249 -875 -6215
rect -891 -6265 -841 -6249
rect -798 -6293 -782 -6259
rect -606 -6293 -590 -6259
rect -3326 -6333 -3191 -6317
rect -3326 -6368 -3225 -6333
rect -1600 -6333 -1465 -6317
rect -3326 -6384 -3191 -6368
rect -3157 -6397 -3141 -6363
rect -2765 -6397 -2749 -6363
rect -1600 -6368 -1499 -6333
rect -1600 -6384 -1465 -6368
rect -1431 -6397 -1415 -6363
rect -1039 -6397 -1023 -6363
rect -3153 -6507 -3126 -6433
rect -2791 -6507 -2753 -6433
rect -1427 -6507 -1400 -6433
rect -1065 -6507 -1027 -6433
<< viali >>
rect -3197 3874 -2957 3921
rect -1356 3874 -1116 3921
rect 485 3874 725 3921
rect 2326 3874 2566 3921
rect -2538 3838 -2532 3872
rect -2532 3838 -2459 3872
rect -3399 3766 -3365 3772
rect -3399 3692 -3365 3766
rect -3303 3576 -3269 3650
rect -3303 3570 -3269 3576
rect -3207 3766 -3173 3772
rect -3207 3692 -3173 3766
rect -3111 3576 -3077 3650
rect -3111 3570 -3077 3576
rect -3015 3766 -2981 3772
rect -3015 3692 -2981 3766
rect -2919 3576 -2885 3650
rect -2919 3570 -2885 3576
rect -2823 3766 -2789 3772
rect -2823 3692 -2789 3766
rect -2625 3598 -2591 3824
rect -697 3838 -691 3872
rect -691 3838 -618 3872
rect -2415 3742 -2338 3776
rect -1558 3766 -1524 3772
rect -1558 3692 -1524 3766
rect -2538 3646 -2532 3680
rect -2532 3646 -2459 3680
rect -3333 3482 -3299 3517
rect -3044 3482 -3010 3517
rect -3249 3358 -3215 3393
rect -3165 3388 -2789 3422
rect -2415 3550 -2338 3584
rect -1462 3576 -1428 3650
rect -1462 3570 -1428 3576
rect -1366 3766 -1332 3772
rect -1366 3692 -1332 3766
rect -1270 3576 -1236 3650
rect -1270 3570 -1236 3576
rect -1174 3766 -1140 3772
rect -1174 3692 -1140 3766
rect -1078 3576 -1044 3650
rect -1078 3570 -1044 3576
rect -982 3766 -948 3772
rect -982 3692 -948 3766
rect -784 3598 -750 3824
rect 1144 3838 1150 3872
rect 1150 3838 1223 3872
rect -574 3742 -497 3776
rect 283 3766 317 3772
rect 283 3692 317 3766
rect -697 3646 -691 3680
rect -691 3646 -618 3680
rect -1492 3482 -1458 3517
rect -1203 3482 -1169 3517
rect -2532 3388 -2356 3422
rect -2625 3344 -2591 3378
rect -2532 3300 -2356 3334
rect -1408 3358 -1374 3393
rect -1324 3388 -948 3422
rect -574 3550 -497 3584
rect 379 3576 413 3650
rect 379 3570 413 3576
rect 475 3766 509 3772
rect 475 3692 509 3766
rect 571 3576 605 3650
rect 571 3570 605 3576
rect 667 3766 701 3772
rect 667 3692 701 3766
rect 763 3576 797 3650
rect 763 3570 797 3576
rect 859 3766 893 3772
rect 859 3692 893 3766
rect 1057 3598 1091 3824
rect 2985 3838 2991 3872
rect 2991 3838 3064 3872
rect 1267 3742 1344 3776
rect 2124 3766 2158 3772
rect 2124 3692 2158 3766
rect 1144 3646 1150 3680
rect 1150 3646 1223 3680
rect 349 3482 383 3517
rect 638 3482 672 3517
rect -691 3388 -515 3422
rect -784 3344 -750 3378
rect -691 3300 -515 3334
rect 433 3358 467 3393
rect 517 3388 893 3422
rect 1267 3550 1344 3584
rect 2220 3576 2254 3650
rect 2220 3570 2254 3576
rect 2316 3766 2350 3772
rect 2316 3692 2350 3766
rect 2412 3576 2446 3650
rect 2412 3570 2446 3576
rect 2508 3766 2542 3772
rect 2508 3692 2542 3766
rect 2604 3576 2638 3650
rect 2604 3570 2638 3576
rect 2700 3766 2734 3772
rect 2700 3692 2734 3766
rect 2898 3598 2932 3824
rect 3108 3742 3185 3776
rect 2985 3646 2991 3680
rect 2991 3646 3064 3680
rect 2190 3482 2224 3517
rect 2479 3482 2513 3517
rect 1150 3388 1326 3422
rect 1057 3344 1091 3378
rect 1150 3300 1326 3334
rect 2274 3358 2308 3393
rect 2358 3388 2734 3422
rect 3108 3550 3185 3584
rect 2991 3388 3167 3422
rect 2898 3344 2932 3378
rect 2991 3300 3167 3334
rect -3165 3196 -2789 3230
rect -1324 3196 -948 3230
rect 517 3196 893 3230
rect 2358 3196 2734 3230
rect -3150 3086 -2815 3155
rect -1309 3086 -974 3155
rect 532 3086 867 3155
rect 2373 3086 2708 3155
rect -3173 2102 -2933 2149
rect -1447 2102 -1207 2149
rect -2514 2066 -2508 2100
rect -2508 2066 -2435 2100
rect -3375 1994 -3341 2000
rect -3375 1920 -3341 1994
rect -3279 1804 -3245 1878
rect -3279 1798 -3245 1804
rect -3183 1994 -3149 2000
rect -3183 1920 -3149 1994
rect -3087 1804 -3053 1878
rect -3087 1798 -3053 1804
rect -2991 1994 -2957 2000
rect -2991 1920 -2957 1994
rect -2895 1804 -2861 1878
rect -2895 1798 -2861 1804
rect -2799 1994 -2765 2000
rect -2799 1920 -2765 1994
rect -2601 1826 -2567 2052
rect -788 2066 -782 2100
rect -782 2066 -709 2100
rect -2391 1970 -2314 2004
rect -1649 1994 -1615 2000
rect -1649 1920 -1615 1994
rect -2514 1874 -2508 1908
rect -2508 1874 -2435 1908
rect -3309 1710 -3275 1745
rect -3020 1710 -2986 1745
rect -3225 1586 -3191 1621
rect -3141 1616 -2765 1650
rect -2391 1778 -2314 1812
rect -1553 1804 -1519 1878
rect -1553 1798 -1519 1804
rect -1457 1994 -1423 2000
rect -1457 1920 -1423 1994
rect -1361 1804 -1327 1878
rect -1361 1798 -1327 1804
rect -1265 1994 -1231 2000
rect -1265 1920 -1231 1994
rect -1169 1804 -1135 1878
rect -1169 1798 -1135 1804
rect -1073 1994 -1039 2000
rect -1073 1920 -1039 1994
rect -875 1826 -841 2052
rect -665 1970 -588 2004
rect -788 1874 -782 1908
rect -782 1874 -709 1908
rect -1583 1710 -1549 1745
rect -1294 1710 -1260 1745
rect -2508 1616 -2332 1650
rect -2601 1572 -2567 1606
rect -2508 1528 -2332 1562
rect -1499 1586 -1465 1621
rect -1415 1616 -1039 1650
rect -665 1778 -588 1812
rect -782 1616 -606 1650
rect -875 1572 -841 1606
rect -782 1528 -606 1562
rect -3141 1424 -2765 1458
rect -1415 1424 -1039 1458
rect -3126 1314 -2791 1383
rect -1400 1314 -1065 1383
rect -3173 810 -2933 857
rect -1447 810 -1207 857
rect -2514 774 -2508 808
rect -2508 774 -2435 808
rect -3375 702 -3341 708
rect -3375 628 -3341 702
rect -3279 512 -3245 586
rect -3279 506 -3245 512
rect -3183 702 -3149 708
rect -3183 628 -3149 702
rect -3087 512 -3053 586
rect -3087 506 -3053 512
rect -2991 702 -2957 708
rect -2991 628 -2957 702
rect -2895 512 -2861 586
rect -2895 506 -2861 512
rect -2799 702 -2765 708
rect -2799 628 -2765 702
rect -2601 534 -2567 760
rect -788 774 -782 808
rect -782 774 -709 808
rect -2391 678 -2314 712
rect -1649 702 -1615 708
rect -1649 628 -1615 702
rect -2514 582 -2508 616
rect -2508 582 -2435 616
rect -3309 418 -3275 453
rect -3020 418 -2986 453
rect -3225 294 -3191 329
rect -3141 324 -2765 358
rect -2391 486 -2314 520
rect -1553 512 -1519 586
rect -1553 506 -1519 512
rect -1457 702 -1423 708
rect -1457 628 -1423 702
rect -1361 512 -1327 586
rect -1361 506 -1327 512
rect -1265 702 -1231 708
rect -1265 628 -1231 702
rect -1169 512 -1135 586
rect -1169 506 -1135 512
rect -1073 702 -1039 708
rect -1073 628 -1039 702
rect -875 534 -841 760
rect -665 678 -588 712
rect -788 582 -782 616
rect -782 582 -709 616
rect -1583 418 -1549 453
rect -1294 418 -1260 453
rect -2508 324 -2332 358
rect -2601 280 -2567 314
rect -2508 236 -2332 270
rect -1499 294 -1465 329
rect -1415 324 -1039 358
rect -665 486 -588 520
rect -782 324 -606 358
rect -875 280 -841 314
rect -782 236 -606 270
rect -3141 132 -2765 166
rect -1415 132 -1039 166
rect -3126 22 -2791 91
rect -1400 22 -1065 91
rect -3173 -1163 -2933 -1116
rect -1447 -1163 -1207 -1116
rect -2514 -1199 -2508 -1165
rect -2508 -1199 -2435 -1165
rect -3375 -1271 -3341 -1265
rect -3375 -1345 -3341 -1271
rect -3279 -1461 -3245 -1387
rect -3279 -1467 -3245 -1461
rect -3183 -1271 -3149 -1265
rect -3183 -1345 -3149 -1271
rect -3087 -1461 -3053 -1387
rect -3087 -1467 -3053 -1461
rect -2991 -1271 -2957 -1265
rect -2991 -1345 -2957 -1271
rect -2895 -1461 -2861 -1387
rect -2895 -1467 -2861 -1461
rect -2799 -1271 -2765 -1265
rect -2799 -1345 -2765 -1271
rect -2601 -1439 -2567 -1213
rect -788 -1199 -782 -1165
rect -782 -1199 -709 -1165
rect -2391 -1295 -2314 -1261
rect -1649 -1271 -1615 -1265
rect -1649 -1345 -1615 -1271
rect -2514 -1391 -2508 -1357
rect -2508 -1391 -2435 -1357
rect -3309 -1555 -3275 -1520
rect -3020 -1555 -2986 -1520
rect -3225 -1679 -3191 -1644
rect -3141 -1649 -2765 -1615
rect -2391 -1487 -2314 -1453
rect -1553 -1461 -1519 -1387
rect -1553 -1467 -1519 -1461
rect -1457 -1271 -1423 -1265
rect -1457 -1345 -1423 -1271
rect -1361 -1461 -1327 -1387
rect -1361 -1467 -1327 -1461
rect -1265 -1271 -1231 -1265
rect -1265 -1345 -1231 -1271
rect -1169 -1461 -1135 -1387
rect -1169 -1467 -1135 -1461
rect -1073 -1271 -1039 -1265
rect -1073 -1345 -1039 -1271
rect -875 -1439 -841 -1213
rect -665 -1295 -588 -1261
rect -788 -1391 -782 -1357
rect -782 -1391 -709 -1357
rect -1583 -1555 -1549 -1520
rect -1294 -1555 -1260 -1520
rect -2508 -1649 -2332 -1615
rect -2601 -1693 -2567 -1659
rect -2508 -1737 -2332 -1703
rect -1499 -1679 -1465 -1644
rect -1415 -1649 -1039 -1615
rect -665 -1487 -588 -1453
rect -782 -1649 -606 -1615
rect -875 -1693 -841 -1659
rect -782 -1737 -606 -1703
rect -3141 -1841 -2765 -1807
rect -1415 -1841 -1039 -1807
rect -3126 -1951 -2791 -1882
rect -1400 -1951 -1065 -1882
rect -3173 -2455 -2933 -2408
rect -1447 -2455 -1207 -2408
rect -2514 -2491 -2508 -2457
rect -2508 -2491 -2435 -2457
rect -3375 -2563 -3341 -2557
rect -3375 -2637 -3341 -2563
rect -3279 -2753 -3245 -2679
rect -3279 -2759 -3245 -2753
rect -3183 -2563 -3149 -2557
rect -3183 -2637 -3149 -2563
rect -3087 -2753 -3053 -2679
rect -3087 -2759 -3053 -2753
rect -2991 -2563 -2957 -2557
rect -2991 -2637 -2957 -2563
rect -2895 -2753 -2861 -2679
rect -2895 -2759 -2861 -2753
rect -2799 -2563 -2765 -2557
rect -2799 -2637 -2765 -2563
rect -2601 -2731 -2567 -2505
rect -788 -2491 -782 -2457
rect -782 -2491 -709 -2457
rect -2391 -2587 -2314 -2553
rect -1649 -2563 -1615 -2557
rect -1649 -2637 -1615 -2563
rect -2514 -2683 -2508 -2649
rect -2508 -2683 -2435 -2649
rect -3309 -2847 -3275 -2812
rect -3020 -2847 -2986 -2812
rect -3225 -2971 -3191 -2936
rect -3141 -2941 -2765 -2907
rect -2391 -2779 -2314 -2745
rect -1553 -2753 -1519 -2679
rect -1553 -2759 -1519 -2753
rect -1457 -2563 -1423 -2557
rect -1457 -2637 -1423 -2563
rect -1361 -2753 -1327 -2679
rect -1361 -2759 -1327 -2753
rect -1265 -2563 -1231 -2557
rect -1265 -2637 -1231 -2563
rect -1169 -2753 -1135 -2679
rect -1169 -2759 -1135 -2753
rect -1073 -2563 -1039 -2557
rect -1073 -2637 -1039 -2563
rect -875 -2731 -841 -2505
rect -665 -2587 -588 -2553
rect -788 -2683 -782 -2649
rect -782 -2683 -709 -2649
rect -1583 -2847 -1549 -2812
rect -1294 -2847 -1260 -2812
rect -2508 -2941 -2332 -2907
rect -2601 -2985 -2567 -2951
rect -2508 -3029 -2332 -2995
rect -1499 -2971 -1465 -2936
rect -1415 -2941 -1039 -2907
rect -665 -2779 -588 -2745
rect -782 -2941 -606 -2907
rect -875 -2985 -841 -2951
rect -782 -3029 -606 -2995
rect -3141 -3133 -2765 -3099
rect -1415 -3133 -1039 -3099
rect -3126 -3243 -2791 -3174
rect -1400 -3243 -1065 -3174
rect -3173 -4427 -2933 -4380
rect -1447 -4427 -1207 -4380
rect -2514 -4463 -2508 -4429
rect -2508 -4463 -2435 -4429
rect -3375 -4535 -3341 -4529
rect -3375 -4609 -3341 -4535
rect -3279 -4725 -3245 -4651
rect -3279 -4731 -3245 -4725
rect -3183 -4535 -3149 -4529
rect -3183 -4609 -3149 -4535
rect -3087 -4725 -3053 -4651
rect -3087 -4731 -3053 -4725
rect -2991 -4535 -2957 -4529
rect -2991 -4609 -2957 -4535
rect -2895 -4725 -2861 -4651
rect -2895 -4731 -2861 -4725
rect -2799 -4535 -2765 -4529
rect -2799 -4609 -2765 -4535
rect -2601 -4703 -2567 -4477
rect -788 -4463 -782 -4429
rect -782 -4463 -709 -4429
rect -2391 -4559 -2314 -4525
rect -1649 -4535 -1615 -4529
rect -1649 -4609 -1615 -4535
rect -2514 -4655 -2508 -4621
rect -2508 -4655 -2435 -4621
rect -3309 -4819 -3275 -4784
rect -3020 -4819 -2986 -4784
rect -3225 -4943 -3191 -4908
rect -3141 -4913 -2765 -4879
rect -2391 -4751 -2314 -4717
rect -1553 -4725 -1519 -4651
rect -1553 -4731 -1519 -4725
rect -1457 -4535 -1423 -4529
rect -1457 -4609 -1423 -4535
rect -1361 -4725 -1327 -4651
rect -1361 -4731 -1327 -4725
rect -1265 -4535 -1231 -4529
rect -1265 -4609 -1231 -4535
rect -1169 -4725 -1135 -4651
rect -1169 -4731 -1135 -4725
rect -1073 -4535 -1039 -4529
rect -1073 -4609 -1039 -4535
rect -875 -4703 -841 -4477
rect -665 -4559 -588 -4525
rect -788 -4655 -782 -4621
rect -782 -4655 -709 -4621
rect -1583 -4819 -1549 -4784
rect -1294 -4819 -1260 -4784
rect -2508 -4913 -2332 -4879
rect -2601 -4957 -2567 -4923
rect -2508 -5001 -2332 -4967
rect -1499 -4943 -1465 -4908
rect -1415 -4913 -1039 -4879
rect -665 -4751 -588 -4717
rect -782 -4913 -606 -4879
rect -875 -4957 -841 -4923
rect -782 -5001 -606 -4967
rect -3141 -5105 -2765 -5071
rect -1415 -5105 -1039 -5071
rect -3126 -5215 -2791 -5146
rect -1400 -5215 -1065 -5146
rect -3173 -5719 -2933 -5672
rect -1447 -5719 -1207 -5672
rect -2514 -5755 -2508 -5721
rect -2508 -5755 -2435 -5721
rect -3375 -5827 -3341 -5821
rect -3375 -5901 -3341 -5827
rect -3279 -6017 -3245 -5943
rect -3279 -6023 -3245 -6017
rect -3183 -5827 -3149 -5821
rect -3183 -5901 -3149 -5827
rect -3087 -6017 -3053 -5943
rect -3087 -6023 -3053 -6017
rect -2991 -5827 -2957 -5821
rect -2991 -5901 -2957 -5827
rect -2895 -6017 -2861 -5943
rect -2895 -6023 -2861 -6017
rect -2799 -5827 -2765 -5821
rect -2799 -5901 -2765 -5827
rect -2601 -5995 -2567 -5769
rect -788 -5755 -782 -5721
rect -782 -5755 -709 -5721
rect -2391 -5851 -2314 -5817
rect -1649 -5827 -1615 -5821
rect -1649 -5901 -1615 -5827
rect -2514 -5947 -2508 -5913
rect -2508 -5947 -2435 -5913
rect -3309 -6111 -3275 -6076
rect -3020 -6111 -2986 -6076
rect -3225 -6235 -3191 -6200
rect -3141 -6205 -2765 -6171
rect -2391 -6043 -2314 -6009
rect -1553 -6017 -1519 -5943
rect -1553 -6023 -1519 -6017
rect -1457 -5827 -1423 -5821
rect -1457 -5901 -1423 -5827
rect -1361 -6017 -1327 -5943
rect -1361 -6023 -1327 -6017
rect -1265 -5827 -1231 -5821
rect -1265 -5901 -1231 -5827
rect -1169 -6017 -1135 -5943
rect -1169 -6023 -1135 -6017
rect -1073 -5827 -1039 -5821
rect -1073 -5901 -1039 -5827
rect -875 -5995 -841 -5769
rect -665 -5851 -588 -5817
rect -788 -5947 -782 -5913
rect -782 -5947 -709 -5913
rect -1583 -6111 -1549 -6076
rect -1294 -6111 -1260 -6076
rect -2508 -6205 -2332 -6171
rect -2601 -6249 -2567 -6215
rect -2508 -6293 -2332 -6259
rect -1499 -6235 -1465 -6200
rect -1415 -6205 -1039 -6171
rect -665 -6043 -588 -6009
rect -782 -6205 -606 -6171
rect -875 -6249 -841 -6215
rect -782 -6293 -606 -6259
rect -3141 -6397 -2765 -6363
rect -1415 -6397 -1039 -6363
rect -3126 -6507 -2791 -6438
rect -1400 -6507 -1065 -6438
<< metal1 >>
rect -3271 3921 -2934 3933
rect -3271 3874 -3197 3921
rect -2957 3874 -2934 3921
rect -1430 3921 -1093 3933
rect -3271 3814 -2934 3874
rect -2548 3872 -2326 3920
rect -2548 3868 -2538 3872
rect -2658 3824 -2575 3840
rect -3412 3778 -2778 3814
rect -3412 3772 -2777 3778
rect -3412 3692 -3399 3772
rect -3365 3692 -3207 3772
rect -3173 3692 -3015 3772
rect -2981 3692 -2823 3772
rect -2789 3692 -2777 3772
rect -3412 3686 -2777 3692
rect -3412 3685 -2778 3686
rect -2658 3656 -2625 3824
rect -3319 3650 -2625 3656
rect -3319 3570 -3303 3650
rect -3269 3570 -3111 3650
rect -3077 3570 -2919 3650
rect -2885 3598 -2625 3650
rect -2591 3598 -2575 3824
rect -2544 3838 -2538 3868
rect -2459 3868 -2326 3872
rect -1430 3874 -1356 3921
rect -1116 3874 -1093 3921
rect 411 3921 748 3933
rect -2459 3838 -2453 3868
rect -2544 3680 -2453 3838
rect -2544 3646 -2538 3680
rect -2459 3646 -2453 3680
rect -2544 3630 -2453 3646
rect -2421 3776 -2268 3840
rect -1430 3814 -1093 3874
rect -707 3872 -485 3920
rect -707 3868 -697 3872
rect -817 3824 -734 3840
rect -2421 3742 -2415 3776
rect -2338 3742 -2268 3776
rect -2885 3570 -2575 3598
rect -2421 3584 -2268 3742
rect -1571 3778 -937 3814
rect -1571 3772 -936 3778
rect -1571 3692 -1558 3772
rect -1524 3692 -1366 3772
rect -1332 3692 -1174 3772
rect -1140 3692 -982 3772
rect -948 3692 -936 3772
rect -1571 3686 -936 3692
rect -1571 3685 -937 3686
rect -817 3656 -784 3824
rect -3319 3564 -2575 3570
rect -3447 3517 -3283 3535
rect -3447 3515 -3333 3517
rect -3447 3405 -3422 3515
rect -3299 3482 -3283 3517
rect -3327 3405 -3283 3482
rect -3447 3400 -3283 3405
rect -3255 3517 -2995 3536
rect -3255 3482 -3044 3517
rect -3010 3482 -2995 3517
rect -3255 3462 -2995 3482
rect -3255 3393 -3205 3462
rect -2919 3434 -2575 3564
rect -3544 3371 -3354 3372
rect -3255 3371 -3249 3393
rect -3544 3358 -3249 3371
rect -3215 3358 -3205 3393
rect -3177 3422 -2575 3434
rect -3177 3388 -3165 3422
rect -2789 3388 -2575 3422
rect -3177 3382 -2575 3388
rect -2544 3550 -2415 3584
rect -2338 3550 -2268 3584
rect -1478 3650 -784 3656
rect -1478 3570 -1462 3650
rect -1428 3570 -1270 3650
rect -1236 3570 -1078 3650
rect -1044 3598 -784 3650
rect -750 3598 -734 3824
rect -703 3838 -697 3868
rect -618 3868 -485 3872
rect 411 3874 485 3921
rect 725 3874 748 3921
rect 2252 3921 2589 3933
rect -618 3838 -612 3868
rect -703 3680 -612 3838
rect -703 3646 -697 3680
rect -618 3646 -612 3680
rect -703 3630 -612 3646
rect -580 3776 -427 3840
rect 411 3814 748 3874
rect 1134 3872 1356 3920
rect 1134 3868 1144 3872
rect 1024 3824 1107 3840
rect -580 3742 -574 3776
rect -497 3742 -427 3776
rect -1044 3570 -734 3598
rect -580 3584 -427 3742
rect 270 3778 904 3814
rect 270 3772 905 3778
rect 270 3692 283 3772
rect 317 3692 475 3772
rect 509 3692 667 3772
rect 701 3692 859 3772
rect 893 3692 905 3772
rect 270 3686 905 3692
rect 270 3685 904 3686
rect 1024 3656 1057 3824
rect -1478 3564 -734 3570
rect -2544 3515 -2268 3550
rect -1606 3517 -1442 3535
rect -1606 3515 -1492 3517
rect -2544 3422 -2205 3515
rect -2544 3388 -2532 3422
rect -2356 3388 -2205 3422
rect -1606 3405 -1581 3515
rect -1458 3482 -1442 3517
rect -1486 3405 -1442 3482
rect -1606 3400 -1442 3405
rect -1414 3517 -1154 3536
rect -1414 3482 -1203 3517
rect -1169 3482 -1154 3517
rect -1414 3462 -1154 3482
rect -2544 3382 -2344 3388
rect -3544 3244 -3205 3358
rect -2658 3378 -2575 3382
rect -2658 3344 -2625 3378
rect -2591 3344 -2575 3378
rect -2658 3327 -2575 3344
rect -2544 3334 -2344 3341
rect -2544 3300 -2532 3334
rect -2356 3300 -2344 3334
rect -2316 3327 -2205 3388
rect -1414 3393 -1364 3462
rect -1078 3434 -734 3564
rect -1414 3371 -1408 3393
rect -1748 3358 -1408 3371
rect -1374 3358 -1364 3393
rect -1336 3422 -734 3434
rect -1336 3388 -1324 3422
rect -948 3388 -734 3422
rect -1336 3382 -734 3388
rect -703 3550 -574 3584
rect -497 3550 -427 3584
rect 363 3650 1057 3656
rect 363 3570 379 3650
rect 413 3570 571 3650
rect 605 3570 763 3650
rect 797 3598 1057 3650
rect 1091 3598 1107 3824
rect 1138 3838 1144 3868
rect 1223 3868 1356 3872
rect 2252 3874 2326 3921
rect 2566 3874 2589 3921
rect 1223 3838 1229 3868
rect 1138 3680 1229 3838
rect 1138 3646 1144 3680
rect 1223 3646 1229 3680
rect 1138 3630 1229 3646
rect 1261 3776 1414 3840
rect 2252 3814 2589 3874
rect 2975 3872 3197 3920
rect 2975 3868 2985 3872
rect 2865 3824 2948 3840
rect 1261 3742 1267 3776
rect 1344 3742 1414 3776
rect 797 3570 1107 3598
rect 1261 3584 1414 3742
rect 2111 3778 2745 3814
rect 2111 3772 2746 3778
rect 2111 3692 2124 3772
rect 2158 3692 2316 3772
rect 2350 3692 2508 3772
rect 2542 3692 2700 3772
rect 2734 3692 2746 3772
rect 2111 3686 2746 3692
rect 2111 3685 2745 3686
rect 2865 3656 2898 3824
rect 363 3564 1107 3570
rect -703 3515 -427 3550
rect 235 3517 399 3535
rect 235 3515 349 3517
rect -703 3422 -364 3515
rect -703 3388 -691 3422
rect -515 3388 -364 3422
rect 235 3405 260 3515
rect 383 3482 399 3517
rect 355 3405 399 3482
rect 235 3400 399 3405
rect 427 3517 687 3536
rect 427 3482 638 3517
rect 672 3482 687 3517
rect 427 3462 687 3482
rect -703 3382 -503 3388
rect -2544 3299 -2344 3300
rect -2548 3252 -2340 3299
rect -3544 3218 -3506 3244
rect -3542 3066 -3506 3218
rect -3384 3235 -3205 3244
rect -3384 3066 -3354 3235
rect -3177 3230 -2777 3236
rect -3177 3196 -3165 3230
rect -2789 3196 -2777 3230
rect -3177 3155 -2777 3196
rect -3177 3086 -3150 3155
rect -2815 3086 -2777 3155
rect -3177 3067 -2777 3086
rect -1748 3235 -1364 3358
rect -817 3378 -734 3382
rect -817 3344 -784 3378
rect -750 3344 -734 3378
rect -817 3327 -734 3344
rect -703 3334 -503 3341
rect -703 3300 -691 3334
rect -515 3300 -503 3334
rect -475 3327 -364 3388
rect 427 3393 477 3462
rect 763 3434 1107 3564
rect 427 3371 433 3393
rect 100 3358 433 3371
rect 467 3358 477 3393
rect 505 3422 1107 3434
rect 505 3388 517 3422
rect 893 3388 1107 3422
rect 505 3382 1107 3388
rect 1138 3550 1267 3584
rect 1344 3550 1414 3584
rect 2204 3650 2898 3656
rect 2204 3570 2220 3650
rect 2254 3570 2412 3650
rect 2446 3570 2604 3650
rect 2638 3598 2898 3650
rect 2932 3598 2948 3824
rect 2979 3838 2985 3868
rect 3064 3868 3197 3872
rect 3064 3838 3070 3868
rect 2979 3680 3070 3838
rect 2979 3646 2985 3680
rect 3064 3646 3070 3680
rect 2979 3630 3070 3646
rect 3102 3776 3255 3840
rect 3102 3742 3108 3776
rect 3185 3742 3255 3776
rect 2638 3570 2948 3598
rect 3102 3584 3255 3742
rect 2204 3564 2948 3570
rect 1138 3515 1414 3550
rect 2076 3517 2240 3535
rect 2076 3515 2190 3517
rect 1138 3422 1477 3515
rect 1138 3388 1150 3422
rect 1326 3388 1477 3422
rect 2076 3405 2101 3515
rect 2224 3482 2240 3517
rect 2196 3405 2240 3482
rect 2076 3400 2240 3405
rect 2268 3517 2528 3536
rect 2268 3482 2479 3517
rect 2513 3482 2528 3517
rect 2268 3462 2528 3482
rect 1138 3382 1338 3388
rect -703 3299 -503 3300
rect -707 3252 -499 3299
rect -1748 3215 -1549 3235
rect -3542 3044 -3354 3066
rect -1748 3043 -1722 3215
rect -1584 3043 -1549 3215
rect -1336 3230 -936 3236
rect -1336 3196 -1324 3230
rect -948 3196 -936 3230
rect -1336 3155 -936 3196
rect -1336 3086 -1309 3155
rect -974 3086 -936 3155
rect -1336 3067 -936 3086
rect 100 3235 477 3358
rect 1024 3378 1107 3382
rect 1024 3344 1057 3378
rect 1091 3344 1107 3378
rect 1024 3327 1107 3344
rect 1138 3334 1338 3341
rect 1138 3300 1150 3334
rect 1326 3300 1338 3334
rect 1366 3327 1477 3388
rect 2268 3393 2318 3462
rect 2604 3434 2948 3564
rect 2268 3371 2274 3393
rect 2001 3358 2274 3371
rect 2308 3358 2318 3393
rect 2346 3422 2948 3434
rect 2346 3388 2358 3422
rect 2734 3388 2948 3422
rect 2346 3382 2948 3388
rect 2979 3550 3108 3584
rect 3185 3550 3255 3584
rect 2979 3515 3255 3550
rect 2979 3422 3318 3515
rect 2979 3388 2991 3422
rect 3167 3388 3318 3422
rect 2979 3382 3179 3388
rect 2001 3323 2318 3358
rect 2865 3378 2948 3382
rect 2865 3344 2898 3378
rect 2932 3344 2948 3378
rect 2865 3327 2948 3344
rect 2979 3334 3179 3341
rect 1138 3299 1338 3300
rect 1134 3252 1342 3299
rect 1752 3297 2318 3323
rect 2979 3300 2991 3334
rect 3167 3300 3179 3334
rect 3207 3327 3318 3388
rect 2979 3299 3179 3300
rect 100 3189 320 3235
rect 100 3066 127 3189
rect 303 3066 320 3189
rect 505 3230 905 3236
rect 505 3196 517 3230
rect 893 3196 905 3230
rect 505 3155 905 3196
rect 505 3086 532 3155
rect 867 3086 905 3155
rect 1752 3144 1803 3297
rect 2001 3235 2318 3297
rect 2975 3252 3183 3299
rect 2001 3144 2150 3235
rect 1752 3116 2150 3144
rect 2346 3230 2746 3236
rect 2346 3196 2358 3230
rect 2734 3196 2746 3230
rect 2346 3155 2746 3196
rect 505 3067 905 3086
rect 2346 3086 2373 3155
rect 2708 3086 2746 3155
rect 2346 3067 2746 3086
rect 100 3045 320 3066
rect -1748 3013 -1549 3043
rect -2226 2840 -3 2924
rect -3817 2215 -3534 2234
rect -3818 2167 -3534 2215
rect -3818 1894 -3763 2167
rect -3574 1894 -3534 2167
rect -3247 2149 -2910 2161
rect -3247 2102 -3173 2149
rect -2933 2102 -2910 2149
rect -3247 2042 -2910 2102
rect -2524 2100 -2302 2148
rect -2524 2096 -2514 2100
rect -2634 2052 -2551 2068
rect -3388 2006 -2754 2042
rect -3388 2000 -2753 2006
rect -3388 1920 -3375 2000
rect -3341 1920 -3183 2000
rect -3149 1920 -2991 2000
rect -2957 1920 -2799 2000
rect -2765 1920 -2753 2000
rect -3388 1914 -2753 1920
rect -3388 1913 -2754 1914
rect -3818 1852 -3534 1894
rect -2634 1884 -2601 2052
rect -3295 1878 -2601 1884
rect -3818 1763 -3652 1852
rect -3295 1798 -3279 1878
rect -3245 1798 -3087 1878
rect -3053 1798 -2895 1878
rect -2861 1826 -2601 1878
rect -2567 1826 -2551 2052
rect -2520 2066 -2514 2096
rect -2435 2096 -2302 2100
rect -2435 2066 -2429 2096
rect -2226 2068 -2113 2840
rect -2520 1908 -2429 2066
rect -2520 1874 -2514 1908
rect -2435 1874 -2429 1908
rect -2520 1858 -2429 1874
rect -2397 2004 -2113 2068
rect -2397 1970 -2391 2004
rect -2314 1970 -2113 2004
rect -2397 1938 -2113 1970
rect -2044 2693 -3 2777
rect -2861 1798 -2551 1826
rect -2397 1812 -2244 1938
rect -3295 1792 -2551 1798
rect -3818 1745 -3259 1763
rect -3818 1710 -3309 1745
rect -3275 1710 -3259 1745
rect -3818 1628 -3259 1710
rect -3231 1745 -2971 1764
rect -3231 1710 -3020 1745
rect -2986 1710 -2971 1745
rect -3231 1690 -2971 1710
rect -3818 -1502 -3652 1628
rect -3231 1621 -3181 1690
rect -2895 1662 -2551 1792
rect -3231 1599 -3225 1621
rect -3423 1586 -3225 1599
rect -3191 1586 -3181 1621
rect -3153 1650 -2551 1662
rect -3153 1616 -3141 1650
rect -2765 1616 -2551 1650
rect -3153 1610 -2551 1616
rect -2520 1778 -2391 1812
rect -2314 1778 -2244 1812
rect -2520 1650 -2244 1778
rect -2520 1616 -2508 1650
rect -2332 1616 -2244 1650
rect -2520 1610 -2320 1616
rect -3423 1578 -3181 1586
rect -3423 1477 -3392 1578
rect -3260 1477 -3181 1578
rect -2634 1606 -2551 1610
rect -2634 1572 -2601 1606
rect -2567 1572 -2551 1606
rect -2634 1555 -2551 1572
rect -2520 1562 -2320 1569
rect -2520 1528 -2508 1562
rect -2332 1528 -2320 1562
rect -2292 1555 -2244 1616
rect -2520 1527 -2320 1528
rect -2524 1480 -2316 1527
rect -3423 1463 -3181 1477
rect -3153 1458 -2753 1464
rect -3153 1424 -3141 1458
rect -2765 1424 -2753 1458
rect -3153 1383 -2753 1424
rect -3153 1314 -3126 1383
rect -2791 1314 -2753 1383
rect -3153 1295 -2753 1314
rect -3247 857 -2910 869
rect -3247 810 -3173 857
rect -2933 810 -2910 857
rect -3247 750 -2910 810
rect -2524 808 -2302 856
rect -2524 804 -2514 808
rect -2634 760 -2551 776
rect -3388 714 -2754 750
rect -3388 708 -2753 714
rect -3388 628 -3375 708
rect -3341 628 -3183 708
rect -3149 628 -2991 708
rect -2957 628 -2799 708
rect -2765 628 -2753 708
rect -3388 622 -2753 628
rect -3388 621 -2754 622
rect -2634 592 -2601 760
rect -3295 586 -2601 592
rect -3295 506 -3279 586
rect -3245 506 -3087 586
rect -3053 506 -2895 586
rect -2861 534 -2601 586
rect -2567 534 -2551 760
rect -2520 774 -2514 804
rect -2435 804 -2302 808
rect -2435 774 -2429 804
rect -2520 616 -2429 774
rect -2520 582 -2514 616
rect -2435 582 -2429 616
rect -2520 566 -2429 582
rect -2397 712 -2244 776
rect -2397 678 -2391 712
rect -2314 678 -2244 712
rect -2861 506 -2551 534
rect -2397 520 -2244 678
rect -3295 500 -2551 506
rect -3423 453 -3259 471
rect -3423 451 -3309 453
rect -3423 341 -3398 451
rect -3275 418 -3259 453
rect -3303 341 -3259 418
rect -3423 336 -3259 341
rect -3231 453 -2971 472
rect -3231 418 -3020 453
rect -2986 418 -2971 453
rect -3231 398 -2971 418
rect -3231 329 -3181 398
rect -2895 370 -2551 500
rect -3231 307 -3225 329
rect -3593 294 -3225 307
rect -3191 294 -3181 329
rect -3153 358 -2551 370
rect -3153 324 -3141 358
rect -2765 324 -2551 358
rect -3153 318 -2551 324
rect -2520 486 -2391 520
rect -2314 486 -2244 520
rect -2520 451 -2244 486
rect -2044 451 -1907 2693
rect -215 2545 -3 2629
rect -1521 2149 -1184 2161
rect -1521 2102 -1447 2149
rect -1207 2102 -1184 2149
rect -1521 2042 -1184 2102
rect -798 2100 -576 2148
rect -798 2096 -788 2100
rect -908 2052 -825 2068
rect -1662 2006 -1028 2042
rect -1662 2000 -1027 2006
rect -1662 1920 -1649 2000
rect -1615 1920 -1457 2000
rect -1423 1920 -1265 2000
rect -1231 1920 -1073 2000
rect -1039 1920 -1027 2000
rect -1662 1914 -1027 1920
rect -1662 1913 -1028 1914
rect -908 1884 -875 2052
rect -1569 1878 -875 1884
rect -1569 1798 -1553 1878
rect -1519 1798 -1361 1878
rect -1327 1798 -1169 1878
rect -1135 1826 -875 1878
rect -841 1826 -825 2052
rect -794 2066 -788 2096
rect -709 2096 -576 2100
rect -709 2066 -703 2096
rect -794 1908 -703 2066
rect -794 1874 -788 1908
rect -709 1874 -703 1908
rect -794 1858 -703 1874
rect -671 2004 -518 2068
rect -671 1970 -665 2004
rect -588 1970 -518 2004
rect -1135 1798 -825 1826
rect -671 1812 -518 1970
rect -1569 1792 -825 1798
rect -1697 1745 -1533 1763
rect -1697 1735 -1583 1745
rect -1697 1658 -1676 1735
rect -1549 1710 -1533 1745
rect -1571 1658 -1533 1710
rect -1697 1628 -1533 1658
rect -1505 1745 -1245 1764
rect -1505 1710 -1294 1745
rect -1260 1710 -1245 1745
rect -1505 1690 -1245 1710
rect -1505 1621 -1455 1690
rect -1169 1662 -825 1792
rect -1505 1599 -1499 1621
rect -1697 1586 -1499 1599
rect -1465 1586 -1455 1621
rect -1427 1650 -825 1662
rect -1427 1616 -1415 1650
rect -1039 1616 -825 1650
rect -1427 1610 -825 1616
rect -794 1778 -665 1812
rect -588 1778 -518 1812
rect -794 1702 -518 1778
rect -215 1702 -84 2545
rect -794 1650 -84 1702
rect -794 1616 -782 1650
rect -606 1616 -84 1650
rect -794 1610 -594 1616
rect -1697 1584 -1455 1586
rect -1697 1480 -1681 1584
rect -1564 1480 -1455 1584
rect -908 1606 -825 1610
rect -908 1572 -875 1606
rect -841 1572 -825 1606
rect -908 1555 -825 1572
rect -794 1562 -594 1569
rect -794 1528 -782 1562
rect -606 1528 -594 1562
rect -566 1555 -84 1616
rect -794 1527 -594 1528
rect -798 1480 -590 1527
rect -1697 1463 -1455 1480
rect -1427 1458 -1027 1464
rect -1427 1424 -1415 1458
rect -1039 1424 -1027 1458
rect -1427 1383 -1027 1424
rect -1427 1314 -1400 1383
rect -1065 1314 -1027 1383
rect -1427 1295 -1027 1314
rect -1521 857 -1184 869
rect -1521 810 -1447 857
rect -1207 810 -1184 857
rect -1521 750 -1184 810
rect -798 808 -576 856
rect -798 804 -788 808
rect -908 760 -825 776
rect -1662 714 -1028 750
rect -1662 708 -1027 714
rect -1662 628 -1649 708
rect -1615 628 -1457 708
rect -1423 628 -1265 708
rect -1231 628 -1073 708
rect -1039 628 -1027 708
rect -1662 622 -1027 628
rect -1662 621 -1028 622
rect -908 592 -875 760
rect -1569 586 -875 592
rect -1569 506 -1553 586
rect -1519 506 -1361 586
rect -1327 506 -1169 586
rect -1135 534 -875 586
rect -841 534 -825 760
rect -794 774 -788 804
rect -709 804 -576 808
rect -709 774 -703 804
rect -794 616 -703 774
rect -794 582 -788 616
rect -709 582 -703 616
rect -794 566 -703 582
rect -671 712 -518 776
rect -671 678 -665 712
rect -588 678 -518 712
rect -1135 506 -825 534
rect -671 528 -518 678
rect -671 526 -433 528
rect -671 520 -262 526
rect -1569 500 -825 506
rect -2520 358 -1907 451
rect -2520 324 -2508 358
rect -2332 324 -1907 358
rect -1697 453 -1533 471
rect -1697 351 -1682 453
rect -1606 418 -1583 453
rect -1549 418 -1533 453
rect -1606 351 -1533 418
rect -1697 336 -1533 351
rect -1505 453 -1245 472
rect -1505 418 -1294 453
rect -1260 418 -1245 453
rect -1505 398 -1245 418
rect -2520 318 -2320 324
rect -3593 182 -3181 294
rect -2634 314 -2551 318
rect -2634 280 -2601 314
rect -2567 280 -2551 314
rect -2634 263 -2551 280
rect -2520 270 -2320 277
rect -2520 236 -2508 270
rect -2332 236 -2320 270
rect -2292 265 -1907 324
rect -1505 329 -1455 398
rect -1169 370 -825 500
rect -1505 307 -1499 329
rect -1697 294 -1499 307
rect -1465 294 -1455 329
rect -1427 358 -825 370
rect -1427 324 -1415 358
rect -1039 324 -825 358
rect -1427 318 -825 324
rect -794 486 -665 520
rect -588 486 -262 520
rect -794 480 -262 486
rect -794 358 -521 480
rect -794 324 -782 358
rect -606 324 -521 358
rect -794 318 -594 324
rect -1697 286 -1455 294
rect -2292 263 -1968 265
rect -2520 235 -2320 236
rect -2524 188 -2316 235
rect -1697 197 -1680 286
rect -1553 197 -1455 286
rect -908 314 -825 318
rect -908 280 -875 314
rect -841 280 -825 314
rect -908 263 -825 280
rect -566 298 -521 324
rect -311 298 -262 480
rect -794 270 -594 277
rect -794 236 -782 270
rect -606 236 -594 270
rect -566 263 -262 298
rect -794 235 -594 236
rect -3593 -16 -3568 182
rect -3422 171 -3181 182
rect -3422 -16 -3332 171
rect -3153 166 -2753 172
rect -1697 171 -1455 197
rect -798 188 -590 235
rect -3153 132 -3141 166
rect -2765 132 -2753 166
rect -3153 91 -2753 132
rect -3153 22 -3126 91
rect -2791 22 -2753 91
rect -3153 3 -2753 22
rect -1427 166 -1027 172
rect -1427 132 -1415 166
rect -1039 132 -1027 166
rect -1427 91 -1027 132
rect -1427 22 -1400 91
rect -1065 22 -1027 91
rect -1427 3 -1027 22
rect -3593 -31 -3332 -16
rect -2226 -425 -3 -341
rect -3247 -1116 -2910 -1104
rect -3247 -1163 -3173 -1116
rect -2933 -1163 -2910 -1116
rect -3247 -1223 -2910 -1163
rect -2524 -1165 -2302 -1117
rect -2524 -1169 -2514 -1165
rect -2634 -1213 -2551 -1197
rect -3388 -1259 -2754 -1223
rect -3388 -1265 -2753 -1259
rect -3388 -1345 -3375 -1265
rect -3341 -1345 -3183 -1265
rect -3149 -1345 -2991 -1265
rect -2957 -1345 -2799 -1265
rect -2765 -1345 -2753 -1265
rect -3388 -1351 -2753 -1345
rect -3388 -1352 -2754 -1351
rect -2634 -1381 -2601 -1213
rect -3295 -1387 -2601 -1381
rect -3295 -1467 -3279 -1387
rect -3245 -1467 -3087 -1387
rect -3053 -1467 -2895 -1387
rect -2861 -1439 -2601 -1387
rect -2567 -1439 -2551 -1213
rect -2520 -1199 -2514 -1169
rect -2435 -1169 -2302 -1165
rect -2435 -1199 -2429 -1169
rect -2226 -1197 -2113 -425
rect -2520 -1357 -2429 -1199
rect -2520 -1391 -2514 -1357
rect -2435 -1391 -2429 -1357
rect -2520 -1407 -2429 -1391
rect -2397 -1261 -2113 -1197
rect -2397 -1295 -2391 -1261
rect -2314 -1295 -2113 -1261
rect -2397 -1327 -2113 -1295
rect -2044 -572 -3 -488
rect -2861 -1467 -2551 -1439
rect -2397 -1453 -2244 -1327
rect -3295 -1473 -2551 -1467
rect -3818 -1520 -3259 -1502
rect -3818 -1555 -3309 -1520
rect -3275 -1555 -3259 -1520
rect -3818 -1637 -3259 -1555
rect -3231 -1520 -2971 -1501
rect -3231 -1555 -3020 -1520
rect -2986 -1555 -2971 -1520
rect -3231 -1575 -2971 -1555
rect -3818 -4766 -3652 -1637
rect -3231 -1644 -3181 -1575
rect -2895 -1603 -2551 -1473
rect -3231 -1666 -3225 -1644
rect -3423 -1679 -3225 -1666
rect -3191 -1679 -3181 -1644
rect -3153 -1615 -2551 -1603
rect -3153 -1649 -3141 -1615
rect -2765 -1649 -2551 -1615
rect -3153 -1655 -2551 -1649
rect -2520 -1487 -2391 -1453
rect -2314 -1487 -2244 -1453
rect -2520 -1615 -2244 -1487
rect -2520 -1649 -2508 -1615
rect -2332 -1649 -2244 -1615
rect -2520 -1655 -2320 -1649
rect -3423 -1687 -3181 -1679
rect -3423 -1788 -3392 -1687
rect -3260 -1788 -3181 -1687
rect -2634 -1659 -2551 -1655
rect -2634 -1693 -2601 -1659
rect -2567 -1693 -2551 -1659
rect -2634 -1710 -2551 -1693
rect -2520 -1703 -2320 -1696
rect -2520 -1737 -2508 -1703
rect -2332 -1737 -2320 -1703
rect -2292 -1710 -2244 -1649
rect -2520 -1738 -2320 -1737
rect -2524 -1785 -2316 -1738
rect -3423 -1802 -3181 -1788
rect -3153 -1807 -2753 -1801
rect -3153 -1841 -3141 -1807
rect -2765 -1841 -2753 -1807
rect -3153 -1882 -2753 -1841
rect -3153 -1951 -3126 -1882
rect -2791 -1951 -2753 -1882
rect -3153 -1970 -2753 -1951
rect -3247 -2408 -2910 -2396
rect -3247 -2455 -3173 -2408
rect -2933 -2455 -2910 -2408
rect -3247 -2515 -2910 -2455
rect -2524 -2457 -2302 -2409
rect -2524 -2461 -2514 -2457
rect -2634 -2505 -2551 -2489
rect -3388 -2551 -2754 -2515
rect -3388 -2557 -2753 -2551
rect -3388 -2637 -3375 -2557
rect -3341 -2637 -3183 -2557
rect -3149 -2637 -2991 -2557
rect -2957 -2637 -2799 -2557
rect -2765 -2637 -2753 -2557
rect -3388 -2643 -2753 -2637
rect -3388 -2644 -2754 -2643
rect -2634 -2673 -2601 -2505
rect -3295 -2679 -2601 -2673
rect -3295 -2759 -3279 -2679
rect -3245 -2759 -3087 -2679
rect -3053 -2759 -2895 -2679
rect -2861 -2731 -2601 -2679
rect -2567 -2731 -2551 -2505
rect -2520 -2491 -2514 -2461
rect -2435 -2461 -2302 -2457
rect -2435 -2491 -2429 -2461
rect -2520 -2649 -2429 -2491
rect -2520 -2683 -2514 -2649
rect -2435 -2683 -2429 -2649
rect -2520 -2699 -2429 -2683
rect -2397 -2553 -2244 -2489
rect -2397 -2587 -2391 -2553
rect -2314 -2587 -2244 -2553
rect -2861 -2759 -2551 -2731
rect -2397 -2745 -2244 -2587
rect -3295 -2765 -2551 -2759
rect -3423 -2812 -3259 -2794
rect -3423 -2814 -3309 -2812
rect -3423 -2924 -3398 -2814
rect -3275 -2847 -3259 -2812
rect -3303 -2924 -3259 -2847
rect -3423 -2929 -3259 -2924
rect -3231 -2812 -2971 -2793
rect -3231 -2847 -3020 -2812
rect -2986 -2847 -2971 -2812
rect -3231 -2867 -2971 -2847
rect -3231 -2936 -3181 -2867
rect -2895 -2895 -2551 -2765
rect -3231 -2958 -3225 -2936
rect -3593 -2971 -3225 -2958
rect -3191 -2971 -3181 -2936
rect -3153 -2907 -2551 -2895
rect -3153 -2941 -3141 -2907
rect -2765 -2941 -2551 -2907
rect -3153 -2947 -2551 -2941
rect -2520 -2779 -2391 -2745
rect -2314 -2779 -2244 -2745
rect -2520 -2814 -2244 -2779
rect -2044 -2814 -1907 -572
rect -215 -720 -3 -636
rect -1521 -1116 -1184 -1104
rect -1521 -1163 -1447 -1116
rect -1207 -1163 -1184 -1116
rect -1521 -1223 -1184 -1163
rect -798 -1165 -576 -1117
rect -798 -1169 -788 -1165
rect -908 -1213 -825 -1197
rect -1662 -1259 -1028 -1223
rect -1662 -1265 -1027 -1259
rect -1662 -1345 -1649 -1265
rect -1615 -1345 -1457 -1265
rect -1423 -1345 -1265 -1265
rect -1231 -1345 -1073 -1265
rect -1039 -1345 -1027 -1265
rect -1662 -1351 -1027 -1345
rect -1662 -1352 -1028 -1351
rect -908 -1381 -875 -1213
rect -1569 -1387 -875 -1381
rect -1569 -1467 -1553 -1387
rect -1519 -1467 -1361 -1387
rect -1327 -1467 -1169 -1387
rect -1135 -1439 -875 -1387
rect -841 -1439 -825 -1213
rect -794 -1199 -788 -1169
rect -709 -1169 -576 -1165
rect -709 -1199 -703 -1169
rect -794 -1357 -703 -1199
rect -794 -1391 -788 -1357
rect -709 -1391 -703 -1357
rect -794 -1407 -703 -1391
rect -671 -1261 -518 -1197
rect -671 -1295 -665 -1261
rect -588 -1295 -518 -1261
rect -1135 -1467 -825 -1439
rect -671 -1453 -518 -1295
rect -1569 -1473 -825 -1467
rect -1697 -1520 -1533 -1502
rect -1697 -1530 -1583 -1520
rect -1697 -1607 -1676 -1530
rect -1549 -1555 -1533 -1520
rect -1571 -1607 -1533 -1555
rect -1697 -1637 -1533 -1607
rect -1505 -1520 -1245 -1501
rect -1505 -1555 -1294 -1520
rect -1260 -1555 -1245 -1520
rect -1505 -1575 -1245 -1555
rect -1505 -1644 -1455 -1575
rect -1169 -1603 -825 -1473
rect -1505 -1666 -1499 -1644
rect -1697 -1679 -1499 -1666
rect -1465 -1679 -1455 -1644
rect -1427 -1615 -825 -1603
rect -1427 -1649 -1415 -1615
rect -1039 -1649 -825 -1615
rect -1427 -1655 -825 -1649
rect -794 -1487 -665 -1453
rect -588 -1487 -518 -1453
rect -794 -1563 -518 -1487
rect -215 -1563 -84 -720
rect -794 -1615 -84 -1563
rect -794 -1649 -782 -1615
rect -606 -1649 -84 -1615
rect -794 -1655 -594 -1649
rect -1697 -1681 -1455 -1679
rect -1697 -1785 -1681 -1681
rect -1564 -1785 -1455 -1681
rect -908 -1659 -825 -1655
rect -908 -1693 -875 -1659
rect -841 -1693 -825 -1659
rect -908 -1710 -825 -1693
rect -794 -1703 -594 -1696
rect -794 -1737 -782 -1703
rect -606 -1737 -594 -1703
rect -566 -1710 -84 -1649
rect -794 -1738 -594 -1737
rect -798 -1785 -590 -1738
rect -1697 -1802 -1455 -1785
rect -1427 -1807 -1027 -1801
rect -1427 -1841 -1415 -1807
rect -1039 -1841 -1027 -1807
rect -1427 -1882 -1027 -1841
rect -1427 -1951 -1400 -1882
rect -1065 -1951 -1027 -1882
rect -1427 -1970 -1027 -1951
rect -1521 -2408 -1184 -2396
rect -1521 -2455 -1447 -2408
rect -1207 -2455 -1184 -2408
rect -1521 -2515 -1184 -2455
rect -798 -2457 -576 -2409
rect -798 -2461 -788 -2457
rect -908 -2505 -825 -2489
rect -1662 -2551 -1028 -2515
rect -1662 -2557 -1027 -2551
rect -1662 -2637 -1649 -2557
rect -1615 -2637 -1457 -2557
rect -1423 -2637 -1265 -2557
rect -1231 -2637 -1073 -2557
rect -1039 -2637 -1027 -2557
rect -1662 -2643 -1027 -2637
rect -1662 -2644 -1028 -2643
rect -908 -2673 -875 -2505
rect -1569 -2679 -875 -2673
rect -1569 -2759 -1553 -2679
rect -1519 -2759 -1361 -2679
rect -1327 -2759 -1169 -2679
rect -1135 -2731 -875 -2679
rect -841 -2731 -825 -2505
rect -794 -2491 -788 -2461
rect -709 -2461 -576 -2457
rect -709 -2491 -703 -2461
rect -794 -2649 -703 -2491
rect -794 -2683 -788 -2649
rect -709 -2683 -703 -2649
rect -794 -2699 -703 -2683
rect -671 -2553 -518 -2489
rect -671 -2587 -665 -2553
rect -588 -2587 -518 -2553
rect -1135 -2759 -825 -2731
rect -671 -2737 -518 -2587
rect -671 -2739 -433 -2737
rect -671 -2745 -262 -2739
rect -1569 -2765 -825 -2759
rect -2520 -2907 -1907 -2814
rect -2520 -2941 -2508 -2907
rect -2332 -2941 -1907 -2907
rect -1697 -2812 -1533 -2794
rect -1697 -2914 -1682 -2812
rect -1606 -2847 -1583 -2812
rect -1549 -2847 -1533 -2812
rect -1606 -2914 -1533 -2847
rect -1697 -2929 -1533 -2914
rect -1505 -2812 -1245 -2793
rect -1505 -2847 -1294 -2812
rect -1260 -2847 -1245 -2812
rect -1505 -2867 -1245 -2847
rect -2520 -2947 -2320 -2941
rect -3593 -3083 -3181 -2971
rect -2634 -2951 -2551 -2947
rect -2634 -2985 -2601 -2951
rect -2567 -2985 -2551 -2951
rect -2634 -3002 -2551 -2985
rect -2520 -2995 -2320 -2988
rect -2520 -3029 -2508 -2995
rect -2332 -3029 -2320 -2995
rect -2292 -3000 -1907 -2941
rect -1505 -2936 -1455 -2867
rect -1169 -2895 -825 -2765
rect -1505 -2958 -1499 -2936
rect -1697 -2971 -1499 -2958
rect -1465 -2971 -1455 -2936
rect -1427 -2907 -825 -2895
rect -1427 -2941 -1415 -2907
rect -1039 -2941 -825 -2907
rect -1427 -2947 -825 -2941
rect -794 -2779 -665 -2745
rect -588 -2779 -262 -2745
rect -794 -2785 -262 -2779
rect -794 -2907 -521 -2785
rect -794 -2941 -782 -2907
rect -606 -2941 -521 -2907
rect -794 -2947 -594 -2941
rect -1697 -2979 -1455 -2971
rect -2292 -3002 -1968 -3000
rect -2520 -3030 -2320 -3029
rect -2524 -3077 -2316 -3030
rect -1697 -3068 -1680 -2979
rect -1553 -3068 -1455 -2979
rect -908 -2951 -825 -2947
rect -908 -2985 -875 -2951
rect -841 -2985 -825 -2951
rect -908 -3002 -825 -2985
rect -566 -2967 -521 -2941
rect -311 -2967 -262 -2785
rect -794 -2995 -594 -2988
rect -794 -3029 -782 -2995
rect -606 -3029 -594 -2995
rect -566 -3002 -262 -2967
rect -794 -3030 -594 -3029
rect -3593 -3281 -3568 -3083
rect -3422 -3094 -3181 -3083
rect -3422 -3281 -3332 -3094
rect -3153 -3099 -2753 -3093
rect -1697 -3094 -1455 -3068
rect -798 -3077 -590 -3030
rect -3153 -3133 -3141 -3099
rect -2765 -3133 -2753 -3099
rect -3153 -3174 -2753 -3133
rect -3153 -3243 -3126 -3174
rect -2791 -3243 -2753 -3174
rect -3153 -3262 -2753 -3243
rect -1427 -3099 -1027 -3093
rect -1427 -3133 -1415 -3099
rect -1039 -3133 -1027 -3099
rect -1427 -3174 -1027 -3133
rect -1427 -3243 -1400 -3174
rect -1065 -3243 -1027 -3174
rect -1427 -3262 -1027 -3243
rect -3593 -3296 -3332 -3281
rect -2226 -3689 -3 -3605
rect -3247 -4380 -2910 -4368
rect -3247 -4427 -3173 -4380
rect -2933 -4427 -2910 -4380
rect -3247 -4487 -2910 -4427
rect -2524 -4429 -2302 -4381
rect -2524 -4433 -2514 -4429
rect -2634 -4477 -2551 -4461
rect -3388 -4523 -2754 -4487
rect -3388 -4529 -2753 -4523
rect -3388 -4609 -3375 -4529
rect -3341 -4609 -3183 -4529
rect -3149 -4609 -2991 -4529
rect -2957 -4609 -2799 -4529
rect -2765 -4609 -2753 -4529
rect -3388 -4615 -2753 -4609
rect -3388 -4616 -2754 -4615
rect -2634 -4645 -2601 -4477
rect -3295 -4651 -2601 -4645
rect -3295 -4731 -3279 -4651
rect -3245 -4731 -3087 -4651
rect -3053 -4731 -2895 -4651
rect -2861 -4703 -2601 -4651
rect -2567 -4703 -2551 -4477
rect -2520 -4463 -2514 -4433
rect -2435 -4433 -2302 -4429
rect -2435 -4463 -2429 -4433
rect -2226 -4461 -2113 -3689
rect -2520 -4621 -2429 -4463
rect -2520 -4655 -2514 -4621
rect -2435 -4655 -2429 -4621
rect -2520 -4671 -2429 -4655
rect -2397 -4525 -2113 -4461
rect -2397 -4559 -2391 -4525
rect -2314 -4559 -2113 -4525
rect -2397 -4591 -2113 -4559
rect -2044 -3836 -3 -3752
rect -2861 -4731 -2551 -4703
rect -2397 -4717 -2244 -4591
rect -3295 -4737 -2551 -4731
rect -3818 -4784 -3259 -4766
rect -3818 -4819 -3309 -4784
rect -3275 -4819 -3259 -4784
rect -3818 -4901 -3259 -4819
rect -3231 -4784 -2971 -4765
rect -3231 -4819 -3020 -4784
rect -2986 -4819 -2971 -4784
rect -3231 -4839 -2971 -4819
rect -3231 -4908 -3181 -4839
rect -2895 -4867 -2551 -4737
rect -3231 -4930 -3225 -4908
rect -3423 -4943 -3225 -4930
rect -3191 -4943 -3181 -4908
rect -3153 -4879 -2551 -4867
rect -3153 -4913 -3141 -4879
rect -2765 -4913 -2551 -4879
rect -3153 -4919 -2551 -4913
rect -2520 -4751 -2391 -4717
rect -2314 -4751 -2244 -4717
rect -2520 -4879 -2244 -4751
rect -2520 -4913 -2508 -4879
rect -2332 -4913 -2244 -4879
rect -2520 -4919 -2320 -4913
rect -3423 -4951 -3181 -4943
rect -3423 -5052 -3392 -4951
rect -3260 -5052 -3181 -4951
rect -2634 -4923 -2551 -4919
rect -2634 -4957 -2601 -4923
rect -2567 -4957 -2551 -4923
rect -2634 -4974 -2551 -4957
rect -2520 -4967 -2320 -4960
rect -2520 -5001 -2508 -4967
rect -2332 -5001 -2320 -4967
rect -2292 -4974 -2244 -4913
rect -2520 -5002 -2320 -5001
rect -2524 -5049 -2316 -5002
rect -3423 -5066 -3181 -5052
rect -3153 -5071 -2753 -5065
rect -3153 -5105 -3141 -5071
rect -2765 -5105 -2753 -5071
rect -3153 -5146 -2753 -5105
rect -3153 -5215 -3126 -5146
rect -2791 -5215 -2753 -5146
rect -3153 -5234 -2753 -5215
rect -3247 -5672 -2910 -5660
rect -3247 -5719 -3173 -5672
rect -2933 -5719 -2910 -5672
rect -3247 -5779 -2910 -5719
rect -2524 -5721 -2302 -5673
rect -2524 -5725 -2514 -5721
rect -2634 -5769 -2551 -5753
rect -3388 -5815 -2754 -5779
rect -3388 -5821 -2753 -5815
rect -3388 -5901 -3375 -5821
rect -3341 -5901 -3183 -5821
rect -3149 -5901 -2991 -5821
rect -2957 -5901 -2799 -5821
rect -2765 -5901 -2753 -5821
rect -3388 -5907 -2753 -5901
rect -3388 -5908 -2754 -5907
rect -2634 -5937 -2601 -5769
rect -3295 -5943 -2601 -5937
rect -3295 -6023 -3279 -5943
rect -3245 -6023 -3087 -5943
rect -3053 -6023 -2895 -5943
rect -2861 -5995 -2601 -5943
rect -2567 -5995 -2551 -5769
rect -2520 -5755 -2514 -5725
rect -2435 -5725 -2302 -5721
rect -2435 -5755 -2429 -5725
rect -2520 -5913 -2429 -5755
rect -2520 -5947 -2514 -5913
rect -2435 -5947 -2429 -5913
rect -2520 -5963 -2429 -5947
rect -2397 -5817 -2244 -5753
rect -2397 -5851 -2391 -5817
rect -2314 -5851 -2244 -5817
rect -2861 -6023 -2551 -5995
rect -2397 -6009 -2244 -5851
rect -3295 -6029 -2551 -6023
rect -3423 -6076 -3259 -6058
rect -3423 -6078 -3309 -6076
rect -3423 -6188 -3398 -6078
rect -3275 -6111 -3259 -6076
rect -3303 -6188 -3259 -6111
rect -3423 -6193 -3259 -6188
rect -3231 -6076 -2971 -6057
rect -3231 -6111 -3020 -6076
rect -2986 -6111 -2971 -6076
rect -3231 -6131 -2971 -6111
rect -3231 -6200 -3181 -6131
rect -2895 -6159 -2551 -6029
rect -3231 -6222 -3225 -6200
rect -3593 -6235 -3225 -6222
rect -3191 -6235 -3181 -6200
rect -3153 -6171 -2551 -6159
rect -3153 -6205 -3141 -6171
rect -2765 -6205 -2551 -6171
rect -3153 -6211 -2551 -6205
rect -2520 -6043 -2391 -6009
rect -2314 -6043 -2244 -6009
rect -2520 -6078 -2244 -6043
rect -2044 -6078 -1907 -3836
rect -215 -3984 -3 -3900
rect -1521 -4380 -1184 -4368
rect -1521 -4427 -1447 -4380
rect -1207 -4427 -1184 -4380
rect -1521 -4487 -1184 -4427
rect -798 -4429 -576 -4381
rect -798 -4433 -788 -4429
rect -908 -4477 -825 -4461
rect -1662 -4523 -1028 -4487
rect -1662 -4529 -1027 -4523
rect -1662 -4609 -1649 -4529
rect -1615 -4609 -1457 -4529
rect -1423 -4609 -1265 -4529
rect -1231 -4609 -1073 -4529
rect -1039 -4609 -1027 -4529
rect -1662 -4615 -1027 -4609
rect -1662 -4616 -1028 -4615
rect -908 -4645 -875 -4477
rect -1569 -4651 -875 -4645
rect -1569 -4731 -1553 -4651
rect -1519 -4731 -1361 -4651
rect -1327 -4731 -1169 -4651
rect -1135 -4703 -875 -4651
rect -841 -4703 -825 -4477
rect -794 -4463 -788 -4433
rect -709 -4433 -576 -4429
rect -709 -4463 -703 -4433
rect -794 -4621 -703 -4463
rect -794 -4655 -788 -4621
rect -709 -4655 -703 -4621
rect -794 -4671 -703 -4655
rect -671 -4525 -518 -4461
rect -671 -4559 -665 -4525
rect -588 -4559 -518 -4525
rect -1135 -4731 -825 -4703
rect -671 -4717 -518 -4559
rect -1569 -4737 -825 -4731
rect -1697 -4784 -1533 -4766
rect -1697 -4794 -1583 -4784
rect -1697 -4871 -1676 -4794
rect -1549 -4819 -1533 -4784
rect -1571 -4871 -1533 -4819
rect -1697 -4901 -1533 -4871
rect -1505 -4784 -1245 -4765
rect -1505 -4819 -1294 -4784
rect -1260 -4819 -1245 -4784
rect -1505 -4839 -1245 -4819
rect -1505 -4908 -1455 -4839
rect -1169 -4867 -825 -4737
rect -1505 -4930 -1499 -4908
rect -1697 -4943 -1499 -4930
rect -1465 -4943 -1455 -4908
rect -1427 -4879 -825 -4867
rect -1427 -4913 -1415 -4879
rect -1039 -4913 -825 -4879
rect -1427 -4919 -825 -4913
rect -794 -4751 -665 -4717
rect -588 -4751 -518 -4717
rect -794 -4827 -518 -4751
rect -215 -4827 -84 -3984
rect -794 -4879 -84 -4827
rect -794 -4913 -782 -4879
rect -606 -4913 -84 -4879
rect -794 -4919 -594 -4913
rect -1697 -4945 -1455 -4943
rect -1697 -5049 -1681 -4945
rect -1564 -5049 -1455 -4945
rect -908 -4923 -825 -4919
rect -908 -4957 -875 -4923
rect -841 -4957 -825 -4923
rect -908 -4974 -825 -4957
rect -794 -4967 -594 -4960
rect -794 -5001 -782 -4967
rect -606 -5001 -594 -4967
rect -566 -4974 -84 -4913
rect -794 -5002 -594 -5001
rect -798 -5049 -590 -5002
rect -1697 -5066 -1455 -5049
rect -1427 -5071 -1027 -5065
rect -1427 -5105 -1415 -5071
rect -1039 -5105 -1027 -5071
rect -1427 -5146 -1027 -5105
rect -1427 -5215 -1400 -5146
rect -1065 -5215 -1027 -5146
rect -1427 -5234 -1027 -5215
rect -1521 -5672 -1184 -5660
rect -1521 -5719 -1447 -5672
rect -1207 -5719 -1184 -5672
rect -1521 -5779 -1184 -5719
rect -798 -5721 -576 -5673
rect -798 -5725 -788 -5721
rect -908 -5769 -825 -5753
rect -1662 -5815 -1028 -5779
rect -1662 -5821 -1027 -5815
rect -1662 -5901 -1649 -5821
rect -1615 -5901 -1457 -5821
rect -1423 -5901 -1265 -5821
rect -1231 -5901 -1073 -5821
rect -1039 -5901 -1027 -5821
rect -1662 -5907 -1027 -5901
rect -1662 -5908 -1028 -5907
rect -908 -5937 -875 -5769
rect -1569 -5943 -875 -5937
rect -1569 -6023 -1553 -5943
rect -1519 -6023 -1361 -5943
rect -1327 -6023 -1169 -5943
rect -1135 -5995 -875 -5943
rect -841 -5995 -825 -5769
rect -794 -5755 -788 -5725
rect -709 -5725 -576 -5721
rect -709 -5755 -703 -5725
rect -794 -5913 -703 -5755
rect -794 -5947 -788 -5913
rect -709 -5947 -703 -5913
rect -794 -5963 -703 -5947
rect -671 -5817 -518 -5753
rect -671 -5851 -665 -5817
rect -588 -5851 -518 -5817
rect -1135 -6023 -825 -5995
rect -671 -6001 -518 -5851
rect -671 -6003 -433 -6001
rect -671 -6009 -262 -6003
rect -1569 -6029 -825 -6023
rect -2520 -6171 -1907 -6078
rect -2520 -6205 -2508 -6171
rect -2332 -6205 -1907 -6171
rect -1697 -6076 -1533 -6058
rect -1697 -6178 -1682 -6076
rect -1606 -6111 -1583 -6076
rect -1549 -6111 -1533 -6076
rect -1606 -6178 -1533 -6111
rect -1697 -6193 -1533 -6178
rect -1505 -6076 -1245 -6057
rect -1505 -6111 -1294 -6076
rect -1260 -6111 -1245 -6076
rect -1505 -6131 -1245 -6111
rect -2520 -6211 -2320 -6205
rect -3593 -6347 -3181 -6235
rect -2634 -6215 -2551 -6211
rect -2634 -6249 -2601 -6215
rect -2567 -6249 -2551 -6215
rect -2634 -6266 -2551 -6249
rect -2520 -6259 -2320 -6252
rect -2520 -6293 -2508 -6259
rect -2332 -6293 -2320 -6259
rect -2292 -6264 -1907 -6205
rect -1505 -6200 -1455 -6131
rect -1169 -6159 -825 -6029
rect -1505 -6222 -1499 -6200
rect -1697 -6235 -1499 -6222
rect -1465 -6235 -1455 -6200
rect -1427 -6171 -825 -6159
rect -1427 -6205 -1415 -6171
rect -1039 -6205 -825 -6171
rect -1427 -6211 -825 -6205
rect -794 -6043 -665 -6009
rect -588 -6043 -262 -6009
rect -794 -6049 -262 -6043
rect -794 -6171 -521 -6049
rect -794 -6205 -782 -6171
rect -606 -6205 -521 -6171
rect -794 -6211 -594 -6205
rect -1697 -6243 -1455 -6235
rect -2292 -6266 -1968 -6264
rect -2520 -6294 -2320 -6293
rect -2524 -6341 -2316 -6294
rect -1697 -6332 -1680 -6243
rect -1553 -6332 -1455 -6243
rect -908 -6215 -825 -6211
rect -908 -6249 -875 -6215
rect -841 -6249 -825 -6215
rect -908 -6266 -825 -6249
rect -566 -6231 -521 -6205
rect -311 -6231 -262 -6049
rect -794 -6259 -594 -6252
rect -794 -6293 -782 -6259
rect -606 -6293 -594 -6259
rect -566 -6266 -262 -6231
rect -794 -6294 -594 -6293
rect -3593 -6545 -3568 -6347
rect -3422 -6358 -3181 -6347
rect -3422 -6545 -3332 -6358
rect -3153 -6363 -2753 -6357
rect -1697 -6358 -1455 -6332
rect -798 -6341 -590 -6294
rect -3153 -6397 -3141 -6363
rect -2765 -6397 -2753 -6363
rect -3153 -6438 -2753 -6397
rect -3153 -6507 -3126 -6438
rect -2791 -6507 -2753 -6438
rect -3153 -6526 -2753 -6507
rect -1427 -6363 -1027 -6357
rect -1427 -6397 -1415 -6363
rect -1039 -6397 -1027 -6363
rect -1427 -6438 -1027 -6397
rect -1427 -6507 -1400 -6438
rect -1065 -6507 -1027 -6438
rect -1427 -6526 -1027 -6507
rect -3593 -6560 -3332 -6545
<< via1 >>
rect -3422 3482 -3333 3515
rect -3333 3482 -3327 3515
rect -3422 3405 -3327 3482
rect -1581 3482 -1492 3515
rect -1492 3482 -1486 3515
rect -1581 3405 -1486 3482
rect 260 3482 349 3515
rect 349 3482 355 3515
rect 260 3405 355 3482
rect -3506 3066 -3384 3244
rect 2101 3482 2190 3515
rect 2190 3482 2196 3515
rect 2101 3405 2196 3482
rect -1722 3043 -1584 3215
rect 127 3066 303 3189
rect 1803 3144 2001 3297
rect -3763 1894 -3574 2167
rect -3392 1477 -3260 1578
rect -3398 418 -3309 451
rect -3309 418 -3303 451
rect -3398 341 -3303 418
rect -1676 1710 -1583 1735
rect -1583 1710 -1571 1735
rect -1676 1658 -1571 1710
rect -1681 1480 -1564 1584
rect -1682 351 -1606 453
rect -1680 197 -1553 286
rect -521 298 -311 480
rect -3568 -16 -3422 182
rect -3392 -1788 -3260 -1687
rect -3398 -2847 -3309 -2814
rect -3309 -2847 -3303 -2814
rect -3398 -2924 -3303 -2847
rect -1676 -1555 -1583 -1530
rect -1583 -1555 -1571 -1530
rect -1676 -1607 -1571 -1555
rect -1681 -1785 -1564 -1681
rect -1682 -2914 -1606 -2812
rect -1680 -3068 -1553 -2979
rect -521 -2967 -311 -2785
rect -3568 -3281 -3422 -3083
rect -3392 -5052 -3260 -4951
rect -3398 -6111 -3309 -6078
rect -3309 -6111 -3303 -6078
rect -3398 -6188 -3303 -6111
rect -1676 -4819 -1583 -4794
rect -1583 -4819 -1571 -4794
rect -1676 -4871 -1571 -4819
rect -1681 -5049 -1564 -4945
rect -1682 -6178 -1606 -6076
rect -1680 -6332 -1553 -6243
rect -521 -6231 -311 -6049
rect -3568 -6545 -3422 -6347
<< metal2 >>
rect -3591 4118 2084 4255
rect -3591 3538 -3448 4118
rect -3591 3515 -3296 3538
rect -1749 3536 -1606 4118
rect 92 3540 235 4118
rect -1749 3515 -1441 3536
rect 92 3515 400 3540
rect 1933 3539 2076 4118
rect 1933 3515 2238 3539
rect -3591 3405 -3422 3515
rect -3327 3405 -3296 3515
rect -3591 3399 -3296 3405
rect -3448 3398 -3296 3399
rect -2251 3511 -2177 3515
rect -2251 3324 -2030 3511
rect -1749 3405 -1581 3515
rect -1486 3405 -1441 3515
rect -1749 3400 -1441 3405
rect -364 3511 -244 3515
rect -364 3327 -135 3511
rect 92 3405 260 3515
rect 355 3405 400 3515
rect 92 3400 400 3405
rect 1477 3510 1516 3515
rect 1477 3327 1600 3510
rect 1933 3405 2101 3515
rect 2196 3405 2238 3515
rect 3453 3514 3608 3518
rect 1933 3400 2238 3405
rect 3318 3327 3608 3514
rect -3542 3244 -3356 3284
rect -3542 3066 -3506 3244
rect -3384 3066 -3356 3244
rect -3542 3048 -3356 3066
rect -2216 2727 -2030 3324
rect -1748 3215 -1558 3247
rect -1748 3043 -1722 3215
rect -1584 3158 -1558 3215
rect -1584 3144 -1412 3158
rect -1584 3043 -1563 3144
rect -1748 3022 -1563 3043
rect -1426 3022 -1412 3144
rect -1748 3013 -1412 3022
rect -275 2833 -135 3327
rect 100 3189 318 3210
rect 100 3066 127 3189
rect 303 3066 318 3189
rect 100 3045 318 3066
rect 1505 2985 1600 3327
rect 1752 3297 2032 3323
rect 1752 3144 1803 3297
rect 2001 3144 2032 3297
rect 1752 3116 2032 3144
rect 3453 3186 3608 3327
rect 3453 3064 13159 3186
rect 3458 3036 13159 3064
rect 1505 2984 10159 2985
rect 1505 2876 10170 2984
rect -1285 2727 -968 2736
rect -2216 2666 -968 2727
rect -285 2722 6879 2833
rect -2216 2614 3582 2666
rect -1285 2553 3582 2614
rect -1285 2544 -968 2553
rect -1869 2517 -1700 2527
rect -1869 2489 -1407 2517
rect -1869 2383 -1556 2489
rect -1432 2383 -1407 2489
rect 3458 2408 3581 2553
rect -1869 2354 -1407 2383
rect 6750 2376 6878 2722
rect 10028 2388 10170 2876
rect -3817 2167 -3534 2234
rect -3817 1894 -3763 2167
rect -3574 1894 -3534 2167
rect -3817 1852 -3534 1894
rect -1869 1763 -1700 2354
rect -2166 1751 -1533 1763
rect -2166 1637 -2151 1751
rect -2020 1735 -1533 1751
rect -2020 1658 -1676 1735
rect -1571 1658 -1533 1735
rect -2020 1637 -1533 1658
rect -2166 1628 -1533 1637
rect -3588 1578 -3225 1599
rect -3588 1477 -3392 1578
rect -3260 1477 -3225 1578
rect -3588 1463 -3225 1477
rect -1866 1584 -1547 1599
rect -1866 1480 -1681 1584
rect -1564 1480 -1547 1584
rect -1866 1463 -1547 1480
rect -312 1468 -3 1475
rect -3588 1204 -3412 1463
rect -1866 1204 -1690 1463
rect -3590 1069 -1690 1204
rect -3588 471 -3412 1069
rect -1866 471 -1690 1069
rect -351 1335 -3 1468
rect -518 526 -433 528
rect -351 526 -260 1335
rect -566 480 -260 526
rect -3588 451 -3281 471
rect -3588 341 -3398 451
rect -3303 341 -3281 451
rect -3588 336 -3281 341
rect -1866 453 -1593 471
rect -1866 351 -1682 453
rect -1606 351 -1593 453
rect -1866 336 -1593 351
rect -1867 300 -1528 306
rect -1868 286 -1528 300
rect -1868 236 -1680 286
rect -3593 182 -3395 211
rect -3593 -16 -3568 182
rect -3422 -16 -3395 182
rect -3593 -31 -3395 -16
rect -1868 -210 -1818 236
rect -1729 197 -1680 236
rect -1553 197 -1528 286
rect -566 298 -521 480
rect -311 298 -260 480
rect -566 263 -260 298
rect -1729 171 -1528 197
rect -1729 -108 -1692 171
rect -1729 -210 -1693 -108
rect -1868 -254 -1693 -210
rect 10 -200 287 -196
rect 10 -401 315 -200
rect 3275 -213 3407 -128
rect 6574 -187 6881 -83
rect 3275 -343 3638 -213
rect 3342 -344 3638 -343
rect -3604 -447 -299 -427
rect -3604 -453 -471 -447
rect -3604 -593 -3575 -453
rect -3446 -587 -471 -453
rect -342 -587 -299 -447
rect -3446 -593 -299 -587
rect -3604 -614 -299 -593
rect 171 -822 315 -401
rect 3452 -848 3636 -344
rect 6755 -863 6878 -187
rect 9870 -241 9997 -101
rect 10040 -241 10168 -240
rect 9865 -397 10168 -241
rect 9870 -398 9997 -397
rect 10040 -839 10168 -397
rect -2166 -1512 -1533 -1502
rect -2166 -1626 -2154 -1512
rect -2023 -1514 -1533 -1512
rect -2020 -1530 -1533 -1514
rect -2020 -1607 -1676 -1530
rect -1571 -1607 -1533 -1530
rect -2166 -1628 -2151 -1626
rect -2020 -1628 -1533 -1607
rect -2166 -1637 -1533 -1628
rect -3588 -1687 -3225 -1666
rect -3588 -1788 -3392 -1687
rect -3260 -1788 -3225 -1687
rect -3588 -1802 -3225 -1788
rect -1866 -1681 -1547 -1666
rect -1866 -1785 -1681 -1681
rect -1564 -1785 -1547 -1681
rect -1866 -1802 -1547 -1785
rect -312 -1797 -3 -1790
rect -3588 -2061 -3412 -1802
rect -1866 -2061 -1690 -1802
rect -3590 -2196 -1690 -2061
rect -3588 -2794 -3412 -2196
rect -1866 -2794 -1690 -2196
rect -351 -1930 -3 -1797
rect -518 -2739 -433 -2737
rect -351 -2739 -260 -1930
rect -566 -2785 -260 -2739
rect -3588 -2814 -3281 -2794
rect -3588 -2924 -3398 -2814
rect -3303 -2924 -3281 -2814
rect -3588 -2929 -3281 -2924
rect -1866 -2812 -1593 -2794
rect -1866 -2914 -1682 -2812
rect -1606 -2914 -1593 -2812
rect -1866 -2929 -1593 -2914
rect -1867 -2965 -1528 -2959
rect -1868 -2979 -1528 -2965
rect -1868 -3008 -1680 -2979
rect -3593 -3083 -3395 -3054
rect -3593 -3281 -3568 -3083
rect -3422 -3281 -3395 -3083
rect -3593 -3296 -3395 -3281
rect -1868 -3454 -1822 -3008
rect -1733 -3029 -1680 -3008
rect -1729 -3068 -1680 -3029
rect -1553 -3068 -1528 -2979
rect -566 -2967 -521 -2785
rect -311 -2967 -260 -2785
rect -566 -3002 -260 -2967
rect -1729 -3094 -1528 -3068
rect -1729 -3373 -1692 -3094
rect -1868 -3475 -1818 -3454
rect -1729 -3475 -1693 -3373
rect -1868 -3519 -1693 -3475
rect -11 -3621 314 -3495
rect 3281 -3497 3615 -3375
rect 169 -4142 299 -3621
rect 3456 -4161 3592 -3497
rect 6570 -3532 6886 -3387
rect 9874 -3505 10165 -3369
rect 6744 -4189 6874 -3532
rect 10040 -4161 10164 -3505
rect -2166 -4776 -1533 -4766
rect -2166 -4890 -2154 -4776
rect -2017 -4794 -1533 -4776
rect -2017 -4871 -1676 -4794
rect -1571 -4871 -1533 -4794
rect -2017 -4890 -1533 -4871
rect -2166 -4892 -2151 -4890
rect -2020 -4892 -1533 -4890
rect -2166 -4901 -1533 -4892
rect -3588 -4951 -3225 -4930
rect -3588 -5052 -3392 -4951
rect -3260 -5052 -3225 -4951
rect -3588 -5066 -3225 -5052
rect -1866 -4945 -1547 -4930
rect -1866 -5049 -1681 -4945
rect -1564 -5049 -1547 -4945
rect -1866 -5066 -1547 -5049
rect -312 -5061 -3 -5054
rect -3588 -5325 -3412 -5066
rect -1866 -5325 -1690 -5066
rect -3590 -5460 -1690 -5325
rect -3588 -6058 -3412 -5460
rect -1866 -6058 -1690 -5460
rect -351 -5194 -3 -5061
rect -518 -6003 -433 -6001
rect -351 -6003 -260 -5194
rect -566 -6049 -260 -6003
rect -3588 -6078 -3281 -6058
rect -3588 -6188 -3398 -6078
rect -3303 -6188 -3281 -6078
rect -3588 -6193 -3281 -6188
rect -1866 -6076 -1593 -6058
rect -1866 -6178 -1682 -6076
rect -1606 -6178 -1593 -6076
rect -1866 -6193 -1593 -6178
rect -1867 -6229 -1528 -6223
rect -1868 -6243 -1528 -6229
rect -1868 -6272 -1680 -6243
rect -1868 -6287 -1822 -6272
rect -3593 -6347 -3395 -6318
rect -3593 -6545 -3568 -6347
rect -3422 -6545 -3395 -6347
rect -3593 -6560 -3395 -6545
rect -1868 -6733 -1825 -6287
rect -1733 -6293 -1680 -6272
rect -1729 -6332 -1680 -6293
rect -1553 -6332 -1528 -6243
rect -566 -6231 -521 -6049
rect -311 -6231 -260 -6049
rect -566 -6266 -260 -6231
rect -1729 -6358 -1528 -6332
rect -1729 -6637 -1692 -6358
rect -1868 -6739 -1818 -6733
rect -1729 -6739 -1693 -6637
rect -1868 -6783 -1693 -6739
<< via2 >>
rect -3506 3066 -3384 3244
rect -1563 3022 -1426 3144
rect 127 3066 303 3189
rect 1803 3144 2001 3297
rect -1556 2383 -1432 2489
rect -3763 1894 -3574 2167
rect -2151 1637 -2020 1751
rect -3568 -16 -3422 182
rect -1818 -210 -1729 236
rect -3575 -593 -3446 -453
rect -471 -587 -342 -447
rect -2154 -1514 -2023 -1512
rect -2154 -1626 -2020 -1514
rect -2151 -1628 -2020 -1626
rect -3568 -3281 -3422 -3083
rect -1822 -3029 -1733 -3008
rect -1822 -3454 -1729 -3029
rect -1818 -3475 -1729 -3454
rect -2154 -4890 -2017 -4776
rect -2151 -4892 -2020 -4890
rect -1822 -6287 -1733 -6272
rect -3568 -6545 -3422 -6347
rect -1825 -6293 -1733 -6287
rect -1825 -6733 -1729 -6293
rect -1818 -6739 -1729 -6733
<< metal3 >>
rect -3817 4255 -3635 4259
rect -3817 4090 1969 4255
rect -3817 2234 -3635 4090
rect -3544 3244 -3354 3372
rect -3544 3218 -3506 3244
rect -3542 3066 -3506 3218
rect -3384 3218 -3354 3244
rect 1752 3323 1969 4090
rect 1752 3297 2032 3323
rect -3384 3066 -3358 3218
rect 100 3189 318 3210
rect -3542 2836 -3358 3066
rect -1583 3144 -1415 3161
rect -1583 3022 -1563 3144
rect -1426 3022 -1415 3144
rect 100 3066 127 3189
rect 303 3066 318 3189
rect 1752 3144 1803 3297
rect 2001 3144 2032 3297
rect 1752 3116 2032 3144
rect 100 3052 318 3066
rect -480 3045 318 3052
rect -480 3033 271 3045
rect -3542 2832 -1710 2836
rect -3542 2636 -1708 2832
rect -3817 2167 -3534 2234
rect -3817 1894 -3763 2167
rect -3574 1894 -3534 2167
rect -3817 1852 -3534 1894
rect -2166 1751 -2007 1796
rect -2166 1637 -2151 1751
rect -2020 1637 -2007 1751
rect -3607 211 -3416 332
rect -3607 182 -3395 211
rect -3607 -16 -3568 182
rect -3422 -16 -3395 182
rect -3607 -31 -3395 -16
rect -3607 -453 -3416 -31
rect -3607 -593 -3575 -453
rect -3446 -593 -3416 -453
rect -3607 -3054 -3416 -593
rect -2166 -1512 -2007 1637
rect -2166 -1626 -2154 -1512
rect -2023 -1514 -2007 -1512
rect -2166 -1628 -2151 -1626
rect -2020 -1628 -2007 -1514
rect -3607 -3083 -3395 -3054
rect -3607 -3281 -3568 -3083
rect -3422 -3281 -3395 -3083
rect -3607 -3296 -3395 -3281
rect -3607 -6318 -3416 -3296
rect -2166 -4776 -2007 -1628
rect -2166 -4890 -2154 -4776
rect -2017 -4890 -2007 -4776
rect -2166 -4892 -2151 -4890
rect -2020 -4892 -2007 -4890
rect -2166 -4901 -2007 -4892
rect -1893 236 -1708 2636
rect -1583 2489 -1415 3022
rect -1583 2383 -1556 2489
rect -1432 2383 -1415 2489
rect -1583 2362 -1415 2383
rect -481 2868 271 3033
rect -481 2858 265 2868
rect -1893 -210 -1818 236
rect -1729 -210 -1708 236
rect -1893 -3008 -1708 -210
rect -481 -447 -301 2858
rect -481 -587 -471 -447
rect -342 -587 -301 -447
rect -481 -623 -301 -587
rect -1893 -3454 -1822 -3008
rect -1733 -3029 -1708 -3008
rect -1893 -3475 -1818 -3454
rect -1729 -3475 -1708 -3029
rect -1893 -6272 -1708 -3475
rect -1893 -6287 -1822 -6272
rect -3607 -6347 -3395 -6318
rect -3607 -6545 -3568 -6347
rect -3422 -6545 -3395 -6347
rect -3607 -6560 -3395 -6545
rect -3607 -6772 -3416 -6560
rect -1893 -6733 -1825 -6287
rect -1733 -6293 -1708 -6272
rect -1893 -6739 -1818 -6733
rect -1729 -6739 -1708 -6293
rect -1893 -6782 -1708 -6739
use 4bit_ADDER  4bit_ADDER_0
timestamp 1736606925
transform 1 0 171 0 1 -165
box -174 -146 13189 3089
use 4bit_ADDER  4bit_ADDER_1
timestamp 1736606925
transform 1 0 171 0 1 -3430
box -174 -146 13189 3089
use 4bit_ADDER  4bit_ADDER_2
timestamp 1736606925
transform 1 0 171 0 1 -6694
box -174 -146 13189 3089
<< labels >>
rlabel metal1 -2500 3920 -2500 3920 1 VDD
port 1 n
rlabel metal1 -2268 3471 -2268 3471 3 Y
port 3 e
rlabel metal1 -602 3252 -602 3252 5 VSS
port 4 s
rlabel metal1 -659 3920 -659 3920 1 VDD
port 1 n
rlabel metal1 -427 3471 -427 3471 3 Y
port 3 e
rlabel metal1 1239 3252 1239 3252 5 VSS
port 4 s
rlabel metal1 1182 3920 1182 3920 1 VDD
port 1 n
rlabel metal1 1038 3471 1038 3471 7 A
port 2 e
rlabel metal1 1414 3471 1414 3471 3 Y
port 3 e
rlabel metal1 3080 3252 3080 3252 5 VSS
port 4 s
rlabel metal1 3023 3920 3023 3920 1 VDD
port 1 n
rlabel metal1 2879 3471 2879 3471 7 A
port 2 e
rlabel metal1 3255 3471 3255 3471 3 Y
port 3 e
flabel metal2 -3228 -2190 -3108 -2070 1 FreeSerif 160 0 0 0 B2
port 7 n
flabel metal2 -3584 3886 -3464 4006 1 FreeSerif 160 0 0 0 B0
port 8 n
flabel metal2 -3220 -5452 -3100 -5332 1 FreeSerif 160 0 0 0 B3
port 9 n
flabel metal2 -2952 -576 -2832 -456 1 FreeSerif 160 0 0 0 A1
port 11 n
flabel metal3 -3190 2678 -3070 2798 1 FreeSerif 160 0 0 0 A3
port 12 n
flabel metal2 12820 3054 12940 3174 1 FreeSerif 160 0 0 0 SO
port 13 n
flabel space 13166 -32 13262 54 1 FreeSerif 160 0 0 0 S1
port 14 n
flabel space 13182 -3394 13278 -3308 1 FreeSerif 160 0 0 0 S2
port 15 n
flabel space 6586 -6668 6682 -6582 1 FreeSerif 160 0 0 0 S5
port 16 n
flabel space 9878 -6670 9974 -6584 1 FreeSerif 160 0 0 0 S4
port 17 n
flabel space 13182 -6664 13278 -6578 1 FreeSerif 160 0 0 0 S3
port 18 n
flabel space 54 -6728 150 -6642 1 FreeSerif 160 0 0 0 S7
port 19 n
flabel space 3294 -6664 3390 -6578 1 FreeSerif 160 0 0 0 S6
port 20 n
rlabel metal1 -803 3471 -803 3471 7 A
port 2 e
rlabel metal1 -2644 3471 -2644 3471 7 A
port 2 e
rlabel metal1 -2443 3252 -2443 3252 5 VSS
port 4 s
flabel metal3 -2146 -202 -2026 -82 1 FreeSerif 160 0 0 0 A2
port 10 n
flabel metal2 -3556 1080 -3436 1200 1 FreeSerif 160 0 0 0 B1
port 5 n
flabel metal1 -3794 1646 -3674 1766 1 FreeSerif 160 0 0 0 A0
port 6 n
rlabel metal1 -518 1699 -518 1699 3 Y
port 3 e
rlabel metal1 -894 1699 -894 1699 7 A
port 2 e
rlabel metal1 -750 2148 -750 2148 1 VDD
port 1 n
rlabel metal1 -693 1480 -693 1480 5 VSS
port 4 s
rlabel metal1 -894 407 -894 407 7 A
port 2 e
rlabel metal1 -750 856 -750 856 1 VDD
port 1 n
rlabel metal1 -693 188 -693 188 5 VSS
port 4 s
rlabel metal1 -2244 407 -2244 407 3 Y
port 3 e
rlabel metal1 -2620 407 -2620 407 7 A
port 2 e
rlabel metal1 -2476 856 -2476 856 1 VDD
port 1 n
rlabel metal1 -2419 188 -2419 188 5 VSS
port 4 s
rlabel via1 -518 407 -518 407 3 Y
port 3 e
rlabel metal1 -2244 1699 -2244 1699 3 Y
port 3 e
rlabel metal1 -2620 1699 -2620 1699 7 A
port 2 e
rlabel metal1 -2476 2148 -2476 2148 1 VDD
port 1 n
rlabel metal1 -2419 1480 -2419 1480 5 VSS
port 4 s
rlabel metal1 -518 -1566 -518 -1566 3 Y
port 3 e
rlabel metal1 -894 -1566 -894 -1566 7 A
port 2 e
rlabel metal1 -750 -1117 -750 -1117 1 VDD
port 1 n
rlabel metal1 -693 -1785 -693 -1785 5 VSS
port 4 s
rlabel metal1 -894 -2858 -894 -2858 7 A
port 2 e
rlabel metal1 -750 -2409 -750 -2409 1 VDD
port 1 n
rlabel metal1 -693 -3077 -693 -3077 5 VSS
port 4 s
rlabel metal1 -2244 -2858 -2244 -2858 3 Y
port 3 e
rlabel metal1 -2620 -2858 -2620 -2858 7 A
port 2 e
rlabel metal1 -2476 -2409 -2476 -2409 1 VDD
port 1 n
rlabel metal1 -2419 -3077 -2419 -3077 5 VSS
port 4 s
rlabel via1 -518 -2858 -518 -2858 3 Y
port 3 e
rlabel metal1 -2244 -1566 -2244 -1566 3 Y
port 3 e
rlabel metal1 -2620 -1566 -2620 -1566 7 A
port 2 e
rlabel metal1 -2476 -1117 -2476 -1117 1 VDD
port 1 n
rlabel metal1 -2419 -1785 -2419 -1785 5 VSS
port 4 s
rlabel metal1 -518 -4830 -518 -4830 3 Y
port 3 e
rlabel metal1 -894 -4830 -894 -4830 7 A
port 2 e
rlabel metal1 -750 -4381 -750 -4381 1 VDD
port 1 n
rlabel metal1 -693 -5049 -693 -5049 5 VSS
port 4 s
rlabel metal1 -894 -6122 -894 -6122 7 A
port 2 e
rlabel metal1 -750 -5673 -750 -5673 1 VDD
port 1 n
rlabel metal1 -693 -6341 -693 -6341 5 VSS
port 4 s
rlabel metal1 -2244 -6122 -2244 -6122 3 Y
port 3 e
rlabel metal1 -2620 -6122 -2620 -6122 7 A
port 2 e
rlabel metal1 -2476 -5673 -2476 -5673 1 VDD
port 1 n
rlabel metal1 -2419 -6341 -2419 -6341 5 VSS
port 4 s
rlabel via1 -518 -6122 -518 -6122 3 Y
port 3 e
rlabel metal1 -2244 -4830 -2244 -4830 3 Y
port 3 e
rlabel metal1 -2620 -4830 -2620 -4830 7 A
port 2 e
rlabel metal1 -2476 -4381 -2476 -4381 1 VDD
port 1 n
rlabel metal1 -2419 -5049 -2419 -5049 5 VSS
port 4 s
<< end >>
