magic
tech sky130B
magscale 1 2
timestamp 1732912614
<< nwell >>
rect -353 -261 353 223
<< pmos >>
rect -255 -161 -225 161
rect -159 -161 -129 161
rect -63 -161 -33 161
rect 33 -161 63 161
rect 129 -161 159 161
rect 225 -161 255 161
<< pdiff >>
rect -317 149 -255 161
rect -317 -149 -305 149
rect -271 -149 -255 149
rect -317 -161 -255 -149
rect -225 149 -159 161
rect -225 -149 -209 149
rect -175 -149 -159 149
rect -225 -161 -159 -149
rect -129 149 -63 161
rect -129 -149 -113 149
rect -79 -149 -63 149
rect -129 -161 -63 -149
rect -33 149 33 161
rect -33 -149 -17 149
rect 17 -149 33 149
rect -33 -161 33 -149
rect 63 149 129 161
rect 63 -149 79 149
rect 113 -149 129 149
rect 63 -161 129 -149
rect 159 149 225 161
rect 159 -149 175 149
rect 209 -149 225 149
rect 159 -161 225 -149
rect 255 149 317 161
rect 255 -149 271 149
rect 305 -149 317 149
rect 255 -161 317 -149
<< pdiffc >>
rect -305 -149 -271 149
rect -209 -149 -175 149
rect -113 -149 -79 149
rect -17 -149 17 149
rect 79 -149 113 149
rect 175 -149 209 149
rect 271 -149 305 149
<< poly >>
rect -255 161 -225 187
rect -159 161 -129 187
rect -63 161 -33 187
rect 33 161 63 187
rect 129 161 159 187
rect 225 161 255 187
rect -255 -192 -225 -161
rect -159 -192 -129 -161
rect -63 -187 -33 -161
rect 33 -187 63 -161
rect -63 -192 63 -187
rect 129 -192 159 -161
rect 225 -192 255 -161
rect -273 -208 -129 -192
rect -273 -242 -257 -208
rect -223 -242 -129 -208
rect -273 -258 -129 -242
rect -81 -208 63 -192
rect -81 -242 -65 -208
rect -31 -242 63 -208
rect -81 -258 63 -242
rect 111 -208 255 -192
rect 111 -242 127 -208
rect 161 -242 255 -208
rect 111 -258 255 -242
<< polycont >>
rect -257 -242 -223 -208
rect -65 -242 -31 -208
rect 127 -242 161 -208
<< locali >>
rect -305 155 -271 165
rect -305 -165 -271 -149
rect -209 149 -175 165
rect -209 -165 -175 -155
rect -113 155 -79 165
rect -113 -165 -79 -149
rect -17 149 17 165
rect -17 -165 17 -155
rect 79 155 113 165
rect 79 -165 113 -149
rect 175 149 209 165
rect 175 -165 209 -155
rect 271 155 305 165
rect 271 -165 305 -149
rect -273 -242 -257 -208
rect -223 -242 -207 -208
rect -81 -242 -65 -208
rect -31 -242 -15 -208
rect 111 -242 127 -208
rect 161 -242 177 -208
<< viali >>
rect -305 149 -271 155
rect -305 23 -271 149
rect -209 -149 -175 -23
rect -209 -155 -175 -149
rect -113 149 -79 155
rect -113 23 -79 149
rect -17 -149 17 -23
rect -17 -155 17 -149
rect 79 149 113 155
rect 79 23 113 149
rect 175 -149 209 -23
rect 175 -155 209 -149
rect 271 149 305 155
rect 271 23 305 149
<< metal1 >>
rect -317 155 317 161
rect -317 23 -305 155
rect -271 23 -113 155
rect -79 23 79 155
rect 113 23 271 155
rect 305 23 317 155
rect -317 15 317 23
rect -225 -21 409 -15
rect -225 -23 410 -21
rect -225 -155 -209 -23
rect -175 -155 -17 -23
rect 17 -155 175 -23
rect 209 -155 410 -23
rect -225 -161 410 -155
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.605 l 0.15 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
