magic
tech sky130B
magscale 1 2
timestamp 1735985840
<< metal1 >>
rect 6 1844 78 1924
rect 178 1852 234 1924
rect 1318 1836 1390 1924
rect 1490 1846 1544 1924
rect 2618 1842 2690 1924
rect 2790 1844 2844 1922
rect 3826 1840 3898 1922
rect 3994 1846 4052 1922
rect 5024 1850 5072 1924
rect 5190 1848 5238 1922
rect 6150 1846 6198 1920
rect 6308 1850 6356 1924
rect 7358 1852 7406 1926
rect 7518 1850 7566 1924
rect 8540 1848 8588 1922
rect 8706 1848 8754 1922
rect 1012 -466 1081 70
rect 2318 -276 2387 50
rect 3625 -112 3694 70
rect 4821 -64 4890 66
rect 3582 -181 3694 -112
rect 4042 -133 4890 -64
rect 2318 -345 3191 -276
rect 1012 -535 2711 -466
rect 2642 -1081 2711 -535
rect 3122 -1072 3191 -345
rect 3582 -1078 3651 -181
rect 4042 -1072 4111 -133
rect 6005 -192 6074 56
rect 4522 -261 6074 -192
rect 4522 -1096 4591 -261
rect 7117 -304 7186 90
rect 5022 -373 7186 -304
rect 5022 -1094 5091 -373
rect 8313 -410 8382 78
rect 5502 -479 8382 -410
rect 5502 -1088 5571 -479
rect 9515 -598 9584 70
rect 6002 -667 9584 -598
rect 6002 -1081 6071 -667
rect 3012 -2650 3048 -2618
rect 3492 -2650 3528 -2618
rect 3952 -2650 3988 -2618
rect 4412 -2650 4448 -2618
rect 4892 -2650 4928 -2618
rect 5392 -2650 5428 -2618
rect 5872 -2646 5908 -2614
rect 6372 -2650 6408 -2618
use NAND8  NAND8_0 ~/Desktop/vlsi_sky130b/design/mag/NAND8
timestamp 1735984326
transform 1 0 5260 0 1 734
box -5260 -734 4324 1197
use NOT8  NOT8_0 ~/Desktop/vlsi_sky130b/design/mag/NOT
timestamp 1735843251
transform 1 0 2718 0 1 -2155
box -110 -501 3853 1143
<< labels >>
rlabel metal1 6 1844 78 1924 1 A0
port 1 n
rlabel metal1 178 1852 234 1924 1 B0
port 2 n
rlabel metal1 1318 1836 1390 1924 1 A1
port 3 n
rlabel metal1 1490 1846 1544 1924 1 B1
port 4 n
rlabel metal1 2790 1844 2844 1922 1 B2
port 5 n
rlabel metal1 2618 1842 2690 1924 1 A2
port 6 n
rlabel metal1 3826 1840 3898 1922 1 A3
port 7 n
rlabel metal1 3994 1846 4052 1922 1 B3
port 8 n
rlabel metal1 5190 1848 5238 1922 1 B4
port 9 n
rlabel metal1 5024 1850 5072 1924 1 A4
port 10 n
rlabel metal1 6150 1846 6198 1920 1 A5
port 11 n
rlabel metal1 6308 1850 6356 1924 1 B5
port 12 n
rlabel metal1 7518 1850 7566 1924 1 B6
port 13 n
rlabel metal1 7358 1852 7406 1926 1 A6
port 14 n
rlabel metal1 8540 1848 8588 1922 1 A7
port 15 n
rlabel metal1 8706 1848 8754 1922 1 B7
port 16 n
rlabel metal1 3012 -2650 3048 -2618 5 S0
port 17 s
rlabel metal1 3492 -2650 3528 -2618 5 S1
port 18 s
rlabel metal1 3952 -2650 3988 -2618 5 S2
port 19 s
rlabel metal1 4412 -2650 4448 -2618 5 S3
port 20 s
rlabel metal1 4892 -2650 4928 -2618 5 S4
port 21 s
rlabel metal1 5392 -2650 5428 -2618 5 S5
port 22 s
rlabel metal1 5872 -2646 5908 -2614 5 S6
port 23 s
rlabel metal1 6372 -2650 6408 -2618 5 S7
port 24 s
<< end >>
