magic
tech sky130B
magscale 1 2
timestamp 1735226356
<< error_s >>
rect 123 265 6842 684
rect 223 139 423 197
rect 602 139 802 197
rect 1075 139 1275 197
rect 1454 139 1654 197
rect 1927 139 2127 197
rect 2306 139 2506 197
rect 2779 139 2979 197
rect 3158 139 3358 197
rect 3631 139 3831 197
rect 4010 139 4210 197
rect 4483 139 4683 197
rect 4862 139 5062 197
rect 5335 140 5535 198
rect 5714 140 5914 198
rect 6187 140 6387 198
rect 6566 140 6766 198
rect 223 51 423 109
rect 602 51 802 109
rect 1075 51 1275 109
rect 1454 51 1654 109
rect 1927 51 2127 109
rect 2306 51 2506 109
rect 2779 51 2979 109
rect 3158 51 3358 109
rect 3631 51 3831 109
rect 4010 51 4210 109
rect 4483 51 4683 109
rect 4862 51 5062 109
rect 5335 52 5535 110
rect 5714 52 5914 110
rect 6187 52 6387 110
rect 6566 52 6766 110
rect 348 18 668 42
rect 1200 18 1520 42
rect 2052 18 2372 42
rect 2904 18 3224 42
rect 3756 18 4076 42
rect 4608 18 4928 42
rect 5460 19 5780 43
rect 6312 19 6632 43
rect 348 -254 372 18
rect 1200 -254 1224 18
rect 2052 -254 2076 18
rect 2904 -254 2928 18
rect 3756 -254 3780 18
rect 4608 -254 4632 18
rect 5460 -253 5484 19
rect 6312 -253 6336 19
rect 348 -278 668 -254
rect 1200 -278 1520 -254
rect 2052 -278 2372 -254
rect 2904 -278 3224 -254
rect 3756 -278 4076 -254
rect 4608 -278 4928 -254
rect 5460 -277 5780 -253
rect 6312 -277 6632 -253
<< nwell >>
rect 123 265 6842 684
<< metal1 >>
rect 26 683 192 858
rect 878 683 1044 858
rect 1730 683 1896 858
rect 2582 683 2748 858
rect 3434 683 3600 858
rect 4286 684 4452 859
rect 123 603 192 683
rect 975 603 1044 683
rect 122 -278 288 15
rect 878 6 947 603
rect 1827 602 1896 683
rect 2679 602 2748 683
rect 3531 602 3600 683
rect 4383 602 4452 684
rect 5138 683 5304 858
rect 6087 857 6156 858
rect 5235 602 5304 683
rect 5990 682 6156 857
rect 6087 602 6156 682
rect 878 -278 1044 6
rect 1730 -2 1799 595
rect 2582 5 2651 602
rect 3434 5 3503 602
rect 4286 5 4355 602
rect 5138 5 5207 602
rect 5990 5 6059 602
rect 6842 5 6911 602
rect 1730 -278 1896 -2
rect 2582 -279 2748 5
rect 3434 -279 3600 5
rect 4286 -279 4452 5
rect 5138 -279 5304 5
rect 5990 -279 6156 5
rect 6842 -279 7008 5
use buffer  buffer_0 ~/Documents/Dersler/VLSI/vlsi_sky130b/design/mag/inv
timestamp 1735226356
transform 1 0 4615 0 1 313
box 1472 -590 2227 547
use buffer  buffer_1
timestamp 1735226356
transform 1 0 -1349 0 1 312
box 1472 -590 2227 547
use buffer  buffer_2
timestamp 1735226356
transform 1 0 -497 0 1 312
box 1472 -590 2227 547
use buffer  buffer_3
timestamp 1735226356
transform 1 0 355 0 1 312
box 1472 -590 2227 547
use buffer  buffer_4
timestamp 1735226356
transform 1 0 1207 0 1 312
box 1472 -590 2227 547
use buffer  buffer_5
timestamp 1735226356
transform 1 0 2059 0 1 312
box 1472 -590 2227 547
use buffer  buffer_6
timestamp 1735226356
transform 1 0 2911 0 1 312
box 1472 -590 2227 547
use buffer  buffer_7
timestamp 1735226356
transform 1 0 3763 0 1 313
box 1472 -590 2227 547
<< end >>
