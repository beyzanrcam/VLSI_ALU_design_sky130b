magic
tech sky130B
magscale 1 2
timestamp 1736693491
<< nwell >>
rect 1282 2682 1443 2683
rect -168 1782 4600 2682
rect 5760 1946 6094 1969
rect 5742 1916 6278 1946
rect 5733 1844 6278 1916
rect 5742 1542 6278 1844
rect 5770 1537 6278 1542
rect 5802 1536 6278 1537
<< poly >>
rect -282 1715 -59 1725
rect -282 1626 -266 1715
rect -177 1626 -59 1715
rect -282 1616 -59 1626
rect 1332 1715 1547 1725
rect 1332 1626 1348 1715
rect 1437 1626 1547 1715
rect 1332 1616 1547 1626
rect 3016 1713 3251 1723
rect 3016 1624 3032 1713
rect 3121 1624 3251 1713
rect 3016 1614 3251 1624
<< polycont >>
rect -266 1626 -177 1715
rect 1348 1626 1437 1715
rect 3032 1624 3121 1713
<< locali >>
rect -275 1715 -166 1770
rect -275 1626 -266 1715
rect -177 1626 -166 1715
rect -275 1616 -166 1626
rect 1338 1715 1447 1743
rect 3022 1745 3131 1888
rect 3022 1723 3138 1745
rect 1338 1626 1348 1715
rect 1437 1626 1447 1715
rect 1338 1616 1447 1626
rect 3016 1713 3138 1723
rect 3016 1624 3032 1713
rect 3121 1624 3138 1713
rect -266 1610 -177 1616
rect 1348 1610 1437 1616
rect 3016 1613 3138 1624
rect 3032 1610 3121 1613
<< viali >>
rect 3022 1888 3131 1985
rect -275 1770 -166 1867
rect 1338 1743 1447 1840
<< metal1 >>
rect -463 1604 -355 2700
rect -274 2297 -165 2690
rect -274 1873 -165 2185
rect -287 1867 -154 1873
rect -287 1770 -275 1867
rect -166 1770 -154 1867
rect 1338 1846 1447 2742
rect 2890 1913 2982 2720
rect 3022 2296 3131 2720
rect 4446 2316 6187 2637
rect 3022 2187 3034 2296
rect 3022 1991 3131 2187
rect -287 1764 -154 1770
rect 1326 1840 1459 1846
rect 1326 1743 1338 1840
rect 1447 1743 1459 1840
rect 2890 1844 2899 1913
rect 2968 1844 2982 1913
rect 3010 1985 3143 1991
rect 3010 1888 3022 1985
rect 3131 1888 3143 1985
rect 5261 1916 6184 2316
rect 5261 1898 5733 1916
rect 3010 1882 3143 1888
rect 5281 1848 5733 1898
rect 5965 1898 6184 1916
rect 5965 1848 6181 1898
rect 2890 1810 2982 1844
rect 1326 1737 1459 1743
rect 2759 1610 2872 1656
rect -481 1461 -47 1604
rect 1187 1461 1559 1604
rect 2759 1531 2857 1610
rect 2759 1519 2987 1531
rect 2850 955 2987 1519
rect 3114 1459 3120 1602
rect 3189 1459 3269 1602
rect 4473 1549 4916 1608
rect 4473 1494 5178 1549
rect 5760 1542 5908 1692
rect 5735 1536 5908 1542
rect 4802 1435 5178 1494
rect 5760 1418 5908 1536
rect 6209 1428 6251 1453
rect 5064 955 5200 1406
rect 5485 1180 5594 1250
rect 5475 1174 5602 1180
rect 5475 1065 5484 1174
rect 5594 1065 5602 1174
rect 5475 1056 5602 1065
rect 5971 1174 6080 1300
rect 5971 1059 6080 1065
rect 2850 818 5200 955
<< via1 >>
rect -274 2185 -165 2297
rect 3034 2187 3131 2296
rect 2899 1844 2968 1913
rect 3120 1459 3189 1602
rect 5484 1065 5594 1174
rect 5971 1065 6080 1174
<< metal2 >>
rect -280 2297 -160 2304
rect -280 2185 -274 2297
rect -165 2296 -160 2297
rect -165 2187 3034 2296
rect 3131 2187 3137 2296
rect -165 2185 -160 2187
rect -280 2179 -160 2185
rect 2899 1913 2968 1919
rect 2899 1565 2968 1844
rect 3120 1602 3189 1608
rect 2899 1496 3120 1565
rect 3120 1453 3189 1459
rect 3744 1174 3853 1251
rect 5474 1174 5605 1184
rect 3744 1065 5484 1174
rect 5594 1065 5971 1174
rect 6080 1065 6086 1174
rect 5474 1055 5605 1065
<< metal4 >>
rect -52 2509 4453 2657
<< metal5 >>
rect 181 989 4352 1346
use inv  inv_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/inv
timestamp 1736620191
transform 1 0 5870 0 1 1461
box 0 -311 412 486
use NAND2  NAND2_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NAND/NAND2
timestamp 1736620191
transform 1 0 4708 0 1 1165
box 356 -17 1062 804
use XOR2  XOR2_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/XOR
timestamp 1736689398
transform 1 0 3229 0 1 917
box -109 77 1371 1764
use XOR2  XOR2_1
timestamp 1736689398
transform 1 0 -81 0 1 919
box -109 77 1371 1764
use XOR2  XOR2_2
timestamp 1736689398
transform 1 0 1525 0 1 919
box -109 77 1371 1764
<< labels >>
flabel metal1 -237 2635 -190 2673 0 FreeSans 160 0 0 0 A_MSB
port 1 nsew
flabel metal1 -432 2633 -385 2671 0 FreeSans 160 0 0 0 B_MSB
port 2 nsew
flabel metal1 1367 2683 1414 2721 0 FreeSans 160 0 0 0 OPCODE3
port 3 nsew
flabel metal1 2920 2675 2962 2700 0 FreeSans 160 0 0 0 Y_MSB
port 4 nsew
flabel metal1 6209 1428 6251 1453 0 FreeSans 160 0 0 0 V
port 5 nsew
<< end >>
