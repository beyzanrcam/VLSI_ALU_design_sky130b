magic
tech sky130B
magscale 1 2
timestamp 1736187666
<< metal1 >>
rect 3113 953 3316 1044
rect 6404 953 6607 1044
rect 9695 953 9898 1044
rect 12986 953 13189 1044
rect 16277 953 16480 1044
rect 19567 953 19770 1044
rect 22858 953 23061 1044
rect 26149 953 26352 1044
use FULL_ADDER_XORED  FULL_ADDER_XORED_0
timestamp 1736187666
transform 1 0 118 0 1 1114
box -292 -1260 3108 3309
use FULL_ADDER_XORED  FULL_ADDER_XORED_1
timestamp 1736187666
transform 1 0 3409 0 1 1114
box -292 -1260 3108 3309
use FULL_ADDER_XORED  FULL_ADDER_XORED_2
timestamp 1736187666
transform 1 0 6700 0 1 1114
box -292 -1260 3108 3309
use FULL_ADDER_XORED  FULL_ADDER_XORED_3
timestamp 1736187666
transform 1 0 9991 0 1 1114
box -292 -1260 3108 3309
use FULL_ADDER_XORED  FULL_ADDER_XORED_4
timestamp 1736187666
transform 1 0 13282 0 1 1114
box -292 -1260 3108 3309
use FULL_ADDER_XORED  FULL_ADDER_XORED_5
timestamp 1736187666
transform 1 0 16572 0 1 1114
box -292 -1260 3108 3309
use FULL_ADDER_XORED  FULL_ADDER_XORED_6
timestamp 1736187666
transform 1 0 19863 0 1 1114
box -292 -1260 3108 3309
use FULL_ADDER_XORED  FULL_ADDER_XORED_7
timestamp 1736187666
transform 1 0 23154 0 1 1114
box -292 -1260 3108 3309
<< end >>
