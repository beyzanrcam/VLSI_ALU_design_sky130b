magic
tech sky130B
magscale 1 2
timestamp 1736096163
<< nwell >>
rect 10 444 908 571
rect 45 414 872 444
<< psubdiff >>
rect 206 -335 268 -311
rect 240 -683 268 -335
rect 206 -735 268 -683
rect 240 -1086 268 -735
rect 206 -1111 268 -1086
<< nsubdiff >>
rect 46 510 872 526
rect 46 475 297 510
rect 585 489 872 510
rect 585 475 871 489
rect 46 472 871 475
<< psubdiffcont >>
rect 206 -683 240 -335
rect 206 -1086 240 -735
<< nsubdiffcont >>
rect 297 475 585 510
<< poly >>
rect 146 -248 176 42
rect 340 2 370 42
rect 282 -1 402 2
rect 522 -1 552 32
rect 726 -1 756 40
rect 282 -68 426 -1
rect 492 -26 552 -1
rect 282 -206 456 -68
rect 146 -278 360 -248
rect 330 -287 360 -278
rect 426 -311 456 -206
rect 498 -288 552 -26
rect 666 -131 756 -1
rect 522 -311 552 -288
rect 618 -161 756 -131
rect 618 -311 648 -161
<< locali >>
rect 281 475 297 510
rect 585 475 611 510
rect 206 -335 311 -304
rect 241 -1086 311 -335
rect 206 -1115 311 -1086
<< viali >>
rect 297 475 585 510
rect 206 -683 240 -335
rect 240 -683 241 -335
rect 206 -735 241 -683
rect 206 -1086 240 -735
rect 240 -1086 241 -735
<< metal1 >>
rect 45 510 872 526
rect 45 475 297 510
rect 585 475 872 510
rect 45 414 872 475
rect 809 109 909 230
rect 10 -1 156 65
rect 212 -1 349 65
rect 212 -29 278 -1
rect 10 -95 278 -29
rect 399 -2 540 64
rect 569 -1 733 65
rect 399 -38 465 -2
rect 502 -3 536 -2
rect 317 -123 465 -38
rect 10 -189 465 -123
rect 569 -217 635 -1
rect 10 -283 635 -217
rect 799 -311 909 109
rect 122 -335 321 -311
rect 122 -1086 206 -335
rect 241 -1086 321 -335
rect 122 -1175 321 -1086
rect 658 -326 909 -311
rect 658 -1111 908 -326
use efenmos2  efenmos2_1
timestamp 1736094670
transform 1 0 489 0 1 -711
box -221 -426 221 426
use pmos4_f2  pmos4_f2_0
timestamp 1735579975
transform 1 0 459 0 1 257
box -449 -261 449 223
<< labels >>
flabel metal1 17 -277 51 -228 0 FreeSans 160 0 0 0 A
port 1 nsew
flabel metal1 20 -177 54 -128 0 FreeSans 160 0 0 0 B
port 2 nsew
flabel metal1 21 -89 55 -40 0 FreeSans 160 0 0 0 C
port 3 nsew
flabel metal1 22 4 56 53 0 FreeSans 160 0 0 0 D
port 4 nsew
flabel metal1 159 -1095 193 -1046 0 FreeSans 160 0 0 0 VSS
port 5 nsew
flabel nwell 422 466 456 515 0 FreeSans 160 0 0 0 VDD
port 6 nsew
flabel metal1 855 -214 889 -165 0 FreeSans 160 0 0 0 Y
port 8 nsew
<< end >>
