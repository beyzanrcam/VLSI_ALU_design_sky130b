magic
tech sky130B
magscale 1 2
timestamp 1736696497
<< metal1 >>
rect -27350 6877 1670 6966
rect -27525 4541 -27436 4547
rect -27350 4541 -27261 6877
rect -21821 6595 -21815 6684
rect -21726 6595 -21720 6684
rect -15130 6664 -15022 6670
rect -27436 4452 -25005 4541
rect -22644 4490 -22532 4500
rect -27525 4446 -27436 4452
rect -22644 4418 -22632 4490
rect -22560 4418 -22532 4490
rect -22644 4398 -22532 4418
rect -21815 4304 -21726 6595
rect -15022 6556 1484 6664
rect -15130 6550 -15022 6556
rect -19318 6376 -19312 6448
rect -19240 6376 -19234 6448
rect -19312 4308 -19240 6376
rect -18534 6279 -18528 6368
rect -18439 6279 -18433 6368
rect -18528 4432 -18439 6279
rect -16025 6124 -16019 6196
rect -15947 6124 -15941 6196
rect -16019 4313 -15947 6124
rect -15236 5884 -15230 5973
rect -15141 5884 -15135 5973
rect -15230 4331 -15141 5884
rect 1376 5818 1484 6556
rect 1581 6130 1670 6877
rect -12748 5681 -12742 5753
rect -12670 5681 -12664 5753
rect -12742 4436 -12670 5681
rect -11946 5537 -11940 5626
rect -11851 5537 -11845 5626
rect -11940 4438 -11851 5537
rect -9445 5385 -9439 5457
rect -9367 5385 -9361 5457
rect 3189 5390 3195 5442
rect 3247 5390 3253 5442
rect -9439 4434 -9367 5385
rect -6173 5339 -6084 5346
rect -8646 5227 -8640 5316
rect -8551 5227 -8545 5316
rect -6173 5269 -6166 5339
rect -6096 5269 -6084 5339
rect -6173 5261 -6084 5269
rect -8640 4490 -8551 5227
rect -6166 4453 -6096 5261
rect -5357 4991 -5351 5080
rect -5262 4991 -5256 5080
rect 8026 5020 8106 5116
rect -5351 4459 -5262 4991
rect -2881 4746 -2875 4818
rect -2803 4746 -2797 4818
rect -2875 4461 -2803 4746
rect 419 4612 425 4684
rect 497 4612 503 4684
rect -2064 4473 -2058 4562
rect -1969 4473 -1963 4562
rect 425 4513 497 4612
rect 2921 4275 2987 4281
rect 4885 4275 4951 4281
rect 2987 4209 4885 4275
rect 4951 4209 4993 4275
rect 2921 4203 2987 4209
rect 4885 4203 4951 4209
rect 5339 4083 5411 4089
rect 5339 3540 5411 4011
rect 605 3365 5411 3540
rect 1922 2519 2013 2538
rect 1922 2453 1934 2519
rect 2000 2453 2013 2519
rect -25060 1117 -24824 1208
rect -25060 -123 -24969 1117
rect -8633 309 -8567 315
rect -15223 296 -15157 302
rect -21801 284 -21735 290
rect -25066 -214 -25060 -123
rect -24969 -214 -24963 -123
rect -21801 -492 -21735 218
rect -18505 -306 -18439 286
rect -18505 -372 -15446 -306
rect -21801 -558 -15583 -492
rect -15649 -1309 -15583 -558
rect -15512 -1138 -15446 -372
rect -15223 -948 -15157 230
rect -11969 223 -11963 289
rect -11897 223 -11891 289
rect -11963 -785 -11897 223
rect -8633 -618 -8567 243
rect -5349 292 -5283 298
rect -5349 -421 -5283 226
rect -2061 261 -1995 267
rect -2061 -232 -1995 195
rect 248 -40 339 -34
rect 1922 -40 2013 2453
rect 6917 2147 6966 2213
rect 7032 2147 7299 2213
rect 13152 1469 13208 1558
rect 6953 1111 7019 1117
rect 7019 1045 7283 1111
rect 6953 1039 7019 1045
rect 339 -131 2013 -40
rect 248 -137 339 -131
rect -2061 -238 5481 -232
rect -2061 -298 5485 -238
rect -5349 -487 5327 -421
rect -8633 -684 5162 -618
rect -11963 -851 5014 -785
rect -15223 -1014 4904 -948
rect -15512 -1204 4639 -1138
rect -15649 -1375 1625 -1309
rect 1691 -1375 4493 -1309
rect 3886 -1551 3970 -1545
rect -7879 -6291 -7873 -6225
rect -7807 -6291 -7801 -6225
rect -7873 -6533 -7807 -6291
rect -5439 -6533 -5373 -6527
rect -7873 -6599 -5439 -6533
rect -5439 -6605 -5373 -6599
rect -7879 -8271 -4977 -8205
rect -24837 -10970 -24748 -10964
rect -24837 -11065 -24748 -11059
rect -5043 -11161 -4977 -8271
rect -5043 -11233 -4977 -11227
rect -7881 -11789 473 -11723
rect -1325 -12387 295 -12321
rect -7799 -12798 -7688 -12792
rect -1325 -12797 -1259 -12387
rect -7799 -12915 -7688 -12909
rect -6359 -12863 -1259 -12797
rect -1209 -12549 125 -12483
rect -6359 -13379 -6293 -12863
rect -1209 -12927 -1143 -12549
rect -11157 -13445 -11151 -13379
rect -11085 -13445 -6293 -13379
rect -6213 -12993 -1143 -12927
rect -1076 -12682 -57 -12623
rect -6213 -13577 -6147 -12993
rect -1076 -13069 -1017 -12682
rect -768 -12818 -684 -12812
rect -684 -12902 -676 -12834
rect -768 -12932 -676 -12902
rect -14449 -13643 -14443 -13577
rect -14377 -13643 -6147 -13577
rect -6088 -13128 -1017 -13069
rect -760 -13066 -676 -12932
rect -6088 -13700 -6029 -13128
rect -760 -13150 -374 -13066
rect -768 -13259 -684 -13258
rect -5292 -13312 -5286 -13259
rect -5233 -13312 -682 -13259
rect -5814 -13408 -5730 -13402
rect -5730 -13492 -850 -13408
rect -5814 -13498 -5730 -13492
rect -17736 -13759 -17730 -13700
rect -17671 -13759 -6029 -13700
rect -1201 -13666 -1117 -13660
rect -4632 -13818 -4626 -13734
rect -4542 -13818 -3436 -13734
rect -1374 -13750 -1201 -13720
rect -1374 -13804 -1117 -13750
rect -14814 -13976 -14808 -13924
rect -14756 -13976 -14750 -13924
rect -21025 -14475 -20959 -14469
rect -20959 -14541 -19311 -14475
rect -21025 -14547 -20959 -14541
rect -24936 -15658 -24916 -15586
rect -24844 -15658 -24818 -15586
rect -24931 -17012 -24925 -16923
rect -24836 -17012 -24830 -16923
rect -24927 -18054 -24921 -17984
rect -24851 -18054 -24845 -17984
rect -20405 -17986 -20399 -17934
rect -20347 -17986 -20341 -17934
rect -20414 -18434 -20362 -18428
rect -20356 -18486 -20350 -18434
rect -20414 -18492 -20362 -18486
rect -19377 -18705 -19311 -14541
rect -17978 -15586 -17880 -15576
rect -17978 -15658 -17966 -15586
rect -17894 -15658 -17880 -15586
rect -17978 -15666 -17880 -15658
rect -18133 -15738 -17893 -15724
rect -18133 -15827 -18123 -15738
rect -18034 -15790 -17893 -15738
rect -18034 -15827 -18005 -15790
rect -18133 -15847 -18005 -15827
rect -18082 -16980 -18010 -16974
rect -18010 -17052 -17892 -16980
rect -18082 -17058 -18010 -17052
rect -18096 -17113 -17992 -17102
rect -18096 -17202 -18089 -17113
rect -18000 -17202 -17830 -17113
rect -18096 -17208 -17992 -17202
rect -14806 -17799 -14758 -13976
rect -10855 -14032 -10779 -13897
rect -5376 -13928 -5370 -13876
rect -5318 -13880 -5312 -13876
rect -5174 -13880 -3570 -13860
rect -5318 -13924 -3570 -13880
rect -5318 -13928 -5312 -13924
rect -5174 -13944 -3570 -13924
rect -14708 -14088 -14656 -14082
rect -5969 -14065 -5963 -13983
rect -5881 -14065 -3716 -13983
rect -10855 -14114 -10779 -14108
rect -14708 -14146 -14656 -14140
rect -6954 -14142 -6902 -14136
rect -14808 -17863 -14756 -17799
rect -14706 -18307 -14658 -14146
rect -10850 -14331 -10795 -14325
rect -12730 -15586 -12656 -15570
rect -12730 -15658 -12724 -15586
rect -12652 -15658 -12512 -15586
rect -12730 -15666 -12656 -15658
rect -12566 -15738 -12440 -15728
rect -12566 -15837 -12555 -15738
rect -12456 -15837 -12440 -15738
rect -12566 -15848 -12440 -15837
rect -14618 -16016 -14612 -15964
rect -14560 -16016 -14554 -15964
rect -14806 -18355 -14658 -18307
rect -18065 -18385 -17995 -18379
rect -17995 -18455 -17893 -18385
rect -18065 -18461 -17995 -18455
rect -18099 -18515 -18010 -18509
rect -18010 -18604 -17834 -18515
rect -18099 -18610 -18010 -18604
rect -19383 -18771 -19377 -18705
rect -19311 -18771 -19305 -18705
rect -14610 -18787 -14562 -16016
rect -14496 -16186 -14444 -16180
rect -14496 -16244 -14444 -16238
rect -14806 -18835 -14562 -18787
rect -20406 -18914 -20340 -18908
rect -20406 -18966 -20399 -18914
rect -20347 -18966 -20340 -18914
rect -20406 -18972 -20340 -18966
rect -24876 -19175 -24870 -19103
rect -24798 -19175 -24792 -19103
rect -14494 -19287 -14446 -16244
rect -10850 -16457 -10795 -14386
rect -10307 -14771 -10252 -14765
rect -10849 -16751 -10797 -16457
rect -10307 -16774 -10252 -14826
rect -6954 -15246 -6902 -14194
rect -6966 -15298 -6902 -15246
rect -6834 -14490 -6782 -14484
rect -8690 -15496 -8594 -15486
rect -8690 -15568 -8676 -15496
rect -8604 -15568 -8594 -15496
rect -8690 -15586 -8594 -15568
rect -8690 -15588 -8476 -15586
rect -8676 -15658 -8476 -15588
rect -6834 -15746 -6782 -14542
rect -5020 -14494 -4926 -14484
rect -5020 -14566 -5008 -14494
rect -4936 -14566 -4926 -14494
rect -3899 -14491 -3833 -14485
rect -3798 -14556 -3716 -14065
rect -3899 -14563 -3833 -14557
rect -5020 -14576 -4926 -14566
rect -6662 -14860 -6614 -14850
rect -6674 -14870 -6600 -14860
rect -6674 -14922 -6664 -14870
rect -6612 -14922 -6600 -14870
rect -6674 -14930 -6600 -14922
rect -6970 -15798 -6782 -15746
rect -8554 -16140 -8482 -16087
rect -8570 -16152 -8470 -16140
rect -8570 -16224 -8554 -16152
rect -8482 -16224 -8470 -16152
rect -8570 -16236 -8470 -16224
rect -6662 -16228 -6614 -14930
rect -3654 -15182 -3570 -13944
rect -4044 -15266 -3570 -15182
rect -4974 -15306 -4880 -15294
rect -4974 -15378 -4966 -15306
rect -4894 -15378 -4880 -15306
rect -4044 -15334 -3960 -15266
rect -4974 -15386 -4880 -15378
rect -3520 -16069 -3436 -13818
rect -934 -14539 -850 -13492
rect -1336 -14623 -850 -14539
rect -768 -15358 -684 -13312
rect -1344 -15442 -684 -15358
rect -4044 -16153 -3436 -16069
rect -458 -16177 -374 -13150
rect -6960 -16276 -6614 -16228
rect -1356 -16261 -368 -16177
rect -8551 -16685 -8482 -16571
rect -116 -16706 -57 -12682
rect 59 -16557 125 -12549
rect 229 -16409 295 -12387
rect 407 -15427 473 -11789
rect 407 -15499 473 -15493
rect 229 -16475 1433 -16409
rect 59 -16623 1287 -16557
rect -8551 -16760 -8482 -16754
rect -12666 -18396 -12594 -18390
rect -12594 -18468 -12550 -18396
rect -12666 -18474 -12594 -18468
rect -12633 -18573 -12544 -18567
rect -12544 -18662 -12494 -18573
rect -12633 -18668 -12544 -18662
rect -14812 -19335 -14446 -19287
rect -20410 -19466 -20404 -19414
rect -20352 -19466 -20346 -19414
rect -18024 -19622 -17942 -19614
rect -10328 -19622 -10233 -16774
rect -6958 -16776 -5186 -16728
rect -116 -16765 1137 -16706
rect -8549 -17188 -8480 -17071
rect -5397 -17149 -5307 -17148
rect -5407 -17154 -5288 -17149
rect -8560 -17205 -8464 -17188
rect -8560 -17274 -8549 -17205
rect -8480 -17274 -8464 -17205
rect -6958 -17256 -5536 -17208
rect -5407 -17243 -5397 -17154
rect -5307 -17243 -5288 -17154
rect -5407 -17252 -5288 -17243
rect -8560 -17286 -8464 -17274
rect -8554 -17615 -8485 -17551
rect -8554 -17690 -8485 -17684
rect -6972 -17716 -5652 -17668
rect -8554 -18097 -8485 -18011
rect -8554 -18172 -8485 -18166
rect -6958 -18176 -5804 -18128
rect -8554 -18567 -8485 -18471
rect -8554 -18642 -8485 -18636
rect -6958 -18656 -5982 -18608
rect -8584 -19098 -8512 -18948
rect -8590 -19170 -8584 -19098
rect -8512 -19170 -8506 -19098
rect -18024 -19685 -18016 -19622
rect -17953 -19685 -17942 -19622
rect -18024 -19692 -17942 -19685
rect -18016 -19847 -17953 -19692
rect -10874 -19717 -10233 -19622
rect -14808 -19866 -14760 -19767
rect -20324 -19894 -20272 -19888
rect -20397 -19944 -20324 -19896
rect -20324 -19952 -20272 -19946
rect -17994 -19907 -17906 -19898
rect -17994 -19978 -17986 -19907
rect -17915 -19978 -17906 -19907
rect -14814 -19918 -14808 -19866
rect -14756 -19918 -14750 -19866
rect -17994 -19986 -17906 -19978
rect -14806 -20275 -12700 -20227
rect -24956 -20291 -24844 -20290
rect -24956 -20363 -24936 -20291
rect -24864 -20363 -24844 -20291
rect -24956 -20364 -24844 -20363
rect -20405 -20406 -20399 -20354
rect -20347 -20406 -20341 -20354
rect -24940 -20444 -24792 -20436
rect -24940 -20533 -24902 -20444
rect -24811 -20533 -24792 -20444
rect -24940 -20534 -24792 -20533
rect -14806 -20735 -12822 -20687
rect -18578 -20816 -18572 -20814
rect -20414 -20864 -18572 -20816
rect -18578 -20866 -18572 -20864
rect -18520 -20866 -18514 -20814
rect -18053 -21176 -17992 -21170
rect -17992 -21237 -17900 -21176
rect -14820 -21215 -12966 -21167
rect -18053 -21243 -17992 -21237
rect -18692 -21294 -18640 -21288
rect -20408 -21344 -18692 -21296
rect -17968 -21322 -17904 -21274
rect -18692 -21352 -18640 -21346
rect -17974 -21340 -17886 -21322
rect -17974 -21404 -17968 -21340
rect -17904 -21404 -17886 -21340
rect -17974 -21410 -17886 -21404
rect -18067 -22666 -18061 -22600
rect -17995 -22666 -17898 -22600
rect -18080 -22745 -17952 -22724
rect -18080 -22834 -18071 -22745
rect -17982 -22834 -17876 -22745
rect -18080 -22846 -17952 -22834
rect -18050 -23986 -17962 -23978
rect -18050 -24058 -18042 -23986
rect -17970 -24058 -17900 -23986
rect -18050 -24066 -17962 -24058
rect -18084 -24131 -17958 -24102
rect -18084 -24220 -18063 -24131
rect -17974 -24220 -17880 -24131
rect -18084 -24246 -17958 -24220
rect -24934 -24261 -24778 -24252
rect -24934 -24350 -24907 -24261
rect -24813 -24350 -24778 -24261
rect -24934 -24360 -24778 -24350
rect -13014 -25106 -12966 -21215
rect -12870 -22284 -12822 -20735
rect -12748 -22092 -12700 -20275
rect -12618 -21367 -12524 -21354
rect -12618 -21437 -12609 -21367
rect -12539 -21437 -12524 -21367
rect -12618 -21448 -12524 -21437
rect -12640 -21527 -12518 -21518
rect -12640 -21616 -12628 -21527
rect -12539 -21616 -12482 -21527
rect -12640 -21624 -12518 -21616
rect -12750 -22098 -12698 -22092
rect -12750 -22156 -12698 -22150
rect -12878 -22336 -12872 -22284
rect -12820 -22336 -12814 -22284
rect -10868 -22334 -10606 -22245
rect -12688 -23951 -12602 -23946
rect -12688 -23952 -12676 -23951
rect -12736 -24014 -12676 -23952
rect -12613 -24014 -12517 -23951
rect -12736 -24016 -12578 -24014
rect -12738 -24092 -12574 -24076
rect -12738 -24163 -12685 -24092
rect -12614 -24163 -12477 -24092
rect -12738 -24164 -12574 -24163
rect -10695 -24593 -10606 -22334
rect -6030 -24356 -5982 -18656
rect -6032 -24362 -5980 -24356
rect -5852 -24358 -5804 -18176
rect -5700 -22398 -5652 -17716
rect -5584 -20422 -5536 -17256
rect -5592 -20474 -5586 -20422
rect -5534 -20474 -5528 -20422
rect -5702 -22404 -5650 -22398
rect -5702 -22462 -5650 -22456
rect -5860 -24410 -5854 -24358
rect -5802 -24410 -5796 -24358
rect -6032 -24420 -5980 -24414
rect -5396 -24593 -5307 -17252
rect -5234 -17314 -5186 -16776
rect -4056 -16942 -3972 -16888
rect -4056 -16980 -3908 -16942
rect -4056 -17064 -2524 -16980
rect 816 -16996 900 -16992
rect -5236 -17320 -5184 -17314
rect -5236 -17378 -5184 -17372
rect -4062 -17791 -2674 -17707
rect -4052 -18610 -2830 -18526
rect -4078 -19429 -2998 -19345
rect -5174 -20056 -5074 -20044
rect -5174 -20128 -5166 -20056
rect -5094 -20128 -5074 -20056
rect -5174 -20134 -5074 -20128
rect -5166 -20202 -5094 -20134
rect -5166 -20274 -4972 -20202
rect -4052 -20248 -3176 -20164
rect -4064 -21046 -3822 -20983
rect -4064 -21067 -3906 -21046
rect -3906 -21136 -3822 -21130
rect -5130 -21525 -5047 -21519
rect -5130 -22437 -5047 -21608
rect -5140 -22520 -5047 -22437
rect -10695 -24682 -5298 -24593
rect -5396 -24688 -5307 -24682
rect -5130 -24796 -5047 -22520
rect -10647 -24879 -5047 -24796
rect -10647 -24987 -10563 -24879
rect -10920 -25070 -10563 -24987
rect -6038 -25036 -6032 -24984
rect -5980 -25036 -5974 -24984
rect -13016 -25112 -12964 -25106
rect -13016 -25170 -12964 -25164
rect -10479 -25107 -10393 -25096
rect -17964 -25350 -17878 -25344
rect -17964 -25422 -17956 -25350
rect -17884 -25422 -17878 -25350
rect -17964 -25428 -17878 -25422
rect -17982 -25553 -17878 -25480
rect -17982 -25642 -17976 -25553
rect -17887 -25642 -17878 -25553
rect -17982 -25650 -17878 -25642
rect -12770 -26744 -12612 -26742
rect -12770 -26805 -12743 -26744
rect -12682 -26805 -12480 -26744
rect -12770 -26806 -12612 -26805
rect -12794 -26998 -12748 -26934
rect -12684 -26998 -12472 -26934
rect -10479 -27674 -10393 -25193
rect -10865 -27760 -10393 -27674
rect -10152 -25530 -10048 -25524
rect -10152 -27954 -10048 -25634
rect -10366 -28058 -10048 -27954
rect -12758 -29446 -12724 -29374
rect -12652 -29446 -12468 -29374
rect -12772 -29537 -12586 -29520
rect -12772 -29626 -12727 -29537
rect -12638 -29626 -12432 -29537
rect -10366 -30233 -10262 -28058
rect -10883 -30337 -10262 -30233
rect -12834 -31918 -12670 -31900
rect -12834 -31990 -12758 -31918
rect -12686 -31990 -12478 -31918
rect -12838 -32087 -12674 -32086
rect -12838 -32176 -12791 -32087
rect -12702 -32176 -12464 -32087
rect -10915 -33009 -9857 -32916
rect -9764 -33009 -9758 -32916
rect -6030 -33110 -5982 -25036
rect -5860 -25086 -5854 -25034
rect -5802 -25086 -5796 -25034
rect -5852 -25742 -5804 -25086
rect -5860 -25794 -5854 -25742
rect -5802 -25794 -5796 -25742
rect -6032 -33116 -5980 -33110
rect -6032 -33174 -5980 -33168
rect -3260 -33272 -3176 -20248
rect -3082 -25874 -2998 -19429
rect -2914 -22526 -2830 -18610
rect -2751 -21748 -2680 -17791
rect -2608 -17980 -2524 -17064
rect -1344 -17080 914 -16996
rect 674 -17086 758 -17080
rect 816 -17812 900 -17080
rect 674 -17815 758 -17812
rect -1302 -17899 758 -17815
rect -2608 -18070 -2524 -18064
rect -1340 -18718 574 -18634
rect -1366 -19537 404 -19453
rect -413 -19617 -347 -19611
rect -2426 -20128 -2420 -20056
rect -2348 -20128 -2342 -20056
rect -2420 -20170 -2348 -20128
rect -2420 -20232 -2320 -20170
rect -2420 -20304 -2266 -20232
rect -1354 -20356 -614 -20272
rect -2751 -21825 -2680 -21819
rect -2914 -22616 -2830 -22610
rect -3082 -25964 -2998 -25958
rect -3260 -33362 -3176 -33356
rect -698 -33494 -614 -20356
rect -698 -33584 -614 -33578
rect -413 -33801 -347 -19683
rect 320 -26064 404 -19537
rect 490 -22696 574 -18718
rect 674 -21872 758 -17899
rect 816 -17902 900 -17896
rect 674 -21962 758 -21956
rect 484 -22780 490 -22696
rect 574 -22780 580 -22696
rect 320 -26154 404 -26148
rect 1078 -29278 1137 -16765
rect 1221 -21389 1287 -16623
rect 1367 -20217 1433 -16475
rect 1367 -20289 1433 -20283
rect 3886 -21046 3970 -1635
rect 4164 -1602 4248 -1596
rect 4164 -13666 4248 -1686
rect 4158 -13750 4164 -13666
rect 4248 -13750 4254 -13666
rect 3880 -21130 3886 -21046
rect 3970 -21130 3976 -21046
rect 1215 -21455 1221 -21389
rect 1287 -21455 1293 -21389
rect 4427 -28308 4493 -1375
rect 4573 -28064 4639 -1204
rect 4838 -17961 4904 -1014
rect 4948 -15747 5014 -851
rect 5096 -13052 5162 -684
rect 5261 -6685 5327 -487
rect 5419 -6437 5485 -298
rect 13190 -2964 15683 -2934
rect 13169 -3000 15683 -2964
rect 13169 -3047 13216 -3000
rect 5413 -6503 5419 -6437
rect 5485 -6503 5491 -6437
rect 5261 -6751 5492 -6685
rect 5426 -11065 5492 -6751
rect 13172 -7413 13219 -7330
rect 13180 -7481 15547 -7415
rect 5426 -11137 5492 -11131
rect 13139 -12012 15435 -11946
rect 13183 -12104 13230 -12021
rect 5096 -13118 5354 -13052
rect 5420 -13118 5426 -13052
rect 4948 -15813 5473 -15747
rect 5407 -17552 5473 -15813
rect 13178 -16518 13225 -16463
rect 13178 -16546 15223 -16518
rect 13193 -16584 15223 -16546
rect 5401 -17619 5407 -17552
rect 5473 -17619 5479 -17552
rect 15157 -17570 15223 -16584
rect 15369 -17476 15435 -12012
rect 15481 -17382 15547 -7481
rect 15617 -17354 15683 -3000
rect 15481 -17448 15683 -17382
rect 15369 -17542 15683 -17476
rect 15157 -17636 15683 -17570
rect 4838 -18027 5471 -17961
rect 4745 -21389 4811 -21383
rect 4811 -21455 5319 -21389
rect 4745 -21461 4811 -21455
rect 5253 -24739 5319 -21455
rect 5405 -24649 5471 -18027
rect 18354 -18573 18391 -18471
rect 15066 -19602 15699 -19536
rect 13181 -21039 13228 -21034
rect 15066 -21039 15132 -19602
rect 13181 -21105 15132 -21039
rect 15261 -19696 15685 -19630
rect 13181 -21117 13228 -21105
rect 5732 -24649 5798 -24643
rect 5405 -24715 5732 -24649
rect 5732 -24721 5798 -24715
rect 5253 -24745 5383 -24739
rect 5253 -24811 5317 -24745
rect 5317 -24817 5383 -24811
rect 15261 -25506 15327 -19696
rect 13186 -25531 15327 -25506
rect 13179 -25572 15327 -25531
rect 15447 -19790 15683 -19724
rect 13179 -25614 13226 -25572
rect 4573 -28130 5520 -28064
rect 4427 -28374 5329 -28308
rect 1078 -29337 4860 -29278
rect 4919 -29337 4925 -29278
rect 5263 -29395 5329 -28374
rect 5454 -29177 5520 -28130
rect 5454 -29249 5520 -29243
rect 5263 -29461 5491 -29395
rect 5425 -33705 5491 -29461
rect 15447 -30040 15513 -19790
rect 13153 -30106 15513 -30040
rect 5425 -33777 5491 -33771
rect 3663 -33801 3729 -33795
rect -413 -33867 3663 -33801
rect 3663 -33873 3729 -33867
rect -12588 -34576 -12582 -34504
rect -12510 -34576 -12504 -34504
rect 15619 -34535 15685 -19818
rect 13156 -34601 15685 -34535
rect -12746 -34671 -12582 -34670
rect -12746 -34760 -12726 -34671
rect -12637 -34760 -12476 -34671
rect 13144 -34776 13232 -34666
rect 13151 -35666 13235 -34780
rect 13035 -36363 13082 -36280
<< via1 >>
rect -21815 6595 -21726 6684
rect -27525 4452 -27436 4541
rect -22632 4418 -22560 4490
rect -15130 6556 -15022 6664
rect -19312 6376 -19240 6448
rect -18528 6279 -18439 6368
rect -16019 6124 -15947 6196
rect -15230 5884 -15141 5973
rect -12742 5681 -12670 5753
rect -11940 5537 -11851 5626
rect -9439 5385 -9367 5457
rect 3195 5390 3247 5442
rect -8640 5227 -8551 5316
rect -6166 5269 -6096 5339
rect -5351 4991 -5262 5080
rect -2875 4746 -2803 4818
rect 425 4612 497 4684
rect -2058 4473 -1969 4562
rect 2921 4209 2987 4275
rect 4885 4209 4951 4275
rect 5339 4011 5411 4083
rect 1934 2453 2000 2519
rect -21801 218 -21735 284
rect -25060 -214 -24969 -123
rect -15223 230 -15157 296
rect -11963 223 -11897 289
rect -8633 243 -8567 309
rect -5349 226 -5283 292
rect -2061 195 -1995 261
rect 6966 2147 7032 2213
rect 6953 1045 7019 1111
rect 248 -131 339 -40
rect 1625 -1375 1691 -1309
rect 3886 -1635 3970 -1551
rect -7873 -6291 -7807 -6225
rect -5439 -6599 -5373 -6533
rect -24837 -11059 -24748 -10970
rect -5043 -11227 -4977 -11161
rect -7799 -12909 -7688 -12798
rect -11151 -13445 -11085 -13379
rect -768 -12902 -684 -12818
rect -14443 -13643 -14377 -13577
rect -5286 -13312 -5233 -13259
rect -5814 -13492 -5730 -13408
rect -17730 -13759 -17671 -13700
rect -4626 -13818 -4542 -13734
rect -1201 -13750 -1117 -13666
rect -14808 -13976 -14756 -13924
rect -21025 -14541 -20959 -14475
rect -24916 -15658 -24844 -15586
rect -24903 -15828 -24812 -15739
rect -24908 -16842 -24836 -16770
rect -24925 -17012 -24836 -16923
rect -24921 -18054 -24851 -17984
rect -20399 -17986 -20347 -17934
rect -24917 -18217 -24824 -18128
rect -20414 -18486 -20356 -18434
rect -17966 -15658 -17894 -15586
rect -18123 -15827 -18034 -15738
rect -18082 -17052 -18010 -16980
rect -18089 -17202 -18000 -17113
rect -5370 -13928 -5318 -13876
rect -14708 -14140 -14656 -14088
rect -10855 -14108 -10779 -14032
rect -5963 -14065 -5881 -13983
rect -6954 -14194 -6902 -14142
rect -10850 -14386 -10795 -14331
rect -12724 -15658 -12652 -15586
rect -12555 -15837 -12456 -15738
rect -14612 -16016 -14560 -15964
rect -18065 -18455 -17995 -18385
rect -18099 -18604 -18010 -18515
rect -19377 -18771 -19311 -18705
rect -14496 -16238 -14444 -16186
rect -20399 -18966 -20347 -18914
rect -24870 -19175 -24798 -19103
rect -24889 -19345 -24796 -19256
rect -10307 -14826 -10252 -14771
rect -6834 -14542 -6782 -14490
rect -8676 -15568 -8604 -15496
rect -5008 -14566 -4936 -14494
rect -3899 -14557 -3833 -14491
rect -6664 -14922 -6612 -14870
rect -8554 -16224 -8482 -16152
rect -4966 -15378 -4894 -15306
rect -2288 -14566 -2216 -14494
rect -2264 -15378 -2192 -15306
rect -4995 -16195 -4925 -16125
rect -2285 -16195 -2215 -16125
rect -8551 -16754 -8482 -16685
rect 407 -15493 473 -15427
rect -12666 -18468 -12594 -18396
rect -12633 -18662 -12544 -18573
rect -20404 -19466 -20352 -19414
rect -8549 -17274 -8480 -17205
rect -5397 -17243 -5307 -17154
rect -8554 -17684 -8485 -17615
rect -8554 -18166 -8485 -18097
rect -8554 -18636 -8485 -18567
rect -8584 -19170 -8512 -19098
rect -18016 -19685 -17953 -19622
rect -20324 -19946 -20272 -19894
rect -17986 -19978 -17915 -19907
rect -14808 -19918 -14756 -19866
rect -24936 -20363 -24864 -20291
rect -20399 -20406 -20347 -20354
rect -24902 -20533 -24811 -20444
rect -18572 -20866 -18520 -20814
rect -18053 -21237 -17992 -21176
rect -18692 -21346 -18640 -21294
rect -17968 -21404 -17904 -21340
rect -24924 -21569 -24852 -21497
rect -24913 -21739 -24823 -21650
rect -18061 -22666 -17995 -22600
rect -24890 -22870 -24818 -22798
rect -18071 -22834 -17982 -22745
rect -24913 -23040 -24819 -22951
rect -18042 -24058 -17970 -23986
rect -24926 -24180 -24854 -24108
rect -18063 -24220 -17974 -24131
rect -24907 -24350 -24813 -24261
rect -12609 -21437 -12539 -21367
rect -12628 -21616 -12539 -21527
rect -12750 -22150 -12698 -22098
rect -12872 -22336 -12820 -22284
rect -12676 -24014 -12613 -23951
rect -12685 -24163 -12614 -24092
rect -5586 -20474 -5534 -20422
rect -5702 -22456 -5650 -22404
rect -6032 -24414 -5980 -24362
rect -5854 -24410 -5802 -24358
rect -5000 -17021 -4937 -16958
rect -2291 -17021 -2228 -16958
rect -5236 -17372 -5184 -17320
rect -4979 -17841 -4918 -17780
rect -5006 -18654 -4934 -18582
rect -5014 -19502 -4942 -19430
rect -5166 -20128 -5094 -20056
rect -3906 -21130 -3822 -21046
rect -5130 -21608 -5047 -21525
rect -6032 -25036 -5980 -24984
rect -13016 -25164 -12964 -25112
rect -10479 -25193 -10393 -25107
rect -17956 -25422 -17884 -25350
rect -17976 -25642 -17887 -25553
rect -12743 -26805 -12682 -26744
rect -12748 -26998 -12684 -26934
rect -10152 -25634 -10048 -25530
rect -12724 -29446 -12652 -29374
rect -12727 -29626 -12638 -29537
rect -12758 -31990 -12686 -31918
rect -12791 -32176 -12702 -32087
rect -9857 -33009 -9764 -32916
rect -5854 -25086 -5802 -25034
rect -5854 -25794 -5802 -25742
rect -6032 -33168 -5980 -33116
rect -2269 -17841 -2208 -17780
rect -2608 -18064 -2524 -17980
rect -2294 -18654 -2222 -18582
rect -2300 -19502 -2228 -19430
rect -413 -19683 -347 -19617
rect -2420 -20128 -2348 -20056
rect -2751 -21819 -2680 -21748
rect -2914 -22610 -2830 -22526
rect -3082 -25958 -2998 -25874
rect -3260 -33356 -3176 -33272
rect -698 -33578 -614 -33494
rect 816 -17896 900 -17812
rect 674 -21956 758 -21872
rect 490 -22780 574 -22696
rect 320 -26148 404 -26064
rect 1367 -20283 1433 -20217
rect 4164 -1686 4248 -1602
rect 4164 -13750 4248 -13666
rect 3886 -21130 3970 -21046
rect 1221 -21455 1287 -21389
rect 5419 -6503 5485 -6437
rect 5426 -11131 5492 -11065
rect 5354 -13118 5420 -13052
rect 5407 -17619 5473 -17552
rect 4745 -21455 4811 -21389
rect 5732 -24715 5798 -24649
rect 5317 -24811 5383 -24745
rect 4860 -29337 4919 -29278
rect 5454 -29243 5520 -29177
rect 5425 -33771 5491 -33705
rect 3663 -33867 3729 -33801
rect -12582 -34576 -12510 -34504
rect -12726 -34760 -12637 -34671
<< metal2 >>
rect -22627 7080 -22565 7084
rect -22632 7075 -22560 7080
rect -22632 7013 -22627 7075
rect -22565 7013 -22560 7075
rect -27531 4452 -27525 4541
rect -27436 4452 -27430 4541
rect -22632 4490 -22560 7013
rect -21840 6812 -17646 6920
rect -21840 6809 -21732 6812
rect -21840 6730 -21811 6809
rect -21840 6700 -21732 6730
rect -21840 6684 -21712 6700
rect -21840 6595 -21815 6684
rect -21726 6595 -21712 6684
rect -17754 6664 -17646 6812
rect -19307 6655 -19245 6659
rect -21840 6592 -21712 6595
rect -19312 6650 -19240 6655
rect -21840 6589 -21726 6592
rect -21840 6544 -21732 6589
rect -19312 6588 -19307 6650
rect -19245 6588 -19240 6650
rect -19312 6448 -19240 6588
rect -17754 6556 -15130 6664
rect -15022 6556 -15016 6664
rect -18524 6501 -18445 6505
rect -19312 6370 -19240 6376
rect -18528 6496 -18439 6501
rect -18528 6417 -18524 6496
rect -18445 6417 -18439 6496
rect -18528 6368 -18439 6417
rect -16019 6304 -15947 6309
rect -18528 6273 -18439 6279
rect -16023 6242 -16014 6304
rect -15952 6242 -15943 6304
rect -16019 6196 -15947 6242
rect -15226 6155 -15147 6159
rect -16019 6118 -15947 6124
rect -15230 6150 -15141 6155
rect -15230 6071 -15226 6150
rect -15147 6071 -15141 6150
rect -15230 5973 -15141 6071
rect -12737 5978 -12675 5982
rect -15230 5878 -15141 5884
rect -12742 5973 -12670 5978
rect -12742 5911 -12737 5973
rect -12675 5911 -12670 5973
rect -12742 5753 -12670 5911
rect -11940 5784 -11851 5789
rect -11945 5705 -11936 5784
rect -11857 5705 -11848 5784
rect -12742 5675 -12670 5681
rect -11940 5626 -11851 5705
rect -9434 5613 -9372 5617
rect -11940 5531 -11851 5537
rect -9439 5608 -9367 5613
rect -9439 5546 -9434 5608
rect -9372 5546 -9367 5608
rect -9439 5457 -9367 5546
rect -8636 5486 -8557 5490
rect -9439 5379 -9367 5385
rect -8640 5481 -8551 5486
rect -8640 5402 -8636 5481
rect -8557 5402 -8551 5481
rect -8640 5316 -8551 5402
rect 3195 5442 3247 5448
rect 3195 5384 3247 5390
rect -6173 5339 -6084 5346
rect -6173 5269 -6166 5339
rect -6096 5269 -6084 5339
rect -6173 5261 -6084 5269
rect -8640 5221 -8551 5227
rect -5363 5202 -5253 5215
rect -5363 5123 -5353 5202
rect -5268 5123 -5253 5202
rect -5363 5113 -5253 5123
rect -5351 5080 -5262 5113
rect -2870 5028 -2808 5032
rect -5351 4985 -5262 4991
rect -2875 5023 -2803 5028
rect -2875 4961 -2870 5023
rect -2808 4961 -2803 5023
rect -2875 4818 -2803 4961
rect -2054 4881 -1975 4885
rect -2875 4740 -2803 4746
rect -2058 4876 -1969 4881
rect -2058 4797 -2054 4876
rect -1975 4797 -1969 4876
rect -2058 4562 -1969 4797
rect 430 4726 492 4730
rect 425 4721 497 4726
rect 425 4684 430 4721
rect 492 4684 497 4721
rect 425 4606 497 4612
rect -2058 4467 -1969 4473
rect -22632 4412 -22560 4418
rect 1625 4209 2921 4275
rect 2987 4209 2993 4275
rect -21807 218 -21801 284
rect -21735 218 -21729 284
rect -15229 230 -15223 296
rect -15157 230 -15151 296
rect -11963 289 -11897 295
rect -8639 243 -8633 309
rect -8567 243 -8561 309
rect -5355 226 -5349 292
rect -5283 226 -5277 292
rect -11963 217 -11897 223
rect -2067 195 -2061 261
rect -1995 195 -1989 261
rect -25060 -123 -24969 -117
rect 242 -123 248 -40
rect -24969 -131 248 -123
rect 339 -131 345 -40
rect -24969 -214 339 -131
rect -25060 -220 -24969 -214
rect 1225 -2009 1291 379
rect 1625 -1298 1691 4209
rect 3198 4128 3243 5384
rect 4922 5187 4978 5188
rect 4885 5060 4978 5187
rect 4885 4275 4951 5060
rect 4879 4209 4885 4275
rect 4951 4209 4957 4275
rect 3198 4083 5411 4128
rect 5333 4011 5339 4083
rect 5411 4011 5417 4083
rect 6436 4022 6445 4081
rect 6504 4022 6513 4081
rect 5339 3863 5411 4011
rect 1934 2519 2000 2525
rect 2000 2453 5811 2519
rect 1934 2447 2000 2453
rect 6576 2215 6642 2423
rect 6576 2149 6683 2215
rect 6617 923 6683 2149
rect 6947 1045 6953 1111
rect 7019 1045 7025 1111
rect 3886 825 5825 891
rect 1618 -1309 1704 -1298
rect 1618 -1375 1625 -1309
rect 1691 -1375 1704 -1309
rect 1618 -1380 1704 -1375
rect 3886 -1551 3970 825
rect 4166 733 5815 770
rect 4164 704 5815 733
rect 3880 -1635 3886 -1551
rect 3970 -1635 3976 -1551
rect 4164 -1602 4248 704
rect 5554 -509 5563 -450
rect 5622 -509 5631 -450
rect 5994 -483 6003 -424
rect 6062 -483 6071 -424
rect 6434 -514 6443 -455
rect 6502 -514 6511 -455
rect 4158 -1686 4164 -1602
rect 4248 -1686 4254 -1602
rect 1225 -2075 5821 -2009
rect -8187 -2171 5798 -2105
rect -25216 -2524 -25155 -2520
rect -25220 -2529 -24499 -2524
rect -25220 -2591 -25216 -2529
rect -25155 -2591 -24499 -2529
rect -25220 -2595 -24499 -2591
rect -25216 -2600 -25155 -2595
rect -8187 -3159 -8121 -2171
rect -6334 -2274 5796 -2226
rect -25512 -5030 -25432 -5026
rect -25060 -5030 -24340 -4997
rect -25512 -5035 -24340 -5030
rect -25512 -5097 -25504 -5035
rect -25442 -5097 -24340 -5035
rect -25512 -5102 -24340 -5097
rect -25512 -5106 -25432 -5102
rect -25060 -5133 -24340 -5102
rect -7873 -6225 -7807 -6219
rect -7873 -6297 -7807 -6291
rect -25655 -6746 -25576 -6742
rect -25659 -6751 -24378 -6746
rect -25659 -6832 -25655 -6751
rect -25576 -6832 -24378 -6751
rect -25659 -6835 -24378 -6832
rect -25655 -6841 -25576 -6835
rect -25809 -8297 -25749 -8293
rect -25814 -8302 -24463 -8297
rect -25814 -8362 -25809 -8302
rect -25749 -8362 -24463 -8302
rect -25814 -8367 -24463 -8362
rect -25809 -8371 -25749 -8367
rect -25990 -10155 -25880 -10146
rect -25305 -10155 -23050 -10101
rect -25990 -10160 -23050 -10155
rect -25990 -10241 -25978 -10160
rect -25899 -10236 -23050 -10160
rect -25899 -10241 -25048 -10236
rect -25990 -10244 -25048 -10241
rect -25990 -10252 -25880 -10244
rect -25369 -10976 -24837 -10970
rect -25374 -11055 -25365 -10976
rect -25286 -11055 -24837 -10976
rect -25369 -11059 -24837 -11055
rect -24748 -11059 -24742 -10970
rect -23185 -10997 -23050 -10236
rect -23185 -11132 -22869 -10997
rect -26164 -11586 -26102 -11582
rect -26169 -11591 -24520 -11586
rect -26169 -11653 -26164 -11591
rect -26102 -11653 -24520 -11591
rect -26169 -11658 -24520 -11653
rect -26164 -11662 -26102 -11658
rect -22912 -13016 -22744 -13010
rect -26340 -13054 -22744 -13016
rect -26340 -13063 -22742 -13054
rect -26340 -13144 -26327 -13063
rect -26248 -13144 -22742 -13063
rect -26340 -13184 -22742 -13144
rect -21025 -14475 -20959 -12899
rect -17730 -13700 -17671 -12825
rect -14443 -13577 -14377 -12821
rect -11151 -13379 -11085 -12783
rect -7805 -12909 -7799 -12798
rect -7688 -12909 -7682 -12798
rect -11151 -13451 -11085 -13445
rect -14443 -13649 -14377 -13643
rect -17730 -13765 -17671 -13759
rect -6334 -13840 -6286 -2274
rect -20148 -13888 -6286 -13840
rect -6254 -2376 5858 -2328
rect -21031 -14541 -21025 -14475
rect -20959 -14541 -20953 -14475
rect -24936 -15658 -24916 -15586
rect -24844 -15658 -24820 -15586
rect -24936 -15739 -24800 -15738
rect -24936 -15828 -24903 -15739
rect -24812 -15828 -24800 -15739
rect -24920 -16842 -24908 -16770
rect -24836 -16842 -24820 -16770
rect -24925 -16923 -24836 -16917
rect -24836 -17012 -24827 -16923
rect -24925 -17018 -24836 -17012
rect -20399 -17934 -20347 -17928
rect -24921 -17982 -24851 -17978
rect -24934 -17984 -24834 -17982
rect -24934 -18054 -24921 -17984
rect -24851 -18054 -24834 -17984
rect -20148 -17936 -20100 -13888
rect -14808 -13920 -14756 -13918
rect -6254 -13920 -6206 -2376
rect -14808 -13924 -6206 -13920
rect -20347 -17984 -20100 -17936
rect -20070 -13988 -14888 -13940
rect -14756 -13968 -6206 -13924
rect -6160 -3486 6238 -3426
rect -14808 -13982 -14756 -13976
rect -20399 -17992 -20347 -17986
rect -24921 -18060 -24851 -18054
rect -24936 -18128 -24806 -18126
rect -24936 -18217 -24917 -18128
rect -24824 -18217 -24806 -18128
rect -24936 -18218 -24806 -18217
rect -20408 -18434 -20356 -18428
rect -20420 -18486 -20414 -18434
rect -20070 -18436 -20022 -13988
rect -14936 -14010 -14888 -13988
rect -20356 -18484 -20022 -18436
rect -19958 -14084 -14970 -14036
rect -14936 -14058 -10918 -14010
rect -6160 -14032 -6100 -3486
rect -6062 -3584 5820 -3536
rect -20408 -18492 -20356 -18486
rect -20406 -18914 -20340 -18908
rect -20406 -18966 -20399 -18914
rect -20347 -18916 -20340 -18914
rect -19958 -18916 -19910 -14084
rect -15018 -14170 -14970 -14084
rect -14714 -14140 -14708 -14088
rect -14656 -14090 -14650 -14088
rect -14656 -14138 -11022 -14090
rect -14656 -14140 -14650 -14138
rect -15018 -14218 -12652 -14170
rect -12700 -15454 -12652 -14218
rect -11070 -14250 -11022 -14138
rect -10966 -14152 -10918 -14058
rect -10861 -14108 -10855 -14032
rect -10779 -14108 -6092 -14032
rect -6062 -14136 -6014 -3584
rect -5959 -3703 5798 -3637
rect -5959 -3793 -5893 -3703
rect -5963 -13983 -5881 -3793
rect -5799 -3824 5799 -3758
rect -5799 -4072 -5733 -3824
rect -5814 -13408 -5730 -4072
rect 5554 -4919 5563 -4860
rect 5622 -4919 5631 -4860
rect 5994 -4939 6003 -4880
rect 6062 -4939 6071 -4880
rect 6433 -4948 6442 -4889
rect 6501 -4948 6510 -4889
rect 5419 -6432 5485 -6431
rect 5412 -6437 5485 -6432
rect 5412 -6503 5419 -6437
rect 5485 -6503 5798 -6437
rect 5412 -6504 5485 -6503
rect -5445 -6599 -5439 -6533
rect -5373 -6599 5819 -6533
rect -5694 -6639 -5646 -6638
rect -5694 -6705 5798 -6639
rect -5820 -13492 -5814 -13408
rect -5730 -13492 -5724 -13408
rect -5963 -14071 -5881 -14065
rect -6958 -14142 -6014 -14136
rect -10966 -14200 -7014 -14152
rect -6960 -14194 -6954 -14142
rect -6902 -14184 -6014 -14142
rect -6902 -14194 -6896 -14184
rect -7062 -14232 -7014 -14200
rect -5694 -14232 -5646 -6705
rect -5615 -6766 5798 -6743
rect -11070 -14298 -7108 -14250
rect -7062 -14280 -5646 -14232
rect -5616 -6809 5798 -6766
rect -7156 -14314 -7108 -14298
rect -5616 -14314 -5568 -6809
rect -5507 -7847 5798 -7845
rect -10856 -14386 -10850 -14331
rect -10795 -14386 -7187 -14331
rect -7156 -14362 -5568 -14314
rect -5536 -7911 5798 -7847
rect -7242 -14402 -7187 -14386
rect -5536 -14402 -5481 -7911
rect -5451 -8033 5798 -7967
rect -12114 -14474 -7308 -14426
rect -7242 -14457 -5481 -14402
rect -12114 -15454 -12066 -14474
rect -7356 -14586 -7308 -14474
rect -5450 -14490 -5398 -8033
rect -5367 -8131 5798 -8065
rect -5366 -13870 -5322 -8131
rect -5286 -8186 -5233 -8180
rect -5286 -8252 5798 -8186
rect -5286 -13259 -5233 -8252
rect 5554 -9582 5563 -9523
rect 5622 -9582 5631 -9523
rect 5994 -9587 6003 -9528
rect 6062 -9587 6071 -9528
rect 6436 -9573 6445 -9514
rect 6504 -9573 6513 -9514
rect 5420 -11131 5426 -11065
rect 5492 -11131 5803 -11065
rect -5049 -11227 -5043 -11161
rect -4977 -11227 5798 -11161
rect -5195 -11276 5798 -11267
rect -5286 -13318 -5233 -13312
rect -5200 -11333 5798 -11276
rect -5200 -13382 -5152 -11333
rect -5115 -11379 5798 -11371
rect -5284 -13430 -5152 -13382
rect -5116 -11437 5798 -11379
rect -5370 -13876 -5318 -13870
rect -5370 -13934 -5318 -13928
rect -5284 -13988 -5236 -13430
rect -5116 -13469 -5061 -11437
rect -6840 -14542 -6834 -14490
rect -6782 -14542 -5398 -14490
rect -5368 -14036 -5236 -13988
rect -5196 -13524 -5061 -13469
rect -5022 -12473 -4974 -12472
rect -5022 -12539 5798 -12473
rect -5368 -14586 -5320 -14036
rect -5196 -14083 -5141 -13524
rect -5022 -13566 -4974 -12539
rect -7356 -14634 -5320 -14586
rect -5284 -14138 -5141 -14083
rect -5108 -13614 -4974 -13566
rect -4796 -12595 -4748 -12592
rect -4796 -12661 5839 -12595
rect -5284 -14685 -5229 -14138
rect -5108 -14180 -5060 -13614
rect -10150 -14690 -5229 -14685
rect -12700 -15502 -12066 -15454
rect -10606 -14738 -5229 -14690
rect -17978 -15586 -17880 -15576
rect -17978 -15658 -17966 -15586
rect -17894 -15658 -17880 -15586
rect -17978 -15666 -17880 -15658
rect -12734 -15586 -12608 -15552
rect -12734 -15658 -12724 -15586
rect -12652 -15658 -12608 -15586
rect -12734 -15672 -12608 -15658
rect -18130 -15738 -18026 -15730
rect -18130 -15827 -18123 -15738
rect -18034 -15827 -18026 -15738
rect -18130 -15836 -18026 -15827
rect -12566 -15738 -12440 -15728
rect -12566 -15837 -12555 -15738
rect -12456 -15837 -12440 -15738
rect -12566 -15848 -12440 -15837
rect -14612 -15964 -14560 -15958
rect -10606 -15966 -10558 -14738
rect -10150 -14740 -5229 -14738
rect -5194 -14228 -5060 -14180
rect -10313 -14826 -10307 -14771
rect -10252 -14778 -6429 -14771
rect -5194 -14778 -5146 -14228
rect -5020 -14494 -4926 -14484
rect -5020 -14566 -5008 -14494
rect -4936 -14566 -4926 -14494
rect -5020 -14576 -4926 -14566
rect -4796 -14726 -4748 -12661
rect -4633 -12759 5798 -12693
rect -4626 -13734 -4542 -12759
rect -774 -12902 -768 -12818
rect -684 -12902 5792 -12818
rect 5354 -13052 5420 -13046
rect 4164 -13666 4248 -13660
rect -1207 -13750 -1201 -13666
rect -1117 -13750 4164 -13666
rect 4164 -13756 4248 -13750
rect -4626 -13824 -4542 -13818
rect -3912 -14491 -3812 -14472
rect -3912 -14557 -3899 -14491
rect -3833 -14557 -3812 -14491
rect -3912 -14574 -3812 -14557
rect -2296 -14494 -2202 -14482
rect -2296 -14566 -2288 -14494
rect -2216 -14566 -2202 -14494
rect -2296 -14574 -2202 -14566
rect -10252 -14826 -5146 -14778
rect -5110 -14774 -4748 -14726
rect -6674 -14870 -6600 -14860
rect -6674 -14922 -6664 -14870
rect -6612 -14872 -6600 -14870
rect -5110 -14872 -5062 -14774
rect -6612 -14920 -5062 -14872
rect -6612 -14922 -6600 -14920
rect -6674 -14930 -6600 -14922
rect -4974 -15306 -4880 -15294
rect -8690 -15496 -8594 -15486
rect -8690 -15568 -8676 -15496
rect -8604 -15568 -8594 -15496
rect -8690 -15588 -8594 -15568
rect -6114 -15533 -6066 -15372
rect -4974 -15378 -4966 -15306
rect -4894 -15378 -4880 -15306
rect -4974 -15386 -4880 -15378
rect -2276 -15306 -2182 -15296
rect -2276 -15378 -2264 -15306
rect -2192 -15378 -2182 -15306
rect -2276 -15388 -2182 -15378
rect 401 -15493 407 -15427
rect 473 -15493 4595 -15427
rect -6114 -15599 4429 -15533
rect -6114 -15644 -6066 -15599
rect -14560 -16014 -10558 -15966
rect -10500 -15692 -6066 -15644
rect -14612 -16022 -14560 -16016
rect -10500 -16086 -10452 -15692
rect -20347 -18964 -19910 -18916
rect -19848 -16134 -10452 -16086
rect -10410 -15772 -5990 -15724
rect -20347 -18966 -20340 -18964
rect -20406 -18972 -20340 -18966
rect -24870 -19102 -24798 -19097
rect -24892 -19103 -24778 -19102
rect -24892 -19175 -24870 -19103
rect -24798 -19175 -24778 -19103
rect -24892 -19176 -24778 -19175
rect -24870 -19181 -24798 -19176
rect -24916 -19345 -24889 -19256
rect -24796 -19345 -24780 -19256
rect -24916 -19346 -24780 -19345
rect -20404 -19414 -20352 -19408
rect -19848 -19416 -19800 -16134
rect -14502 -16238 -14496 -16186
rect -14444 -16188 -14438 -16186
rect -10410 -16188 -10362 -15772
rect -6038 -15930 -5990 -15772
rect 4363 -15795 4429 -15599
rect 4529 -15689 4595 -15493
rect 5354 -15593 5420 -13118
rect 5554 -14109 5563 -14050
rect 5622 -14109 5631 -14050
rect 5994 -14093 6003 -14034
rect 6062 -14093 6071 -14034
rect 6433 -14076 6442 -14017
rect 6501 -14076 6510 -14017
rect 5354 -15659 5798 -15593
rect 4529 -15755 5809 -15689
rect 4363 -15861 5815 -15795
rect -6038 -15952 -3582 -15930
rect 4366 -15952 5918 -15920
rect -6038 -15968 5918 -15952
rect -6038 -15978 4414 -15968
rect -3647 -16000 4414 -15978
rect -5002 -16125 -4908 -16110
rect -14444 -16236 -10362 -16188
rect -8570 -16152 -8470 -16140
rect -8570 -16224 -8554 -16152
rect -8482 -16224 -8470 -16152
rect -5002 -16195 -4995 -16125
rect -4925 -16195 -4908 -16125
rect -5002 -16202 -4908 -16195
rect -2294 -16125 -2200 -16114
rect -2294 -16195 -2285 -16125
rect -2215 -16195 -2200 -16125
rect -2294 -16206 -2200 -16195
rect -8570 -16236 -8470 -16224
rect -14444 -16238 -14438 -16236
rect -8566 -16685 -8470 -16670
rect -8566 -16754 -8551 -16685
rect -8482 -16754 -8470 -16685
rect -8566 -16768 -8470 -16754
rect -5010 -16958 -4916 -16940
rect -18077 -16980 -18015 -16976
rect -18088 -17052 -18082 -16980
rect -18010 -17052 -18004 -16980
rect -5010 -17021 -5000 -16958
rect -4937 -17021 -4916 -16958
rect -5010 -17032 -4916 -17021
rect -2298 -16958 -2204 -16938
rect -2298 -17021 -2291 -16958
rect -2228 -17021 -2204 -16958
rect -2298 -17030 -2204 -17021
rect -18077 -17056 -18015 -17052
rect 1537 -17067 5798 -16982
rect -18096 -17113 -17992 -17102
rect -18096 -17202 -18089 -17113
rect -18000 -17202 -17992 -17113
rect -5407 -17154 -5288 -17149
rect 1537 -17154 1622 -17067
rect -18096 -17208 -17992 -17202
rect -8560 -17205 -8464 -17188
rect -8560 -17274 -8549 -17205
rect -8480 -17274 -8464 -17205
rect -5414 -17243 -5397 -17154
rect -5307 -17243 1624 -17154
rect 1680 -17178 6618 -17130
rect -5407 -17252 -5288 -17243
rect -8560 -17286 -8464 -17274
rect -5242 -17372 -5236 -17320
rect -5184 -17372 -5178 -17320
rect -5234 -17548 -5186 -17372
rect 1680 -17548 1728 -17178
rect 1799 -17224 5799 -17221
rect -5234 -17596 1728 -17548
rect 1794 -17287 5799 -17224
rect -8570 -17615 -8474 -17598
rect -8570 -17684 -8554 -17615
rect -8485 -17684 -8474 -17615
rect 1794 -17648 1878 -17287
rect 1941 -17408 5831 -17342
rect -8570 -17696 -8474 -17684
rect -926 -17732 1878 -17648
rect -4988 -17780 -4894 -17758
rect -4988 -17841 -4979 -17780
rect -4918 -17841 -4894 -17780
rect -4988 -17850 -4894 -17841
rect -2280 -17780 -2186 -17760
rect -2280 -17841 -2269 -17780
rect -2208 -17841 -2186 -17780
rect -2280 -17852 -2186 -17841
rect -926 -17980 -842 -17732
rect 1942 -17812 2026 -17408
rect 810 -17896 816 -17812
rect 900 -17896 2026 -17812
rect 5407 -17552 5473 -17546
rect -2614 -18064 -2608 -17980
rect -2524 -18064 -842 -17980
rect -8568 -18097 -8472 -18080
rect -8568 -18166 -8554 -18097
rect -8485 -18166 -8472 -18097
rect -8568 -18178 -8472 -18166
rect -18060 -18385 -18000 -18381
rect -18071 -18455 -18065 -18385
rect -17995 -18455 -17989 -18385
rect -12661 -18396 -12599 -18392
rect -18060 -18459 -18000 -18455
rect -12672 -18468 -12666 -18396
rect -12594 -18468 -12588 -18396
rect -12661 -18472 -12599 -18468
rect -18094 -18515 -18015 -18511
rect -18105 -18604 -18099 -18515
rect -18010 -18604 -18004 -18515
rect -8564 -18567 -8468 -18548
rect -12628 -18573 -12549 -18569
rect -18094 -18608 -18015 -18604
rect -12639 -18662 -12633 -18573
rect -12544 -18662 -12538 -18573
rect -8564 -18636 -8554 -18567
rect -8485 -18636 -8468 -18567
rect -8564 -18646 -8468 -18636
rect -5014 -18582 -4920 -18572
rect -5014 -18654 -5006 -18582
rect -4934 -18654 -4920 -18582
rect -12628 -18666 -12549 -18662
rect -5014 -18664 -4920 -18654
rect -2302 -18582 -2208 -18572
rect -2302 -18654 -2294 -18582
rect -2222 -18654 -2208 -18582
rect -2302 -18664 -2208 -18654
rect -19377 -18705 -19311 -18699
rect -19311 -18771 -14471 -18705
rect -19377 -18777 -19311 -18771
rect -20352 -19464 -19800 -19416
rect -20404 -19472 -20352 -19466
rect -18024 -19622 -17942 -19614
rect -18024 -19685 -18016 -19622
rect -17953 -19685 -17942 -19622
rect -14537 -19617 -14471 -18771
rect -8584 -19098 -8512 -19092
rect -8584 -19176 -8512 -19170
rect -5026 -19430 -4932 -19420
rect -5026 -19502 -5014 -19430
rect -4942 -19502 -4932 -19430
rect -5026 -19512 -4932 -19502
rect -2308 -19430 -2214 -19420
rect -2308 -19502 -2300 -19430
rect -2228 -19502 -2214 -19430
rect -2308 -19512 -2214 -19502
rect -14537 -19683 -413 -19617
rect -347 -19683 -341 -19617
rect -18024 -19692 -17942 -19685
rect -20317 -19762 -10635 -19753
rect -20322 -19819 -10635 -19762
rect -20322 -19894 -20274 -19819
rect -14808 -19866 -14756 -19860
rect -20330 -19946 -20324 -19894
rect -20272 -19946 -20266 -19894
rect -17994 -19907 -17906 -19898
rect -17994 -19978 -17986 -19907
rect -17915 -19978 -17906 -19907
rect -14756 -19916 -10766 -19868
rect -14808 -19924 -14756 -19918
rect -17994 -19986 -17906 -19978
rect -10814 -20290 -10766 -19916
rect -10701 -20195 -10635 -19819
rect -5174 -20056 -5074 -20044
rect -5174 -20128 -5166 -20056
rect -5094 -20128 -5074 -20056
rect -2420 -20056 -2348 -20050
rect -2424 -20123 -2420 -20061
rect -2348 -20123 -2344 -20061
rect 5407 -20121 5473 -17619
rect 5554 -18615 5563 -18556
rect 5622 -18615 5631 -18556
rect 5994 -18633 6003 -18574
rect 6062 -18633 6071 -18574
rect 6431 -18626 6440 -18567
rect 6499 -18626 6508 -18567
rect -5174 -20134 -5074 -20128
rect -2420 -20134 -2348 -20128
rect 5407 -20187 5798 -20121
rect -10701 -20261 -337 -20195
rect -24956 -20291 -24844 -20290
rect -24956 -20363 -24936 -20291
rect -24864 -20363 -24844 -20291
rect -10814 -20338 -446 -20290
rect -24956 -20364 -24844 -20363
rect -20399 -20354 -20347 -20348
rect -20347 -20360 -18426 -20356
rect -20347 -20404 -18421 -20360
rect -20399 -20412 -20347 -20406
rect -24940 -20444 -24792 -20436
rect -24940 -20533 -24902 -20444
rect -24811 -20533 -24792 -20444
rect -24940 -20534 -24792 -20533
rect -18572 -20814 -18520 -20808
rect -18572 -20872 -18520 -20866
rect -18698 -21346 -18692 -21294
rect -18640 -21346 -18634 -21294
rect -24936 -21497 -24812 -21464
rect -24936 -21569 -24924 -21497
rect -24852 -21569 -24812 -21497
rect -24936 -21574 -24812 -21569
rect -24936 -21650 -24812 -21638
rect -24936 -21739 -24913 -21650
rect -24823 -21739 -24812 -21650
rect -24936 -21748 -24812 -21739
rect -18690 -21784 -18642 -21346
rect -18570 -21672 -18522 -20872
rect -18466 -21596 -18421 -20404
rect -5586 -20422 -5534 -20416
rect -5586 -20480 -5534 -20474
rect -494 -20430 -446 -20338
rect -403 -20323 -337 -20261
rect 1361 -20283 1367 -20217
rect 1433 -20283 5803 -20217
rect -403 -20389 5798 -20323
rect -494 -20478 5912 -20430
rect -18051 -21176 -17995 -21170
rect -18059 -21237 -18053 -21176
rect -17992 -21237 -17986 -21176
rect -18051 -21244 -17995 -21237
rect -17974 -21340 -17886 -21322
rect -17974 -21404 -17968 -21340
rect -17904 -21404 -17886 -21340
rect -17974 -21410 -17886 -21404
rect -12618 -21367 -12524 -21354
rect -12618 -21437 -12609 -21367
rect -12539 -21437 -12524 -21367
rect -12618 -21448 -12524 -21437
rect -12640 -21527 -12518 -21518
rect -18466 -21641 -16235 -21596
rect -12640 -21616 -12628 -21527
rect -12539 -21616 -12518 -21527
rect -12640 -21624 -12518 -21616
rect -18570 -21720 -16310 -21672
rect -18690 -21832 -16420 -21784
rect -16468 -22230 -16420 -21832
rect -16358 -22116 -16310 -21720
rect -16280 -22020 -16235 -21641
rect -5584 -21664 -5536 -20480
rect 3886 -21046 3970 -21040
rect -3912 -21130 -3906 -21046
rect -3822 -21130 3886 -21046
rect 3886 -21136 3970 -21130
rect 1221 -21389 1287 -21383
rect 1287 -21455 4745 -21389
rect 4811 -21455 4817 -21389
rect 1221 -21461 1287 -21455
rect -5136 -21608 -5130 -21525
rect -5047 -21608 6237 -21525
rect -5584 -21712 6004 -21664
rect -2757 -21819 -2751 -21748
rect -2680 -21819 6679 -21748
rect 668 -21956 674 -21872
rect 758 -21956 5966 -21872
rect -16280 -22065 5277 -22020
rect -16358 -22164 -12790 -22116
rect -12756 -22150 -12750 -22098
rect -12698 -22100 -12692 -22098
rect -12698 -22148 5166 -22100
rect -12698 -22150 -12692 -22148
rect -12838 -22182 -12790 -22164
rect -12838 -22230 -10534 -22182
rect -16468 -22278 -12972 -22230
rect -13020 -22400 -12972 -22278
rect -12872 -22284 -12820 -22278
rect -12820 -22334 -10620 -22286
rect -12872 -22342 -12820 -22336
rect -13020 -22448 -10720 -22400
rect -18074 -22600 -17972 -22582
rect -18074 -22666 -18061 -22600
rect -17995 -22666 -17972 -22600
rect -18074 -22678 -17972 -22666
rect -18080 -22745 -17952 -22724
rect -24900 -22798 -24806 -22786
rect -24900 -22870 -24890 -22798
rect -24818 -22870 -24806 -22798
rect -18080 -22834 -18071 -22745
rect -17982 -22834 -17952 -22745
rect -18080 -22846 -17952 -22834
rect -24900 -22882 -24806 -22870
rect -24926 -22951 -24808 -22942
rect -24926 -23040 -24913 -22951
rect -24819 -23040 -24808 -22951
rect -24926 -23052 -24808 -23040
rect -12688 -23951 -12602 -23946
rect -12688 -23952 -12676 -23951
rect -18050 -23986 -17962 -23978
rect -18050 -24058 -18042 -23986
rect -17970 -24058 -17962 -23986
rect -12736 -24014 -12676 -23952
rect -12613 -23952 -12602 -23951
rect -12613 -24014 -12578 -23952
rect -12736 -24016 -12578 -24014
rect -18050 -24066 -17962 -24058
rect -12738 -24092 -12574 -24076
rect -24938 -24108 -24848 -24102
rect -24938 -24180 -24926 -24108
rect -24854 -24180 -24848 -24108
rect -24938 -24186 -24848 -24180
rect -18084 -24131 -17958 -24102
rect -18084 -24220 -18063 -24131
rect -17974 -24220 -17958 -24131
rect -12738 -24163 -12685 -24092
rect -12614 -24163 -12574 -24092
rect -12738 -24164 -12574 -24163
rect -18084 -24246 -17958 -24220
rect -24920 -24261 -24800 -24250
rect -24920 -24350 -24907 -24261
rect -24813 -24350 -24800 -24261
rect -24920 -24362 -24800 -24350
rect -13022 -25164 -13016 -25112
rect -12964 -25114 -12958 -25112
rect -12964 -25162 -10844 -25114
rect -12964 -25164 -12958 -25162
rect -17964 -25350 -17878 -25344
rect -17964 -25422 -17956 -25350
rect -17884 -25422 -17878 -25350
rect -17964 -25428 -17878 -25422
rect -17982 -25553 -17878 -25480
rect -17982 -25642 -17976 -25553
rect -17887 -25642 -17878 -25553
rect -17982 -25650 -17878 -25642
rect -10892 -25824 -10844 -25162
rect -10768 -25724 -10720 -22448
rect -10668 -25368 -10620 -22334
rect -10582 -25242 -10534 -22230
rect -10479 -22299 5069 -22213
rect -10479 -25098 -10393 -22299
rect -5708 -22456 -5702 -22404
rect -5650 -22406 -5644 -22404
rect -5650 -22454 4942 -22406
rect -5650 -22456 -5644 -22454
rect -2920 -22610 -2914 -22526
rect -2830 -22529 4836 -22526
rect -2830 -22610 4849 -22529
rect 490 -22696 574 -22690
rect 574 -22705 4656 -22696
rect 574 -22780 4717 -22705
rect 490 -22786 574 -22780
rect -5854 -24358 -5802 -24352
rect -6038 -24414 -6032 -24362
rect -5980 -24414 -5974 -24362
rect -6030 -24978 -5982 -24414
rect -5854 -24416 -5802 -24410
rect -6032 -24984 -5980 -24978
rect -5852 -25028 -5804 -24416
rect -6032 -25042 -5980 -25036
rect -5854 -25034 -5802 -25028
rect -5854 -25092 -5802 -25086
rect -10490 -25107 -10366 -25098
rect -10490 -25193 -10479 -25107
rect -10393 -25193 -10366 -25107
rect -10490 -25206 -10366 -25193
rect -10582 -25290 4462 -25242
rect -10668 -25416 4354 -25368
rect -10158 -25634 -10152 -25530
rect -10048 -25634 4226 -25530
rect -10768 -25772 -5970 -25724
rect -10892 -25872 -6064 -25824
rect -6112 -26420 -6064 -25872
rect -6018 -26332 -5970 -25772
rect -5854 -25742 -5802 -25736
rect -5802 -25792 4004 -25744
rect -5854 -25800 -5802 -25794
rect -3088 -25958 -3082 -25874
rect -2998 -25958 3902 -25874
rect 314 -26148 320 -26064
rect 404 -26148 3740 -26064
rect -6018 -26380 3558 -26332
rect -6112 -26468 3472 -26420
rect -12770 -26744 -12612 -26742
rect -12770 -26805 -12743 -26744
rect -12682 -26805 -12612 -26744
rect -12770 -26806 -12612 -26805
rect -12794 -26998 -12748 -26934
rect -12684 -26998 -12636 -26934
rect -12758 -29446 -12724 -29374
rect -12652 -29446 -12598 -29374
rect -12772 -29537 -12586 -29520
rect -12772 -29626 -12727 -29537
rect -12638 -29626 -12586 -29537
rect -12834 -31918 -12670 -31900
rect -12834 -31990 -12758 -31918
rect -12686 -31990 -12670 -31918
rect -12838 -32087 -12674 -32086
rect -12838 -32176 -12791 -32087
rect -12702 -32176 -12674 -32087
rect -9857 -32916 -9764 -32910
rect -9764 -33009 3112 -32916
rect -9857 -33015 -9764 -33009
rect -6038 -33168 -6032 -33116
rect -5980 -33118 -5974 -33116
rect -5980 -33166 2846 -33118
rect -5980 -33168 -5974 -33166
rect -3266 -33356 -3260 -33272
rect -3176 -33356 2696 -33272
rect -704 -33578 -698 -33494
rect -614 -33578 2428 -33494
rect -12582 -34504 -12510 -34498
rect -12582 -34582 -12510 -34576
rect -12746 -34671 -12582 -34670
rect -12746 -34760 -12726 -34671
rect -12637 -34760 -12582 -34671
rect 2344 -35454 2428 -33578
rect 2612 -35333 2696 -33356
rect 2798 -35235 2846 -33166
rect 3025 -35113 3091 -33009
rect 3424 -34011 3472 -26468
rect 3510 -33907 3558 -26380
rect 3656 -30926 3740 -26148
rect 3818 -30805 3902 -25958
rect 3956 -30722 4004 -25792
rect 4122 -30562 4226 -25634
rect 4306 -29500 4354 -25416
rect 4414 -29390 4462 -25290
rect 4651 -26398 4717 -22780
rect 4783 -26277 4849 -22610
rect 4894 -26179 4942 -22454
rect 4983 -26057 5069 -22299
rect 5118 -24962 5166 -22148
rect 5232 -24861 5277 -22065
rect 5554 -23159 5563 -23100
rect 5622 -23159 5631 -23100
rect 5994 -23149 6003 -23090
rect 6062 -23149 6071 -23090
rect 6439 -23124 6448 -23065
rect 6507 -23124 6516 -23065
rect 5726 -24715 5732 -24649
rect 5798 -24715 5804 -24649
rect 5311 -24811 5317 -24745
rect 5383 -24811 5809 -24745
rect 5232 -24906 5788 -24861
rect 5118 -25010 5808 -24962
rect 4983 -26123 5811 -26057
rect 4894 -26228 5827 -26179
rect 4899 -26245 5827 -26228
rect 4783 -26343 5799 -26277
rect 4651 -26464 5807 -26398
rect 5554 -27699 5563 -27640
rect 5622 -27699 5631 -27640
rect 5994 -27694 6003 -27635
rect 6062 -27694 6071 -27635
rect 6429 -27640 6438 -27581
rect 6497 -27640 6506 -27581
rect 5448 -29243 5454 -29177
rect 5520 -29243 5798 -29177
rect 4860 -29273 4919 -29272
rect 4860 -29278 5798 -29273
rect 4919 -29337 5798 -29278
rect 4860 -29339 5798 -29337
rect 4860 -29343 4919 -29339
rect 4414 -29438 5858 -29390
rect 4306 -29548 5804 -29500
rect 4122 -30666 5856 -30562
rect 3956 -30770 6030 -30722
rect 3818 -30871 5803 -30805
rect 3818 -30874 3902 -30871
rect 3656 -30992 5809 -30926
rect 3656 -30994 3740 -30992
rect 5554 -32208 5563 -32149
rect 5622 -32208 5631 -32149
rect 5994 -32223 6003 -32164
rect 6062 -32223 6071 -32164
rect 5419 -33771 5425 -33705
rect 5491 -33771 5804 -33705
rect 3657 -33867 3663 -33801
rect 3729 -33867 5811 -33801
rect 3510 -33958 5799 -33907
rect 3511 -33973 5799 -33958
rect 3424 -34077 5821 -34011
rect 3424 -34082 3756 -34077
rect 3025 -35179 5807 -35113
rect 2789 -35301 5817 -35235
rect 2612 -35399 5801 -35333
rect 2612 -35400 2696 -35399
rect 2328 -35520 5805 -35454
<< via2 >>
rect -22627 7013 -22565 7075
rect -27520 4457 -27441 4536
rect -21811 6730 -21732 6809
rect -19307 6588 -19245 6650
rect -18524 6417 -18445 6496
rect -16014 6242 -15952 6304
rect -15226 6071 -15147 6150
rect -12737 5911 -12675 5973
rect -11936 5705 -11857 5784
rect -9434 5546 -9372 5608
rect -8636 5402 -8557 5481
rect -6161 5274 -6101 5334
rect -5353 5123 -5268 5202
rect -2870 4961 -2808 5023
rect -2054 4797 -1975 4876
rect 430 4684 492 4721
rect 430 4659 492 4684
rect 5558 4029 5627 4099
rect 5998 4029 6067 4099
rect 6445 4022 6504 4081
rect 5563 -509 5622 -450
rect 6003 -483 6062 -424
rect 6443 -514 6502 -455
rect -25216 -2591 -25155 -2529
rect -25504 -5097 -25442 -5035
rect -25655 -6832 -25576 -6751
rect -25809 -8362 -25749 -8302
rect -25978 -10241 -25899 -10160
rect -25365 -11055 -25286 -10976
rect -26164 -11653 -26102 -11591
rect -26327 -13144 -26248 -13063
rect -24916 -15658 -24844 -15586
rect -24903 -15828 -24812 -15739
rect -24908 -16842 -24836 -16770
rect -24915 -17012 -24836 -16923
rect -24921 -18054 -24851 -17984
rect -24917 -18217 -24824 -18128
rect 5563 -4919 5622 -4860
rect 6003 -4939 6062 -4880
rect 6442 -4948 6501 -4889
rect 5563 -9582 5622 -9523
rect 6003 -9587 6062 -9528
rect 6445 -9573 6504 -9514
rect -17961 -15653 -17899 -15591
rect -12719 -15653 -12657 -15591
rect -18118 -15822 -18039 -15743
rect -12555 -15837 -12456 -15738
rect -5003 -14561 -4941 -14499
rect -2283 -14561 -2221 -14499
rect -8671 -15563 -8609 -15501
rect -4961 -15373 -4899 -15311
rect -2259 -15373 -2197 -15311
rect -24870 -19175 -24798 -19103
rect -24875 -19345 -24796 -19256
rect 5563 -14109 5622 -14050
rect 6003 -14093 6062 -14034
rect 6442 -14076 6501 -14017
rect -8549 -16219 -8487 -16157
rect -4990 -16190 -4930 -16130
rect -2280 -16190 -2220 -16130
rect -8551 -16754 -8482 -16685
rect -18077 -17047 -18015 -16985
rect -4997 -17018 -4941 -16962
rect -2288 -17018 -2232 -16962
rect -18085 -17197 -18005 -17118
rect -8549 -17274 -8480 -17205
rect -8554 -17684 -8485 -17615
rect -4977 -17839 -4921 -17783
rect -2267 -17839 -2211 -17783
rect -8554 -18166 -8485 -18097
rect -18060 -18450 -18000 -18390
rect -12661 -18463 -12599 -18401
rect -18094 -18599 -18015 -18520
rect -12628 -18657 -12549 -18578
rect -8554 -18636 -8485 -18567
rect -5001 -18649 -4939 -18587
rect -2289 -18649 -2227 -18587
rect -18013 -19682 -17957 -19626
rect -8579 -19165 -8517 -19103
rect -5009 -19497 -4947 -19435
rect -2295 -19497 -2233 -19435
rect -17981 -19973 -17920 -19912
rect -5161 -20123 -5099 -20061
rect -2415 -20123 -2353 -20061
rect 5563 -18615 5622 -18556
rect 6003 -18633 6062 -18574
rect 6440 -18626 6499 -18567
rect -24936 -20363 -24864 -20291
rect -24902 -20533 -24811 -20444
rect -24914 -21569 -24852 -21497
rect -24913 -21739 -24823 -21650
rect -18051 -21235 -17995 -21179
rect -17964 -21400 -17908 -21344
rect -12604 -21432 -12544 -21372
rect -12623 -21611 -12544 -21532
rect -18061 -22666 -17995 -22600
rect -24890 -22870 -24818 -22798
rect -18067 -22829 -17987 -22750
rect -24913 -23040 -24819 -22951
rect -18037 -24053 -17975 -23991
rect -12673 -24011 -12617 -23955
rect -24926 -24180 -24864 -24108
rect -18058 -24215 -17979 -24136
rect -12681 -24158 -12619 -24097
rect -24907 -24350 -24813 -24261
rect -17951 -25417 -17889 -25355
rect -17971 -25637 -17892 -25558
rect -12741 -26803 -12685 -26747
rect -12744 -26994 -12688 -26938
rect -12719 -29441 -12657 -29379
rect -12723 -29621 -12643 -29542
rect -12753 -31985 -12691 -31923
rect -12787 -32171 -12707 -32092
rect -12577 -34571 -12515 -34509
rect -12721 -34755 -12642 -34676
rect 5563 -23159 5622 -23100
rect 6003 -23149 6062 -23090
rect 6448 -23124 6507 -23065
rect 5563 -27699 5622 -27640
rect 6003 -27694 6062 -27635
rect 6438 -27640 6497 -27581
rect 5563 -32208 5622 -32149
rect 6003 -32223 6062 -32164
rect 6438 -32201 6507 -32131
<< metal3 >>
rect -27376 7075 -22560 7080
rect -27376 7013 -22627 7075
rect -22565 7013 -22560 7075
rect -27376 7008 -22560 7013
rect -27525 4536 -27436 4541
rect -27525 4457 -27520 4536
rect -27441 4457 -27436 4536
rect -27525 -24260 -27436 4457
rect -27376 -24108 -27304 7008
rect -27210 6809 -21727 6814
rect -27210 6730 -21811 6809
rect -21732 6730 -21727 6809
rect -27210 6725 -21727 6730
rect -27210 6717 -27121 6725
rect -27210 -22950 -27131 6717
rect -27070 6650 -19240 6655
rect -27070 6588 -19307 6650
rect -19245 6588 -19240 6650
rect -27070 6583 -19240 6588
rect -27070 -22798 -26998 6583
rect -26921 6496 -18440 6501
rect -26921 6417 -18524 6496
rect -18445 6417 -18440 6496
rect -26921 6412 -18440 6417
rect -26921 6411 -26832 6412
rect -26921 -21642 -26842 6411
rect -26782 6304 -15947 6309
rect -26782 6242 -16014 6304
rect -15952 6242 -15947 6304
rect -26782 6237 -15947 6242
rect -26782 -21497 -26710 6237
rect -26650 6150 -15142 6155
rect -26650 6071 -15226 6150
rect -15147 6071 -15142 6150
rect -26650 6066 -15142 6071
rect -26650 -20443 -26564 6066
rect -26500 5973 -12670 5978
rect -26500 5911 -12737 5973
rect -12675 5911 -12670 5973
rect -26500 5906 -12670 5911
rect -26500 -20291 -26428 5906
rect -26332 5784 -11852 5789
rect -26332 5705 -11936 5784
rect -11857 5705 -11852 5784
rect -26332 5700 -11852 5705
rect -26332 -13063 -26243 5700
rect -26332 -13144 -26327 -13063
rect -26248 -13144 -26243 -13063
rect -26332 -19255 -26243 -13144
rect -26169 5608 -9367 5613
rect -26169 5546 -9434 5608
rect -9372 5546 -9367 5608
rect -26169 5541 -9367 5546
rect -26169 -11591 -26097 5541
rect -9298 5481 -8552 5486
rect -9298 5479 -8636 5481
rect -26169 -11653 -26164 -11591
rect -26102 -11653 -26097 -11591
rect -26169 -19103 -26097 -11653
rect -25983 5402 -8636 5479
rect -8557 5402 -8552 5481
rect -25983 5397 -8552 5402
rect -25983 -10160 -25894 5397
rect -8489 5336 -6096 5339
rect -25983 -10241 -25978 -10160
rect -25899 -10241 -25894 -10160
rect -25983 -18127 -25894 -10241
rect -25814 5334 -6096 5336
rect -25814 5274 -6161 5334
rect -6101 5274 -6096 5334
rect -25814 5269 -6096 5274
rect -25814 -8302 -25744 5269
rect -25814 -8362 -25809 -8302
rect -25749 -8362 -25744 -8302
rect -25814 -17984 -25744 -8362
rect -25660 5202 -5263 5207
rect -25660 5123 -5353 5202
rect -5268 5123 -5263 5202
rect -25660 5118 -5263 5123
rect -25660 -6751 -25571 5118
rect -25660 -6832 -25655 -6751
rect -25576 -6832 -25571 -6751
rect -25660 -16922 -25571 -6832
rect -25509 5023 -2803 5028
rect -25509 4961 -2870 5023
rect -2808 4961 -2803 5023
rect -25509 4956 -2803 4961
rect -25509 -5035 -25437 4956
rect -25509 -5097 -25504 -5035
rect -25442 -5097 -25437 -5035
rect -25509 -16770 -25437 -5097
rect -25370 4876 -1970 4881
rect -25370 4797 -2054 4876
rect -1975 4797 -1970 4876
rect -25370 4792 -1970 4797
rect -25370 -10976 -25281 4792
rect -25370 -11055 -25365 -10976
rect -25286 -11055 -25281 -10976
rect -25370 -15738 -25281 -11055
rect -25221 4721 497 4726
rect -25221 4659 430 4721
rect 492 4659 497 4721
rect -25221 4654 497 4659
rect -25221 -2529 -25150 4654
rect 5553 4099 5632 4104
rect 5553 4029 5558 4099
rect 5627 4029 5632 4099
rect 5553 4024 5632 4029
rect 5993 4099 6072 4104
rect 5993 4029 5998 4099
rect 6067 4029 6072 4099
rect 5993 4024 6072 4029
rect 6440 4081 6509 4086
rect -25221 -2591 -25216 -2529
rect -25155 -2591 -25150 -2529
rect -25221 -15586 -25150 -2591
rect 5558 -450 5627 4024
rect 5558 -509 5563 -450
rect 5622 -509 5627 -450
rect 5558 -4860 5627 -509
rect 5558 -4919 5563 -4860
rect 5622 -4919 5627 -4860
rect 5558 -9523 5627 -4919
rect 5558 -9582 5563 -9523
rect 5622 -9582 5627 -9523
rect 5558 -14050 5627 -9582
rect 5558 -14109 5563 -14050
rect 5622 -14109 5627 -14050
rect -6212 -14496 -2216 -14494
rect -6780 -14499 -2216 -14496
rect -6780 -14561 -5003 -14499
rect -4941 -14561 -2283 -14499
rect -2221 -14561 -2216 -14499
rect -6780 -14566 -2216 -14561
rect -6780 -14568 -6124 -14566
rect -8676 -15501 -8604 -15496
rect -8676 -15563 -8671 -15501
rect -8609 -15563 -8604 -15501
rect -24921 -15586 -24839 -15581
rect -12730 -15586 -12656 -15570
rect -25221 -15658 -24916 -15586
rect -24844 -15591 -9810 -15586
rect -24844 -15653 -17961 -15591
rect -17899 -15653 -12719 -15591
rect -12657 -15632 -9810 -15591
rect -8676 -15632 -8604 -15563
rect -6780 -15632 -6708 -14568
rect -6596 -15311 -2184 -15306
rect -6596 -15373 -4961 -15311
rect -4899 -15373 -2259 -15311
rect -2197 -15373 -2184 -15311
rect -6596 -15378 -2184 -15373
rect -12657 -15653 -6688 -15632
rect -24844 -15658 -6688 -15653
rect -24921 -15663 -24839 -15658
rect -12730 -15666 -12656 -15658
rect -9882 -15704 -6688 -15658
rect -9882 -15708 -9810 -15704
rect -24908 -15738 -24807 -15734
rect -12560 -15738 -12451 -15733
rect -25370 -15739 -12555 -15738
rect -25370 -15827 -24903 -15739
rect -24908 -15828 -24903 -15827
rect -24812 -15743 -12555 -15739
rect -24812 -15822 -18118 -15743
rect -18039 -15822 -12555 -15743
rect -24812 -15827 -12555 -15822
rect -24812 -15828 -24807 -15827
rect -24908 -15833 -24807 -15828
rect -12560 -15837 -12555 -15827
rect -12456 -15827 -10774 -15738
rect -12456 -15837 -12451 -15827
rect -12560 -15842 -12451 -15837
rect -6596 -16152 -6524 -15378
rect -6209 -16130 -2203 -16125
rect -10052 -16157 -6510 -16152
rect -10052 -16219 -8549 -16157
rect -8487 -16219 -6510 -16157
rect -10052 -16224 -6510 -16219
rect -6209 -16190 -4990 -16130
rect -4930 -16190 -2280 -16130
rect -2220 -16190 -2203 -16130
rect -6209 -16195 -2203 -16190
rect -24913 -16770 -24831 -16765
rect -25509 -16842 -24908 -16770
rect -24836 -16842 -18526 -16770
rect -24913 -16847 -24831 -16842
rect -24920 -16922 -24831 -16918
rect -25660 -16923 -18736 -16922
rect -25660 -17011 -24915 -16923
rect -24920 -17012 -24915 -17011
rect -24836 -17011 -18736 -16923
rect -24836 -17012 -24831 -17011
rect -24920 -17017 -24831 -17012
rect -18825 -17113 -18736 -17011
rect -18598 -16980 -18526 -16842
rect -18598 -16985 -13076 -16980
rect -18598 -17047 -18077 -16985
rect -18015 -17047 -13076 -16985
rect -18598 -17052 -13076 -17047
rect -18825 -17118 -17178 -17113
rect -18825 -17197 -18085 -17118
rect -18005 -17155 -17178 -17118
rect -18005 -17197 -13292 -17155
rect -18825 -17202 -13292 -17197
rect -17304 -17244 -13292 -17202
rect -22395 -17977 -18413 -17907
rect -24926 -17984 -24846 -17979
rect -22395 -17984 -22325 -17977
rect -25814 -18054 -24921 -17984
rect -24851 -18054 -22325 -17984
rect -24926 -18059 -24846 -18054
rect -24922 -18127 -24819 -18123
rect -25983 -18128 -22118 -18127
rect -25983 -18216 -24917 -18128
rect -24922 -18217 -24917 -18216
rect -24824 -18216 -22118 -18128
rect -24824 -18217 -24819 -18216
rect -24922 -18222 -24819 -18217
rect -22207 -18315 -22118 -18216
rect -22207 -18404 -18592 -18315
rect -18681 -18515 -18592 -18404
rect -18483 -18385 -18413 -17977
rect -16571 -18301 -13459 -18231
rect -16571 -18385 -16501 -18301
rect -18483 -18390 -16501 -18385
rect -18483 -18450 -18060 -18390
rect -18000 -18450 -16501 -18390
rect -18483 -18455 -16501 -18450
rect -18681 -18520 -16570 -18515
rect -18681 -18599 -18094 -18520
rect -18015 -18599 -16570 -18520
rect -18681 -18604 -16570 -18599
rect -16659 -18695 -16570 -18604
rect -16659 -18784 -13618 -18695
rect -13707 -18903 -13618 -18784
rect -13529 -18769 -13459 -18301
rect -13381 -18573 -13292 -17244
rect -13148 -18396 -13076 -17052
rect -10052 -18396 -9980 -16224
rect -8556 -16685 -8477 -16680
rect -8556 -16687 -8551 -16685
rect -13148 -18401 -9980 -18396
rect -13148 -18463 -12661 -18401
rect -12599 -18463 -9980 -18401
rect -13148 -18468 -9980 -18463
rect -9825 -16754 -8551 -16687
rect -8482 -16687 -8477 -16685
rect -6209 -16687 -6139 -16195
rect -8482 -16754 -6139 -16687
rect -9825 -16757 -6139 -16754
rect -13381 -18578 -12544 -18573
rect -13381 -18657 -12628 -18578
rect -12549 -18657 -12544 -18578
rect -13381 -18662 -12544 -18657
rect -13529 -18839 -12679 -18769
rect -22106 -18980 -18438 -18908
rect -24875 -19103 -24793 -19098
rect -22106 -19103 -22034 -18980
rect -26169 -19175 -24870 -19103
rect -24798 -19175 -22034 -19103
rect -24875 -19180 -24793 -19175
rect -24880 -19255 -24791 -19251
rect -26332 -19256 -22060 -19255
rect -26332 -19344 -24875 -19256
rect -24880 -19345 -24875 -19344
rect -24796 -19344 -22060 -19256
rect -24796 -19345 -24791 -19344
rect -24880 -19350 -24791 -19345
rect -22149 -19385 -22060 -19344
rect -22149 -19474 -18636 -19385
rect -18725 -19907 -18636 -19474
rect -18506 -19780 -18442 -18980
rect -13707 -18992 -12844 -18903
rect -18018 -19626 -17952 -19621
rect -18018 -19682 -18013 -19626
rect -17957 -19682 -17952 -19626
rect -18018 -19687 -17952 -19682
rect -18017 -19780 -17954 -19687
rect -18506 -19843 -13041 -19780
rect -18506 -19844 -18442 -19843
rect -18725 -19912 -16507 -19907
rect -18725 -19973 -17981 -19912
rect -17920 -19973 -16507 -19912
rect -18725 -19978 -16507 -19973
rect -16578 -20132 -16507 -19978
rect -16578 -20203 -13191 -20132
rect -24941 -20291 -24859 -20286
rect -26500 -20363 -24936 -20291
rect -24864 -20363 -18314 -20291
rect -24941 -20368 -24859 -20363
rect -24907 -20443 -24806 -20439
rect -26650 -20444 -22144 -20443
rect -26650 -20532 -24902 -20444
rect -24907 -20533 -24902 -20532
rect -24811 -20532 -22144 -20444
rect -24811 -20533 -24806 -20532
rect -24907 -20538 -24806 -20533
rect -22233 -20717 -22144 -20532
rect -22233 -20806 -18498 -20717
rect -18587 -21340 -18498 -20806
rect -18380 -21177 -18319 -20363
rect -18056 -21177 -17990 -21174
rect -16037 -21177 -13362 -21120
rect -18380 -21179 -13362 -21177
rect -18380 -21235 -18051 -21179
rect -17995 -21181 -13362 -21179
rect -17995 -21235 -15976 -21181
rect -18380 -21238 -15976 -21235
rect -18056 -21240 -17990 -21238
rect -17969 -21340 -17903 -21339
rect -18587 -21344 -16574 -21340
rect -18587 -21350 -17964 -21344
rect -18574 -21400 -17964 -21350
rect -17908 -21400 -16574 -21344
rect -18574 -21404 -16574 -21400
rect -17969 -21405 -17903 -21404
rect -24919 -21497 -24847 -21492
rect -26782 -21569 -24914 -21497
rect -24852 -21569 -22110 -21497
rect -24919 -21574 -24847 -21569
rect -26921 -21649 -26832 -21642
rect -24918 -21649 -24818 -21645
rect -26921 -21650 -22298 -21649
rect -26921 -21738 -24913 -21650
rect -24918 -21739 -24913 -21738
rect -24823 -21738 -22298 -21650
rect -24823 -21739 -24818 -21738
rect -24918 -21744 -24818 -21739
rect -22387 -22745 -22298 -21738
rect -22182 -22586 -22110 -21569
rect -16638 -21578 -16574 -21404
rect -16638 -21642 -13506 -21578
rect -22182 -22600 -13654 -22586
rect -22182 -22658 -18061 -22600
rect -18066 -22666 -18061 -22658
rect -17995 -22658 -13654 -22600
rect -17995 -22666 -17990 -22658
rect -18066 -22671 -17990 -22666
rect -22387 -22750 -13824 -22745
rect -24895 -22798 -24813 -22793
rect -27070 -22870 -24890 -22798
rect -24818 -22870 -22488 -22798
rect -22387 -22829 -18067 -22750
rect -17987 -22829 -13824 -22750
rect -22387 -22834 -13824 -22829
rect -24895 -22875 -24813 -22870
rect -24918 -22950 -24814 -22946
rect -27210 -22951 -22674 -22950
rect -27210 -23039 -24913 -22951
rect -24918 -23040 -24913 -23039
rect -24819 -23039 -22674 -22951
rect -24819 -23040 -24814 -23039
rect -24918 -23045 -24814 -23040
rect -24931 -24108 -24859 -24103
rect -27376 -24180 -24926 -24108
rect -24864 -24180 -22986 -24108
rect -24931 -24185 -24859 -24180
rect -24934 -24260 -24778 -24252
rect -27525 -24261 -23124 -24260
rect -27525 -24349 -24907 -24261
rect -24934 -24350 -24907 -24349
rect -24813 -24349 -23124 -24261
rect -24813 -24350 -24778 -24349
rect -24934 -24360 -24778 -24350
rect -23213 -25553 -23124 -24349
rect -23058 -25350 -22986 -24180
rect -22763 -24131 -22674 -23039
rect -22560 -23986 -22488 -22870
rect -22560 -23991 -14032 -23986
rect -22560 -24053 -18037 -23991
rect -17975 -24053 -14032 -23991
rect -22560 -24058 -14032 -24053
rect -22763 -24136 -14178 -24131
rect -22763 -24215 -18058 -24136
rect -17979 -24215 -14178 -24136
rect -22763 -24220 -14178 -24215
rect -23058 -25355 -14392 -25350
rect -23058 -25417 -17951 -25355
rect -17889 -25417 -14392 -25355
rect -23058 -25422 -14392 -25417
rect -23213 -25558 -14534 -25553
rect -23213 -25637 -17971 -25558
rect -17892 -25637 -14534 -25558
rect -23213 -25642 -14534 -25637
rect -14623 -34671 -14534 -25642
rect -14464 -34504 -14392 -25422
rect -14267 -32087 -14178 -24220
rect -14104 -31918 -14032 -24058
rect -13913 -29537 -13824 -22834
rect -13726 -29374 -13654 -22658
rect -13570 -26934 -13506 -21642
rect -13423 -26745 -13362 -21181
rect -13262 -24092 -13191 -20203
rect -13104 -23952 -13041 -19843
rect -12933 -21527 -12844 -18992
rect -12749 -21367 -12679 -18839
rect -12749 -21372 -9935 -21367
rect -12749 -21432 -12604 -21372
rect -12544 -21385 -9935 -21372
rect -9825 -21385 -9755 -16757
rect -8556 -16759 -8477 -16757
rect -5002 -16959 -4936 -16957
rect -2293 -16959 -2227 -16957
rect -5941 -16962 -2195 -16959
rect -5941 -17018 -4997 -16962
rect -4941 -17018 -2288 -16962
rect -2232 -17018 -2195 -16962
rect -5941 -17022 -2195 -17018
rect -8554 -17205 -8475 -17200
rect -8554 -17209 -8549 -17205
rect -12544 -21432 -9755 -21385
rect -12749 -21437 -9755 -21432
rect -10035 -21455 -9755 -21437
rect -9648 -17272 -8549 -17209
rect -12933 -21532 -12486 -21527
rect -12933 -21611 -12623 -21532
rect -12544 -21611 -12486 -21532
rect -12933 -21616 -12486 -21611
rect -12688 -23952 -12602 -23946
rect -9648 -23952 -9585 -17272
rect -8554 -17274 -8549 -17272
rect -8480 -17209 -8475 -17205
rect -5941 -17209 -5878 -17022
rect -5002 -17023 -4936 -17022
rect -2293 -17023 -2227 -17022
rect -8480 -17272 -5875 -17209
rect -8480 -17274 -8475 -17272
rect -8554 -17279 -8475 -17274
rect -8559 -17615 -8480 -17610
rect -8559 -17616 -8554 -17615
rect -13104 -23955 -9585 -23952
rect -13104 -24011 -12673 -23955
rect -12617 -24011 -9585 -23955
rect -13104 -24015 -9585 -24011
rect -9457 -17677 -8554 -17616
rect -12678 -24016 -12612 -24015
rect -12738 -24092 -12574 -24076
rect -13262 -24097 -12523 -24092
rect -13262 -24158 -12681 -24097
rect -12619 -24158 -12523 -24097
rect -13262 -24163 -12523 -24158
rect -12738 -24164 -12574 -24163
rect -12770 -26745 -12612 -26742
rect -9457 -26745 -9396 -17677
rect -8559 -17684 -8554 -17677
rect -8485 -17616 -8480 -17615
rect -8485 -17677 -5420 -17616
rect -8485 -17684 -8480 -17677
rect -8559 -17689 -8480 -17684
rect -5481 -17781 -5420 -17677
rect -4982 -17781 -4916 -17778
rect -2272 -17781 -2206 -17778
rect -5481 -17783 -2196 -17781
rect -5481 -17839 -4977 -17783
rect -4921 -17839 -2267 -17783
rect -2211 -17839 -2196 -17783
rect -5481 -17842 -2196 -17839
rect -4982 -17844 -4916 -17842
rect -2272 -17844 -2206 -17842
rect -8559 -18094 -8480 -18092
rect -13423 -26747 -9396 -26745
rect -13423 -26803 -12741 -26747
rect -12685 -26803 -9396 -26747
rect -13423 -26806 -9396 -26803
rect -9308 -18097 -5472 -18094
rect -9308 -18166 -8554 -18097
rect -8485 -18166 -5472 -18097
rect -12746 -26808 -12680 -26806
rect -12749 -26934 -12683 -26933
rect -13570 -26938 -12532 -26934
rect -13570 -26994 -12744 -26938
rect -12688 -26994 -12532 -26938
rect -13570 -26998 -12532 -26994
rect -12749 -26999 -12683 -26998
rect -9308 -29374 -9236 -18166
rect -8559 -18171 -8480 -18166
rect -13726 -29379 -9236 -29374
rect -13726 -29441 -12719 -29379
rect -12657 -29441 -9236 -29379
rect -13726 -29446 -9236 -29441
rect -9076 -18567 -5782 -18562
rect -9076 -18634 -8554 -18567
rect -13913 -29542 -12094 -29537
rect -13913 -29621 -12723 -29542
rect -12643 -29621 -12094 -29542
rect -13913 -29626 -12094 -29621
rect -12834 -31918 -12670 -31900
rect -9076 -31918 -9004 -18634
rect -8559 -18636 -8554 -18634
rect -8485 -18634 -5782 -18567
rect -8485 -18636 -8480 -18634
rect -8559 -18641 -8480 -18636
rect -14104 -31923 -9004 -31918
rect -14104 -31985 -12753 -31923
rect -12691 -31985 -9004 -31923
rect -14104 -31990 -9004 -31985
rect -8828 -19103 -5924 -19098
rect -8828 -19165 -8579 -19103
rect -8517 -19165 -5924 -19103
rect -8828 -19170 -5924 -19165
rect -14267 -32092 -12460 -32087
rect -14267 -32171 -12787 -32092
rect -12707 -32171 -12460 -32092
rect -14267 -32176 -12460 -32171
rect -8828 -34504 -8756 -19170
rect -5996 -20056 -5924 -19170
rect -5854 -19430 -5782 -18634
rect -5544 -18582 -5472 -18166
rect 5558 -18556 5627 -14109
rect -5544 -18587 -2222 -18582
rect -5544 -18649 -5001 -18587
rect -4939 -18649 -2289 -18587
rect -2227 -18649 -2222 -18587
rect -5544 -18654 -2222 -18649
rect 5558 -18615 5563 -18556
rect 5622 -18615 5627 -18556
rect -5854 -19435 -2216 -19430
rect -5854 -19497 -5009 -19435
rect -4947 -19497 -2295 -19435
rect -2233 -19497 -2216 -19435
rect -5854 -19502 -2216 -19497
rect -5996 -20061 -2348 -20056
rect -5996 -20123 -5161 -20061
rect -5099 -20123 -2415 -20061
rect -2353 -20123 -2348 -20061
rect -5996 -20128 -2348 -20123
rect 5558 -23100 5627 -18615
rect 5558 -23159 5563 -23100
rect 5622 -23159 5627 -23100
rect 5558 -27640 5627 -23159
rect 5558 -27699 5563 -27640
rect 5622 -27699 5627 -27640
rect 5558 -32149 5627 -27699
rect 5558 -32208 5563 -32149
rect 5622 -32208 5627 -32149
rect 5558 -32279 5627 -32208
rect 5998 -424 6067 4024
rect 6440 4022 6445 4081
rect 6504 4022 6509 4081
rect 6440 3020 6509 4022
rect 6144 2951 6509 3020
rect 6144 302 6213 2951
rect 6144 233 6507 302
rect 5998 -483 6003 -424
rect 6062 -483 6067 -424
rect 5998 -4880 6067 -483
rect 6438 -455 6507 233
rect 6438 -514 6443 -455
rect 6502 -514 6507 -455
rect 6438 -1465 6507 -514
rect 6168 -1534 6507 -1465
rect 6168 -4240 6237 -1534
rect 6168 -4309 6506 -4240
rect 5998 -4939 6003 -4880
rect 6062 -4939 6067 -4880
rect 5998 -9528 6067 -4939
rect 6437 -4889 6506 -4309
rect 6437 -4948 6442 -4889
rect 6501 -4948 6506 -4889
rect 6437 -5912 6506 -4948
rect 6165 -5981 6506 -5912
rect 6165 -9037 6234 -5981
rect 6165 -9106 6509 -9037
rect 5998 -9587 6003 -9528
rect 6062 -9587 6067 -9528
rect 5998 -14034 6067 -9587
rect 6440 -9514 6509 -9106
rect 6440 -9573 6445 -9514
rect 6504 -9573 6509 -9514
rect 6440 -10527 6509 -9573
rect 6166 -10596 6509 -10527
rect 6166 -13281 6235 -10596
rect 6166 -13350 6506 -13281
rect 5998 -14093 6003 -14034
rect 6062 -14093 6067 -14034
rect 5998 -18574 6067 -14093
rect 6437 -14017 6506 -13350
rect 6437 -14076 6442 -14017
rect 6501 -14076 6506 -14017
rect 6437 -15089 6506 -14076
rect 6155 -15158 6506 -15089
rect 6155 -17862 6224 -15158
rect 6155 -17931 6504 -17862
rect 5998 -18633 6003 -18574
rect 6062 -18633 6067 -18574
rect 5998 -23090 6067 -18633
rect 6435 -18567 6504 -17931
rect 6435 -18626 6440 -18567
rect 6499 -18626 6504 -18567
rect 6435 -19597 6504 -18626
rect 6166 -19666 6504 -19597
rect 6166 -22390 6235 -19666
rect 6166 -22459 6512 -22390
rect 5998 -23149 6003 -23090
rect 6062 -23149 6067 -23090
rect 5998 -27635 6067 -23149
rect 6443 -23065 6512 -22459
rect 6443 -23124 6448 -23065
rect 6507 -23124 6512 -23065
rect 6443 -24122 6512 -23124
rect 6155 -24191 6512 -24122
rect 6155 -26902 6224 -24191
rect 6155 -26971 6502 -26902
rect 5998 -27694 6003 -27635
rect 6062 -27694 6067 -27635
rect 5998 -32164 6067 -27694
rect 6433 -27581 6502 -26971
rect 6433 -27640 6438 -27581
rect 6497 -27640 6502 -27581
rect 6433 -28684 6502 -27640
rect 6145 -28753 6502 -28684
rect 6145 -31454 6214 -28753
rect 6145 -31523 6507 -31454
rect 6438 -32126 6507 -31523
rect 5998 -32223 6003 -32164
rect 6062 -32223 6067 -32164
rect 6433 -32131 6512 -32126
rect 6433 -32201 6438 -32131
rect 6507 -32201 6512 -32131
rect 6433 -32206 6512 -32201
rect 5998 -32228 6067 -32223
rect -14464 -34509 -8756 -34504
rect -14464 -34571 -12577 -34509
rect -12515 -34571 -8756 -34509
rect -14464 -34576 -8756 -34571
rect -14623 -34676 -12520 -34671
rect -14623 -34755 -12721 -34676
rect -12642 -34755 -12520 -34676
rect -14623 -34760 -12520 -34755
<< metal4 >>
rect -208 6040 6474 6352
rect -22644 4398 -22532 4500
rect -208 4367 104 6040
rect 6162 4462 6474 6040
rect 5006 4200 6474 4462
rect 5006 3668 6834 4200
rect -20361 -2211 -20271 1010
rect 5006 -428 5318 3668
rect 12166 2634 13912 2970
rect 13576 208 13912 2634
rect 11816 -104 13912 208
rect 12066 -128 13912 -104
rect 5006 -740 6890 -428
rect 5006 -1450 5318 -740
rect 12098 -1450 12410 -128
rect 5006 -1538 12410 -1450
rect 5006 -1730 12502 -1538
rect 13576 -1730 13912 -128
rect 5006 -1762 13912 -1730
rect 5006 -4832 5318 -1762
rect 12098 -2030 13912 -1762
rect 12166 -2066 13912 -2030
rect 13576 -4328 13912 -2066
rect 11866 -4664 13912 -4328
rect 5006 -5144 6820 -4832
rect 5006 -9450 5318 -5144
rect 13576 -6000 13912 -4664
rect 12028 -6336 13912 -6000
rect 13576 -8750 13912 -6336
rect 11866 -9086 13912 -8750
rect 5006 -9762 7020 -9450
rect -21095 -15679 -20762 -11843
rect -5026 -13504 -2152 -13388
rect -5026 -14485 -4910 -13504
rect -2268 -14530 -2152 -13504
rect 5006 -13946 5318 -9762
rect 13576 -10584 13912 -9086
rect 12014 -10920 13912 -10584
rect 13576 -13326 13912 -10920
rect 11842 -13662 13912 -13326
rect 5006 -14258 6904 -13946
rect -8554 -14870 -4983 -14707
rect -24936 -15865 -17965 -15679
rect -8554 -15766 -8391 -14870
rect -24936 -15949 -8473 -15865
rect -21891 -21721 -21621 -15949
rect -18235 -16135 -8473 -15949
rect 5006 -18520 5318 -14258
rect 13576 -15146 13912 -13662
rect 12214 -15482 13912 -15146
rect 11738 -18112 12264 -17878
rect 13576 -18112 13912 -15482
rect 11738 -18214 13912 -18112
rect 11928 -18448 13912 -18214
rect 13576 -18480 13912 -18448
rect 17292 -18212 17830 -17876
rect 17292 -18480 17628 -18212
rect 5006 -18832 6920 -18520
rect 13576 -18816 17628 -18480
rect 5006 -22982 5318 -18832
rect 13576 -19756 13912 -18816
rect 12162 -20092 13912 -19756
rect 13576 -22544 13912 -20092
rect 11814 -22880 13912 -22544
rect 5006 -23294 6904 -22982
rect 5006 -27658 5318 -23294
rect 13576 -24278 13912 -22880
rect 12224 -24614 13912 -24278
rect 13576 -26858 13912 -24614
rect 11852 -27194 13912 -26858
rect 5006 -27970 6774 -27658
rect 5006 -32178 5318 -27970
rect 13576 -28748 13912 -27194
rect 12120 -29084 13912 -28748
rect 13576 -31544 13912 -29084
rect 11824 -31880 13912 -31544
rect 5006 -32490 6962 -32178
rect 5006 -32698 5318 -32490
rect 13576 -33282 13912 -31880
rect 12158 -33618 14308 -33282
rect 13972 -35856 14308 -33618
rect 11918 -36352 12254 -36052
rect 13480 -36192 14308 -35856
rect 13972 -36352 14308 -36192
rect 11918 -36688 14308 -36352
<< metal5 >>
rect -27804 -37316 20350 6916
use 8bit_ADDER  8bit_ADDER_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/ADDER
timestamp 1736693491
transform 1 0 -24940 0 1 164
box -180 -380 26456 4515
use AND8  AND8_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/AND8
timestamp 1736693803
transform 0 -1 -23005 1 0 -24350
box 0 -2656 9584 1931
use buffer  buffer_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/inv
timestamp 1736620191
transform 0 1 12838 -1 0 -35620
box -5 -422 786 852
use left_shifter  left_shifter_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/SHIFTER
timestamp 1736620191
transform 0 -1 -3884 1 0 -22631
box 1467 -110 8528 1164
use MULT  MULT_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/MULT
timestamp 1736693491
transform 1 0 -21044 0 1 -6231
box -3818 -7001 13360 4259
use mux8  mux8_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/MUX
timestamp 1736674958
transform 1 0 7400 0 1 784
box -1848 -1184 5835 3344
use mux8  mux8_1
timestamp 1736674958
transform 1 0 7400 0 1 -3744
box -1848 -1184 5835 3344
use mux8  mux8_2
timestamp 1736674958
transform 1 0 7400 0 1 -8172
box -1848 -1184 5835 3344
use mux8  mux8_3
timestamp 1736674958
transform 1 0 7400 0 1 -12800
box -1848 -1184 5835 3344
use mux8  mux8_4
timestamp 1736674958
transform 1 0 7400 0 1 -17328
box -1848 -1184 5835 3344
use mux8  mux8_5
timestamp 1736674958
transform 1 0 7400 0 1 -21856
box -1848 -1184 5835 3344
use mux8  mux8_6
timestamp 1736674958
transform 1 0 7400 0 1 -35440
box -1848 -1184 5835 3344
use mux8  mux8_7
timestamp 1736674958
transform 1 0 7400 0 1 -26384
box -1848 -1184 5835 3344
use mux8  mux8_8
timestamp 1736674958
transform 1 0 7400 0 1 -30912
box -1848 -1184 5835 3344
use NOT8  NOT8_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NOT
timestamp 1736694824
transform 0 -1 -7411 1 0 -18944
box -110 -501 3853 1143
use OR8  OR8_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/OR
timestamp 1736694850
transform 0 -1 -18638 1 0 -27353
box 1807 -3880 12892 -390
use right_shifter  right_shifter_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/SHIFTER
timestamp 1736620191
transform 0 -1 -1168 1 0 -21808
box 1124 -110 8185 1164
use V_FLAG  V_FLAG_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/ZV_FLAG
timestamp 1736693491
transform 1 0 1839 0 1 3628
box -481 818 6282 2742
use XOR8  XOR8_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/XOR
timestamp 1736693491
transform 0 -1 -10856 1 0 -34519
box -239 -77 20622 1756
use ZFLAG  ZFLAG_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/ZV_FLAG
timestamp 1736620191
transform 1 0 15545 0 1 -20424
box -7 -79 2863 3814
<< labels >>
flabel metal3 -24908 -15649 -24849 -15604 0 FreeSans 800 0 0 0 B0
port 0 nsew
flabel metal3 -24899 -16827 -24840 -16782 0 FreeSans 800 0 0 0 B1
port 1 nsew
flabel metal3 -24910 -18036 -24851 -17991 0 FreeSans 800 0 0 0 B2
port 2 nsew
flabel metal3 -24840 -19162 -24781 -19117 0 FreeSans 800 0 0 0 B3
port 3 nsew
flabel metal3 -24887 -20352 -24828 -20307 0 FreeSans 800 0 0 0 B4
port 4 nsew
flabel metal3 -24879 -21556 -24820 -21511 0 FreeSans 800 0 0 0 B5
port 5 nsew
flabel metal3 -24879 -22857 -24820 -22812 0 FreeSans 800 0 0 0 B6
port 6 nsew
flabel metal3 -24878 -15812 -24819 -15767 0 FreeSans 800 0 0 0 A0
port 8 nsew
flabel metal3 -24898 -16988 -24839 -16943 0 FreeSans 800 0 0 0 A1
port 9 nsew
flabel metal3 -24905 -18196 -24846 -18151 0 FreeSans 800 0 0 0 A2
port 10 nsew
flabel metal3 -24846 -19319 -24787 -19274 0 FreeSans 800 0 0 0 A3
port 11 nsew
flabel metal3 -24884 -20512 -24825 -20467 0 FreeSans 800 0 0 0 A4
port 12 nsew
flabel metal3 -24902 -21706 -24843 -21661 0 FreeSans 800 0 0 0 A5
port 13 nsew
flabel metal3 -24888 -23019 -24829 -22974 0 FreeSans 800 0 0 0 A6
port 15 nsew
flabel metal3 -24885 -24327 -24826 -24282 0 FreeSans 800 0 0 0 A7
port 16 nsew
flabel metal1 13169 -3047 13216 -2964 0 FreeSans 800 0 0 0 Y0
port 17 nsew
flabel metal1 13172 -7413 13219 -7330 0 FreeSans 800 0 0 0 Y1
port 18 nsew
flabel metal1 13183 -12104 13230 -12021 0 FreeSans 800 0 0 0 Y2
port 20 nsew
flabel metal1 13178 -16546 13225 -16463 0 FreeSans 800 0 0 0 Y3
port 21 nsew
flabel metal1 13181 -21117 13228 -21034 0 FreeSans 800 0 0 0 Y4
port 22 nsew
flabel metal1 13179 -25614 13226 -25531 0 FreeSans 800 0 0 0 Y5
port 23 nsew
flabel metal1 13178 -30106 13225 -30058 0 FreeSans 800 0 0 0 Y6
port 24 nsew
flabel metal1 13035 -36363 13082 -36280 0 FreeSans 800 0 0 0 S
port 26 nsew
flabel metal1 18354 -18573 18391 -18471 0 FreeSans 800 0 0 0 Z
port 27 nsew
flabel metal1 13152 1469 13208 1558 0 FreeSans 800 0 0 0 C
port 28 nsew
flabel metal1 8026 5020 8106 5116 0 FreeSans 1600 0 0 0 V
port 29 nsew
flabel metal4 5732 4158 5880 4280 0 FreeSans 1600 0 0 0 VDD
port 30 nsew
flabel metal5 8982 4290 9670 4732 0 FreeSans 1600 0 0 0 VSS
port 32 nsew
flabel metal1 13172 -34752 13202 -34724 0 FreeSans 1600 0 0 0 Y7
port 34 nsew
flabel metal1 -9072 -16096 -8778 -16087 0 FreeSans 1600 0 0 0 VDD
flabel metal1 -9072 -16096 -8778 -16087 0 FreeSans 1600 0 0 0 VDD
flabel metal3 -25060 -24176 -24986 -24108 0 FreeSans 1600 0 0 0 B7
port 36 nsew
<< end >>
