magic
tech sky130B
magscale 1 2
timestamp 1736596529
<< metal1 >>
rect 1807 -1356 1873 -467
rect 1927 -1251 1993 -467
rect 1927 -1317 2066 -1251
rect 1807 -1422 2066 -1356
rect 2986 -2245 3055 -1586
rect 5726 -2126 5795 -1586
rect 6905 -2126 6974 -1606
rect 8325 -1886 8394 -1586
rect 9965 -1866 10034 -1546
rect 5726 -2195 6323 -2126
rect 2986 -2314 5843 -2245
rect 6254 -2305 6323 -2195
rect 6714 -2195 6974 -2126
rect 7174 -1955 8394 -1886
rect 8445 -1935 10034 -1866
rect 6714 -2305 6783 -2195
rect 7174 -2305 7243 -1955
rect 8445 -2026 8514 -1935
rect 11385 -1986 11454 -1566
rect 7654 -2095 8514 -2026
rect 8634 -2055 11454 -1986
rect 7654 -2305 7723 -2095
rect 8634 -2305 8703 -2055
rect 12705 -2146 12774 -1586
rect 9134 -2215 12774 -2146
rect 9134 -2305 9203 -2215
use nor2  nor2_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NOR/NOR2
timestamp 1736020690
transform 1 0 11800 0 1 -1320
box 0 -480 1090 580
use nor2  nor2_1
timestamp 1736020690
transform 1 0 2000 0 1 -1320
box 0 -480 1090 580
use nor2  nor2_2
timestamp 1736020690
transform 1 0 3400 0 1 -1320
box 0 -480 1090 580
use nor2  nor2_3
timestamp 1736020690
transform 1 0 4800 0 1 -1320
box 0 -480 1090 580
use nor2  nor2_4
timestamp 1736020690
transform 1 0 6200 0 1 -1320
box 0 -480 1090 580
use nor2  nor2_5
timestamp 1736020690
transform 1 0 7600 0 1 -1320
box 0 -480 1090 580
use nor2  nor2_6
timestamp 1736020690
transform 1 0 9000 0 1 -1320
box 0 -480 1090 580
use nor2  nor2_7
timestamp 1736020690
transform 1 0 10400 0 1 -1320
box 0 -480 1090 580
use NOT8  NOT8_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NOT
timestamp 1736595726
transform 1 0 5850 0 1 -3379
box -110 -501 3853 1143
<< end >>
