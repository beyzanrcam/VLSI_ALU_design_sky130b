magic
tech sky130B
magscale 1 2
timestamp 1736680159
<< nwell >>
rect -292 625 2999 1536
rect -292 -679 2999 -159
<< poly >>
rect -118 660 74 717
rect -118 550 -99 660
rect -52 550 74 660
rect -118 458 74 550
rect 1413 615 1729 630
rect 1413 475 1458 615
rect 1531 475 1729 615
rect 1413 458 1729 475
<< polycont >>
rect -99 550 -52 660
rect 1458 475 1531 615
<< locali >>
rect -117 660 -32 683
rect -117 550 -99 660
rect -52 550 -32 660
rect -117 530 -32 550
rect 1358 608 1392 625
rect 1439 615 1548 630
rect 1358 511 1383 608
rect 1358 495 1392 511
rect 1439 475 1458 615
rect 1531 475 1548 615
rect 1439 458 1548 475
<< viali >>
rect -99 550 -52 660
rect 1458 512 1531 615
<< metal1 >>
rect -117 660 18 684
rect -117 550 -99 660
rect -3 552 18 660
rect 1357 625 1548 630
rect -52 550 18 552
rect -117 530 18 550
rect 1356 615 1548 625
rect 1356 608 1458 615
rect 1531 608 1548 615
rect 1356 511 1383 608
rect 1533 511 1548 608
rect 1356 495 1548 511
rect 1519 420 1724 446
rect 1519 323 1559 420
rect 1675 323 1724 420
rect 1519 303 1724 323
rect 2862 316 3108 525
rect 2999 129 3108 316
rect 2999 43 3008 129
rect 3099 43 3108 129
rect 2999 31 3108 43
rect -93 -86 1135 -70
rect -93 -155 1020 -86
rect 1119 -155 1135 -86
rect -93 -161 1135 -155
rect 1518 -82 2995 -70
rect 1518 -148 1532 -82
rect 1603 -148 2995 -82
rect 1518 -161 2995 -148
rect 401 -277 675 -268
rect 401 -349 410 -277
rect 666 -349 675 -277
rect 401 -358 675 -349
rect 1690 -277 1964 -268
rect 1690 -349 1699 -277
rect 1955 -349 1964 -277
rect 1690 -358 1964 -349
rect 2407 -277 2681 -268
rect 2407 -349 2416 -277
rect 2672 -349 2681 -277
rect 2407 -358 2681 -349
rect 189 -673 353 -646
rect 189 -753 221 -673
rect 319 -753 353 -673
rect 189 -781 353 -753
rect 1298 -674 1462 -651
rect 1298 -754 1332 -674
rect 1430 -754 1462 -674
rect 1298 -781 1462 -754
rect 1826 -759 2243 -669
rect -7 -866 384 -809
rect -7 -932 12 -866
rect 265 -932 384 -866
rect -7 -946 384 -932
rect 477 -1023 830 -1010
rect 1722 -1016 1784 -997
rect 477 -1075 486 -1023
rect 821 -1075 830 -1023
rect 477 -1084 830 -1075
rect 1711 -1028 1795 -1016
rect 1711 -1090 1722 -1028
rect 1784 -1090 1795 -1028
rect 1711 -1101 1795 -1090
rect 2576 -1055 2654 -1042
rect 2576 -1107 2589 -1055
rect 2641 -1107 2654 -1055
rect 2576 -1120 2654 -1107
<< via1 >>
rect -93 552 -52 660
rect -52 552 -3 660
rect 1383 512 1458 608
rect 1458 512 1531 608
rect 1531 512 1533 608
rect 1383 511 1533 512
rect 4 319 80 427
rect 1559 323 1675 420
rect 3008 43 3099 129
rect 1020 -155 1119 -86
rect 1532 -148 1603 -82
rect 410 -349 666 -277
rect 1699 -349 1955 -277
rect 2416 -349 2672 -277
rect 221 -753 319 -673
rect 776 -760 859 -612
rect 1332 -754 1430 -674
rect 2753 -742 2873 -662
rect 12 -932 265 -866
rect 1322 -937 1507 -877
rect 2194 -903 2339 -828
rect 486 -1075 821 -1023
rect 1722 -1090 1784 -1028
rect 2589 -1107 2641 -1055
<< metal2 >>
rect -292 440 -183 1536
rect -117 683 -3 1536
rect -117 660 286 683
rect -117 552 -93 660
rect -3 552 286 660
rect -117 530 286 552
rect -117 529 -3 530
rect -292 439 65 440
rect -292 427 94 439
rect -292 327 4 427
rect -18 319 4 327
rect 80 319 94 427
rect -18 -846 83 319
rect 190 -646 286 530
rect 1299 608 1571 624
rect 1299 511 1383 608
rect 1533 511 1571 608
rect 1299 476 1571 511
rect 1004 -86 1135 -70
rect 1004 -155 1020 -86
rect 1119 -155 1135 -86
rect 401 -277 675 -268
rect 401 -349 410 -277
rect 666 -349 675 -277
rect 401 -358 675 -349
rect 763 -612 872 -597
rect 189 -673 353 -646
rect 189 -753 221 -673
rect 319 -753 353 -673
rect 189 -781 353 -753
rect 763 -760 776 -612
rect 859 -760 872 -612
rect 763 -772 872 -760
rect -18 -866 353 -846
rect -18 -932 12 -866
rect 265 -932 353 -866
rect -18 -945 353 -932
rect 477 -1019 830 -1010
rect 477 -1075 486 -1019
rect 821 -1075 830 -1019
rect 477 -1084 830 -1075
rect 1004 -1158 1135 -155
rect 1299 -651 1395 476
rect 1518 420 1724 446
rect 1518 323 1559 420
rect 1675 323 1724 420
rect 1518 303 1724 323
rect 1518 -82 1613 303
rect 1518 -148 1532 -82
rect 1603 -148 1613 -82
rect 1298 -674 1462 -651
rect 1298 -754 1332 -674
rect 1430 -754 1462 -674
rect 1298 -781 1462 -754
rect 1518 -862 1613 -148
rect 2999 129 3108 138
rect 2999 43 3008 129
rect 3099 43 3108 129
rect 1690 -277 1964 -268
rect 1690 -349 1699 -277
rect 1955 -349 1964 -277
rect 1690 -358 1964 -349
rect 2407 -277 2681 -268
rect 2407 -349 2416 -277
rect 2672 -349 2681 -277
rect 2407 -358 2681 -349
rect 2708 -662 2886 -611
rect 2708 -742 2753 -662
rect 2873 -742 2886 -662
rect 2708 -759 2886 -742
rect 1298 -877 1613 -862
rect 1298 -937 1322 -877
rect 1507 -937 1613 -877
rect 2182 -828 2357 -817
rect 2182 -903 2194 -828
rect 2339 -903 2357 -828
rect 2182 -915 2357 -903
rect 1298 -947 1613 -937
rect 1711 -1028 1795 -1016
rect 1711 -1090 1722 -1028
rect 1784 -1090 1795 -1028
rect 1711 -1101 1795 -1090
rect 2576 -1053 2654 -1042
rect 2576 -1109 2587 -1053
rect 2643 -1109 2654 -1053
rect 2576 -1120 2654 -1109
rect 2708 -1158 2828 -759
rect 2999 -1099 3108 43
rect 1004 -1260 2828 -1158
<< via2 >>
rect 410 -349 666 -277
rect 776 -760 859 -612
rect 486 -1023 821 -1019
rect 486 -1075 821 -1023
rect 1699 -349 1955 -277
rect 2416 -349 2672 -277
rect 2194 -903 2339 -828
rect 1722 -1090 1784 -1028
rect 2587 -1055 2643 -1053
rect 2587 -1107 2589 -1055
rect 2589 -1107 2641 -1055
rect 2641 -1107 2643 -1055
rect 2587 -1109 2643 -1107
<< metal3 >>
rect 401 -277 675 -268
rect 401 -349 410 -277
rect 666 -349 675 -277
rect 401 -358 675 -349
rect 1690 -277 1964 -268
rect 1690 -349 1699 -277
rect 1955 -349 1964 -277
rect 1690 -358 1964 -349
rect 2407 -277 2681 -268
rect 2407 -349 2416 -277
rect 2672 -349 2681 -277
rect 2407 -358 2681 -349
rect 759 -612 881 -579
rect 759 -760 776 -612
rect 859 -760 881 -612
rect 759 -813 881 -760
rect 759 -828 2360 -813
rect 759 -903 2194 -828
rect 2339 -903 2360 -828
rect 759 -915 2360 -903
rect 477 -1011 830 -1010
rect 477 -1075 486 -1011
rect 821 -1075 830 -1011
rect 477 -1084 830 -1075
rect 1697 -1023 1809 -1009
rect 1697 -1095 1717 -1023
rect 1789 -1095 1809 -1023
rect 1697 -1106 1809 -1095
rect 2564 -1048 2667 -1034
rect 2564 -1114 2582 -1048
rect 2648 -1114 2667 -1048
rect 2564 -1132 2667 -1114
<< via3 >>
rect 410 -349 666 -277
rect 1699 -349 1955 -277
rect 2416 -349 2672 -277
rect 486 -1019 821 -1011
rect 486 -1075 821 -1019
rect 1717 -1028 1789 -1023
rect 1717 -1090 1722 -1028
rect 1722 -1090 1784 -1028
rect 1784 -1090 1789 -1028
rect 1717 -1095 1789 -1090
rect 2582 -1053 2648 -1048
rect 2582 -1109 2587 -1053
rect 2587 -1109 2643 -1053
rect 2643 -1109 2648 -1053
rect 2582 -1114 2648 -1109
<< metal4 >>
rect 597 1497 723 1536
rect 597 1371 2272 1497
rect 1418 -268 1596 1371
rect 401 -277 2681 -268
rect 401 -349 410 -277
rect 666 -349 1699 -277
rect 1955 -349 2416 -277
rect 2672 -349 2681 -277
rect 401 -358 2681 -349
rect 477 -1075 486 -1010
rect 821 -1075 830 -1010
rect 477 -1084 830 -1075
<< via4 >>
rect 486 -1011 821 -821
rect 486 -1057 821 -1011
rect 1617 -1023 1889 -923
rect 1617 -1095 1717 -1023
rect 1717 -1095 1789 -1023
rect 1789 -1095 1889 -1023
rect 1617 -1195 1889 -1095
rect 2479 -1048 2751 -945
rect 2479 -1114 2582 -1048
rect 2582 -1114 2648 -1048
rect 2648 -1114 2751 -1048
rect 2479 -1217 2751 -1114
<< metal5 >>
rect -166 -821 2994 1536
rect -166 -1057 486 -821
rect 821 -923 2994 -821
rect 821 -1057 1617 -923
rect -166 -1195 1617 -1057
rect 1889 -945 2994 -923
rect 1889 -1195 2479 -945
rect -166 -1217 2479 -1195
rect 2751 -1217 2994 -945
rect -166 -1421 2994 -1217
use NAND2  NAND2_0 ~/Desktop/vlsi_sky130b/design/mag/NAND/NAND2
timestamp 1736620191
transform 1 0 -167 0 1 -1051
box 356 -17 1062 804
use NAND2  NAND2_1
timestamp 1736620191
transform 1 0 942 0 1 -1051
box 356 -17 1062 804
use NAND2  NAND2_2
timestamp 1736620191
transform 1 0 1824 0 1 -1051
box 356 -17 1062 804
use XOR2  XOR2_0 ~/Desktop/vlsi_sky130b/design/mag/XOR
timestamp 1736620191
transform 1 0 69 0 1 -239
box -109 77 1371 1764
use XOR2  XOR2_1
timestamp 1736620191
transform 1 0 1628 0 1 -239
box -109 77 1371 1764
<< labels >>
rlabel metal1 -80 -152 -44 -82 5 COUT
port 4 s
rlabel metal2 3014 -1066 3094 -986 5 OUT
port 5 s
rlabel metal1 2808 -144 2958 -100 5 CIN
port 6 s
rlabel metal5 433 -1321 834 -1244 5 VSS
port 8 s
rlabel metal2 -279 1470 -199 1529 5 A
port 9 s
rlabel metal2 -102 1470 -22 1529 5 B
port 10 s
rlabel metal4 1355 1383 1610 1485 5 VDD
port 11 s
<< end >>
