magic
tech sky130A
magscale 1 2
timestamp 1736606925
<< nwell >>
rect 6413 2450 6512 2634
rect 9708 2491 9799 2635
<< metal1 >>
rect -174 3005 9807 3089
rect -174 2858 6517 2942
rect -174 2710 3226 2794
rect 3117 2633 3226 2710
rect 3117 2538 3129 2633
rect 3218 2538 3226 2633
rect 3117 2527 3226 2538
rect 6407 2634 6517 2858
rect 6407 2450 6413 2634
rect 6512 2450 6517 2634
rect 9699 2635 9807 3005
rect 9699 2491 9708 2635
rect 9799 2491 9807 2635
rect 9699 2480 9807 2491
rect 6407 2443 6517 2450
rect -160 1063 49 1083
rect -160 961 -130 1063
rect -12 961 49 1063
rect -160 931 49 961
rect 3113 953 3316 1044
rect 6404 953 6607 1044
rect 9695 953 9898 1044
rect 12934 91 12983 1042
rect 12986 953 13189 1044
rect 12441 1 12992 91
rect 12934 -3 12983 1
<< via1 >>
rect 3129 2538 3218 2633
rect 6413 2450 6512 2634
rect 9708 2491 9799 2635
rect -130 961 -12 1063
<< metal2 >>
rect -174 1500 -96 1640
rect -166 1063 19 1079
rect -166 961 -130 1063
rect -12 961 19 1063
rect -166 -125 19 961
rect 12985 16 13185 127
use FULL_ADDER  FULL_ADDER_0
timestamp 1736606925
transform 1 0 118 0 1 1114
box -292 -1260 3108 1536
use FULL_ADDER  FULL_ADDER_1
timestamp 1736606925
transform 1 0 3409 0 1 1114
box -292 -1260 3108 1536
use FULL_ADDER  FULL_ADDER_2
timestamp 1736606925
transform 1 0 6700 0 1 1114
box -292 -1260 3108 1536
use FULL_ADDER  FULL_ADDER_3
timestamp 1736606925
transform 1 0 9991 0 1 1114
box -292 -1260 3108 1536
<< end >>
