magic
tech sky130B
magscale 1 2
timestamp 1736187666
<< nwell >>
rect -292 625 2999 1536
rect -292 -679 2999 -159
<< poly >>
rect 2110 2501 2361 2506
rect 1704 2489 2361 2501
rect 1704 2269 2142 2489
rect 2334 2269 2361 2489
rect 1704 2243 2361 2269
rect 1704 2242 2351 2243
rect -118 660 74 717
rect -118 550 -99 660
rect -52 550 74 660
rect -118 458 74 550
rect 1413 615 1729 630
rect 1413 475 1458 615
rect 1531 475 1729 615
rect 1413 458 1729 475
<< polycont >>
rect 2142 2269 2334 2489
rect -99 550 -52 660
rect 1458 475 1531 615
<< locali >>
rect 2110 2489 2361 2506
rect 2110 2269 2142 2489
rect 2334 2269 2361 2489
rect 2110 2243 2361 2269
rect -117 660 -32 683
rect -117 550 -99 660
rect -52 550 -32 660
rect -117 530 -32 550
rect 1358 608 1392 625
rect 1439 615 1548 630
rect 1358 511 1383 608
rect 1358 495 1392 511
rect 1439 475 1458 615
rect 1531 475 1548 615
rect 1439 458 1548 475
<< viali >>
rect 2185 2346 2305 2488
rect -99 550 -52 660
rect 1458 512 1531 615
<< metal1 >>
rect 2166 2489 2324 3297
rect 2142 2488 2334 2489
rect 2142 2346 2185 2488
rect 2305 2346 2334 2488
rect -3 2271 656 2309
rect -3 2131 31 2271
rect 625 2131 656 2271
rect 2142 2269 2334 2346
rect 2391 2230 2566 3281
rect -3 2100 656 2131
rect 1931 2087 2566 2230
rect -117 660 18 684
rect -117 550 -99 660
rect -3 552 18 660
rect 1357 625 1548 630
rect -52 550 18 552
rect -117 530 18 550
rect 1356 615 1548 625
rect 1356 608 1458 615
rect 1531 608 1548 615
rect 1356 511 1383 608
rect 1533 511 1548 608
rect 1356 495 1548 511
rect 1519 420 1724 446
rect 1519 323 1559 420
rect 1675 323 1724 420
rect 1519 303 1724 323
rect 2862 316 3108 525
rect 2999 129 3108 316
rect 2999 43 3008 129
rect 3099 43 3108 129
rect 2999 31 3108 43
rect -93 -86 1135 -70
rect -93 -155 1020 -86
rect 1119 -155 1135 -86
rect -93 -161 1135 -155
rect 1518 -82 2995 -70
rect 1518 -148 1532 -82
rect 1603 -148 2995 -82
rect 1518 -161 2995 -148
rect 189 -673 353 -646
rect 189 -753 221 -673
rect 319 -753 353 -673
rect 189 -781 353 -753
rect 1298 -674 1462 -651
rect 1298 -754 1332 -674
rect 1430 -754 1462 -674
rect 1298 -781 1462 -754
rect 1826 -759 2243 -669
rect -7 -866 384 -809
rect -7 -932 12 -866
rect 265 -932 384 -866
rect -7 -946 384 -932
<< via1 >>
rect 31 2131 625 2271
rect -93 552 -52 660
rect -52 552 -3 660
rect 1383 512 1458 608
rect 1458 512 1531 608
rect 1531 512 1533 608
rect 1383 511 1533 512
rect 4 319 80 427
rect 1559 323 1675 420
rect 3008 43 3099 129
rect 1020 -155 1119 -86
rect 1532 -148 1603 -82
rect 221 -753 319 -673
rect 776 -760 859 -612
rect 1332 -754 1430 -674
rect 2753 -742 2873 -662
rect 12 -932 265 -866
rect 1322 -937 1507 -877
rect 2194 -903 2339 -828
<< metal2 >>
rect -292 440 -183 2731
rect -117 2271 656 2309
rect -117 2131 31 2271
rect 625 2131 656 2271
rect -117 2100 656 2131
rect -117 683 -3 2100
rect -117 660 286 683
rect -117 552 -93 660
rect -3 552 286 660
rect -117 530 286 552
rect -117 529 -3 530
rect -292 439 65 440
rect -292 427 94 439
rect -292 327 4 427
rect -7 319 4 327
rect 80 319 94 427
rect -7 -846 94 319
rect 190 -646 286 530
rect 1299 608 1571 624
rect 1299 511 1383 608
rect 1533 511 1571 608
rect 1299 476 1571 511
rect 1004 -86 1135 -70
rect 1004 -155 1020 -86
rect 1119 -155 1135 -86
rect 763 -612 872 -597
rect 189 -673 353 -646
rect 189 -753 221 -673
rect 319 -753 353 -673
rect 189 -781 353 -753
rect 763 -760 776 -612
rect 859 -760 872 -612
rect 763 -772 872 -760
rect -7 -866 353 -846
rect -7 -932 12 -866
rect 265 -932 353 -866
rect -7 -945 353 -932
rect 1004 -1158 1135 -155
rect 1299 -651 1395 476
rect 1518 420 1724 446
rect 1518 323 1559 420
rect 1675 323 1724 420
rect 1518 303 1724 323
rect 1518 -82 1613 303
rect 1518 -148 1532 -82
rect 1603 -148 1613 -82
rect 1298 -674 1462 -651
rect 1298 -754 1332 -674
rect 1430 -754 1462 -674
rect 1298 -781 1462 -754
rect 1518 -862 1613 -148
rect 2999 129 3108 138
rect 2999 43 3008 129
rect 3099 43 3108 129
rect 2708 -662 2886 -611
rect 2708 -742 2753 -662
rect 2873 -742 2886 -662
rect 2708 -759 2886 -742
rect 1298 -877 1613 -862
rect 1298 -937 1322 -877
rect 1507 -937 1613 -877
rect 2182 -828 2357 -817
rect 2182 -903 2194 -828
rect 2339 -903 2357 -828
rect 2182 -915 2357 -903
rect 1298 -947 1613 -937
rect 2708 -1158 2828 -759
rect 2999 -1099 3108 43
rect 1004 -1260 2828 -1158
<< via2 >>
rect 776 -760 859 -612
rect 2194 -903 2339 -828
<< metal3 >>
rect 759 -612 881 -579
rect 759 -760 776 -612
rect 859 -760 881 -612
rect 759 -813 881 -760
rect 759 -828 2360 -813
rect 759 -903 2194 -828
rect 2339 -903 2360 -828
rect 759 -915 2360 -903
use NAND2  NAND2_0
timestamp 1736181444
transform 1 0 -167 0 1 -1051
box 356 -63 1062 892
use NAND2  NAND2_1
timestamp 1736181444
transform 1 0 942 0 1 -1051
box 356 -63 1062 892
use NAND2  NAND2_2
timestamp 1736181444
transform 1 0 1824 0 1 -1051
box 356 -63 1062 892
use XOR2  XOR2_0
timestamp 1736181444
transform 1 0 69 0 1 -239
box -109 222 1371 1764
use XOR2  XOR2_1
timestamp 1736181444
transform 1 0 1628 0 1 -239
box -109 222 1371 1764
use XOR2  XOR2_2
timestamp 1736181444
transform -1 0 2027 0 1 1545
box -109 222 1371 1764
<< end >>
