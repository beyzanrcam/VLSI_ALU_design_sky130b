magic
tech sky130B
magscale 1 2
timestamp 1736020054
<< nwell >>
rect -602 991 790 1966
<< nmos >>
rect -10 429 20 629
rect 86 429 116 629
rect 182 429 212 629
rect 278 429 308 629
<< pmos >>
rect -394 1047 -364 1903
rect -298 1047 -268 1903
rect -202 1047 -172 1903
rect -106 1047 -76 1903
rect -10 1047 20 1903
rect 86 1047 116 1903
rect 182 1047 212 1903
rect 278 1047 308 1903
rect 374 1047 404 1903
rect 470 1047 500 1903
rect 566 1047 596 1903
rect 662 1047 692 1903
<< ndiff >>
rect -72 617 -10 629
rect -72 441 -60 617
rect -26 441 -10 617
rect -72 429 -10 441
rect 20 617 86 629
rect 20 441 36 617
rect 70 441 86 617
rect 20 429 86 441
rect 116 617 182 629
rect 116 441 132 617
rect 166 441 182 617
rect 116 429 182 441
rect 212 617 278 629
rect 212 441 228 617
rect 262 441 278 617
rect 212 429 278 441
rect 308 617 370 629
rect 308 441 324 617
rect 358 441 370 617
rect 308 429 370 441
<< pdiff >>
rect -456 1891 -394 1903
rect -456 1059 -444 1891
rect -410 1059 -394 1891
rect -456 1047 -394 1059
rect -364 1891 -298 1903
rect -364 1059 -348 1891
rect -314 1059 -298 1891
rect -364 1047 -298 1059
rect -268 1891 -202 1903
rect -268 1059 -252 1891
rect -218 1059 -202 1891
rect -268 1047 -202 1059
rect -172 1891 -106 1903
rect -172 1059 -156 1891
rect -122 1059 -106 1891
rect -172 1047 -106 1059
rect -76 1891 -10 1903
rect -76 1059 -60 1891
rect -26 1059 -10 1891
rect -76 1047 -10 1059
rect 20 1891 86 1903
rect 20 1059 36 1891
rect 70 1059 86 1891
rect 20 1047 86 1059
rect 116 1891 182 1903
rect 116 1059 132 1891
rect 166 1059 182 1891
rect 116 1047 182 1059
rect 212 1891 278 1903
rect 212 1059 228 1891
rect 262 1059 278 1891
rect 212 1047 278 1059
rect 308 1891 374 1903
rect 308 1059 324 1891
rect 358 1059 374 1891
rect 308 1047 374 1059
rect 404 1891 470 1903
rect 404 1059 420 1891
rect 454 1059 470 1891
rect 404 1047 470 1059
rect 500 1891 566 1903
rect 500 1059 516 1891
rect 550 1059 566 1891
rect 500 1047 566 1059
rect 596 1891 662 1903
rect 596 1059 612 1891
rect 646 1059 662 1891
rect 596 1047 662 1059
rect 692 1891 754 1903
rect 692 1059 708 1891
rect 742 1059 754 1891
rect 692 1047 754 1059
<< ndiffc >>
rect -60 441 -26 617
rect 36 441 70 617
rect 132 441 166 617
rect 228 441 262 617
rect 324 441 358 617
<< pdiffc >>
rect -444 1059 -410 1891
rect -348 1059 -314 1891
rect -252 1059 -218 1891
rect -156 1059 -122 1891
rect -60 1059 -26 1891
rect 36 1059 70 1891
rect 132 1059 166 1891
rect 228 1059 262 1891
rect 324 1059 358 1891
rect 420 1059 454 1891
rect 516 1059 550 1891
rect 612 1059 646 1891
rect 708 1059 742 1891
<< psubdiff >>
rect -72 307 370 375
rect -72 194 -8 307
rect 322 194 370 307
rect -72 118 370 194
<< nsubdiff >>
rect -566 1413 -456 1903
rect -566 1059 -516 1413
rect -482 1059 -456 1413
rect -566 1047 -456 1059
<< psubdiffcont >>
rect -8 194 322 307
<< nsubdiffcont >>
rect -516 1059 -482 1413
<< poly >>
rect -394 1903 -364 1929
rect -298 1903 -268 1929
rect -202 1903 -172 1929
rect -106 1903 -76 1929
rect -10 1903 20 1929
rect 86 1903 116 1929
rect 182 1903 212 1929
rect 278 1903 308 1929
rect 374 1903 404 1929
rect 470 1903 500 1929
rect 566 1903 596 1929
rect 662 1903 692 1929
rect -394 1021 -364 1047
rect -298 1021 -268 1047
rect -202 1021 -172 1047
rect -394 1000 -172 1021
rect -394 991 -222 1000
rect -238 966 -222 991
rect -188 966 -172 1000
rect -106 1021 -76 1047
rect -10 1021 20 1047
rect 86 1021 116 1047
rect -106 1000 116 1021
rect -106 991 66 1000
rect -238 950 -172 966
rect 50 966 66 991
rect 100 966 116 1000
rect 50 950 116 966
rect -202 674 -172 950
rect -202 644 20 674
rect -10 629 20 644
rect 86 629 116 950
rect 182 1021 212 1047
rect 278 1021 308 1047
rect 374 1021 404 1047
rect 182 1000 404 1021
rect 182 966 198 1000
rect 232 991 404 1000
rect 470 1021 500 1047
rect 566 1021 596 1047
rect 662 1021 692 1047
rect 470 991 692 1021
rect 232 966 248 991
rect 182 950 248 966
rect 182 629 212 950
rect 470 734 500 991
rect 434 718 500 734
rect 434 697 450 718
rect 278 684 450 697
rect 484 684 500 718
rect 278 667 500 684
rect 278 629 308 667
rect -10 403 20 429
rect 86 403 116 429
rect 182 403 212 429
rect 278 403 308 429
<< polycont >>
rect -222 966 -188 1000
rect 66 966 100 1000
rect 198 966 232 1000
rect 450 684 484 718
<< locali >>
rect -444 1891 -410 1907
rect -516 1413 -482 1429
rect -516 1043 -482 1059
rect -444 1043 -410 1059
rect -348 1891 -314 1907
rect -348 1043 -314 1059
rect -252 1891 -218 1907
rect -252 1043 -218 1059
rect -156 1891 -122 1907
rect -156 1043 -122 1059
rect -60 1891 -26 1907
rect -60 1043 -26 1059
rect 36 1891 70 1907
rect 36 1043 70 1059
rect 132 1891 166 1907
rect 132 1043 166 1059
rect 228 1891 262 1907
rect 228 1043 262 1059
rect 324 1891 358 1907
rect 324 1043 358 1059
rect 420 1891 454 1907
rect 420 1043 454 1059
rect 516 1891 550 1907
rect 516 1043 550 1059
rect 612 1891 646 1907
rect 612 1043 646 1059
rect 708 1891 742 1907
rect 708 1043 742 1059
rect -238 966 -222 1000
rect -188 966 -172 1000
rect 50 966 66 1000
rect 100 966 116 1000
rect 182 966 198 1000
rect 232 966 248 1000
rect 434 684 450 718
rect 484 684 500 718
rect -60 617 -26 633
rect -60 375 -26 441
rect 36 617 70 633
rect 36 425 70 441
rect 132 617 166 633
rect 132 375 166 441
rect 228 617 262 633
rect 228 425 262 441
rect 324 617 358 633
rect 324 375 358 441
rect -60 307 358 375
rect -60 194 -8 307
rect 322 194 358 307
rect -60 146 358 194
<< viali >>
rect -516 1059 -482 1413
rect -444 1059 -410 1413
rect -348 1535 -314 1891
rect -252 1059 -218 1413
rect -156 1535 -122 1891
rect -60 1059 -26 1413
rect 36 1535 70 1891
rect 132 1059 166 1413
rect 228 1535 262 1891
rect 324 1059 358 1413
rect 420 1535 454 1891
rect 516 1059 550 1413
rect 612 1535 646 1891
rect 708 1059 742 1413
rect -222 966 -188 1000
rect 66 966 100 1000
rect 198 966 232 1000
rect 450 684 484 718
rect 36 441 70 617
rect 228 441 262 617
rect -8 194 322 307
<< metal1 >>
rect -354 1891 76 1903
rect -354 1535 -348 1891
rect -314 1535 -156 1891
rect -122 1535 36 1891
rect 70 1535 76 1891
rect -354 1523 76 1535
rect 222 1891 652 1903
rect 222 1535 228 1891
rect 262 1535 420 1891
rect 454 1535 612 1891
rect 646 1535 652 1891
rect 222 1523 652 1535
rect -531 1413 -212 1425
rect -531 1059 -516 1413
rect -482 1059 -444 1413
rect -410 1059 -252 1413
rect -218 1059 -212 1413
rect -531 1047 -212 1059
rect -66 1413 364 1425
rect -66 1059 -60 1413
rect -26 1059 132 1413
rect 166 1059 324 1413
rect 358 1059 364 1413
rect -66 1047 364 1059
rect 510 1413 748 1425
rect 510 1059 516 1413
rect 550 1059 708 1413
rect 742 1059 748 1413
rect 510 1047 748 1059
rect 611 1016 748 1047
rect -602 1000 -172 1016
rect -602 966 -222 1000
rect -188 966 -172 1000
rect -602 950 -172 966
rect -141 1000 116 1016
rect -141 966 66 1000
rect 100 966 116 1000
rect -141 950 116 966
rect 182 1000 248 1016
rect 182 966 198 1000
rect 232 966 248 1000
rect -141 922 -75 950
rect 182 922 248 966
rect -602 856 -75 922
rect -42 856 248 922
rect 611 950 790 1016
rect -42 828 25 856
rect -602 762 25 828
rect -602 718 500 734
rect -602 684 450 718
rect 484 684 500 718
rect -602 668 500 684
rect 611 629 748 950
rect 30 617 748 629
rect 30 441 36 617
rect 70 441 228 617
rect 262 441 748 617
rect 30 429 748 441
rect -20 307 334 317
rect -20 194 -8 307
rect 322 194 334 307
rect -20 187 334 194
<< labels >>
rlabel metal1 -602 981 -602 981 3 A
port 6 e
rlabel metal1 -602 889 -602 889 3 B
port 7 e
rlabel metal1 -602 793 -602 793 3 C
port 8 e
rlabel metal1 -602 698 -602 698 3 D
port 9 e
rlabel metal1 158 187 158 187 5 VSS
port 10 s
rlabel metal1 -531 1235 -531 1235 5 VDD
port 11 s
rlabel metal1 790 982 790 982 3 Y
port 12 e
<< end >>
