magic
tech sky130B
magscale 1 2
timestamp 1736019897
<< error_p >>
rect -641 -484 641 491
<< nwell >>
rect -641 -484 641 491
<< pmos >>
rect -543 -428 -513 428
rect -447 -428 -417 428
rect -351 -428 -321 428
rect -255 -428 -225 428
rect -159 -428 -129 428
rect -63 -428 -33 428
rect 33 -428 63 428
rect 129 -428 159 428
rect 225 -428 255 428
rect 321 -428 351 428
rect 417 -428 447 428
rect 513 -428 543 428
<< pdiff >>
rect -605 416 -543 428
rect -605 -416 -593 416
rect -559 -416 -543 416
rect -605 -428 -543 -416
rect -513 416 -447 428
rect -513 -416 -497 416
rect -463 -416 -447 416
rect -513 -428 -447 -416
rect -417 416 -351 428
rect -417 -416 -401 416
rect -367 -416 -351 416
rect -417 -428 -351 -416
rect -321 416 -255 428
rect -321 -416 -305 416
rect -271 -416 -255 416
rect -321 -428 -255 -416
rect -225 416 -159 428
rect -225 -416 -209 416
rect -175 -416 -159 416
rect -225 -428 -159 -416
rect -129 416 -63 428
rect -129 -416 -113 416
rect -79 -416 -63 416
rect -129 -428 -63 -416
rect -33 416 33 428
rect -33 -416 -17 416
rect 17 -416 33 416
rect -33 -428 33 -416
rect 63 416 129 428
rect 63 -416 79 416
rect 113 -416 129 416
rect 63 -428 129 -416
rect 159 416 225 428
rect 159 -416 175 416
rect 209 -416 225 416
rect 159 -428 225 -416
rect 255 416 321 428
rect 255 -416 271 416
rect 305 -416 321 416
rect 255 -428 321 -416
rect 351 416 417 428
rect 351 -416 367 416
rect 401 -416 417 416
rect 351 -428 417 -416
rect 447 416 513 428
rect 447 -416 463 416
rect 497 -416 513 416
rect 447 -428 513 -416
rect 543 416 605 428
rect 543 -416 559 416
rect 593 -416 605 416
rect 543 -428 605 -416
<< pdiffc >>
rect -593 -416 -559 416
rect -497 -416 -463 416
rect -401 -416 -367 416
rect -305 -416 -271 416
rect -209 -416 -175 416
rect -113 -416 -79 416
rect -17 -416 17 416
rect 79 -416 113 416
rect 175 -416 209 416
rect 271 -416 305 416
rect 367 -416 401 416
rect 463 -416 497 416
rect 559 -416 593 416
<< poly >>
rect -543 428 -513 454
rect -447 428 -417 454
rect -351 428 -321 454
rect -255 428 -225 454
rect -159 428 -129 454
rect -63 428 -33 454
rect 33 428 63 454
rect 129 428 159 454
rect 225 428 255 454
rect 321 428 351 454
rect 417 428 447 454
rect 513 428 543 454
rect -543 -454 -513 -428
rect -447 -454 -417 -428
rect -351 -454 -321 -428
rect -543 -484 -321 -454
rect -255 -454 -225 -428
rect -159 -454 -129 -428
rect -63 -454 -33 -428
rect -255 -484 -33 -454
rect 33 -454 63 -428
rect 129 -454 159 -428
rect 225 -454 255 -428
rect 33 -484 255 -454
rect 321 -454 351 -428
rect 417 -454 447 -428
rect 513 -454 543 -428
rect 321 -484 543 -454
<< locali >>
rect -593 416 -559 432
rect -593 -432 -559 -416
rect -497 416 -463 432
rect -497 -432 -463 -416
rect -401 416 -367 432
rect -401 -432 -367 -416
rect -305 416 -271 432
rect -305 -432 -271 -416
rect -209 416 -175 432
rect -209 -432 -175 -416
rect -113 416 -79 432
rect -113 -432 -79 -416
rect -17 416 17 432
rect -17 -432 17 -416
rect 79 416 113 432
rect 79 -432 113 -416
rect 175 416 209 432
rect 175 -432 209 -416
rect 271 416 305 432
rect 271 -432 305 -416
rect 367 416 401 432
rect 367 -432 401 -416
rect 463 416 497 432
rect 463 -432 497 -416
rect 559 416 593 432
rect 559 -432 593 -416
<< viali >>
rect -593 -416 -559 -62
rect -497 60 -463 416
rect -401 -416 -367 -62
rect -305 60 -271 416
rect -209 -416 -175 -62
rect -113 60 -79 416
rect -17 -416 17 -62
rect 79 60 113 416
rect 175 -416 209 -62
rect 271 60 305 416
rect 367 -416 401 -62
rect 463 60 497 416
rect 559 -416 593 -62
<< metal1 >>
rect -503 416 -457 428
rect -503 60 -497 416
rect -463 60 -457 416
rect -503 48 -457 60
rect -311 416 -265 428
rect -311 60 -305 416
rect -271 60 -265 416
rect -311 48 -265 60
rect -119 416 -73 428
rect -119 60 -113 416
rect -79 60 -73 416
rect -119 48 -73 60
rect 73 416 119 428
rect 73 60 79 416
rect 113 60 119 416
rect 73 48 119 60
rect 265 416 311 428
rect 265 60 271 416
rect 305 60 311 416
rect 265 48 311 60
rect 457 416 503 428
rect 457 60 463 416
rect 497 60 503 416
rect 457 48 503 60
rect -599 -62 -553 -50
rect -599 -416 -593 -62
rect -559 -416 -553 -62
rect -599 -428 -553 -416
rect -407 -62 -361 -50
rect -407 -416 -401 -62
rect -367 -416 -361 -62
rect -407 -428 -361 -416
rect -215 -62 -169 -50
rect -215 -416 -209 -62
rect -175 -416 -169 -62
rect -215 -428 -169 -416
rect -23 -62 23 -50
rect -23 -416 -17 -62
rect 17 -416 23 -62
rect -23 -428 23 -416
rect 169 -62 215 -50
rect 169 -416 175 -62
rect 209 -416 215 -62
rect 169 -428 215 -416
rect 361 -62 407 -50
rect 361 -416 367 -62
rect 401 -416 407 -62
rect 361 -428 407 -416
rect 553 -62 599 -50
rect 553 -416 559 -62
rect 593 -416 599 -62
rect 553 -428 599 -416
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.28 l 0.15 m 1 nf 12 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
