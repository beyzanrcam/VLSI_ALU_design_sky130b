magic
tech sky130B
magscale 1 2
timestamp 1734801607
<< error_s >>
rect 786 866 6191 867
rect 20 449 6191 866
rect 6192 449 7131 867
rect 20 448 5425 449
rect 120 322 320 380
rect 510 322 710 380
rect 1011 322 1211 380
rect 1401 322 1601 380
rect 1923 322 2123 380
rect 2313 322 2513 380
rect 2815 323 3015 381
rect 3205 323 3405 381
rect 3707 323 3907 381
rect 4097 323 4297 381
rect 4606 323 4806 381
rect 4996 323 5196 381
rect 5525 323 5725 381
rect 5915 323 6115 381
rect 6465 323 6665 381
rect 6855 323 7055 381
rect 120 234 320 292
rect 510 234 710 292
rect 1011 234 1211 292
rect 1401 234 1601 292
rect 1923 234 2123 292
rect 2313 234 2513 292
rect 2815 235 3015 293
rect 3205 235 3405 293
rect 3707 235 3907 293
rect 4097 235 4297 293
rect 4606 235 4806 293
rect 4996 235 5196 293
rect 5525 235 5725 293
rect 5915 235 6115 293
rect 6465 235 6665 293
rect 6855 235 7055 293
rect 257 209 577 233
rect 88 15 89 198
rect 116 22 117 198
rect 257 -63 281 209
rect 979 15 980 187
rect 1007 22 1008 215
rect 1148 209 1468 233
rect 2060 209 2380 233
rect 2952 210 3272 234
rect 3844 210 4164 234
rect 4743 210 5063 234
rect 5662 210 5982 234
rect 6602 210 6922 234
rect 1148 -63 1172 209
rect 2060 -63 2084 209
rect 2952 -62 2976 210
rect 3844 -62 3868 210
rect 4743 -62 4767 210
rect 5662 -62 5686 210
rect 6602 -62 6626 210
rect 257 -87 577 -63
rect 1148 -87 1468 -63
rect 2060 -87 2380 -63
rect 2952 -86 3272 -62
rect 3844 -86 4164 -62
rect 4743 -86 5063 -62
rect 5662 -86 5982 -62
rect 6602 -86 6922 -62
<< metal1 >>
rect 6 198 116 245
rect 6 15 89 198
rect 786 187 869 199
rect 1677 187 1760 199
rect 2589 187 2672 199
rect 3481 188 3564 199
rect 4373 188 4456 199
rect 5272 188 5355 199
rect 6191 188 6274 199
rect 786 113 980 187
rect 1677 113 1871 187
rect 2589 113 2783 187
rect 3481 113 3675 188
rect 4373 113 4567 188
rect 5272 113 5466 188
rect 6191 113 6385 188
rect 897 15 980 113
rect 1788 15 1871 113
rect 2700 15 2783 113
rect 3592 16 3675 113
rect 4484 16 4567 113
rect 5383 16 5466 113
rect 6302 16 6385 113
rect 7131 27 7214 199
use shifter  shifter_0
timestamp 1734801607
transform 1 0 -106 0 1 183
box 112 -270 7320 829
<< end >>
