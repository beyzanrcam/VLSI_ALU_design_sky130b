magic
tech sky130B
magscale 1 2
timestamp 1736600897
<< metal1 >>
rect 2212 -554 2310 -542
rect 2212 -628 2224 -554
rect 2298 -628 2310 -554
rect 2212 -640 2310 -628
rect 3592 -548 3690 -536
rect 3592 -622 3604 -548
rect 3678 -622 3690 -548
rect 3592 -634 3690 -622
rect 4994 -550 5092 -538
rect 4994 -624 5006 -550
rect 5080 -624 5092 -550
rect 1807 -1356 1873 -674
rect 1927 -1251 1993 -674
rect 2224 -868 2298 -640
rect 1927 -1317 2066 -1251
rect 3191 -1356 3257 -674
rect 3300 -1257 3353 -674
rect 3604 -812 3678 -634
rect 4994 -636 5092 -624
rect 6398 -548 6496 -536
rect 6398 -622 6410 -548
rect 6484 -622 6496 -548
rect 6398 -634 6496 -622
rect 7792 -552 7890 -540
rect 7792 -626 7804 -552
rect 7878 -626 7890 -552
rect 3300 -1310 3460 -1257
rect 4581 -1356 4647 -674
rect 4687 -1251 4753 -674
rect 5006 -814 5080 -636
rect 4687 -1317 4866 -1251
rect 6013 -1356 6079 -674
rect 6109 -1251 6175 -674
rect 6410 -816 6484 -634
rect 7792 -638 7890 -626
rect 9198 -550 9296 -538
rect 9198 -624 9210 -550
rect 9284 -624 9296 -550
rect 9198 -636 9296 -624
rect 10584 -554 10682 -542
rect 10584 -628 10596 -554
rect 10670 -628 10682 -554
rect 6109 -1317 6266 -1251
rect 7389 -1356 7455 -674
rect 7507 -1251 7573 -674
rect 7804 -816 7878 -638
rect 7507 -1317 7669 -1251
rect 8773 -1356 8839 -674
rect 8891 -1251 8957 -674
rect 9210 -812 9284 -636
rect 10584 -640 10682 -628
rect 11986 -566 12084 -554
rect 11986 -640 11998 -566
rect 12072 -640 12084 -566
rect 8891 -1317 9079 -1251
rect 10175 -1356 10241 -674
rect 10299 -1251 10365 -674
rect 10596 -814 10670 -640
rect 11986 -652 12084 -640
rect 10299 -1317 10477 -1251
rect 11563 -1356 11629 -674
rect 11697 -1251 11763 -674
rect 11998 -816 12072 -652
rect 11697 -1317 11866 -1251
rect 1807 -1422 2066 -1356
rect 3191 -1422 3466 -1356
rect 4581 -1422 4871 -1356
rect 6013 -1422 6277 -1356
rect 7389 -1422 7666 -1356
rect 8773 -1422 9073 -1356
rect 10175 -1422 10487 -1356
rect 11563 -1422 11893 -1356
rect 2986 -1640 3055 -1586
rect 2504 -1934 2578 -1782
rect 2488 -1950 2594 -1934
rect 2488 -2024 2504 -1950
rect 2578 -2024 2594 -1950
rect 2488 -2040 2594 -2024
rect 2986 -2245 3070 -1640
rect 4311 -1642 4363 -1530
rect 3908 -1932 3986 -1758
rect 3894 -1950 4004 -1932
rect 3894 -2028 3908 -1950
rect 3986 -2028 4004 -1950
rect 3894 -2042 4004 -2028
rect 4310 -2114 4400 -1642
rect 5306 -1900 5370 -1748
rect 5292 -1912 5384 -1900
rect 5292 -1976 5306 -1912
rect 5370 -1976 5384 -1912
rect 5292 -1992 5384 -1976
rect 5726 -1991 5795 -1586
rect 6262 -1722 6358 -1708
rect 6262 -1784 6278 -1722
rect 6340 -1784 6656 -1722
rect 6262 -1802 6358 -1784
rect 5726 -2060 6590 -1991
rect 6521 -2107 6590 -2060
rect 6905 -2087 6974 -1606
rect 7664 -1717 7744 -1704
rect 7664 -1769 7679 -1717
rect 7731 -1720 7744 -1717
rect 7731 -1766 8052 -1720
rect 7731 -1769 7744 -1766
rect 7664 -1784 7744 -1769
rect 8325 -1857 8394 -1586
rect 9116 -1602 9202 -1584
rect 9116 -1654 9134 -1602
rect 9186 -1654 9202 -1602
rect 9116 -1670 9202 -1654
rect 9142 -1722 9178 -1670
rect 9142 -1766 9448 -1722
rect 7656 -1926 8394 -1857
rect 9965 -1866 10034 -1546
rect 10546 -1732 10636 -1714
rect 10546 -1786 10564 -1732
rect 10618 -1786 10840 -1732
rect 10546 -1804 10636 -1786
rect 4310 -2196 6322 -2114
rect 6521 -2176 6780 -2107
rect 6905 -2156 7240 -2087
rect 6254 -2208 6322 -2196
rect 6711 -2208 6780 -2176
rect 7171 -2208 7240 -2156
rect 7656 -2208 7725 -1926
rect 8472 -1935 10034 -1866
rect 8472 -2067 8541 -1935
rect 11385 -1986 11454 -1566
rect 11952 -1733 12042 -1714
rect 11952 -1785 11971 -1733
rect 12023 -1736 12042 -1733
rect 12023 -1782 12240 -1736
rect 12023 -1785 12042 -1782
rect 11952 -1802 12042 -1785
rect 2986 -2314 5843 -2245
rect 6254 -2305 6323 -2208
rect 6711 -2248 6783 -2208
rect 6714 -2305 6783 -2248
rect 7171 -2260 7243 -2208
rect 7174 -2305 7243 -2260
rect 7654 -2268 7725 -2208
rect 8156 -2136 8541 -2067
rect 8634 -2055 11454 -1986
rect 7654 -2305 7723 -2268
rect 8156 -2350 8225 -2136
rect 8634 -2305 8703 -2055
rect 12705 -2146 12774 -1586
rect 9134 -2215 12774 -2146
rect 9134 -2305 9203 -2215
rect 6140 -3878 6184 -3836
rect 6620 -3878 6664 -3836
rect 7080 -3878 7124 -3836
rect 7540 -3878 7584 -3836
rect 8020 -3878 8064 -3836
rect 8520 -3878 8564 -3836
rect 9000 -3878 9044 -3836
rect 9500 -3878 9544 -3836
<< via1 >>
rect 2224 -628 2298 -554
rect 3604 -622 3678 -548
rect 5006 -624 5080 -550
rect 6410 -622 6484 -548
rect 7804 -626 7878 -552
rect 9210 -624 9284 -550
rect 10596 -628 10670 -554
rect 11998 -640 12072 -566
rect 2504 -2024 2578 -1950
rect 3908 -2028 3986 -1950
rect 5306 -1976 5370 -1912
rect 6278 -1784 6340 -1722
rect 7679 -1769 7731 -1717
rect 9134 -1654 9186 -1602
rect 10564 -1786 10618 -1732
rect 11971 -1785 12023 -1733
<< metal2 >>
rect 2212 -554 2310 -542
rect 2212 -628 2224 -554
rect 2298 -628 2310 -554
rect 2212 -640 2310 -628
rect 3592 -548 3690 -536
rect 3592 -622 3604 -548
rect 3678 -622 3690 -548
rect 3592 -634 3690 -622
rect 4994 -550 5092 -538
rect 4994 -624 5006 -550
rect 5080 -624 5092 -550
rect 4994 -636 5092 -624
rect 6398 -548 6496 -536
rect 6398 -622 6410 -548
rect 6484 -622 6496 -548
rect 6398 -634 6496 -622
rect 7792 -552 7890 -540
rect 7792 -626 7804 -552
rect 7878 -626 7890 -552
rect 7792 -638 7890 -626
rect 9198 -550 9296 -538
rect 9198 -624 9210 -550
rect 9284 -624 9296 -550
rect 9198 -636 9296 -624
rect 10584 -554 10682 -542
rect 10584 -628 10596 -554
rect 10670 -628 10682 -554
rect 10584 -640 10682 -628
rect 11986 -566 12084 -554
rect 11986 -640 11998 -566
rect 12072 -640 12084 -566
rect 11986 -652 12084 -640
rect 9116 -1598 9202 -1584
rect 9116 -1658 9130 -1598
rect 9190 -1658 9202 -1598
rect 9116 -1670 9202 -1658
rect 6262 -1722 6358 -1708
rect 6262 -1784 6278 -1722
rect 6340 -1784 6358 -1722
rect 7664 -1713 7744 -1704
rect 7664 -1773 7675 -1713
rect 7735 -1773 7744 -1713
rect 7664 -1784 7744 -1773
rect 10546 -1729 10636 -1714
rect 6262 -1802 6358 -1784
rect 10546 -1789 10561 -1729
rect 10621 -1789 10636 -1729
rect 10546 -1804 10636 -1789
rect 11952 -1729 12042 -1714
rect 11952 -1789 11967 -1729
rect 12027 -1789 12042 -1729
rect 11952 -1802 12042 -1789
rect 5292 -1912 5384 -1900
rect 2488 -1950 2594 -1934
rect 2488 -2024 2504 -1950
rect 2578 -2024 2594 -1950
rect 2488 -2040 2594 -2024
rect 3894 -1950 4004 -1932
rect 3894 -2028 3908 -1950
rect 3986 -2028 4004 -1950
rect 5292 -1976 5306 -1912
rect 5370 -1976 5384 -1912
rect 5292 -1992 5384 -1976
rect 3894 -2042 4004 -2028
<< via2 >>
rect 2224 -628 2298 -554
rect 3604 -622 3678 -548
rect 5006 -624 5080 -550
rect 6410 -622 6484 -548
rect 7804 -626 7878 -552
rect 9210 -624 9284 -550
rect 10596 -628 10670 -554
rect 11998 -640 12072 -566
rect 9130 -1602 9190 -1598
rect 9130 -1654 9134 -1602
rect 9134 -1654 9186 -1602
rect 9186 -1654 9190 -1602
rect 9130 -1658 9190 -1654
rect 6278 -1784 6340 -1722
rect 7675 -1717 7735 -1713
rect 7675 -1769 7679 -1717
rect 7679 -1769 7731 -1717
rect 7731 -1769 7735 -1717
rect 7675 -1773 7735 -1769
rect 10561 -1732 10621 -1729
rect 10561 -1786 10564 -1732
rect 10564 -1786 10618 -1732
rect 10618 -1786 10621 -1732
rect 10561 -1789 10621 -1786
rect 11967 -1733 12027 -1729
rect 11967 -1785 11971 -1733
rect 11971 -1785 12023 -1733
rect 12023 -1785 12027 -1733
rect 11967 -1789 12027 -1785
rect 2504 -2024 2578 -1950
rect 3908 -2028 3986 -1950
rect 5306 -1976 5370 -1912
<< metal3 >>
rect 2212 -549 2310 -542
rect 2212 -633 2219 -549
rect 2303 -633 2310 -549
rect 2212 -640 2310 -633
rect 3592 -543 3690 -536
rect 3592 -627 3599 -543
rect 3683 -627 3690 -543
rect 3592 -634 3690 -627
rect 4994 -545 5092 -538
rect 4994 -629 5001 -545
rect 5085 -629 5092 -545
rect 4994 -636 5092 -629
rect 6398 -543 6496 -536
rect 6398 -627 6405 -543
rect 6489 -627 6496 -543
rect 6398 -634 6496 -627
rect 7792 -547 7890 -540
rect 7792 -631 7799 -547
rect 7883 -631 7890 -547
rect 7792 -638 7890 -631
rect 9198 -545 9296 -538
rect 9198 -629 9205 -545
rect 9289 -629 9296 -545
rect 9198 -636 9296 -629
rect 10584 -549 10682 -542
rect 10584 -633 10591 -549
rect 10675 -633 10682 -549
rect 10584 -640 10682 -633
rect 11986 -561 12084 -554
rect 11986 -645 11993 -561
rect 12077 -645 12084 -561
rect 11986 -652 12084 -645
rect 9098 -1593 9220 -1564
rect 9098 -1663 9125 -1593
rect 9195 -1663 9220 -1593
rect 6254 -1717 6364 -1700
rect 6254 -1789 6273 -1717
rect 6345 -1789 6364 -1717
rect 6254 -1808 6364 -1789
rect 7650 -1708 7764 -1686
rect 9098 -1690 9220 -1663
rect 7650 -1778 7670 -1708
rect 7740 -1778 7764 -1708
rect 7650 -1800 7764 -1778
rect 10532 -1724 10654 -1700
rect 10532 -1794 10556 -1724
rect 10626 -1794 10654 -1724
rect 10532 -1816 10654 -1794
rect 11936 -1724 12058 -1700
rect 11936 -1794 11962 -1724
rect 12032 -1794 12058 -1724
rect 11936 -1816 12058 -1794
rect 5288 -1907 5386 -1894
rect 2488 -1945 2594 -1934
rect 2488 -2029 2499 -1945
rect 2583 -2029 2594 -1945
rect 2488 -2040 2594 -2029
rect 3894 -1945 4004 -1932
rect 3894 -2033 3903 -1945
rect 3991 -2033 4004 -1945
rect 5288 -1981 5301 -1907
rect 5375 -1981 5386 -1907
rect 5288 -1994 5386 -1981
rect 3894 -2042 4004 -2033
<< via3 >>
rect 2219 -554 2303 -549
rect 2219 -628 2224 -554
rect 2224 -628 2298 -554
rect 2298 -628 2303 -554
rect 2219 -633 2303 -628
rect 3599 -548 3683 -543
rect 3599 -622 3604 -548
rect 3604 -622 3678 -548
rect 3678 -622 3683 -548
rect 3599 -627 3683 -622
rect 5001 -550 5085 -545
rect 5001 -624 5006 -550
rect 5006 -624 5080 -550
rect 5080 -624 5085 -550
rect 5001 -629 5085 -624
rect 6405 -548 6489 -543
rect 6405 -622 6410 -548
rect 6410 -622 6484 -548
rect 6484 -622 6489 -548
rect 6405 -627 6489 -622
rect 7799 -552 7883 -547
rect 7799 -626 7804 -552
rect 7804 -626 7878 -552
rect 7878 -626 7883 -552
rect 7799 -631 7883 -626
rect 9205 -550 9289 -545
rect 9205 -624 9210 -550
rect 9210 -624 9284 -550
rect 9284 -624 9289 -550
rect 9205 -629 9289 -624
rect 10591 -554 10675 -549
rect 10591 -628 10596 -554
rect 10596 -628 10670 -554
rect 10670 -628 10675 -554
rect 10591 -633 10675 -628
rect 11993 -566 12077 -561
rect 11993 -640 11998 -566
rect 11998 -640 12072 -566
rect 12072 -640 12077 -566
rect 11993 -645 12077 -640
rect 9125 -1598 9195 -1593
rect 9125 -1658 9130 -1598
rect 9130 -1658 9190 -1598
rect 9190 -1658 9195 -1598
rect 9125 -1663 9195 -1658
rect 6273 -1722 6345 -1717
rect 6273 -1784 6278 -1722
rect 6278 -1784 6340 -1722
rect 6340 -1784 6345 -1722
rect 6273 -1789 6345 -1784
rect 7670 -1713 7740 -1708
rect 7670 -1773 7675 -1713
rect 7675 -1773 7735 -1713
rect 7735 -1773 7740 -1713
rect 7670 -1778 7740 -1773
rect 10556 -1729 10626 -1724
rect 10556 -1789 10561 -1729
rect 10561 -1789 10621 -1729
rect 10621 -1789 10626 -1729
rect 10556 -1794 10626 -1789
rect 11962 -1729 12032 -1724
rect 11962 -1789 11967 -1729
rect 11967 -1789 12027 -1729
rect 12027 -1789 12032 -1729
rect 11962 -1794 12032 -1789
rect 2499 -1950 2583 -1945
rect 2499 -2024 2504 -1950
rect 2504 -2024 2578 -1950
rect 2578 -2024 2583 -1950
rect 2499 -2029 2583 -2024
rect 3903 -1950 3991 -1945
rect 3903 -2028 3908 -1950
rect 3908 -2028 3986 -1950
rect 3986 -2028 3991 -1950
rect 3903 -2033 3991 -2028
rect 5301 -1912 5375 -1907
rect 5301 -1976 5306 -1912
rect 5306 -1976 5370 -1912
rect 5370 -1976 5375 -1912
rect 5301 -1981 5375 -1976
<< metal4 >>
rect 2042 -543 12300 -390
rect 2042 -549 3599 -543
rect 2042 -633 2219 -549
rect 2303 -627 3599 -549
rect 3683 -545 6405 -543
rect 3683 -627 5001 -545
rect 2303 -629 5001 -627
rect 5085 -627 6405 -545
rect 6489 -545 12300 -543
rect 6489 -547 9205 -545
rect 6489 -627 7799 -547
rect 5085 -629 7799 -627
rect 2303 -631 7799 -629
rect 7883 -629 9205 -547
rect 9289 -549 12300 -545
rect 9289 -629 10591 -549
rect 7883 -631 10591 -629
rect 2303 -633 10591 -631
rect 10675 -561 12300 -549
rect 10675 -633 11993 -561
rect 2042 -645 11993 -633
rect 12077 -645 12300 -561
rect 2042 -778 12300 -645
rect 6918 -2392 7198 -778
<< via4 >>
rect 6149 -1717 6469 -1593
rect 2381 -1945 2701 -1827
rect 2381 -2029 2499 -1945
rect 2499 -2029 2583 -1945
rect 2583 -2029 2701 -1945
rect 2381 -2147 2701 -2029
rect 3787 -1945 4107 -1829
rect 3787 -2033 3903 -1945
rect 3903 -2033 3991 -1945
rect 3991 -2033 4107 -1945
rect 3787 -2149 4107 -2033
rect 5178 -1907 5498 -1784
rect 5178 -1981 5301 -1907
rect 5301 -1981 5375 -1907
rect 5375 -1981 5498 -1907
rect 6149 -1789 6273 -1717
rect 6273 -1789 6345 -1717
rect 6345 -1789 6469 -1717
rect 6149 -1913 6469 -1789
rect 5178 -2104 5498 -1981
rect 7545 -1708 7865 -1583
rect 7545 -1778 7670 -1708
rect 7670 -1778 7740 -1708
rect 7740 -1778 7865 -1708
rect 7545 -1903 7865 -1778
rect 9000 -1593 9320 -1468
rect 9000 -1663 9125 -1593
rect 9125 -1663 9195 -1593
rect 9195 -1663 9320 -1593
rect 9000 -1788 9320 -1663
rect 10431 -1724 10751 -1599
rect 10431 -1794 10556 -1724
rect 10556 -1794 10626 -1724
rect 10626 -1794 10751 -1724
rect 10431 -1919 10751 -1794
rect 11837 -1724 12157 -1599
rect 11837 -1794 11962 -1724
rect 11962 -1794 12032 -1724
rect 12032 -1794 12157 -1724
rect 11837 -1919 12157 -1794
<< metal5 >>
rect 1940 -1468 12892 -898
rect 1940 -1583 9000 -1468
rect 1940 -1593 7545 -1583
rect 1940 -1784 6149 -1593
rect 1940 -1827 5178 -1784
rect 1940 -2147 2381 -1827
rect 2701 -1829 5178 -1827
rect 2701 -2147 3787 -1829
rect 1940 -2149 3787 -2147
rect 4107 -2104 5178 -1829
rect 5498 -1913 6149 -1784
rect 6469 -1903 7545 -1593
rect 7865 -1788 9000 -1583
rect 9320 -1599 12892 -1468
rect 9320 -1788 10431 -1599
rect 7865 -1903 10431 -1788
rect 6469 -1913 10431 -1903
rect 5498 -1919 10431 -1913
rect 10751 -1919 11837 -1599
rect 12157 -1919 12892 -1599
rect 5498 -2104 12892 -1919
rect 4107 -2149 12892 -2104
rect 1940 -3874 12892 -2149
rect 12154 -3878 12892 -3874
use NOT8  NOT8_0 ~/Desktop/vlsi_sky130b/design/mag/NOT
timestamp 1736598171
transform 1 0 5850 0 1 -3379
box -110 -501 3853 1143
use nor2  nor2_0 ~/Desktop/vlsi_sky130b/design/mag/NOR/NOR2
timestamp 1736600368
transform 1 0 11800 0 1 -1320
box 0 -480 1090 580
use nor2  nor2_1
timestamp 1736600368
transform 1 0 2000 0 1 -1320
box 0 -480 1090 580
use nor2  nor2_2
timestamp 1736600368
transform 1 0 3400 0 1 -1320
box 0 -480 1090 580
use nor2  nor2_3
timestamp 1736600368
transform 1 0 4800 0 1 -1320
box 0 -480 1090 580
use nor2  nor2_4
timestamp 1736600368
transform 1 0 6200 0 1 -1320
box 0 -480 1090 580
use nor2  nor2_5
timestamp 1736600368
transform 1 0 7600 0 1 -1320
box 0 -480 1090 580
use nor2  nor2_6
timestamp 1736600368
transform 1 0 9000 0 1 -1320
box 0 -480 1090 580
use nor2  nor2_7
timestamp 1736600368
transform 1 0 10400 0 1 -1320
box 0 -480 1090 580
<< labels >>
flabel metal1 1936 -718 1978 -690 0 FreeSans 160 0 0 0 A7
port 0 nsew
flabel metal1 3308 -714 3350 -686 0 FreeSans 160 0 0 0 A6
port 1 nsew
flabel metal1 4698 -722 4740 -694 0 FreeSans 160 0 0 0 A5
port 2 nsew
flabel metal1 6120 -718 6162 -690 0 FreeSans 160 0 0 0 A4
port 3 nsew
flabel metal1 7516 -722 7558 -694 0 FreeSans 160 0 0 0 A3
port 4 nsew
flabel metal1 8904 -722 8946 -694 0 FreeSans 160 0 0 0 A2
port 5 nsew
flabel metal1 10312 -716 10354 -688 0 FreeSans 160 0 0 0 A1
port 6 nsew
flabel metal1 11708 -718 11750 -690 0 FreeSans 160 0 0 0 A0
port 7 nsew
flabel metal1 11574 -716 11616 -688 0 FreeSans 160 0 0 0 B0
port 8 nsew
flabel metal1 10182 -716 10224 -688 0 FreeSans 160 0 0 0 B1
port 9 nsew
flabel metal1 8784 -722 8826 -694 0 FreeSans 160 0 0 0 B2
port 10 nsew
flabel metal1 7402 -722 7444 -694 0 FreeSans 160 0 0 0 B3
port 11 nsew
flabel metal1 6026 -718 6068 -690 0 FreeSans 160 0 0 0 B4
port 12 nsew
flabel metal1 4592 -722 4634 -694 0 FreeSans 160 0 0 0 B5
port 13 nsew
flabel metal1 3200 -714 3242 -686 0 FreeSans 160 0 0 0 B6
port 14 nsew
flabel metal1 1822 -718 1864 -690 0 FreeSans 160 0 0 0 B7
port 15 nsew
flabel metal1 9504 -3874 9538 -3842 0 FreeSans 160 0 0 0 S0
port 23 nsew
flabel metal1 9004 -3876 9038 -3844 0 FreeSans 160 0 0 0 S1
port 22 nsew
flabel metal1 8524 -3874 8558 -3842 0 FreeSans 160 0 0 0 S2
port 21 nsew
flabel metal1 8024 -3874 8058 -3842 0 FreeSans 160 0 0 0 S3
port 20 nsew
flabel metal1 7544 -3874 7578 -3842 0 FreeSans 160 0 0 0 S4
port 19 nsew
flabel metal1 7084 -3874 7118 -3842 0 FreeSans 160 0 0 0 S5
port 18 nsew
flabel metal1 6624 -3874 6658 -3842 0 FreeSans 160 0 0 0 S6
port 17 nsew
flabel metal1 6144 -3874 6178 -3842 0 FreeSans 160 0 0 0 S7
port 16 nsew
flabel metal4 2218 -634 2302 -548 0 FreeSans 1600 0 0 0 VDD
port 24 nsew
flabel metal5 5966 -3670 6066 -3568 0 FreeSans 1600 0 0 0 VSS
port 25 nsew
<< end >>
