magic
tech sky130B
magscale 1 2
timestamp 1733615364
<< error_p >>
rect -545 169 641 207
rect -641 -169 641 169
rect -641 -207 545 -169
<< nwell >>
rect -545 169 641 207
rect -641 -169 641 169
rect -641 -207 545 -169
<< pmos >>
rect -543 -107 -513 107
rect -447 -107 -417 107
rect -351 -107 -321 107
rect -255 -107 -225 107
rect -159 -107 -129 107
rect -63 -107 -33 107
rect 33 -107 63 107
rect 129 -107 159 107
rect 225 -107 255 107
rect 321 -107 351 107
rect 417 -107 447 107
rect 513 -107 543 107
<< pdiff >>
rect -605 95 -543 107
rect -605 -95 -593 95
rect -559 -95 -543 95
rect -605 -107 -543 -95
rect -513 95 -447 107
rect -513 -95 -497 95
rect -463 -95 -447 95
rect -513 -107 -447 -95
rect -417 95 -351 107
rect -417 -95 -401 95
rect -367 -95 -351 95
rect -417 -107 -351 -95
rect -321 95 -255 107
rect -321 -95 -305 95
rect -271 -95 -255 95
rect -321 -107 -255 -95
rect -225 95 -159 107
rect -225 -95 -209 95
rect -175 -95 -159 95
rect -225 -107 -159 -95
rect -129 95 -63 107
rect -129 -95 -113 95
rect -79 -95 -63 95
rect -129 -107 -63 -95
rect -33 95 33 107
rect -33 -95 -17 95
rect 17 -95 33 95
rect -33 -107 33 -95
rect 63 95 129 107
rect 63 -95 79 95
rect 113 -95 129 95
rect 63 -107 129 -95
rect 159 95 225 107
rect 159 -95 175 95
rect 209 -95 225 95
rect 159 -107 225 -95
rect 255 95 321 107
rect 255 -95 271 95
rect 305 -95 321 95
rect 255 -107 321 -95
rect 351 95 417 107
rect 351 -95 367 95
rect 401 -95 417 95
rect 351 -107 417 -95
rect 447 95 513 107
rect 447 -95 463 95
rect 497 -95 513 95
rect 447 -107 513 -95
rect 543 95 605 107
rect 543 -95 559 95
rect 593 -95 605 95
rect 543 -107 605 -95
<< pdiffc >>
rect -593 -95 -559 95
rect -497 -95 -463 95
rect -401 -95 -367 95
rect -305 -95 -271 95
rect -209 -95 -175 95
rect -113 -95 -79 95
rect -17 -95 17 95
rect 79 -95 113 95
rect 175 -95 209 95
rect 271 -95 305 95
rect 367 -95 401 95
rect 463 -95 497 95
rect 559 -95 593 95
<< poly >>
rect -465 188 -399 204
rect -465 154 -449 188
rect -415 154 -399 188
rect -465 138 -399 154
rect -273 188 -207 204
rect -273 154 -257 188
rect -223 154 -207 188
rect -273 138 -207 154
rect -81 188 -15 204
rect -81 154 -65 188
rect -31 154 -15 188
rect -81 138 -15 154
rect 111 188 177 204
rect 111 154 127 188
rect 161 154 177 188
rect 111 138 177 154
rect 303 188 369 204
rect 303 154 319 188
rect 353 154 369 188
rect 303 138 369 154
rect 495 188 561 204
rect 495 154 511 188
rect 545 154 561 188
rect 495 138 561 154
rect -543 107 -513 133
rect -447 107 -417 138
rect -351 107 -321 133
rect -255 107 -225 138
rect -159 107 -129 133
rect -63 107 -33 138
rect 33 107 63 133
rect 129 107 159 138
rect 225 107 255 133
rect 321 107 351 138
rect 417 107 447 133
rect 513 107 543 138
rect -543 -138 -513 -107
rect -447 -133 -417 -107
rect -351 -138 -321 -107
rect -255 -133 -225 -107
rect -159 -138 -129 -107
rect -63 -133 -33 -107
rect 33 -138 63 -107
rect 129 -133 159 -107
rect 225 -138 255 -107
rect 321 -133 351 -107
rect 417 -138 447 -107
rect 513 -133 543 -107
rect -561 -154 -495 -138
rect -561 -188 -545 -154
rect -511 -188 -495 -154
rect -561 -204 -495 -188
rect -369 -154 -303 -138
rect -369 -188 -353 -154
rect -319 -188 -303 -154
rect -369 -204 -303 -188
rect -177 -154 -111 -138
rect -177 -188 -161 -154
rect -127 -188 -111 -154
rect -177 -204 -111 -188
rect 15 -154 81 -138
rect 15 -188 31 -154
rect 65 -188 81 -154
rect 15 -204 81 -188
rect 207 -154 273 -138
rect 207 -188 223 -154
rect 257 -188 273 -154
rect 207 -204 273 -188
rect 399 -154 465 -138
rect 399 -188 415 -154
rect 449 -188 465 -154
rect 399 -204 465 -188
<< polycont >>
rect -449 154 -415 188
rect -257 154 -223 188
rect -65 154 -31 188
rect 127 154 161 188
rect 319 154 353 188
rect 511 154 545 188
rect -545 -188 -511 -154
rect -353 -188 -319 -154
rect -161 -188 -127 -154
rect 31 -188 65 -154
rect 223 -188 257 -154
rect 415 -188 449 -154
<< locali >>
rect -465 154 -449 188
rect -415 154 -399 188
rect -273 154 -257 188
rect -223 154 -207 188
rect -81 154 -65 188
rect -31 154 -15 188
rect 111 154 127 188
rect 161 154 177 188
rect 303 154 319 188
rect 353 154 369 188
rect 495 154 511 188
rect 545 154 561 188
rect -593 95 -559 111
rect -593 -111 -559 -95
rect -497 95 -463 111
rect -497 -111 -463 -95
rect -401 95 -367 111
rect -401 -111 -367 -95
rect -305 95 -271 111
rect -305 -111 -271 -95
rect -209 95 -175 111
rect -209 -111 -175 -95
rect -113 95 -79 111
rect -113 -111 -79 -95
rect -17 95 17 111
rect -17 -111 17 -95
rect 79 95 113 111
rect 79 -111 113 -95
rect 175 95 209 111
rect 175 -111 209 -95
rect 271 95 305 111
rect 271 -111 305 -95
rect 367 95 401 111
rect 367 -111 401 -95
rect 463 95 497 111
rect 463 -111 497 -95
rect 559 95 593 111
rect 559 -111 593 -95
rect -561 -188 -545 -154
rect -511 -188 -495 -154
rect -369 -188 -353 -154
rect -319 -188 -303 -154
rect -177 -188 -161 -154
rect -127 -188 -111 -154
rect 15 -188 31 -154
rect 65 -188 81 -154
rect 207 -188 223 -154
rect 257 -188 273 -154
rect 399 -188 415 -154
rect 449 -188 465 -154
<< viali >>
rect -449 154 -415 188
rect -257 154 -223 188
rect -65 154 -31 188
rect 127 154 161 188
rect 319 154 353 188
rect 511 154 545 188
rect -593 -95 -559 95
rect -497 -95 -463 95
rect -401 -95 -367 95
rect -305 -95 -271 95
rect -209 -95 -175 95
rect -113 -95 -79 95
rect -17 -95 17 95
rect 79 -95 113 95
rect 175 -95 209 95
rect 271 -95 305 95
rect 367 -95 401 95
rect 463 -95 497 95
rect 559 -95 593 95
rect -545 -188 -511 -154
rect -353 -188 -319 -154
rect -161 -188 -127 -154
rect 31 -188 65 -154
rect 223 -188 257 -154
rect 415 -188 449 -154
<< metal1 >>
rect -461 188 -403 194
rect -461 154 -449 188
rect -415 154 -403 188
rect -461 148 -403 154
rect -269 188 -211 194
rect -269 154 -257 188
rect -223 154 -211 188
rect -269 148 -211 154
rect -77 188 -19 194
rect -77 154 -65 188
rect -31 154 -19 188
rect -77 148 -19 154
rect 115 188 173 194
rect 115 154 127 188
rect 161 154 173 188
rect 115 148 173 154
rect 307 188 365 194
rect 307 154 319 188
rect 353 154 365 188
rect 307 148 365 154
rect 499 188 557 194
rect 499 154 511 188
rect 545 154 557 188
rect 499 148 557 154
rect -599 95 -553 107
rect -599 -95 -593 95
rect -559 -95 -553 95
rect -599 -107 -553 -95
rect -503 95 -457 107
rect -503 -95 -497 95
rect -463 -95 -457 95
rect -503 -107 -457 -95
rect -407 95 -361 107
rect -407 -95 -401 95
rect -367 -95 -361 95
rect -407 -107 -361 -95
rect -311 95 -265 107
rect -311 -95 -305 95
rect -271 -95 -265 95
rect -311 -107 -265 -95
rect -215 95 -169 107
rect -215 -95 -209 95
rect -175 -95 -169 95
rect -215 -107 -169 -95
rect -119 95 -73 107
rect -119 -95 -113 95
rect -79 -95 -73 95
rect -119 -107 -73 -95
rect -23 95 23 107
rect -23 -95 -17 95
rect 17 -95 23 95
rect -23 -107 23 -95
rect 73 95 119 107
rect 73 -95 79 95
rect 113 -95 119 95
rect 73 -107 119 -95
rect 169 95 215 107
rect 169 -95 175 95
rect 209 -95 215 95
rect 169 -107 215 -95
rect 265 95 311 107
rect 265 -95 271 95
rect 305 -95 311 95
rect 265 -107 311 -95
rect 361 95 407 107
rect 361 -95 367 95
rect 401 -95 407 95
rect 361 -107 407 -95
rect 457 95 503 107
rect 457 -95 463 95
rect 497 -95 503 95
rect 457 -107 503 -95
rect 553 95 599 107
rect 553 -95 559 95
rect 593 -95 599 95
rect 553 -107 599 -95
rect -557 -154 -499 -148
rect -557 -188 -545 -154
rect -511 -188 -499 -154
rect -557 -194 -499 -188
rect -365 -154 -307 -148
rect -365 -188 -353 -154
rect -319 -188 -307 -154
rect -365 -194 -307 -188
rect -173 -154 -115 -148
rect -173 -188 -161 -154
rect -127 -188 -115 -154
rect -173 -194 -115 -188
rect 19 -154 77 -148
rect 19 -188 31 -154
rect 65 -188 77 -154
rect 19 -194 77 -188
rect 211 -154 269 -148
rect 211 -188 223 -154
rect 257 -188 269 -154
rect 211 -194 269 -188
rect 403 -154 461 -148
rect 403 -188 415 -154
rect 449 -188 461 -154
rect 403 -194 461 -188
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.07 l 0.15 m 1 nf 12 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 1 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
