* NGSPICE file created from ALU.ext - technology: sky130B

.subckt sky130_fd_pr__pfet_01v8_64A2S3 a_n33_n428# a_447_n428# a_n605_n428# a_321_n484#
+ a_n543_n484# a_543_n428# a_159_n428# a_33_n484# a_n255_n484# a_255_n428# w_n641_n484#
+ a_351_n428# a_n417_n428# a_n513_n428# a_n129_n428# a_63_n428# a_n225_n428# a_n321_n428#
X0 a_447_n428# a_321_n484# a_351_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X1 a_n513_n428# a_n543_n484# a_n605_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=1.3268 ps=9.18 w=4.28 l=0.15
X2 a_63_n428# a_33_n484# a_n33_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X3 a_n129_n428# a_n255_n484# a_n225_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X4 a_n417_n428# a_n543_n484# a_n513_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X5 a_n33_n428# a_n255_n484# a_n129_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X6 a_351_n428# a_321_n484# a_255_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X7 a_255_n428# a_33_n484# a_159_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X8 a_n321_n428# a_n543_n484# a_n417_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X9 a_543_n428# a_321_n484# a_447_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=1.3268 pd=9.18 as=0.7062 ps=4.61 w=4.28 l=0.15
X10 a_159_n428# a_33_n484# a_63_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X11 a_n225_n428# a_n255_n484# a_n321_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_S9NJ5Q a_159_n100# a_n159_n126# a_33_n126# a_n129_n100#
+ a_n221_n100# a_63_n100# a_n63_n126# a_n33_n100# a_129_n126# VSUBS
X0 a_n129_n100# a_n159_n126# a_n221_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1 a_63_n100# a_33_n126# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2 a_n33_n100# a_n63_n126# a_n129_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_159_n100# a_129_n126# a_63_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt nor4 A B C D VSS Y VDD
Xsky130_fd_pr__pfet_01v8_64A2S3_0 m1_n20_1047# m1_268_1523# VDD D A Y m1_n20_1047#
+ C B m1_268_1523# VDD Y VDD m1_n308_1523# m1_n308_1523# m1_268_1523# m1_n20_1047#
+ m1_n308_1523# sky130_fd_pr__pfet_01v8_64A2S3
Xsky130_fd_pr__nfet_01v8_S9NJ5Q_0 VSS A C Y VSS Y B VSS D VSS sky130_fd_pr__nfet_01v8_S9NJ5Q
.ends

.subckt sky130_fd_pr__nfet_01v8_6H9P4D a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt efepmos_W107-L15-F3 a_n129_n204# a_n173_n107# w_n209_n207# a_n81_n107#
X0 a_n81_n107# a_n129_n204# a_n173_n107# w_n209_n207# sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1 a_n81_n107# a_n129_n204# a_n173_n107# w_n209_n207# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2 a_n173_n107# a_n129_n204# a_n81_n107# w_n209_n207# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
.ends

.subckt inv A VSS Y VDD
Xsky130_fd_pr__nfet_01v8_6H9P4D_0 Y VSS A VSS sky130_fd_pr__nfet_01v8_6H9P4D
Xefepmos_W107-L15-F3_0 A VDD VDD Y efepmos_W107-L15-F3
.ends

.subckt nmos_2shared_W200-L015-F1 a_63_n200# a_n63_n226# a_n33_n200# a_33_n226# a_n125_n200#
+ VSUBS
X0 a_n33_n200# a_n63_n226# a_n125_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1 a_63_n200# a_33_n226# a_n33_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
.ends

.subckt pmos_p2-w321-L015-f3 a_n317_n107# w_n353_n143# a_n225_n107# a_33_n138# a_n255_n138#
X0 a_n225_n107# a_33_n138# a_n317_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1 a_n225_n107# a_n255_n138# a_n317_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2 a_n317_n107# a_33_n138# a_n225_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3 a_n317_n107# a_n255_n138# a_n225_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4 a_n225_n107# a_n255_n138# a_n317_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X5 a_n317_n107# a_33_n138# a_n225_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
.ends

.subckt NAND2 A B VSS VDD Y
Xnmos_2shared_W200-L015-F1_0 VSS B a_994_146# A Y VSS nmos_2shared_W200-L015-F1
Xpmos_p2-w321-L015-f3_0 VDD VDD Y B A pmos_p2-w321-L015-f3
.ends

.subckt ZFLAG A0 A1 A2 A3 A4 A5 A6 A7 Z VDD VSS
Xnor4_0 A3 A2 A1 A0 VSS nor4_0/Y VDD nor4
Xnor4_1 A4 A5 A6 A7 VSS nor4_1/Y VDD nor4
Xinv_0 inv_0/A VSS Z VDD inv
XNAND2_0 nor4_0/Y nor4_1/Y VSS VDD inv_0/A NAND2
.ends

.subckt buffer VDD Y A VSS
Xinv_0 A VSS inv_1/A VDD inv
Xinv_1 inv_1/A VSS Y VDD inv
.ends

.subckt left_shifter A0 A1 A2 A3 A4 A5 A6 A7 S0 S1 S2 S3 S4 S5 S6 S7 C VDD VSS
Xbuffer_0 VDD S3 A2 VSS buffer
Xbuffer_1 VDD C A7 VSS buffer
Xbuffer_2 VDD S7 A6 VSS buffer
Xbuffer_3 VDD S6 A5 VSS buffer
Xbuffer_4 VDD S5 A4 VSS buffer
Xinv_0 VDD VSS S0 VDD inv
Xbuffer_5 VDD S4 A3 VSS buffer
Xbuffer_6 VDD S1 A0 VSS buffer
Xbuffer_7 VDD S2 A1 VSS buffer
.ends

.subckt right_shifter A0 A1 A2 A3 A4 A5 A6 A7 C S0 S1 S2 S3 S4 S5 S6 S7 VDD VSS
Xbuffer_0 VDD S1 A2 VSS buffer
Xbuffer_1 VDD S6 A7 VSS buffer
Xbuffer_2 VDD S5 A6 VSS buffer
Xbuffer_3 VDD S4 A5 VSS buffer
Xbuffer_4 VDD S3 A4 VSS buffer
Xinv_0 VDD VSS S7 VDD inv
Xbuffer_5 VDD S2 A3 VSS buffer
Xbuffer_6 VDD C A0 VSS buffer
Xbuffer_7 VDD S0 A1 VSS buffer
.ends

.subckt XOR2 A B VSS VDD Y a_99_341#
X0 VDD A a_129_987# VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1 a_129_987# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2 a_129_987# a_n51_367# Y VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3 Y a_99_341# a_129_987# VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X4 Y a_n51_367# a_129_987# VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X5 Y a_n51_367# a_129_987# VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X6 a_129_987# a_99_341# Y VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X7 a_129_987# a_99_341# Y VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X8 VDD B a_129_987# VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X9 a_129_367# a_99_341# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X10 a_99_341# B VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X11 a_129_987# B VDD VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X12 VDD B a_129_987# VDD sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X13 VSS A a_n51_367# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X14 a_129_987# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X15 a_99_341# B VDD VDD sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X16 VDD A a_n51_367# VDD sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X17 VSS a_99_341# a_129_367# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X18 a_129_367# a_99_341# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X19 a_129_367# a_n51_367# Y VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X20 Y A a_705_367# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X21 Y a_n51_367# a_129_367# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X22 Y a_n51_367# a_129_367# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X23 a_705_367# A Y VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X24 a_705_367# A Y VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X25 VSS B a_705_367# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X26 a_705_367# B VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X27 VSS B a_705_367# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt V_FLAG A_MSB B_MSB OPCODE3 Y_MSB V VDD VSS
Xinv_0 inv_0/A VSS V VDD inv
XNAND2_0 XOR2_0/Y XOR2_2/Y VSS VDD inv_0/A NAND2
XXOR2_0 A_MSB Y_MSB VSS VDD XOR2_0/Y XOR2_0/a_99_341# XOR2
XXOR2_1 A_MSB B_MSB VSS VDD XOR2_2/B XOR2_1/a_99_341# XOR2
XXOR2_2 OPCODE3 XOR2_2/B VSS VDD XOR2_2/Y XOR2_2/a_99_341# XOR2
.ends

.subckt FULL_ADDER_XORED A K COUT CIN B VDD VSS OUT
XNAND2_0 XOR2_2/Y A VSS VDD NAND2_2/B NAND2
XNAND2_1 XOR2_1/A CIN VSS VDD NAND2_2/A NAND2
XNAND2_2 NAND2_2/A NAND2_2/B VSS VDD COUT NAND2
XXOR2_0 XOR2_2/Y A VSS VDD XOR2_1/A li_1358_495# XOR2
XXOR2_1 XOR2_1/A CIN VSS VDD OUT XOR2_1/a_99_341# XOR2
XXOR2_2 B K VSS VDD XOR2_2/Y XOR2_2/a_99_341# XOR2
.ends

.subckt x8bit_ADDER K B0 B1 B2 B3 B5 B6 B7 A0 A1 A2 A3 A4 A5 A6 A7 S0 S1 S2 S3 S4
+ S5 S6 S7 C B4 VDD VSS
XFULL_ADDER_XORED_0 A7 K C FULL_ADDER_XORED_0/CIN B7 VDD VSS S7 FULL_ADDER_XORED
XFULL_ADDER_XORED_1 A6 K FULL_ADDER_XORED_0/CIN FULL_ADDER_XORED_1/CIN B6 VDD VSS
+ S6 FULL_ADDER_XORED
XFULL_ADDER_XORED_2 A5 K FULL_ADDER_XORED_1/CIN FULL_ADDER_XORED_2/CIN B5 VDD VSS
+ S5 FULL_ADDER_XORED
XFULL_ADDER_XORED_3 A4 K FULL_ADDER_XORED_2/CIN FULL_ADDER_XORED_3/CIN B4 VDD VSS
+ S4 FULL_ADDER_XORED
XFULL_ADDER_XORED_4 A3 K FULL_ADDER_XORED_3/CIN FULL_ADDER_XORED_4/CIN B3 VDD VSS
+ S3 FULL_ADDER_XORED
XFULL_ADDER_XORED_5 A2 K FULL_ADDER_XORED_4/CIN FULL_ADDER_XORED_5/CIN B2 VDD VSS
+ S2 FULL_ADDER_XORED
XFULL_ADDER_XORED_6 A1 K FULL_ADDER_XORED_5/CIN FULL_ADDER_XORED_6/CIN B1 VDD VSS
+ S1 FULL_ADDER_XORED
XFULL_ADDER_XORED_7 A0 K FULL_ADDER_XORED_6/CIN K B0 VDD VSS S0 FULL_ADDER_XORED
.ends

.subckt NOT8 A7 A6 A5 A4 A3 A2 A1 A0 S0 S1 S2 S3 S4 S5 S6 S7 VDD VSS
Xinv_0 A3 VSS S3 VDD inv
Xinv_1 A7 VSS S7 VDD inv
Xinv_2 A6 VSS S6 VDD inv
Xinv_3 A5 VSS S5 VDD inv
Xinv_4 A4 VSS S4 VDD inv
Xinv_5 A2 VSS S2 VDD inv
Xinv_6 A1 VSS S1 VDD inv
Xinv_7 A0 VSS S0 VDD inv
.ends

.subckt NAND8 A0 B0 A1 B1 A2 B2 A3 B3 A4 B4 A5 B5 A6 B6 A7 B7 P0 P1 P2 P3 P4 P5 P6
+ P7 NAND2_9/VDD VSUBS
XNAND2_7 B6 A6 VSUBS NAND2_9/VDD P6 NAND2
XNAND2_8 B1 A1 VSUBS NAND2_9/VDD P1 NAND2
XNAND2_9 B2 A2 VSUBS NAND2_9/VDD P2 NAND2
XNAND2_0 B7 A7 VSUBS NAND2_9/VDD P7 NAND2
XNAND2_1 B4 A4 VSUBS NAND2_9/VDD P4 NAND2
XNAND2_2 B3 A3 VSUBS NAND2_9/VDD P3 NAND2
XNAND2_4 B0 A0 VSUBS NAND2_9/VDD P0 NAND2
XNAND2_6 B5 A5 VSUBS NAND2_9/VDD P5 NAND2
.ends

.subckt AND8 A7 B7 A6 B6 A5 B5 A4 B4 A3 B3 A2 B2 A1 B1 A0 B0 S0 S1 S2 S3 S4 S5 S6
+ S7 NAND8_0/NAND2_9/VDD NOT8_0/VDD VSUBS
XNOT8_0 NOT8_0/A7 NOT8_0/A6 NOT8_0/A5 NOT8_0/A4 NOT8_0/A3 NOT8_0/A2 NOT8_0/A1 NOT8_0/A0
+ S0 S1 S2 S3 S4 S5 S6 S7 NOT8_0/VDD VSUBS NOT8
XNAND8_0 A7 B7 A6 B6 A5 B5 A4 B4 A3 B3 A2 B2 A1 B1 A0 B0 NOT8_0/A7 NOT8_0/A6 NOT8_0/A5
+ NOT8_0/A4 NOT8_0/A3 NOT8_0/A2 NOT8_0/A1 NOT8_0/A0 NAND8_0/NAND2_9/VDD VSUBS NAND8
.ends

.subckt pmos4_f2 a_n177_n258# a_n413_n161# a_207_n258# w_n449_n261# a_n369_n258# a_n321_n161#
+ a_15_n258#
X0 a_n321_n161# a_207_n258# a_n413_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1 a_n321_n161# a_n369_n258# a_n413_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2 a_n413_n161# a_15_n258# a_n321_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3 a_n413_n161# a_n369_n258# a_n321_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4 a_n321_n161# a_15_n258# a_n413_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X5 a_n321_n161# a_n177_n258# a_n413_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X6 a_n413_n161# a_n177_n258# a_n321_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X7 a_n413_n161# a_207_n258# a_n321_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
.ends

.subckt efenmos2 a_n159_n426# a_33_n426# a_n221_n400# a_n63_n426# a_129_n426# a_159_n400#
+ VSUBS
X0 a_63_n400# a_33_n426# a_n33_n400# VSUBS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1 a_n129_n400# a_n159_n426# a_n221_n400# VSUBS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2 a_n33_n400# a_n63_n426# a_n129_n400# VSUBS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3 a_159_n400# a_129_n426# a_63_n400# VSUBS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
.ends

.subckt NAND4F A B C D VSS VDD Y
Xpmos4_f2_0 C VDD A VDD D Y B pmos4_f2
Xefenmos2_1 D B VSS C A Y VSS efenmos2
.ends

.subckt sky130_fd_pr__pfet_01v8_UFBY79 a_n33_n128# a_n509_n128# a_447_n128# a_159_n128#
+ a_255_n128# a_351_n128# a_n417_n128# a_n447_n225# a_n129_n128# a_63_n128# a_n225_n128#
+ a_33_n225# w_n545_n228# a_n321_n128#
X0 a_63_n128# a_33_n225# a_n33_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1 a_n129_n128# a_n447_n225# a_n225_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2 a_n417_n128# a_n447_n225# a_n509_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X3 a_351_n128# a_33_n225# a_255_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X4 a_n33_n128# a_n447_n225# a_n129_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X5 a_255_n128# a_33_n225# a_159_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X6 a_n321_n128# a_n447_n225# a_n417_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X7 a_159_n128# a_33_n225# a_63_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X8 a_n225_n128# a_n447_n225# a_n321_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X9 a_447_n128# a_33_n225# a_351_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_LZEQWH a_33_n126# a_n125_n100# a_63_n100# a_n63_n126#
+ a_n33_n100# VSUBS
X0 a_63_n100# a_33_n126# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X1 a_n33_n100# a_n63_n126# a_n125_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
.ends

.subckt nor2 A B VSS VDD Y
Xsky130_fd_pr__pfet_01v8_UFBY79_0 m1_760_245# VDD Y m1_760_245# Y m1_760_245# m1_760_245#
+ A VDD Y m1_760_245# B VDD VDD sky130_fd_pr__pfet_01v8_UFBY79
Xsky130_fd_pr__nfet_01v8_LZEQWH_0 A VSS VSS B Y VSS sky130_fd_pr__nfet_01v8_LZEQWH
.ends

.subckt mux8 A0 A1 A2 A5 A6 A7 SEL0 A3 SEL1 Y VDD A4 VSS SEL2
XNAND4F_3 A0 inv_2/Y inv_1/Y inv_3/Y VSS VDD NAND4F_8/C NAND4F
XNAND4F_4 A2 inv_2/Y SEL1 inv_3/Y VSS VDD NAND4F_8/A NAND4F
XNAND4F_5 A6 inv_2/Y SEL1 SEL2 VSS VDD NAND4F_9/A NAND4F
XNAND4F_6 A7 SEL0 SEL1 SEL2 VSS VDD NAND4F_9/B NAND4F
XNAND4F_8 NAND4F_8/A NAND4F_8/B NAND4F_8/C NAND4F_8/D VSS VDD nor2_0/A NAND4F
XNAND4F_7 A5 SEL0 inv_1/Y SEL2 VSS VDD NAND4F_9/D NAND4F
XNAND4F_9 NAND4F_9/A NAND4F_9/B NAND4F_9/C NAND4F_9/D VSS VDD nor2_0/B NAND4F
Xnor2_0 nor2_0/A nor2_0/B VSS VDD inv_0/A nor2
Xinv_0 inv_0/A VSS Y VDD inv
Xinv_1 SEL1 VSS inv_1/Y VDD inv
Xinv_2 SEL0 VSS inv_2/Y VDD inv
Xinv_3 SEL2 VSS inv_3/Y VDD inv
XNAND4F_0 A1 SEL0 inv_1/Y inv_3/Y VSS VDD NAND4F_8/D NAND4F
XNAND4F_1 A4 inv_2/Y inv_1/Y SEL2 VSS VDD NAND4F_9/C NAND4F
XNAND4F_2 A3 SEL0 SEL1 inv_3/Y VSS VDD NAND4F_8/B NAND4F
.ends

.subckt XOR8 B7 A7 A6 A5 A4 A3 A2 A1 A0 B0 B1 B2 B3 B4 B5 B6 S7 S6 S5 S4 S3 S2 S1
+ S0 XOR2_7/VDD VSUBS
XXOR2_3 A5 B5 VSUBS XOR2_7/VDD S5 XOR2_3/a_99_341# XOR2
XXOR2_4 A4 B4 VSUBS XOR2_7/VDD S4 XOR2_4/a_99_341# XOR2
XXOR2_5 A3 B3 VSUBS XOR2_7/VDD S3 XOR2_5/a_99_341# XOR2
XXOR2_6 A2 B2 VSUBS XOR2_7/VDD S2 XOR2_6/a_99_341# XOR2
XXOR2_7 A1 B1 VSUBS XOR2_7/VDD S1 XOR2_7/a_99_341# XOR2
XXOR2_0 A0 B0 VSUBS XOR2_7/VDD S0 XOR2_0/a_99_341# XOR2
XXOR2_1 A7 B7 VSUBS XOR2_7/VDD S7 XOR2_1/a_99_341# XOR2
XXOR2_2 A6 B6 VSUBS XOR2_7/VDD S6 XOR2_2/a_99_341# XOR2
.ends

.subckt OR8 A7 A6 A5 A4 A3 A2 A1 A0 B0 B1 B2 B3 B4 B5 B6 B7 S7 S6 S5 S4 S3 S2 S1 S0
+ VDD VSS
Xnor2_0 A0 B0 VSS VDD nor2_0/Y nor2
Xnor2_1 A7 B7 VSS VDD nor2_1/Y nor2
Xnor2_2 A6 B6 VSS VDD nor2_2/Y nor2
Xnor2_3 A5 B5 VSS VDD nor2_3/Y nor2
Xnor2_4 A4 B4 VSS VDD nor2_4/Y nor2
Xnor2_5 A3 B3 VSS VDD nor2_5/Y nor2
Xnor2_6 A2 B2 VSS VDD nor2_6/Y nor2
Xnor2_7 A1 B1 VSS VDD nor2_7/Y nor2
XNOT8_0 nor2_1/Y nor2_2/Y nor2_3/Y nor2_4/Y nor2_5/Y nor2_6/Y nor2_7/Y nor2_0/Y S0
+ S1 S2 S3 S4 S5 S6 S7 VDD VSS NOT8
.ends

.subckt FULL_ADDER COUT A B CIN VDD VSS OUT
XNAND2_0 B A VSS VDD NAND2_2/B NAND2
XNAND2_1 XOR2_1/A CIN VSS VDD NAND2_2/A NAND2
XNAND2_2 NAND2_2/A NAND2_2/B VSS VDD COUT NAND2
XXOR2_0 B A VSS VDD XOR2_1/A li_1358_495# XOR2
XXOR2_1 XOR2_1/A CIN VSS VDD OUT XOR2_1/a_99_341# XOR2
.ends

.subckt x4bit_ADDER A2 A1 A0 B0 B1 B2 S0 S1 S2 S3 C Cout A3 B3 VDD VSS
XFULL_ADDER_0 Cout A3 B3 FULL_ADDER_0/CIN VDD VSS S3 FULL_ADDER
XFULL_ADDER_1 FULL_ADDER_0/CIN A2 B2 FULL_ADDER_1/CIN VDD VSS S2 FULL_ADDER
XFULL_ADDER_2 FULL_ADDER_1/CIN A1 B1 FULL_ADDER_2/CIN VDD VSS S1 FULL_ADDER
XFULL_ADDER_3 FULL_ADDER_2/CIN A0 B0 C VDD VSS S0 FULL_ADDER
.ends

.subckt MULT A0 B2 B0 B3 A2 A1 SO S1 S2 S5 S4 S3 S7 S6 VDD B1 A3 VSS
XNAND2_13 B2 A3 VSS VDD inv_13/A NAND2
XNAND2_7 B2 A1 VSS VDD inv_7/A NAND2
XNAND2_8 A0 B3 VSS VDD inv_8/A NAND2
XNAND2_14 A2 B3 VSS VDD inv_14/A NAND2
XNAND2_15 B3 A3 VSS VDD inv_15/A NAND2
XNAND2_9 B3 A1 VSS VDD inv_9/A NAND2
Xinv_10 inv_10/A VSS inv_10/Y VDD inv
Xinv_11 inv_11/A VSS inv_11/Y VDD inv
Xinv_12 inv_12/A VSS inv_12/Y VDD inv
Xinv_13 inv_13/A VSS inv_13/Y VDD inv
Xinv_14 inv_14/A VSS inv_14/Y VDD inv
Xinv_15 inv_15/A VSS inv_15/Y VDD inv
Xinv_0 inv_0/A VSS inv_0/Y VDD inv
Xinv_1 inv_1/A VSS inv_1/Y VDD inv
X4bit_ADDER_0 inv_10/Y inv_4/Y inv_5/Y inv_2/Y inv_1/Y inv_0/Y S1 4bit_ADDER_1/B0
+ 4bit_ADDER_1/B1 4bit_ADDER_1/B2 VSS 4bit_ADDER_1/B3 inv_11/Y VSS VDD VSS x4bit_ADDER
Xinv_2 inv_2/A VSS inv_2/Y VDD inv
X4bit_ADDER_1 inv_12/Y inv_7/Y inv_6/Y 4bit_ADDER_1/B0 4bit_ADDER_1/B1 4bit_ADDER_1/B2
+ S2 4bit_ADDER_2/B0 4bit_ADDER_2/B1 4bit_ADDER_2/B2 VSS 4bit_ADDER_2/B3 inv_13/Y
+ 4bit_ADDER_1/B3 VDD VSS x4bit_ADDER
Xinv_3 inv_3/A VSS SO VDD inv
X4bit_ADDER_2 inv_14/Y inv_9/Y inv_8/Y 4bit_ADDER_2/B0 4bit_ADDER_2/B1 4bit_ADDER_2/B2
+ S3 S4 S5 S6 VSS S7 inv_15/Y 4bit_ADDER_2/B3 VDD VSS x4bit_ADDER
Xinv_4 inv_4/A VSS inv_4/Y VDD inv
Xinv_5 inv_5/A VSS inv_5/Y VDD inv
Xinv_7 inv_7/A VSS inv_7/Y VDD inv
Xinv_6 inv_6/A VSS inv_6/Y VDD inv
XNAND2_1 B0 A2 VSS VDD inv_1/A NAND2
XNAND2_0 B0 A3 VSS VDD inv_0/A NAND2
Xinv_8 inv_8/A VSS inv_8/Y VDD inv
XNAND2_2 B0 A1 VSS VDD inv_2/A NAND2
Xinv_9 inv_9/A VSS inv_9/Y VDD inv
XNAND2_3 B0 A0 VSS VDD inv_3/A NAND2
XNAND2_10 A2 B1 VSS VDD inv_10/A NAND2
XNAND2_4 A0 B1 VSS VDD inv_5/A NAND2
XNAND2_11 B1 A3 VSS VDD inv_11/A NAND2
XNAND2_5 B1 A1 VSS VDD inv_4/A NAND2
XNAND2_12 A2 B2 VSS VDD inv_12/A NAND2
XNAND2_6 A0 B2 VSS VDD inv_6/A NAND2
.ends

.subckt ALU B0 B1 B2 B3 B4 B5 B6 A0 A1 A2 A3 A4 A5 A6 A7 Y0 Y1 Y2 Y3 Y4 Y5 Y6 S Z
+ C V VSS Y7 B7 SEL0 SEL1 SEL2 SEL3 VDD
XZFLAG_0 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 Z VDD VSS ZFLAG
Xleft_shifter_0 B0 B1 B2 B3 B4 B5 B6 B7 mux8_1/A6 mux8_2/A6 mux8_3/A6 mux8_4/A6 mux8_5/A6
+ mux8_7/A6 mux8_8/A6 mux8_6/A6 mux8_0/A6 VDD VSS left_shifter
Xright_shifter_0 B0 B1 B2 B3 B4 B5 B6 B7 mux8_0/A7 mux8_1/A7 mux8_2/A7 mux8_3/A7 mux8_4/A7
+ mux8_5/A7 mux8_7/A7 mux8_8/A7 mux8_6/A7 VDD VSS right_shifter
XV_FLAG_0 A7 B7 SEL3 mux8_6/A0 V VDD VSS V_FLAG
X8bit_ADDER_0 SEL3 B0 B1 B2 B3 B5 B6 B7 A0 A1 A2 A3 A4 A5 A6 A7 mux8_1/A0 mux8_2/A0
+ mux8_3/A0 mux8_4/A0 mux8_5/A0 mux8_7/A0 mux8_8/A0 mux8_6/A0 mux8_0/A0 B4 VDD VSS
+ x8bit_ADDER
XAND8_0 A7 B7 A6 B6 A5 B5 A4 B4 A3 B3 A2 B2 A1 B1 A0 B0 mux8_1/A2 mux8_2/A2 mux8_3/A2
+ mux8_4/A2 mux8_5/A2 mux8_7/A2 mux8_8/A2 mux8_6/A2 VDD VDD VSS AND8
Xmux8_1 mux8_1/A0 mux8_1/A1 mux8_1/A2 mux8_1/A5 mux8_1/A6 mux8_1/A7 SEL0 OR8_0/S0
+ SEL1 Y0 VDD mux8_1/A4 VSS SEL2 mux8
Xmux8_0 mux8_0/A0 VSS VSS VSS mux8_0/A6 mux8_0/A7 SEL0 VSS SEL1 C VDD VSS VSS SEL2
+ mux8
XNOT8_0 B7 B6 B5 B4 B3 B2 B1 B0 mux8_1/A5 mux8_2/A5 mux8_3/A5 mux8_4/A5 mux8_5/A5
+ mux8_7/A5 mux8_8/A5 mux8_6/A5 VDD VSS NOT8
Xmux8_2 mux8_2/A0 mux8_2/A1 mux8_2/A2 mux8_2/A5 mux8_2/A6 mux8_2/A7 SEL0 OR8_0/S1
+ SEL1 Y1 VDD mux8_2/A4 VSS SEL2 mux8
Xmux8_3 mux8_3/A0 mux8_3/A1 mux8_3/A2 mux8_3/A5 mux8_3/A6 mux8_3/A7 SEL0 OR8_0/S2
+ SEL1 Y2 VDD mux8_3/A4 VSS SEL2 mux8
Xbuffer_0 VDD S Y7 VSS buffer
Xmux8_4 mux8_4/A0 mux8_4/A1 mux8_4/A2 mux8_4/A5 mux8_4/A6 mux8_4/A7 SEL0 OR8_0/S3
+ SEL1 Y3 VDD mux8_4/A4 VSS SEL2 mux8
Xmux8_5 mux8_5/A0 mux8_5/A1 mux8_5/A2 mux8_5/A5 mux8_5/A6 mux8_5/A7 SEL0 OR8_0/S4
+ SEL1 Y4 VDD mux8_5/A4 VSS SEL2 mux8
Xmux8_6 mux8_6/A0 mux8_6/A1 mux8_6/A2 mux8_6/A5 mux8_6/A6 mux8_6/A7 SEL0 OR8_0/S7
+ SEL1 Y7 VDD mux8_6/A4 VSS SEL2 mux8
Xmux8_7 mux8_7/A0 mux8_7/A1 mux8_7/A2 mux8_7/A5 mux8_7/A6 mux8_7/A7 SEL0 OR8_0/S5
+ SEL1 Y5 VDD mux8_7/A4 VSS SEL2 mux8
Xmux8_8 mux8_8/A0 mux8_8/A1 mux8_8/A2 mux8_8/A5 mux8_8/A6 mux8_8/A7 SEL0 OR8_0/S6
+ SEL1 Y6 VDD mux8_8/A4 VSS SEL2 mux8
XXOR8_0 A7 B7 B6 B5 B4 B3 B2 B1 B0 A0 A1 A2 A3 A4 A5 A6 mux8_6/A4 mux8_8/A4 mux8_7/A4
+ mux8_5/A4 mux8_4/A4 mux8_3/A4 mux8_2/A4 mux8_1/A4 VDD VSS XOR8
XOR8_0 B7 B6 B5 B4 B3 B2 B1 B0 A0 A1 A2 A3 A4 A5 A6 A7 OR8_0/S7 OR8_0/S6 OR8_0/S5
+ OR8_0/S4 OR8_0/S3 OR8_0/S2 OR8_0/S1 OR8_0/S0 VDD VSS OR8
XMULT_0 A0 B2 B0 B3 A2 A1 mux8_1/A1 mux8_2/A1 mux8_3/A1 mux8_7/A1 mux8_5/A1 mux8_4/A1
+ mux8_6/A1 mux8_8/A1 VDD B1 A3 VSS MULT
.ends

