magic
tech sky130B
magscale 1 2
timestamp 1735576878
<< nwell >>
rect 2355 900 7564 1048
rect 8019 900 8088 1048
rect 2355 562 7528 900
<< locali >>
rect 3121 900 3171 901
rect 3940 900 3990 901
rect 4759 900 4809 901
rect 5578 900 5628 901
rect 6397 900 6447 901
rect 7216 900 7266 901
rect 8035 900 8085 901
<< metal1 >>
rect 2286 980 2452 1164
rect 3105 980 3271 1164
rect 3924 980 4090 1164
rect 4743 980 4909 1164
rect 5562 980 5728 1164
rect 6381 980 6547 1164
rect 7200 980 7366 1164
rect 8019 980 8185 1164
rect 2286 900 2355 980
rect 3105 900 3174 980
rect 3924 900 3993 980
rect 4743 900 4812 980
rect 5562 900 5631 980
rect 6381 900 6450 980
rect 7200 900 7269 980
rect 8019 900 8088 980
rect 3271 387 3286 448
rect 1564 74 1648 387
rect 2383 74 2467 387
rect 3202 74 3286 387
rect 4021 74 4105 387
rect 4840 74 4924 387
rect 5659 74 5743 387
rect 6478 74 6562 387
rect 7297 74 7381 387
rect 7988 251 8103 348
rect 8019 74 8103 251
rect 1467 -110 1648 74
rect 2286 -110 2467 74
rect 3105 -110 3286 74
rect 3924 -110 4105 74
rect 4743 -110 4924 74
rect 5562 -110 5743 74
rect 6381 -110 6562 74
rect 7200 -110 7381 74
rect 7922 -110 8103 74
use buffer  buffer_0 ~/Documents/Dersler/VLSI/vlsi_sky130b/design/mag/inv
timestamp 1735575029
transform -1 0 6445 0 1 312
box -5 -422 786 852
use buffer  buffer_1
timestamp 1735575029
transform -1 0 2350 0 1 312
box -5 -422 786 852
use buffer  buffer_2
timestamp 1735575029
transform -1 0 3169 0 1 312
box -5 -422 786 852
use buffer  buffer_3
timestamp 1735575029
transform -1 0 3988 0 1 312
box -5 -422 786 852
use buffer  buffer_4
timestamp 1735575029
transform -1 0 4807 0 1 312
box -5 -422 786 852
use buffer  buffer_5
timestamp 1735575029
transform -1 0 5626 0 1 312
box -5 -422 786 852
use buffer  buffer_6
timestamp 1735575029
transform -1 0 8083 0 1 312
box -5 -422 786 852
use buffer  buffer_7
timestamp 1735575029
transform -1 0 7264 0 1 312
box -5 -422 786 852
<< labels >>
rlabel metal1 8104 1164 8104 1164 5 A0
port 1 s
rlabel metal1 7282 1164 7282 1164 5 A1
port 2 s
rlabel metal1 6468 1164 6468 1164 5 A2
port 3 s
rlabel metal1 5646 1164 5646 1164 5 A3
port 4 s
rlabel metal1 4822 1164 4822 1164 5 A4
port 5 s
rlabel metal1 4003 1164 4003 1164 5 A5
port 6 s
rlabel metal1 3187 1164 3187 1164 5 A6
port 7 s
rlabel metal1 2373 1164 2373 1164 5 A7
port 8 s
rlabel metal1 8003 -110 8003 -110 5 S0
port 9 s
rlabel metal1 7289 -110 7289 -110 5 S1
port 10 s
rlabel metal1 6472 -110 6472 -110 5 S2
port 11 s
rlabel metal1 5653 -110 5653 -110 5 S3
port 12 s
rlabel metal1 4836 -110 4836 -110 5 S4
port 13 s
rlabel metal1 4017 -110 4017 -110 5 S5
port 14 s
rlabel metal1 3180 -110 3180 -110 5 S6
port 15 s
rlabel metal1 2385 -110 2385 -110 5 S7
port 16 s
rlabel metal1 1566 -110 1566 -110 5 C
port 17 s
<< end >>
