magic
tech sky130B
magscale 1 2
timestamp 1733171533
<< nwell >>
rect 113 573 1412 2357
<< nmos >>
rect 445 -34 505 166
rect 563 -34 623 166
rect 681 -34 741 166
rect 799 -34 859 166
rect 917 -34 977 166
rect 1035 -34 1095 166
<< pmos >>
rect 269 726 329 2010
rect 387 726 447 2010
rect 505 726 565 2010
rect 623 726 683 2010
rect 741 726 801 2010
rect 859 726 919 2010
rect 977 726 1037 2010
rect 1095 726 1155 2010
rect 1213 726 1273 2010
<< ndiff >>
rect 387 154 445 166
rect 387 -22 399 154
rect 433 -22 445 154
rect 387 -34 445 -22
rect 505 154 563 166
rect 505 -22 517 154
rect 551 -22 563 154
rect 505 -34 563 -22
rect 623 154 681 166
rect 623 -22 635 154
rect 669 -22 681 154
rect 623 -34 681 -22
rect 741 154 799 166
rect 741 -22 753 154
rect 787 -22 799 154
rect 741 -34 799 -22
rect 859 154 917 166
rect 859 -22 871 154
rect 905 -22 917 154
rect 859 -34 917 -22
rect 977 154 1035 166
rect 977 -22 989 154
rect 1023 -22 1035 154
rect 977 -34 1035 -22
rect 1095 154 1153 166
rect 1095 -22 1107 154
rect 1141 -22 1153 154
rect 1095 -34 1153 -22
<< pdiff >>
rect 211 1998 269 2010
rect 211 738 223 1998
rect 257 738 269 1998
rect 211 726 269 738
rect 329 1998 387 2010
rect 329 738 341 1998
rect 375 738 387 1998
rect 329 726 387 738
rect 447 1998 505 2010
rect 447 738 459 1998
rect 493 738 505 1998
rect 447 726 505 738
rect 565 1998 623 2010
rect 565 738 577 1998
rect 611 738 623 1998
rect 565 726 623 738
rect 683 1998 741 2010
rect 683 738 695 1998
rect 729 738 741 1998
rect 683 726 741 738
rect 801 1998 859 2010
rect 801 738 813 1998
rect 847 738 859 1998
rect 801 726 859 738
rect 919 1998 977 2010
rect 919 738 931 1998
rect 965 738 977 1998
rect 919 726 977 738
rect 1037 1998 1095 2010
rect 1037 738 1049 1998
rect 1083 738 1095 1998
rect 1037 726 1095 738
rect 1155 1998 1213 2010
rect 1155 738 1167 1998
rect 1201 738 1213 1998
rect 1155 726 1213 738
rect 1273 1998 1331 2010
rect 1273 738 1285 1998
rect 1319 738 1331 1998
rect 1273 726 1331 738
<< ndiffc >>
rect 399 -22 433 154
rect 517 -22 551 154
rect 635 -22 669 154
rect 753 -22 787 154
rect 871 -22 905 154
rect 989 -22 1023 154
rect 1107 -22 1141 154
<< pdiffc >>
rect 223 738 257 1998
rect 341 738 375 1998
rect 459 738 493 1998
rect 577 738 611 1998
rect 695 738 729 1998
rect 813 738 847 1998
rect 931 738 965 1998
rect 1049 738 1083 1998
rect 1167 738 1201 1998
rect 1285 738 1319 1998
<< psubdiff >>
rect 387 -128 1151 -88
rect 387 -186 637 -128
rect 909 -186 1151 -128
rect 387 -262 1151 -186
<< nsubdiff >>
rect 175 2209 500 2284
rect 175 2146 259 2209
rect 401 2146 500 2209
rect 175 2072 500 2146
<< psubdiffcont >>
rect 637 -186 909 -128
<< nsubdiffcont >>
rect 259 2146 401 2209
<< poly >>
rect 269 2010 329 2036
rect 387 2010 447 2036
rect 505 2010 565 2036
rect 623 2010 683 2036
rect 741 2010 801 2036
rect 859 2010 919 2036
rect 977 2010 1037 2036
rect 1095 2010 1155 2036
rect 1213 2010 1273 2036
rect 269 695 329 726
rect 387 695 447 726
rect 505 695 565 726
rect 623 695 683 726
rect 741 695 801 726
rect 859 695 919 726
rect 977 695 1037 726
rect 1095 695 1155 726
rect 1213 695 1273 726
rect 266 679 332 695
rect 266 645 282 679
rect 316 645 332 679
rect 266 629 332 645
rect 384 679 450 695
rect 384 645 400 679
rect 434 645 450 679
rect 384 629 450 645
rect 502 679 568 695
rect 502 645 518 679
rect 552 645 568 679
rect 502 629 568 645
rect 620 679 686 695
rect 620 645 636 679
rect 670 645 686 679
rect 620 629 686 645
rect 738 679 804 695
rect 738 645 754 679
rect 788 645 804 679
rect 738 629 804 645
rect 856 679 922 695
rect 856 645 872 679
rect 906 645 922 679
rect 856 629 922 645
rect 974 679 1040 695
rect 974 645 990 679
rect 1024 645 1040 679
rect 974 629 1040 645
rect 1092 679 1158 695
rect 1092 645 1108 679
rect 1142 645 1158 679
rect 1092 629 1158 645
rect 1210 679 1276 695
rect 1210 645 1226 679
rect 1260 645 1276 679
rect 1210 629 1276 645
rect 442 238 508 254
rect 442 204 458 238
rect 492 204 508 238
rect 442 188 508 204
rect 560 238 626 254
rect 560 204 576 238
rect 610 204 626 238
rect 560 188 626 204
rect 678 238 744 254
rect 678 204 694 238
rect 728 204 744 238
rect 678 188 744 204
rect 796 238 862 254
rect 796 204 812 238
rect 846 204 862 238
rect 796 188 862 204
rect 914 238 980 254
rect 914 204 930 238
rect 964 204 980 238
rect 914 188 980 204
rect 1032 238 1098 254
rect 1032 204 1048 238
rect 1082 204 1098 238
rect 1032 188 1098 204
rect 445 166 505 188
rect 563 166 623 188
rect 681 166 741 188
rect 799 166 859 188
rect 917 166 977 188
rect 1035 166 1095 188
rect 445 -60 505 -34
rect 563 -60 623 -34
rect 681 -60 741 -34
rect 799 -60 859 -34
rect 917 -60 977 -34
rect 1035 -60 1095 -34
<< polycont >>
rect 282 645 316 679
rect 400 645 434 679
rect 518 645 552 679
rect 636 645 670 679
rect 754 645 788 679
rect 872 645 906 679
rect 990 645 1024 679
rect 1108 645 1142 679
rect 1226 645 1260 679
rect 458 204 492 238
rect 576 204 610 238
rect 694 204 728 238
rect 812 204 846 238
rect 930 204 964 238
rect 1048 204 1082 238
<< locali >>
rect 175 2210 500 2218
rect 175 2145 258 2210
rect 402 2145 500 2210
rect 175 2137 500 2145
rect 223 1998 257 2014
rect 223 722 257 738
rect 341 1998 375 2014
rect 341 722 375 738
rect 459 1998 493 2014
rect 459 722 493 738
rect 577 1998 611 2014
rect 577 722 611 738
rect 695 1998 729 2014
rect 695 722 729 738
rect 813 1998 847 2014
rect 813 722 847 738
rect 931 1998 965 2014
rect 931 722 965 738
rect 1049 1998 1083 2014
rect 1049 722 1083 738
rect 1167 1998 1201 2014
rect 1167 722 1201 738
rect 1285 1998 1319 2014
rect 1285 722 1319 738
rect 266 645 282 679
rect 316 645 400 679
rect 434 645 518 679
rect 552 645 568 679
rect 620 645 636 679
rect 670 645 754 679
rect 788 645 872 679
rect 906 645 922 679
rect 974 645 990 679
rect 1024 645 1108 679
rect 1142 645 1226 679
rect 1260 645 1276 679
rect 518 306 552 645
rect 754 447 788 645
rect 787 413 788 447
rect 518 238 552 272
rect 754 238 788 413
rect 990 552 1024 645
rect 990 238 1024 518
rect 442 204 458 238
rect 492 204 576 238
rect 610 204 626 238
rect 678 204 694 238
rect 728 204 812 238
rect 846 204 862 238
rect 914 204 930 238
rect 964 204 1048 238
rect 1082 204 1098 238
rect 399 154 433 170
rect 399 -105 433 -22
rect 517 154 551 170
rect 517 -38 551 -22
rect 635 154 669 170
rect 635 -105 669 -22
rect 753 154 787 170
rect 753 -38 787 -22
rect 871 154 905 170
rect 871 -105 905 -22
rect 989 154 1023 170
rect 989 -38 1023 -22
rect 1107 154 1141 170
rect 1107 -105 1141 -22
rect 387 -128 1151 -105
rect 387 -186 637 -128
rect 909 -186 1151 -128
rect 387 -204 1151 -186
<< viali >>
rect 258 2209 402 2210
rect 258 2146 259 2209
rect 259 2146 401 2209
rect 401 2146 402 2209
rect 258 2145 402 2146
rect 223 1425 257 1998
rect 341 738 375 1350
rect 459 1425 493 1998
rect 577 738 611 1350
rect 695 1425 729 1998
rect 813 738 847 1350
rect 931 1425 965 1998
rect 1049 738 1083 1350
rect 1167 1425 1201 1998
rect 1285 738 1319 1350
rect 753 413 787 447
rect 518 272 552 306
rect 990 518 1024 552
rect 517 -22 551 154
rect 753 -22 787 154
rect 989 -22 1023 154
rect 637 -186 909 -128
<< metal1 >>
rect 246 2210 414 2216
rect 246 2145 258 2210
rect 402 2145 414 2210
rect 246 2010 414 2145
rect 217 1998 499 2010
rect 217 1425 223 1998
rect 257 1425 459 1998
rect 493 1425 499 1998
rect 217 1413 499 1425
rect 689 1998 1207 2010
rect 689 1425 695 1998
rect 729 1425 931 1998
rect 965 1425 1167 1998
rect 1201 1425 1207 1998
rect 689 1413 1207 1425
rect 577 1362 853 1363
rect 335 1350 853 1362
rect 335 738 341 1350
rect 375 738 577 1350
rect 611 738 813 1350
rect 847 738 853 1350
rect 335 727 853 738
rect 335 726 617 727
rect 807 726 853 727
rect 1043 1350 1325 1362
rect 1043 738 1049 1350
rect 1083 738 1285 1350
rect 1319 738 1325 1350
rect 1043 726 1325 738
rect 247 552 1036 613
rect 247 518 990 552
rect 1024 518 1036 552
rect 247 515 1036 518
rect 983 511 1036 515
rect 247 447 807 487
rect 247 413 753 447
rect 787 413 807 447
rect 247 389 807 413
rect 246 306 570 353
rect 246 272 518 306
rect 552 272 570 306
rect 246 255 570 272
rect 1167 166 1325 726
rect 511 154 1325 166
rect 511 -22 517 154
rect 551 -22 753 154
rect 787 -22 989 154
rect 1023 -22 1325 154
rect 511 -34 1325 -22
rect 625 -128 921 -120
rect 625 -186 637 -128
rect 909 -186 921 -128
rect 625 -193 921 -186
<< labels >>
flabel metal1 1189 433 1305 551 1 FreeSerif 320 0 0 0 Y
port 1 n
flabel nwell 277 2145 382 2212 1 FreeSerif 320 0 0 0 VDD
port 2 n
flabel metal1 744 -181 804 -134 1 FreeSerif 320 0 0 0 VSS
port 3 n
flabel metal1 253 272 320 340 1 FreeSerif 320 0 0 0 A
port 4 n
flabel metal1 256 405 323 473 1 FreeSerif 320 0 0 0 B
port 5 n
flabel metal1 256 524 323 592 1 FreeSerif 320 0 0 0 C
port 6 n
<< end >>
