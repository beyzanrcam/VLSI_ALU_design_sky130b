magic
tech sky130B
magscale 1 2
timestamp 1735651099
<< nwell >>
rect 1125 562 8088 1048
<< locali >>
rect 1567 900 1617 901
rect 2386 900 2436 901
rect 3205 900 3255 901
rect 4024 900 4074 901
rect 4843 900 4893 901
rect 5662 900 5712 901
rect 6481 900 6531 901
<< metal1 >>
rect 1269 1048 1275 1142
rect 1124 1026 1275 1048
rect 1391 1026 1397 1142
rect 1124 985 1287 1026
rect 1124 899 1193 985
rect 1467 980 1633 1164
rect 2286 980 2452 1164
rect 3105 980 3271 1164
rect 3924 980 4090 1164
rect 4743 980 4909 1164
rect 5562 980 5728 1164
rect 6381 980 6547 1164
rect 7200 980 7366 1164
rect 1564 900 1633 980
rect 2383 900 2452 980
rect 3202 900 3271 980
rect 4021 900 4090 980
rect 4840 900 4909 980
rect 5659 900 5728 980
rect 6478 900 6547 980
rect 7297 900 7366 980
rect 1124 891 1186 899
rect 1271 120 1368 251
rect 1271 17 1368 23
rect 1452 75 1536 471
rect 6366 387 6381 448
rect 1452 74 1549 75
rect 2271 74 2355 387
rect 3090 74 3174 387
rect 3909 74 3993 387
rect 4728 74 4812 387
rect 5547 74 5631 387
rect 6366 74 6450 387
rect 7185 74 7269 387
rect 8004 74 8088 387
rect 1452 -110 1633 74
rect 2271 -110 2452 74
rect 3090 -110 3271 74
rect 3909 -110 4090 74
rect 4728 -110 4909 74
rect 5547 -110 5728 74
rect 6366 -110 6547 74
rect 7185 -110 7366 74
rect 8004 -110 8185 74
<< via1 >>
rect 1275 1026 1391 1142
rect 1271 23 1368 120
<< metal2 >>
rect 1269 1026 1275 1142
rect 1391 1026 1397 1142
rect 1262 23 1271 120
rect 1368 23 1377 120
<< via2 >>
rect 1280 1031 1386 1137
rect 1271 23 1368 120
<< metal3 >>
rect 1276 1142 1390 1147
rect 1275 1141 1391 1142
rect 1275 1027 1276 1141
rect 1390 1027 1391 1141
rect 1275 1026 1391 1027
rect 1276 1021 1390 1026
rect 1266 125 1373 131
rect 1266 12 1373 18
<< via3 >>
rect 1276 1137 1390 1141
rect 1276 1031 1280 1137
rect 1280 1031 1386 1137
rect 1386 1031 1390 1137
rect 1276 1027 1390 1031
rect 1266 120 1373 125
rect 1266 23 1271 120
rect 1271 23 1368 120
rect 1368 23 1373 120
rect 1266 18 1373 23
<< metal4 >>
rect 1275 1141 7751 1142
rect 1275 1027 1276 1141
rect 1390 1027 7751 1141
rect 1275 1026 7751 1027
<< via4 >>
rect 1184 125 1456 208
rect 1184 18 1266 125
rect 1266 18 1373 125
rect 1373 18 1456 125
rect 1184 -64 1456 18
<< metal5 >>
rect 1141 208 7921 251
rect 1141 -64 1184 208
rect 1456 -64 7921 208
rect 1141 -110 7921 -64
use buffer  buffer_0 ~/Documents/Dersler/VLSI/vlsi_sky130b/design/mag/inv
timestamp 1735596573
transform 1 0 5664 0 1 312
box -5 -422 786 852
use buffer  buffer_1
timestamp 1735596573
transform 1 0 1569 0 1 312
box -5 -422 786 852
use buffer  buffer_2
timestamp 1735596573
transform 1 0 2388 0 1 312
box -5 -422 786 852
use buffer  buffer_3
timestamp 1735596573
transform 1 0 3207 0 1 312
box -5 -422 786 852
use buffer  buffer_4
timestamp 1735596573
transform 1 0 4026 0 1 312
box -5 -422 786 852
use buffer  buffer_5
timestamp 1735596573
transform 1 0 4845 0 1 312
box -5 -422 786 852
use buffer  buffer_6
timestamp 1735596573
transform 1 0 7302 0 1 312
box -5 -422 786 852
use buffer  buffer_7
timestamp 1735596573
transform 1 0 6483 0 1 312
box -5 -422 786 852
use inv  inv_0 ~/Documents/Dersler/VLSI/vlsi_sky130b/design/mag/inv
timestamp 1735590487
transform 1 0 1124 0 1 562
box 0 -311 412 486
<< labels >>
rlabel metal1 7281 1164 7281 1164 5 A0
port 1 s
rlabel metal1 6467 1164 6467 1164 5 A1
port 2 s
rlabel metal1 5653 1164 5653 1164 5 A2
port 3 s
rlabel metal1 4826 1164 4826 1164 5 A3
port 4 s
rlabel metal1 4011 1164 4011 1164 5 A4
port 5 s
rlabel metal1 3184 1164 3184 1164 5 A5
port 6 s
rlabel metal1 2366 1164 2366 1164 5 A6
port 7 s
rlabel metal1 1555 1164 1555 1164 5 A7
port 8 s
rlabel metal1 8095 -110 8095 -110 5 C
port 9 s
rlabel metal1 7280 -110 7280 -110 5 S0
port 10 s
rlabel metal1 6461 -110 6461 -110 5 S1
port 11 s
rlabel metal1 5633 -110 5633 -110 5 S2
port 12 s
rlabel metal1 4817 -110 4817 -110 5 S3
port 13 s
rlabel metal1 4000 -110 4000 -110 5 S4
port 14 s
rlabel metal1 3183 -110 3183 -110 5 S5
port 15 s
rlabel metal1 2364 -110 2364 -110 5 S6
port 16 s
rlabel metal1 1546 -110 1546 -110 5 S7
port 17 s
rlabel metal5 4800 -110 4800 -110 5 VSS
port 18 s
rlabel metal4 4826 1142 4826 1142 5 VDD
port 19 s
<< end >>
