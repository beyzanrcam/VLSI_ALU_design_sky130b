magic
tech sky130B
magscale 1 2
timestamp 1736010558
<< nwell >>
rect 3789 899 4035 1429
<< metal1 >>
rect 36 1590 100 1640
rect 518 1588 582 1638
rect 976 1588 1040 1638
rect 1436 1590 1500 1640
rect 1916 1590 1980 1640
rect 2418 1592 2482 1642
rect 2896 1588 2960 1638
rect 3396 1590 3460 1640
rect 4000 1594 4066 1642
rect 4476 1594 4542 1642
rect 4940 1594 5006 1642
rect 5398 1594 5464 1642
rect 5878 1594 5944 1642
rect 6378 1596 6444 1644
rect 6860 1594 6926 1642
rect 7358 1598 7424 1646
rect -691 0 446 48
rect 623 5 926 53
rect -691 -894 -643 0
rect -522 -677 -470 -671
rect -522 -735 -470 -729
rect -520 -911 -472 -735
rect 623 -859 671 5
rect 778 -858 784 -806
rect 836 -858 842 -806
rect 1338 -813 1386 56
rect 1798 -479 1846 60
rect 2278 -397 2326 55
rect 2778 -307 2826 69
rect 3258 -207 3306 69
rect 6739 63 6791 69
rect 3758 -112 3806 51
rect 4353 -2 4359 50
rect 4411 -2 4417 50
rect 4833 6 4839 58
rect 4891 6 4897 58
rect 5299 54 5351 60
rect 5753 2 5759 54
rect 5811 2 5817 54
rect 6239 50 6291 56
rect 5299 -4 5351 2
rect 6739 5 6791 11
rect 7213 -2 7219 50
rect 7271 -2 7277 50
rect 7721 0 8043 48
rect 6239 -8 6291 -2
rect 3758 -160 7879 -112
rect 3258 -255 6702 -207
rect 2778 -355 5503 -307
rect 2278 -445 4359 -397
rect 1798 -527 3178 -479
rect 1338 -861 1970 -813
rect 2080 -867 2086 -815
rect 2138 -867 2144 -815
rect 3130 -984 3178 -527
rect 3289 -863 3295 -811
rect 3347 -863 3353 -811
rect 4311 -1011 4359 -445
rect 4474 -867 4480 -815
rect 4532 -867 4538 -815
rect 5455 -1029 5503 -355
rect 5601 -867 5607 -815
rect 5659 -867 5665 -815
rect 6654 -997 6702 -255
rect 6805 -886 6811 -834
rect 6863 -886 6869 -834
rect 7831 -952 7879 -160
rect 7995 -957 8043 0
rect 322 -2720 354 -2696
rect 1628 -2714 1660 -2690
rect 2930 -2716 2962 -2692
rect 4132 -2714 4164 -2690
rect 5324 -2718 5356 -2694
rect 6424 -2714 6456 -2690
rect 7614 -2724 7668 -2690
rect 8820 -2718 8852 -2694
<< via1 >>
rect -522 -729 -470 -677
rect 784 -858 836 -806
rect 4359 -2 4411 50
rect 4839 6 4891 58
rect 5299 2 5351 54
rect 5759 2 5811 54
rect 6239 -2 6291 50
rect 6739 11 6791 63
rect 7219 -2 7271 50
rect 2086 -867 2138 -815
rect 3295 -863 3347 -811
rect 4480 -867 4532 -815
rect 5607 -867 5659 -815
rect 6811 -886 6863 -834
<< metal2 >>
rect 4839 58 4891 64
rect 4359 50 4411 56
rect -520 0 4359 48
rect -520 -677 -472 0
rect 5759 54 5811 60
rect 4839 0 4891 6
rect 5293 2 5299 54
rect 5351 2 5357 54
rect 4359 -8 4411 -2
rect 4841 -59 4889 0
rect 786 -107 4889 -59
rect -528 -729 -522 -677
rect -470 -729 -464 -677
rect 786 -800 834 -107
rect 5301 -160 5349 2
rect 5759 -4 5811 2
rect 6233 -2 6239 50
rect 6291 -2 6297 50
rect 6733 11 6739 63
rect 6791 11 6797 63
rect 7219 50 7271 56
rect 2088 -208 5349 -160
rect 784 -806 836 -800
rect 2088 -809 2136 -208
rect 5761 -256 5809 -4
rect 3297 -304 5809 -256
rect 3297 -805 3345 -304
rect 6241 -394 6289 -2
rect 4482 -442 6289 -394
rect 784 -864 836 -858
rect 2086 -815 2138 -809
rect 2086 -873 2138 -867
rect 3295 -811 3347 -805
rect 4482 -809 4530 -442
rect 6741 -528 6789 11
rect 7219 -8 7271 -2
rect 5609 -576 6789 -528
rect 5609 -809 5657 -576
rect 7221 -629 7269 -8
rect 6813 -677 7269 -629
rect 3295 -869 3347 -863
rect 4480 -815 4532 -809
rect 4480 -873 4532 -867
rect 5607 -815 5659 -809
rect 6813 -828 6861 -677
rect 5607 -873 5659 -867
rect 6811 -834 6863 -828
rect 6811 -892 6863 -886
<< metal4 >>
rect 3674 1480 4130 1644
use NAND8  NAND8_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NAND8
timestamp 1735984326
transform 1 0 4552 0 1 -1997
box -5260 -734 4324 1197
use NOT8  NOT8_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NOT
timestamp 1735843251
transform 1 0 4073 0 1 501
box -110 -501 3853 1143
use NOT8  NOT8_1
timestamp 1735843251
transform 1 0 110 0 1 501
box -110 -501 3853 1143
<< labels >>
flabel metal1 52 1602 84 1628 0 FreeSans 160 0 0 0 B7
port 1 nsew
flabel metal1 530 1604 562 1630 0 FreeSans 160 0 0 0 B6
port 2 nsew
flabel metal1 992 1600 1024 1626 0 FreeSans 160 0 0 0 B5
port 3 nsew
flabel metal1 1452 1598 1484 1624 0 FreeSans 160 0 0 0 B4
port 4 nsew
flabel metal1 1934 1604 1966 1630 0 FreeSans 160 0 0 0 B3
port 5 nsew
flabel metal1 2436 1604 2468 1630 0 FreeSans 160 0 0 0 B2
port 6 nsew
flabel metal1 2912 1604 2944 1630 0 FreeSans 160 0 0 0 B1
port 7 nsew
flabel metal1 3414 1604 3446 1630 0 FreeSans 160 0 0 0 B0
port 8 nsew
flabel metal1 4012 1602 4044 1628 0 FreeSans 160 0 0 0 A7
port 9 nsew
flabel metal1 4498 1604 4530 1628 0 FreeSans 160 0 0 0 A6
port 10 nsew
flabel metal1 4956 1598 4988 1622 0 FreeSans 160 0 0 0 A5
port 11 nsew
flabel metal1 5418 1604 5450 1628 0 FreeSans 160 0 0 0 A4
port 12 nsew
flabel metal1 5896 1600 5928 1624 0 FreeSans 160 0 0 0 A3
port 13 nsew
flabel metal1 6392 1602 6424 1626 0 FreeSans 160 0 0 0 A2
port 14 nsew
flabel metal1 6876 1606 6908 1630 0 FreeSans 160 0 0 0 A1
port 15 nsew
flabel metal1 7378 1604 7410 1628 0 FreeSans 160 0 0 0 A0
port 16 nsew
flabel metal1 8820 -2718 8852 -2694 0 FreeSans 160 0 0 0 S0
port 17 nsew
flabel metal1 7626 -2718 7658 -2694 0 FreeSans 160 0 0 0 S1
port 18 nsew
flabel metal1 6424 -2714 6456 -2690 0 FreeSans 160 0 0 0 S2
port 19 nsew
flabel metal1 5324 -2718 5356 -2694 0 FreeSans 160 0 0 0 S3
port 20 nsew
flabel metal1 4132 -2714 4164 -2690 0 FreeSans 160 0 0 0 S4
port 21 nsew
flabel metal1 2930 -2716 2962 -2692 0 FreeSans 160 0 0 0 S5
port 22 nsew
flabel metal1 1628 -2714 1660 -2690 0 FreeSans 160 0 0 0 S6
port 23 nsew
flabel metal1 322 -2720 354 -2696 0 FreeSans 160 0 0 0 S7
port 24 nsew
<< end >>
