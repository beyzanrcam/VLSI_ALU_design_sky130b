magic
tech sky130B
magscale 1 2
timestamp 1736276957
<< nwell >>
rect -3447 3502 -2268 4023
rect -1606 3502 -427 4023
rect 235 3502 1414 4023
rect 2076 3502 3255 4023
<< nmos >>
rect -3177 3342 -2777 3372
rect -2544 3346 -2344 3376
rect -1336 3342 -936 3372
rect -703 3346 -503 3376
rect 505 3342 905 3372
rect 1138 3346 1338 3376
rect 2346 3342 2746 3372
rect 2979 3346 3179 3376
rect -3177 3246 -2777 3276
rect -1336 3246 -936 3276
rect 505 3246 905 3276
rect 2346 3246 2746 3276
<< pmos >>
rect -3349 3564 -3319 3778
rect -3253 3564 -3223 3778
rect -3157 3564 -3127 3778
rect -3061 3564 -3031 3778
rect -2965 3564 -2935 3778
rect -2869 3564 -2839 3778
rect -2544 3792 -2330 3822
rect -2544 3696 -2330 3726
rect -2544 3600 -2330 3630
rect -1508 3564 -1478 3778
rect -1412 3564 -1382 3778
rect -1316 3564 -1286 3778
rect -1220 3564 -1190 3778
rect -1124 3564 -1094 3778
rect -1028 3564 -998 3778
rect -703 3792 -489 3822
rect -703 3696 -489 3726
rect -703 3600 -489 3630
rect 333 3564 363 3778
rect 429 3564 459 3778
rect 525 3564 555 3778
rect 621 3564 651 3778
rect 717 3564 747 3778
rect 813 3564 843 3778
rect 1138 3792 1352 3822
rect 1138 3696 1352 3726
rect 1138 3600 1352 3630
rect 2174 3564 2204 3778
rect 2270 3564 2300 3778
rect 2366 3564 2396 3778
rect 2462 3564 2492 3778
rect 2558 3564 2588 3778
rect 2654 3564 2684 3778
rect 2979 3792 3193 3822
rect 2979 3696 3193 3726
rect 2979 3600 3193 3630
<< ndiff >>
rect -3177 3422 -2777 3434
rect -3177 3388 -3165 3422
rect -2789 3388 -2777 3422
rect -2544 3422 -2344 3434
rect -3177 3372 -2777 3388
rect -2544 3388 -2532 3422
rect -2356 3388 -2344 3422
rect -2544 3376 -2344 3388
rect -3177 3276 -2777 3342
rect -2544 3334 -2344 3346
rect -2544 3300 -2532 3334
rect -2356 3300 -2344 3334
rect -2544 3288 -2344 3300
rect -1336 3422 -936 3434
rect -1336 3388 -1324 3422
rect -948 3388 -936 3422
rect -703 3422 -503 3434
rect -1336 3372 -936 3388
rect -703 3388 -691 3422
rect -515 3388 -503 3422
rect -703 3376 -503 3388
rect -1336 3276 -936 3342
rect -703 3334 -503 3346
rect -703 3300 -691 3334
rect -515 3300 -503 3334
rect -703 3288 -503 3300
rect 505 3422 905 3434
rect 505 3388 517 3422
rect 893 3388 905 3422
rect 1138 3422 1338 3434
rect 505 3372 905 3388
rect 1138 3388 1150 3422
rect 1326 3388 1338 3422
rect 1138 3376 1338 3388
rect 505 3276 905 3342
rect 1138 3334 1338 3346
rect 1138 3300 1150 3334
rect 1326 3300 1338 3334
rect 1138 3288 1338 3300
rect 2346 3422 2746 3434
rect 2346 3388 2358 3422
rect 2734 3388 2746 3422
rect 2979 3422 3179 3434
rect 2346 3372 2746 3388
rect 2979 3388 2991 3422
rect 3167 3388 3179 3422
rect 2979 3376 3179 3388
rect 2346 3276 2746 3342
rect 2979 3334 3179 3346
rect 2979 3300 2991 3334
rect 3167 3300 3179 3334
rect 2979 3288 3179 3300
rect -3177 3230 -2777 3246
rect -3177 3196 -3165 3230
rect -2789 3196 -2777 3230
rect -1336 3230 -936 3246
rect -3177 3184 -2777 3196
rect -1336 3196 -1324 3230
rect -948 3196 -936 3230
rect 505 3230 905 3246
rect -1336 3184 -936 3196
rect 505 3196 517 3230
rect 893 3196 905 3230
rect 2346 3230 2746 3246
rect 505 3184 905 3196
rect 2346 3196 2358 3230
rect 2734 3196 2746 3230
rect 2346 3184 2746 3196
<< pdiff >>
rect -2544 3872 -2330 3884
rect -3411 3766 -3349 3778
rect -3411 3576 -3399 3766
rect -3365 3576 -3349 3766
rect -3411 3564 -3349 3576
rect -3319 3766 -3253 3778
rect -3319 3576 -3303 3766
rect -3269 3576 -3253 3766
rect -3319 3564 -3253 3576
rect -3223 3766 -3157 3778
rect -3223 3576 -3207 3766
rect -3173 3576 -3157 3766
rect -3223 3564 -3157 3576
rect -3127 3766 -3061 3778
rect -3127 3576 -3111 3766
rect -3077 3576 -3061 3766
rect -3127 3564 -3061 3576
rect -3031 3766 -2965 3778
rect -3031 3576 -3015 3766
rect -2981 3576 -2965 3766
rect -3031 3564 -2965 3576
rect -2935 3766 -2869 3778
rect -2935 3576 -2919 3766
rect -2885 3576 -2869 3766
rect -2935 3564 -2869 3576
rect -2839 3766 -2777 3778
rect -2839 3576 -2823 3766
rect -2789 3576 -2777 3766
rect -2544 3838 -2532 3872
rect -2342 3838 -2330 3872
rect -2544 3822 -2330 3838
rect -703 3872 -489 3884
rect -2544 3776 -2330 3792
rect -2544 3742 -2532 3776
rect -2338 3742 -2330 3776
rect -2544 3726 -2330 3742
rect -1570 3766 -1508 3778
rect -2544 3680 -2330 3696
rect -2544 3646 -2532 3680
rect -2342 3646 -2330 3680
rect -2544 3630 -2330 3646
rect -2544 3584 -2330 3600
rect -2839 3564 -2777 3576
rect -2544 3550 -2532 3584
rect -2338 3550 -2330 3584
rect -1570 3576 -1558 3766
rect -1524 3576 -1508 3766
rect -1570 3564 -1508 3576
rect -1478 3766 -1412 3778
rect -1478 3576 -1462 3766
rect -1428 3576 -1412 3766
rect -1478 3564 -1412 3576
rect -1382 3766 -1316 3778
rect -1382 3576 -1366 3766
rect -1332 3576 -1316 3766
rect -1382 3564 -1316 3576
rect -1286 3766 -1220 3778
rect -1286 3576 -1270 3766
rect -1236 3576 -1220 3766
rect -1286 3564 -1220 3576
rect -1190 3766 -1124 3778
rect -1190 3576 -1174 3766
rect -1140 3576 -1124 3766
rect -1190 3564 -1124 3576
rect -1094 3766 -1028 3778
rect -1094 3576 -1078 3766
rect -1044 3576 -1028 3766
rect -1094 3564 -1028 3576
rect -998 3766 -936 3778
rect -998 3576 -982 3766
rect -948 3576 -936 3766
rect -703 3838 -691 3872
rect -501 3838 -489 3872
rect -703 3822 -489 3838
rect 1138 3872 1352 3884
rect -703 3776 -489 3792
rect -703 3742 -691 3776
rect -497 3742 -489 3776
rect -703 3726 -489 3742
rect 271 3766 333 3778
rect -703 3680 -489 3696
rect -703 3646 -691 3680
rect -501 3646 -489 3680
rect -703 3630 -489 3646
rect -703 3584 -489 3600
rect -998 3564 -936 3576
rect -2544 3538 -2330 3550
rect -703 3550 -691 3584
rect -497 3550 -489 3584
rect 271 3576 283 3766
rect 317 3576 333 3766
rect 271 3564 333 3576
rect 363 3766 429 3778
rect 363 3576 379 3766
rect 413 3576 429 3766
rect 363 3564 429 3576
rect 459 3766 525 3778
rect 459 3576 475 3766
rect 509 3576 525 3766
rect 459 3564 525 3576
rect 555 3766 621 3778
rect 555 3576 571 3766
rect 605 3576 621 3766
rect 555 3564 621 3576
rect 651 3766 717 3778
rect 651 3576 667 3766
rect 701 3576 717 3766
rect 651 3564 717 3576
rect 747 3766 813 3778
rect 747 3576 763 3766
rect 797 3576 813 3766
rect 747 3564 813 3576
rect 843 3766 905 3778
rect 843 3576 859 3766
rect 893 3576 905 3766
rect 1138 3838 1150 3872
rect 1340 3838 1352 3872
rect 1138 3822 1352 3838
rect 2979 3872 3193 3884
rect 1138 3776 1352 3792
rect 1138 3742 1150 3776
rect 1344 3742 1352 3776
rect 1138 3726 1352 3742
rect 2112 3766 2174 3778
rect 1138 3680 1352 3696
rect 1138 3646 1150 3680
rect 1340 3646 1352 3680
rect 1138 3630 1352 3646
rect 1138 3584 1352 3600
rect 843 3564 905 3576
rect -703 3538 -489 3550
rect 1138 3550 1150 3584
rect 1344 3550 1352 3584
rect 2112 3576 2124 3766
rect 2158 3576 2174 3766
rect 2112 3564 2174 3576
rect 2204 3766 2270 3778
rect 2204 3576 2220 3766
rect 2254 3576 2270 3766
rect 2204 3564 2270 3576
rect 2300 3766 2366 3778
rect 2300 3576 2316 3766
rect 2350 3576 2366 3766
rect 2300 3564 2366 3576
rect 2396 3766 2462 3778
rect 2396 3576 2412 3766
rect 2446 3576 2462 3766
rect 2396 3564 2462 3576
rect 2492 3766 2558 3778
rect 2492 3576 2508 3766
rect 2542 3576 2558 3766
rect 2492 3564 2558 3576
rect 2588 3766 2654 3778
rect 2588 3576 2604 3766
rect 2638 3576 2654 3766
rect 2588 3564 2654 3576
rect 2684 3766 2746 3778
rect 2684 3576 2700 3766
rect 2734 3576 2746 3766
rect 2979 3838 2991 3872
rect 3181 3838 3193 3872
rect 2979 3822 3193 3838
rect 2979 3776 3193 3792
rect 2979 3742 2991 3776
rect 3185 3742 3193 3776
rect 2979 3726 3193 3742
rect 2979 3680 3193 3696
rect 2979 3646 2991 3680
rect 3181 3646 3193 3680
rect 2979 3630 3193 3646
rect 2979 3584 3193 3600
rect 2684 3564 2746 3576
rect 1138 3538 1352 3550
rect 2979 3550 2991 3584
rect 3185 3550 3193 3584
rect 2979 3538 3193 3550
<< ndiffc >>
rect -3165 3388 -2789 3422
rect -2532 3388 -2356 3422
rect -2532 3300 -2356 3334
rect -1324 3388 -948 3422
rect -691 3388 -515 3422
rect -691 3300 -515 3334
rect 517 3388 893 3422
rect 1150 3388 1326 3422
rect 1150 3300 1326 3334
rect 2358 3388 2734 3422
rect 2991 3388 3167 3422
rect 2991 3300 3167 3334
rect -3165 3196 -2789 3230
rect -1324 3196 -948 3230
rect 517 3196 893 3230
rect 2358 3196 2734 3230
<< pdiffc >>
rect -3399 3576 -3365 3766
rect -3303 3576 -3269 3766
rect -3207 3576 -3173 3766
rect -3111 3576 -3077 3766
rect -3015 3576 -2981 3766
rect -2919 3576 -2885 3766
rect -2823 3576 -2789 3766
rect -2532 3838 -2342 3872
rect -2532 3742 -2338 3776
rect -2532 3646 -2342 3680
rect -2532 3550 -2338 3584
rect -1558 3576 -1524 3766
rect -1462 3576 -1428 3766
rect -1366 3576 -1332 3766
rect -1270 3576 -1236 3766
rect -1174 3576 -1140 3766
rect -1078 3576 -1044 3766
rect -982 3576 -948 3766
rect -691 3838 -501 3872
rect -691 3742 -497 3776
rect -691 3646 -501 3680
rect -691 3550 -497 3584
rect 283 3576 317 3766
rect 379 3576 413 3766
rect 475 3576 509 3766
rect 571 3576 605 3766
rect 667 3576 701 3766
rect 763 3576 797 3766
rect 859 3576 893 3766
rect 1150 3838 1340 3872
rect 1150 3742 1344 3776
rect 1150 3646 1340 3680
rect 1150 3550 1344 3584
rect 2124 3576 2158 3766
rect 2220 3576 2254 3766
rect 2316 3576 2350 3766
rect 2412 3576 2446 3766
rect 2508 3576 2542 3766
rect 2604 3576 2638 3766
rect 2700 3576 2734 3766
rect 2991 3838 3181 3872
rect 2991 3742 3185 3776
rect 2991 3646 3181 3680
rect 2991 3550 3185 3584
<< psubdiff >>
rect -3177 3160 -2777 3184
rect -3177 3086 -3150 3160
rect -2815 3086 -2777 3160
rect -3177 3067 -2777 3086
rect -1336 3160 -936 3184
rect -1336 3086 -1309 3160
rect -974 3086 -936 3160
rect -1336 3067 -936 3086
rect 505 3160 905 3184
rect 505 3086 532 3160
rect 867 3086 905 3160
rect 505 3067 905 3086
rect 2346 3160 2746 3184
rect 2346 3086 2373 3160
rect 2708 3086 2746 3160
rect 2346 3067 2746 3086
<< nsubdiff >>
rect -3407 3921 -2790 3982
rect -3407 3874 -3197 3921
rect -2957 3874 -2790 3921
rect -1566 3921 -949 3982
rect -3407 3832 -2790 3874
rect -1566 3874 -1356 3921
rect -1116 3874 -949 3921
rect 275 3921 892 3982
rect -1566 3832 -949 3874
rect 275 3874 485 3921
rect 725 3874 892 3921
rect 2116 3921 2733 3982
rect 275 3832 892 3874
rect 2116 3874 2326 3921
rect 2566 3874 2733 3921
rect 2116 3832 2733 3874
<< psubdiffcont >>
rect -3150 3086 -2815 3160
rect -1309 3086 -974 3160
rect 532 3086 867 3160
rect 2373 3086 2708 3160
<< nsubdiffcont >>
rect -3197 3874 -2957 3921
rect -1356 3874 -1116 3921
rect 485 3874 725 3921
rect 2326 3874 2566 3921
<< poly >>
rect -2641 3824 -2575 3840
rect -3349 3778 -3319 3809
rect -3253 3778 -3223 3809
rect -3157 3778 -3127 3809
rect -3061 3778 -3031 3809
rect -2965 3778 -2935 3809
rect -2869 3778 -2839 3809
rect -2641 3598 -2625 3824
rect -2591 3822 -2575 3824
rect -800 3824 -734 3840
rect -2591 3792 -2544 3822
rect -2330 3792 -2304 3822
rect -2591 3726 -2575 3792
rect -1508 3778 -1478 3809
rect -1412 3778 -1382 3809
rect -1316 3778 -1286 3809
rect -1220 3778 -1190 3809
rect -1124 3778 -1094 3809
rect -1028 3778 -998 3809
rect -2591 3696 -2544 3726
rect -2330 3696 -2304 3726
rect -2591 3630 -2575 3696
rect -2591 3600 -2544 3630
rect -2330 3600 -2304 3630
rect -2591 3598 -2575 3600
rect -2641 3582 -2575 3598
rect -3349 3538 -3319 3564
rect -3253 3538 -3223 3564
rect -3157 3538 -3127 3564
rect -3350 3517 -3127 3538
rect -3350 3482 -3333 3517
rect -3299 3508 -3127 3517
rect -3061 3538 -3031 3564
rect -2965 3538 -2935 3564
rect -2869 3538 -2839 3564
rect -800 3598 -784 3824
rect -750 3822 -734 3824
rect 1041 3824 1107 3840
rect -750 3792 -703 3822
rect -489 3792 -463 3822
rect -750 3726 -734 3792
rect 333 3778 363 3809
rect 429 3778 459 3809
rect 525 3778 555 3809
rect 621 3778 651 3809
rect 717 3778 747 3809
rect 813 3778 843 3809
rect -750 3696 -703 3726
rect -489 3696 -463 3726
rect -750 3630 -734 3696
rect -750 3600 -703 3630
rect -489 3600 -463 3630
rect -750 3598 -734 3600
rect -800 3582 -734 3598
rect -1508 3538 -1478 3564
rect -1412 3538 -1382 3564
rect -1316 3538 -1286 3564
rect -3061 3517 -2839 3538
rect -3299 3482 -3283 3508
rect -3350 3471 -3283 3482
rect -3061 3482 -3044 3517
rect -3010 3508 -2839 3517
rect -1509 3517 -1286 3538
rect -3010 3482 -2994 3508
rect -3061 3471 -2994 3482
rect -1509 3482 -1492 3517
rect -1458 3508 -1286 3517
rect -1220 3538 -1190 3564
rect -1124 3538 -1094 3564
rect -1028 3538 -998 3564
rect 1041 3598 1057 3824
rect 1091 3822 1107 3824
rect 2882 3824 2948 3840
rect 1091 3792 1138 3822
rect 1352 3792 1378 3822
rect 1091 3726 1107 3792
rect 2174 3778 2204 3809
rect 2270 3778 2300 3809
rect 2366 3778 2396 3809
rect 2462 3778 2492 3809
rect 2558 3778 2588 3809
rect 2654 3778 2684 3809
rect 1091 3696 1138 3726
rect 1352 3696 1378 3726
rect 1091 3630 1107 3696
rect 1091 3600 1138 3630
rect 1352 3600 1378 3630
rect 1091 3598 1107 3600
rect 1041 3582 1107 3598
rect 333 3538 363 3564
rect 429 3538 459 3564
rect 525 3538 555 3564
rect -1220 3517 -998 3538
rect -1458 3482 -1442 3508
rect -1509 3471 -1442 3482
rect -1220 3482 -1203 3517
rect -1169 3508 -998 3517
rect 332 3517 555 3538
rect -1169 3482 -1153 3508
rect -1220 3471 -1153 3482
rect 332 3482 349 3517
rect 383 3508 555 3517
rect 621 3538 651 3564
rect 717 3538 747 3564
rect 813 3538 843 3564
rect 2882 3598 2898 3824
rect 2932 3822 2948 3824
rect 2932 3792 2979 3822
rect 3193 3792 3219 3822
rect 2932 3726 2948 3792
rect 2932 3696 2979 3726
rect 3193 3696 3219 3726
rect 2932 3630 2948 3696
rect 2932 3600 2979 3630
rect 3193 3600 3219 3630
rect 2932 3598 2948 3600
rect 2882 3582 2948 3598
rect 2174 3538 2204 3564
rect 2270 3538 2300 3564
rect 2366 3538 2396 3564
rect 621 3517 843 3538
rect 383 3482 399 3508
rect 332 3471 399 3482
rect 621 3482 638 3517
rect 672 3508 843 3517
rect 2173 3517 2396 3538
rect 672 3482 688 3508
rect 621 3471 688 3482
rect 2173 3482 2190 3517
rect 2224 3508 2396 3517
rect 2462 3538 2492 3564
rect 2558 3538 2588 3564
rect 2654 3538 2684 3564
rect 2462 3517 2684 3538
rect 2224 3482 2240 3508
rect 2173 3471 2240 3482
rect 2462 3482 2479 3517
rect 2513 3508 2684 3517
rect 2513 3482 2529 3508
rect 2462 3471 2529 3482
rect -3350 3276 -3307 3471
rect -3265 3393 -3199 3409
rect -3265 3358 -3249 3393
rect -3215 3372 -3199 3393
rect -2641 3378 -2574 3394
rect -3215 3358 -3177 3372
rect -3265 3342 -3177 3358
rect -2777 3342 -2751 3372
rect -2641 3344 -2625 3378
rect -2591 3376 -2574 3378
rect -2591 3346 -2544 3376
rect -2344 3346 -2318 3376
rect -2591 3344 -2574 3346
rect -2641 3328 -2574 3344
rect -1509 3276 -1466 3471
rect -1424 3393 -1358 3409
rect -1424 3358 -1408 3393
rect -1374 3372 -1358 3393
rect -800 3378 -733 3394
rect -1374 3358 -1336 3372
rect -1424 3342 -1336 3358
rect -936 3342 -910 3372
rect -800 3344 -784 3378
rect -750 3376 -733 3378
rect -750 3346 -703 3376
rect -503 3346 -477 3376
rect -750 3344 -733 3346
rect -800 3328 -733 3344
rect 332 3276 375 3471
rect 417 3393 483 3409
rect 417 3358 433 3393
rect 467 3372 483 3393
rect 1041 3378 1108 3394
rect 467 3358 505 3372
rect 417 3342 505 3358
rect 905 3342 931 3372
rect 1041 3344 1057 3378
rect 1091 3376 1108 3378
rect 1091 3346 1138 3376
rect 1338 3346 1364 3376
rect 1091 3344 1108 3346
rect 1041 3328 1108 3344
rect 2173 3276 2216 3471
rect 2258 3393 2324 3409
rect 2258 3358 2274 3393
rect 2308 3372 2324 3393
rect 2882 3378 2949 3394
rect 2308 3358 2346 3372
rect 2258 3342 2346 3358
rect 2746 3342 2772 3372
rect 2882 3344 2898 3378
rect 2932 3376 2949 3378
rect 2932 3346 2979 3376
rect 3179 3346 3205 3376
rect 2932 3344 2949 3346
rect 2882 3328 2949 3344
rect -3350 3260 -3177 3276
rect -3350 3225 -3249 3260
rect -3215 3246 -3177 3260
rect -2777 3246 -2751 3276
rect -1509 3260 -1336 3276
rect -3215 3225 -3199 3246
rect -3350 3209 -3199 3225
rect -1509 3225 -1408 3260
rect -1374 3246 -1336 3260
rect -936 3246 -910 3276
rect 332 3260 505 3276
rect -1374 3225 -1358 3246
rect -1509 3209 -1358 3225
rect 332 3225 433 3260
rect 467 3246 505 3260
rect 905 3246 931 3276
rect 2173 3260 2346 3276
rect 467 3225 483 3246
rect 332 3209 483 3225
rect 2173 3225 2274 3260
rect 2308 3246 2346 3260
rect 2746 3246 2772 3276
rect 2308 3225 2324 3246
rect 2173 3209 2324 3225
<< polycont >>
rect -2625 3598 -2591 3824
rect -3333 3482 -3299 3517
rect -784 3598 -750 3824
rect -3044 3482 -3010 3517
rect -1492 3482 -1458 3517
rect 1057 3598 1091 3824
rect -1203 3482 -1169 3517
rect 349 3482 383 3517
rect 2898 3598 2932 3824
rect 638 3482 672 3517
rect 2190 3482 2224 3517
rect 2479 3482 2513 3517
rect -3249 3358 -3215 3393
rect -2625 3344 -2591 3378
rect -1408 3358 -1374 3393
rect -784 3344 -750 3378
rect 433 3358 467 3393
rect 1057 3344 1091 3378
rect 2274 3358 2308 3393
rect 2898 3344 2932 3378
rect -3249 3225 -3215 3260
rect -1408 3225 -1374 3260
rect 433 3225 467 3260
rect 2274 3225 2308 3260
<< locali >>
rect -3271 3874 -3197 3921
rect -2957 3874 -2857 3921
rect -1430 3874 -1356 3921
rect -1116 3874 -1016 3921
rect 411 3874 485 3921
rect 725 3874 825 3921
rect 2252 3874 2326 3921
rect 2566 3874 2666 3921
rect -2641 3824 -2591 3841
rect -2548 3838 -2538 3872
rect -2342 3838 -2326 3872
rect -3399 3772 -3365 3782
rect -3399 3560 -3365 3576
rect -3303 3766 -3269 3782
rect -3303 3560 -3269 3570
rect -3207 3772 -3173 3782
rect -3207 3560 -3173 3576
rect -3111 3766 -3077 3782
rect -3111 3560 -3077 3570
rect -3015 3772 -2981 3782
rect -3015 3560 -2981 3576
rect -2919 3766 -2885 3782
rect -2919 3560 -2885 3570
rect -2823 3772 -2789 3782
rect -2823 3560 -2789 3576
rect -2641 3598 -2625 3824
rect -800 3824 -750 3841
rect -707 3838 -697 3872
rect -501 3838 -485 3872
rect -2548 3742 -2532 3776
rect -2338 3742 -2320 3776
rect -1558 3772 -1524 3782
rect -2548 3646 -2538 3680
rect -2342 3646 -2326 3680
rect -3350 3482 -3333 3517
rect -3299 3482 -3283 3517
rect -3061 3511 -3044 3517
rect -3249 3482 -3044 3511
rect -3010 3482 -2994 3517
rect -3350 3276 -3307 3482
rect -3249 3477 -2994 3482
rect -3249 3393 -3215 3477
rect -3181 3388 -3165 3422
rect -2789 3388 -2773 3422
rect -3249 3342 -3215 3358
rect -2641 3378 -2591 3598
rect -2548 3550 -2532 3584
rect -2338 3550 -2320 3584
rect -1558 3560 -1524 3576
rect -1462 3766 -1428 3782
rect -1462 3560 -1428 3570
rect -1366 3772 -1332 3782
rect -1366 3560 -1332 3576
rect -1270 3766 -1236 3782
rect -1270 3560 -1236 3570
rect -1174 3772 -1140 3782
rect -1174 3560 -1140 3576
rect -1078 3766 -1044 3782
rect -1078 3560 -1044 3570
rect -982 3772 -948 3782
rect -982 3560 -948 3576
rect -800 3598 -784 3824
rect 1041 3824 1091 3841
rect 1134 3838 1144 3872
rect 1340 3838 1356 3872
rect -707 3742 -691 3776
rect -497 3742 -479 3776
rect 283 3772 317 3782
rect -707 3646 -697 3680
rect -501 3646 -485 3680
rect -1509 3482 -1492 3517
rect -1458 3482 -1442 3517
rect -1220 3511 -1203 3517
rect -1408 3482 -1203 3511
rect -1169 3482 -1153 3517
rect -2548 3388 -2532 3422
rect -2356 3388 -2340 3422
rect -2641 3344 -2625 3378
rect -2641 3328 -2591 3344
rect -2548 3300 -2532 3334
rect -2356 3300 -2340 3334
rect -1509 3276 -1466 3482
rect -1408 3477 -1153 3482
rect -1408 3393 -1374 3477
rect -1340 3388 -1324 3422
rect -948 3388 -932 3422
rect -1408 3342 -1374 3358
rect -800 3378 -750 3598
rect -707 3550 -691 3584
rect -497 3550 -479 3584
rect 283 3560 317 3576
rect 379 3766 413 3782
rect 379 3560 413 3570
rect 475 3772 509 3782
rect 475 3560 509 3576
rect 571 3766 605 3782
rect 571 3560 605 3570
rect 667 3772 701 3782
rect 667 3560 701 3576
rect 763 3766 797 3782
rect 763 3560 797 3570
rect 859 3772 893 3782
rect 859 3560 893 3576
rect 1041 3598 1057 3824
rect 2882 3824 2932 3841
rect 2975 3838 2985 3872
rect 3181 3838 3197 3872
rect 1134 3742 1150 3776
rect 1344 3742 1362 3776
rect 2124 3772 2158 3782
rect 1134 3646 1144 3680
rect 1340 3646 1356 3680
rect 332 3482 349 3517
rect 383 3482 399 3517
rect 621 3511 638 3517
rect 433 3482 638 3511
rect 672 3482 688 3517
rect -707 3388 -691 3422
rect -515 3388 -499 3422
rect -800 3344 -784 3378
rect -800 3328 -750 3344
rect -707 3300 -691 3334
rect -515 3300 -499 3334
rect 332 3276 375 3482
rect 433 3477 688 3482
rect 433 3393 467 3477
rect 501 3388 517 3422
rect 893 3388 909 3422
rect 433 3342 467 3358
rect 1041 3378 1091 3598
rect 1134 3550 1150 3584
rect 1344 3550 1362 3584
rect 2124 3560 2158 3576
rect 2220 3766 2254 3782
rect 2220 3560 2254 3570
rect 2316 3772 2350 3782
rect 2316 3560 2350 3576
rect 2412 3766 2446 3782
rect 2412 3560 2446 3570
rect 2508 3772 2542 3782
rect 2508 3560 2542 3576
rect 2604 3766 2638 3782
rect 2604 3560 2638 3570
rect 2700 3772 2734 3782
rect 2700 3560 2734 3576
rect 2882 3598 2898 3824
rect 2975 3742 2991 3776
rect 3185 3742 3203 3776
rect 2975 3646 2985 3680
rect 3181 3646 3197 3680
rect 2173 3482 2190 3517
rect 2224 3482 2240 3517
rect 2462 3511 2479 3517
rect 2274 3482 2479 3511
rect 2513 3482 2529 3517
rect 1134 3388 1150 3422
rect 1326 3388 1342 3422
rect 1041 3344 1057 3378
rect 1041 3328 1091 3344
rect 1134 3300 1150 3334
rect 1326 3300 1342 3334
rect 2173 3276 2216 3482
rect 2274 3477 2529 3482
rect 2274 3393 2308 3477
rect 2342 3388 2358 3422
rect 2734 3388 2750 3422
rect 2274 3342 2308 3358
rect 2882 3378 2932 3598
rect 2975 3550 2991 3584
rect 3185 3550 3203 3584
rect 2975 3388 2991 3422
rect 3167 3388 3183 3422
rect 2882 3344 2898 3378
rect 2882 3328 2932 3344
rect 2975 3300 2991 3334
rect 3167 3300 3183 3334
rect -3350 3260 -3215 3276
rect -3350 3225 -3249 3260
rect -1509 3260 -1374 3276
rect -3350 3209 -3215 3225
rect -3181 3196 -3165 3230
rect -2789 3196 -2773 3230
rect -1509 3225 -1408 3260
rect 332 3260 467 3276
rect -1509 3209 -1374 3225
rect -1340 3196 -1324 3230
rect -948 3196 -932 3230
rect 332 3225 433 3260
rect 2173 3260 2308 3276
rect 332 3209 467 3225
rect 501 3196 517 3230
rect 893 3196 909 3230
rect 2173 3225 2274 3260
rect 2173 3209 2308 3225
rect 2342 3196 2358 3230
rect 2734 3196 2750 3230
rect -3177 3086 -3150 3160
rect -2815 3086 -2777 3160
rect -1336 3086 -1309 3160
rect -974 3086 -936 3160
rect 505 3086 532 3160
rect 867 3086 905 3160
rect 2346 3086 2373 3160
rect 2708 3086 2746 3160
rect 154 1006 264 1634
rect 154 942 596 1006
<< viali >>
rect -3197 3874 -2957 3921
rect -1356 3874 -1116 3921
rect 485 3874 725 3921
rect 2326 3874 2566 3921
rect -2538 3838 -2532 3872
rect -2532 3838 -2459 3872
rect -3399 3766 -3365 3772
rect -3399 3692 -3365 3766
rect -3303 3576 -3269 3650
rect -3303 3570 -3269 3576
rect -3207 3766 -3173 3772
rect -3207 3692 -3173 3766
rect -3111 3576 -3077 3650
rect -3111 3570 -3077 3576
rect -3015 3766 -2981 3772
rect -3015 3692 -2981 3766
rect -2919 3576 -2885 3650
rect -2919 3570 -2885 3576
rect -2823 3766 -2789 3772
rect -2823 3692 -2789 3766
rect -2625 3598 -2591 3824
rect -697 3838 -691 3872
rect -691 3838 -618 3872
rect -2415 3742 -2338 3776
rect -1558 3766 -1524 3772
rect -1558 3692 -1524 3766
rect -2538 3646 -2532 3680
rect -2532 3646 -2459 3680
rect -3333 3482 -3299 3517
rect -3044 3482 -3010 3517
rect -3249 3358 -3215 3393
rect -3165 3388 -2789 3422
rect -2415 3550 -2338 3584
rect -1462 3576 -1428 3650
rect -1462 3570 -1428 3576
rect -1366 3766 -1332 3772
rect -1366 3692 -1332 3766
rect -1270 3576 -1236 3650
rect -1270 3570 -1236 3576
rect -1174 3766 -1140 3772
rect -1174 3692 -1140 3766
rect -1078 3576 -1044 3650
rect -1078 3570 -1044 3576
rect -982 3766 -948 3772
rect -982 3692 -948 3766
rect -784 3598 -750 3824
rect 1144 3838 1150 3872
rect 1150 3838 1223 3872
rect -574 3742 -497 3776
rect 283 3766 317 3772
rect 283 3692 317 3766
rect -697 3646 -691 3680
rect -691 3646 -618 3680
rect -1492 3482 -1458 3517
rect -1203 3482 -1169 3517
rect -2532 3388 -2356 3422
rect -2625 3344 -2591 3378
rect -2532 3300 -2356 3334
rect -1408 3358 -1374 3393
rect -1324 3388 -948 3422
rect -574 3550 -497 3584
rect 379 3576 413 3650
rect 379 3570 413 3576
rect 475 3766 509 3772
rect 475 3692 509 3766
rect 571 3576 605 3650
rect 571 3570 605 3576
rect 667 3766 701 3772
rect 667 3692 701 3766
rect 763 3576 797 3650
rect 763 3570 797 3576
rect 859 3766 893 3772
rect 859 3692 893 3766
rect 1057 3598 1091 3824
rect 2985 3838 2991 3872
rect 2991 3838 3064 3872
rect 1267 3742 1344 3776
rect 2124 3766 2158 3772
rect 2124 3692 2158 3766
rect 1144 3646 1150 3680
rect 1150 3646 1223 3680
rect 349 3482 383 3517
rect 638 3482 672 3517
rect -691 3388 -515 3422
rect -784 3344 -750 3378
rect -691 3300 -515 3334
rect 433 3358 467 3393
rect 517 3388 893 3422
rect 1267 3550 1344 3584
rect 2220 3576 2254 3650
rect 2220 3570 2254 3576
rect 2316 3766 2350 3772
rect 2316 3692 2350 3766
rect 2412 3576 2446 3650
rect 2412 3570 2446 3576
rect 2508 3766 2542 3772
rect 2508 3692 2542 3766
rect 2604 3576 2638 3650
rect 2604 3570 2638 3576
rect 2700 3766 2734 3772
rect 2700 3692 2734 3766
rect 2898 3598 2932 3824
rect 3108 3742 3185 3776
rect 2985 3646 2991 3680
rect 2991 3646 3064 3680
rect 2190 3482 2224 3517
rect 2479 3482 2513 3517
rect 1150 3388 1326 3422
rect 1057 3344 1091 3378
rect 1150 3300 1326 3334
rect 2274 3358 2308 3393
rect 2358 3388 2734 3422
rect 3108 3550 3185 3584
rect 2991 3388 3167 3422
rect 2898 3344 2932 3378
rect 2991 3300 3167 3334
rect -3165 3196 -2789 3230
rect -1324 3196 -948 3230
rect 517 3196 893 3230
rect 2358 3196 2734 3230
rect -3150 3086 -2815 3155
rect -1309 3086 -974 3155
rect 532 3086 867 3155
rect 2373 3086 2708 3155
<< metal1 >>
rect -3271 3921 -2934 3933
rect -3271 3874 -3197 3921
rect -2957 3874 -2934 3921
rect -1430 3921 -1093 3933
rect -3271 3814 -2934 3874
rect -2548 3872 -2326 3920
rect -2548 3868 -2538 3872
rect -2658 3824 -2575 3840
rect -3412 3778 -2778 3814
rect -3412 3772 -2777 3778
rect -3412 3692 -3399 3772
rect -3365 3692 -3207 3772
rect -3173 3692 -3015 3772
rect -2981 3692 -2823 3772
rect -2789 3692 -2777 3772
rect -3412 3686 -2777 3692
rect -3412 3685 -2778 3686
rect -2658 3656 -2625 3824
rect -3319 3650 -2625 3656
rect -3319 3570 -3303 3650
rect -3269 3570 -3111 3650
rect -3077 3570 -2919 3650
rect -2885 3598 -2625 3650
rect -2591 3598 -2575 3824
rect -2544 3838 -2538 3868
rect -2459 3868 -2326 3872
rect -1430 3874 -1356 3921
rect -1116 3874 -1093 3921
rect 411 3921 748 3933
rect -2459 3838 -2453 3868
rect -2544 3680 -2453 3838
rect -2544 3646 -2538 3680
rect -2459 3646 -2453 3680
rect -2544 3630 -2453 3646
rect -2421 3776 -2268 3840
rect -1430 3814 -1093 3874
rect -707 3872 -485 3920
rect -707 3868 -697 3872
rect -817 3824 -734 3840
rect -2421 3742 -2415 3776
rect -2338 3742 -2268 3776
rect -2885 3570 -2575 3598
rect -2421 3584 -2268 3742
rect -1571 3778 -937 3814
rect -1571 3772 -936 3778
rect -1571 3692 -1558 3772
rect -1524 3692 -1366 3772
rect -1332 3692 -1174 3772
rect -1140 3692 -982 3772
rect -948 3692 -936 3772
rect -1571 3686 -936 3692
rect -1571 3685 -937 3686
rect -817 3656 -784 3824
rect -3319 3564 -2575 3570
rect -3447 3517 -3283 3535
rect -3447 3515 -3333 3517
rect -3447 3405 -3422 3515
rect -3299 3482 -3283 3517
rect -3327 3405 -3283 3482
rect -3447 3400 -3283 3405
rect -3255 3517 -2995 3536
rect -3255 3482 -3044 3517
rect -3010 3482 -2995 3517
rect -3255 3462 -2995 3482
rect -3255 3393 -3205 3462
rect -2919 3434 -2575 3564
rect -3544 3371 -3354 3372
rect -3255 3371 -3249 3393
rect -3544 3358 -3249 3371
rect -3215 3358 -3205 3393
rect -3177 3422 -2575 3434
rect -3177 3388 -3165 3422
rect -2789 3388 -2575 3422
rect -3177 3382 -2575 3388
rect -2544 3550 -2415 3584
rect -2338 3550 -2268 3584
rect -1478 3650 -784 3656
rect -1478 3570 -1462 3650
rect -1428 3570 -1270 3650
rect -1236 3570 -1078 3650
rect -1044 3598 -784 3650
rect -750 3598 -734 3824
rect -703 3838 -697 3868
rect -618 3868 -485 3872
rect 411 3874 485 3921
rect 725 3874 748 3921
rect 2252 3921 2589 3933
rect -618 3838 -612 3868
rect -703 3680 -612 3838
rect -703 3646 -697 3680
rect -618 3646 -612 3680
rect -703 3630 -612 3646
rect -580 3776 -427 3840
rect 411 3814 748 3874
rect 1134 3872 1356 3920
rect 1134 3868 1144 3872
rect 1024 3824 1107 3840
rect -580 3742 -574 3776
rect -497 3742 -427 3776
rect -1044 3570 -734 3598
rect -580 3584 -427 3742
rect 270 3778 904 3814
rect 270 3772 905 3778
rect 270 3692 283 3772
rect 317 3692 475 3772
rect 509 3692 667 3772
rect 701 3692 859 3772
rect 893 3692 905 3772
rect 270 3686 905 3692
rect 270 3685 904 3686
rect 1024 3656 1057 3824
rect -1478 3564 -734 3570
rect -2544 3515 -2268 3550
rect -1606 3517 -1442 3535
rect -1606 3515 -1492 3517
rect -2544 3422 -2205 3515
rect -2544 3388 -2532 3422
rect -2356 3388 -2205 3422
rect -1606 3405 -1581 3515
rect -1458 3482 -1442 3517
rect -1486 3405 -1442 3482
rect -1606 3400 -1442 3405
rect -1414 3517 -1154 3536
rect -1414 3482 -1203 3517
rect -1169 3482 -1154 3517
rect -1414 3462 -1154 3482
rect -2544 3382 -2344 3388
rect -3544 3244 -3205 3358
rect -2658 3378 -2575 3382
rect -2658 3344 -2625 3378
rect -2591 3344 -2575 3378
rect -2658 3327 -2575 3344
rect -2544 3334 -2344 3341
rect -2544 3300 -2532 3334
rect -2356 3300 -2344 3334
rect -2316 3327 -2205 3388
rect -1414 3393 -1364 3462
rect -1078 3434 -734 3564
rect -1414 3371 -1408 3393
rect -1748 3358 -1408 3371
rect -1374 3358 -1364 3393
rect -1336 3422 -734 3434
rect -1336 3388 -1324 3422
rect -948 3388 -734 3422
rect -1336 3382 -734 3388
rect -703 3550 -574 3584
rect -497 3550 -427 3584
rect 363 3650 1057 3656
rect 363 3570 379 3650
rect 413 3570 571 3650
rect 605 3570 763 3650
rect 797 3598 1057 3650
rect 1091 3598 1107 3824
rect 1138 3838 1144 3868
rect 1223 3868 1356 3872
rect 2252 3874 2326 3921
rect 2566 3874 2589 3921
rect 1223 3838 1229 3868
rect 1138 3680 1229 3838
rect 1138 3646 1144 3680
rect 1223 3646 1229 3680
rect 1138 3630 1229 3646
rect 1261 3776 1414 3840
rect 2252 3814 2589 3874
rect 2975 3872 3197 3920
rect 2975 3868 2985 3872
rect 2865 3824 2948 3840
rect 1261 3742 1267 3776
rect 1344 3742 1414 3776
rect 797 3570 1107 3598
rect 1261 3584 1414 3742
rect 2111 3778 2745 3814
rect 2111 3772 2746 3778
rect 2111 3692 2124 3772
rect 2158 3692 2316 3772
rect 2350 3692 2508 3772
rect 2542 3692 2700 3772
rect 2734 3692 2746 3772
rect 2111 3686 2746 3692
rect 2111 3685 2745 3686
rect 2865 3656 2898 3824
rect 363 3564 1107 3570
rect -703 3515 -427 3550
rect 235 3517 399 3535
rect 235 3515 349 3517
rect -703 3422 -364 3515
rect -703 3388 -691 3422
rect -515 3388 -364 3422
rect 235 3405 260 3515
rect 383 3482 399 3517
rect 355 3405 399 3482
rect 235 3400 399 3405
rect 427 3517 687 3536
rect 427 3482 638 3517
rect 672 3482 687 3517
rect 427 3462 687 3482
rect -703 3382 -503 3388
rect -2544 3299 -2344 3300
rect -2548 3252 -2340 3299
rect -3544 3218 -3506 3244
rect -3542 3066 -3506 3218
rect -3384 3235 -3205 3244
rect -3384 3066 -3354 3235
rect -3177 3230 -2777 3236
rect -3177 3196 -3165 3230
rect -2789 3196 -2777 3230
rect -3177 3155 -2777 3196
rect -3177 3086 -3150 3155
rect -2815 3086 -2777 3155
rect -3177 3067 -2777 3086
rect -1748 3235 -1364 3358
rect -817 3378 -734 3382
rect -817 3344 -784 3378
rect -750 3344 -734 3378
rect -817 3327 -734 3344
rect -703 3334 -503 3341
rect -703 3300 -691 3334
rect -515 3300 -503 3334
rect -475 3327 -364 3388
rect 427 3393 477 3462
rect 763 3434 1107 3564
rect 427 3371 433 3393
rect 100 3358 433 3371
rect 467 3358 477 3393
rect 505 3422 1107 3434
rect 505 3388 517 3422
rect 893 3388 1107 3422
rect 505 3382 1107 3388
rect 1138 3550 1267 3584
rect 1344 3550 1414 3584
rect 2204 3650 2898 3656
rect 2204 3570 2220 3650
rect 2254 3570 2412 3650
rect 2446 3570 2604 3650
rect 2638 3598 2898 3650
rect 2932 3598 2948 3824
rect 2979 3838 2985 3868
rect 3064 3868 3197 3872
rect 3064 3838 3070 3868
rect 2979 3680 3070 3838
rect 2979 3646 2985 3680
rect 3064 3646 3070 3680
rect 2979 3630 3070 3646
rect 3102 3776 3255 3840
rect 3102 3742 3108 3776
rect 3185 3742 3255 3776
rect 2638 3570 2948 3598
rect 3102 3584 3255 3742
rect 2204 3564 2948 3570
rect 1138 3515 1414 3550
rect 2076 3517 2240 3535
rect 2076 3515 2190 3517
rect 1138 3422 1477 3515
rect 1138 3388 1150 3422
rect 1326 3388 1477 3422
rect 2076 3405 2101 3515
rect 2224 3482 2240 3517
rect 2196 3405 2240 3482
rect 2076 3400 2240 3405
rect 2268 3517 2528 3536
rect 2268 3482 2479 3517
rect 2513 3482 2528 3517
rect 2268 3462 2528 3482
rect 1138 3382 1338 3388
rect -703 3299 -503 3300
rect -707 3252 -499 3299
rect -1748 3215 -1549 3235
rect -3542 3044 -3354 3066
rect -1748 3043 -1722 3215
rect -1584 3043 -1549 3215
rect -1336 3230 -936 3236
rect -1336 3196 -1324 3230
rect -948 3196 -936 3230
rect -1336 3155 -936 3196
rect -1336 3086 -1309 3155
rect -974 3086 -936 3155
rect -1336 3067 -936 3086
rect 100 3235 477 3358
rect 1024 3378 1107 3382
rect 1024 3344 1057 3378
rect 1091 3344 1107 3378
rect 1024 3327 1107 3344
rect 1138 3334 1338 3341
rect 1138 3300 1150 3334
rect 1326 3300 1338 3334
rect 1366 3327 1477 3388
rect 2268 3393 2318 3462
rect 2604 3434 2948 3564
rect 2268 3371 2274 3393
rect 2001 3358 2274 3371
rect 2308 3358 2318 3393
rect 2346 3422 2948 3434
rect 2346 3388 2358 3422
rect 2734 3388 2948 3422
rect 2346 3382 2948 3388
rect 2979 3550 3108 3584
rect 3185 3550 3255 3584
rect 2979 3515 3255 3550
rect 2979 3422 3318 3515
rect 2979 3388 2991 3422
rect 3167 3388 3318 3422
rect 2979 3382 3179 3388
rect 2001 3323 2318 3358
rect 2865 3378 2948 3382
rect 2865 3344 2898 3378
rect 2932 3344 2948 3378
rect 2865 3327 2948 3344
rect 2979 3334 3179 3341
rect 1138 3299 1338 3300
rect 1134 3252 1342 3299
rect 1752 3297 2318 3323
rect 2979 3300 2991 3334
rect 3167 3300 3179 3334
rect 3207 3327 3318 3388
rect 2979 3299 3179 3300
rect 100 3189 320 3235
rect 100 3066 127 3189
rect 303 3066 320 3189
rect 505 3230 905 3236
rect 505 3196 517 3230
rect 893 3196 905 3230
rect 505 3155 905 3196
rect 505 3086 532 3155
rect 867 3086 905 3155
rect 1752 3144 1803 3297
rect 2001 3235 2318 3297
rect 2975 3252 3183 3299
rect 2001 3144 2150 3235
rect 1752 3116 2150 3144
rect 2346 3230 2746 3236
rect 2346 3196 2358 3230
rect 2734 3196 2746 3230
rect 2346 3155 2746 3196
rect 505 3067 905 3086
rect 2346 3086 2373 3155
rect 2708 3086 2746 3155
rect 2346 3067 2746 3086
rect 100 3045 320 3066
rect -1748 3013 -1549 3043
rect -3817 2215 -3534 2234
rect -3818 2167 -3534 2215
rect -3818 1894 -3763 2167
rect -3574 1894 -3534 2167
rect -3818 1852 -3534 1894
rect -3818 -4901 -3652 1852
<< via1 >>
rect -3422 3482 -3333 3515
rect -3333 3482 -3327 3515
rect -3422 3405 -3327 3482
rect -1581 3482 -1492 3515
rect -1492 3482 -1486 3515
rect -1581 3405 -1486 3482
rect 260 3482 349 3515
rect 349 3482 355 3515
rect 260 3405 355 3482
rect -3506 3066 -3384 3244
rect 2101 3482 2190 3515
rect 2190 3482 2196 3515
rect 2101 3405 2196 3482
rect -1722 3043 -1584 3215
rect 127 3066 303 3189
rect 1803 3144 2001 3297
rect -3763 1894 -3574 2167
<< metal2 >>
rect -3591 4118 2084 4255
rect -3591 3538 -3448 4118
rect -3591 3515 -3296 3538
rect -1749 3536 -1606 4118
rect 92 3540 235 4118
rect -1749 3515 -1441 3536
rect 92 3515 400 3540
rect 1933 3539 2076 4118
rect 1933 3515 2238 3539
rect -3591 3405 -3422 3515
rect -3327 3405 -3296 3515
rect -3591 3399 -3296 3405
rect -3448 3398 -3296 3399
rect -2251 3511 -2177 3515
rect -2251 3324 -2030 3511
rect -1749 3405 -1581 3515
rect -1486 3405 -1441 3515
rect -1749 3400 -1441 3405
rect -364 3511 -244 3515
rect -364 3327 -135 3511
rect 92 3405 260 3515
rect 355 3405 400 3515
rect 92 3400 400 3405
rect 1477 3510 1516 3515
rect 1477 3327 1600 3510
rect 1933 3405 2101 3515
rect 2196 3405 2238 3515
rect 3453 3514 3608 3518
rect 1933 3400 2238 3405
rect 3318 3327 3608 3514
rect -3542 3244 -3356 3284
rect -3542 3066 -3506 3244
rect -3384 3066 -3356 3244
rect -3542 3048 -3356 3066
rect -2216 2727 -2030 3324
rect -1748 3215 -1558 3247
rect -1748 3043 -1722 3215
rect -1584 3158 -1558 3215
rect -1584 3144 -1412 3158
rect -1584 3043 -1563 3144
rect -1748 3022 -1563 3043
rect -1426 3022 -1412 3144
rect -1748 3013 -1412 3022
rect -275 2833 -135 3327
rect 100 3189 318 3210
rect 100 3066 127 3189
rect 303 3066 318 3189
rect 100 3045 318 3066
rect 1505 2985 1600 3327
rect 1752 3297 2032 3323
rect 1752 3144 1803 3297
rect 2001 3144 2032 3297
rect 1752 3116 2032 3144
rect 3453 3186 3608 3327
rect 3453 3064 13159 3186
rect 3458 3036 13159 3064
rect 1505 2984 10159 2985
rect 1505 2876 10170 2984
rect -1285 2727 -968 2736
rect -2216 2666 -968 2727
rect -285 2722 6879 2833
rect -2216 2614 3582 2666
rect -1285 2553 3582 2614
rect -1285 2544 -968 2553
rect -1869 2517 -1700 2527
rect -1869 2489 -1407 2517
rect -1869 2383 -1556 2489
rect -1432 2383 -1407 2489
rect 3458 2408 3581 2553
rect -1869 2354 -1407 2383
rect 6750 2376 6878 2722
rect 10028 2388 10170 2876
rect -3817 2167 -3534 2234
rect -3817 1894 -3763 2167
rect -3574 1894 -3534 2167
rect -3817 1852 -3534 1894
rect -1869 1632 -1700 2354
rect 10 -200 287 -196
rect 10 -401 315 -200
rect 3275 -213 3407 -128
rect 6574 -187 6881 -83
rect 3275 -343 3638 -213
rect 3342 -344 3638 -343
rect -3604 -447 -299 -427
rect -3604 -453 -471 -447
rect -3604 -593 -3575 -453
rect -3446 -587 -471 -453
rect -342 -587 -299 -447
rect -3446 -593 -299 -587
rect -3604 -614 -299 -593
rect 171 -822 315 -401
rect 3452 -848 3636 -344
rect 6755 -863 6878 -187
rect 9870 -241 9997 -101
rect 10040 -241 10168 -240
rect 9865 -397 10168 -241
rect 9870 -398 9997 -397
rect 10040 -839 10168 -397
rect -11 -3621 314 -3495
rect 3281 -3497 3615 -3375
rect 169 -4142 299 -3621
rect 3456 -4161 3592 -3497
rect 6570 -3532 6886 -3387
rect 9874 -3505 10165 -3369
rect 6744 -4189 6874 -3532
rect 10040 -4161 10164 -3505
<< via2 >>
rect -3506 3066 -3384 3244
rect -1563 3022 -1426 3144
rect 127 3066 303 3189
rect 1803 3144 2001 3297
rect -1556 2383 -1432 2489
rect -3763 1894 -3574 2167
rect -2151 1637 -2020 1751
rect -1818 -210 -1729 236
rect -3575 -593 -3446 -453
rect -471 -587 -342 -447
rect -2154 -1626 -2023 -1512
rect -1822 -3454 -1733 -3008
rect -2148 -4890 -2017 -4776
rect -1825 -6733 -1736 -6287
<< metal3 >>
rect -3817 4255 -3635 4259
rect -3817 4090 1969 4255
rect -3817 2234 -3635 4090
rect -3544 3244 -3354 3372
rect -3544 3218 -3506 3244
rect -3542 3066 -3506 3218
rect -3384 3218 -3354 3244
rect 1752 3323 1969 4090
rect 1752 3297 2032 3323
rect -3384 3066 -3358 3218
rect 100 3189 318 3210
rect -3542 2836 -3358 3066
rect -1583 3144 -1415 3161
rect -1583 3022 -1563 3144
rect -1426 3022 -1415 3144
rect 100 3066 127 3189
rect 303 3066 318 3189
rect 1752 3144 1803 3297
rect 2001 3144 2032 3297
rect 1752 3116 2032 3144
rect 100 3052 318 3066
rect -480 3045 318 3052
rect -480 3033 271 3045
rect -3542 2832 -1710 2836
rect -3542 2636 -1708 2832
rect -3817 2167 -3534 2234
rect -3817 1894 -3763 2167
rect -3574 1894 -3534 2167
rect -3817 1852 -3534 1894
rect -2166 1751 -2007 1796
rect -2166 1637 -2151 1751
rect -2020 1637 -2007 1751
rect -3607 -453 -3416 332
rect -3607 -593 -3575 -453
rect -3446 -593 -3416 -453
rect -3607 -6772 -3416 -593
rect -2166 -1512 -2007 1637
rect -2166 -1626 -2154 -1512
rect -2023 -1626 -2007 -1512
rect -2166 -4776 -2007 -1626
rect -2166 -4890 -2148 -4776
rect -2017 -4890 -2007 -4776
rect -2166 -4901 -2007 -4890
rect -1893 236 -1708 2636
rect -1583 2489 -1415 3022
rect -1583 2383 -1556 2489
rect -1432 2383 -1415 2489
rect -1583 2362 -1415 2383
rect -481 2868 271 3033
rect -481 2858 265 2868
rect -1893 -210 -1818 236
rect -1729 -210 -1708 236
rect -1893 -3008 -1708 -210
rect -481 -447 -301 2858
rect -481 -587 -471 -447
rect -342 -587 -301 -447
rect -481 -623 -301 -587
rect -1893 -3454 -1822 -3008
rect -1733 -3454 -1708 -3008
rect -1893 -6287 -1708 -3454
rect -1893 -6733 -1825 -6287
rect -1736 -6733 -1708 -6287
rect -1893 -6782 -1708 -6733
use 4bit_ADDER  4bit_ADDER_0
timestamp 1736273553
transform 1 0 171 0 1 -165
box -3989 -146 13189 3089
use 4bit_ADDER  4bit_ADDER_1
timestamp 1736273553
transform 1 0 171 0 1 -3430
box -3989 -146 13189 3089
use 4bit_ADDER  4bit_ADDER_2
timestamp 1736273553
transform 1 0 171 0 1 -6694
box -3989 -146 13189 3089
<< labels >>
rlabel metal1 -2443 3252 -2443 3252 5 VSS
port 4 s
rlabel metal1 -2500 3920 -2500 3920 1 VDD
port 1 n
rlabel metal1 -2644 3471 -2644 3471 7 A
port 2 e
rlabel metal1 -2268 3471 -2268 3471 3 Y
port 3 e
rlabel metal1 -602 3252 -602 3252 5 VSS
port 4 s
rlabel metal1 -659 3920 -659 3920 1 VDD
port 1 n
rlabel metal1 -803 3471 -803 3471 7 A
port 2 e
rlabel metal1 -427 3471 -427 3471 3 Y
port 3 e
rlabel metal1 1239 3252 1239 3252 5 VSS
port 4 s
rlabel metal1 1182 3920 1182 3920 1 VDD
port 1 n
rlabel metal1 1038 3471 1038 3471 7 A
port 2 e
rlabel metal1 1414 3471 1414 3471 3 Y
port 3 e
rlabel metal1 3080 3252 3080 3252 5 VSS
port 4 s
rlabel metal1 3023 3920 3023 3920 1 VDD
port 1 n
rlabel metal1 2879 3471 2879 3471 7 A
port 2 e
rlabel metal1 3255 3471 3255 3471 3 Y
port 3 e
flabel metal2 -3556 1080 -3436 1200 1 FreeSerif 160 0 0 0 B1
port 5 n
flabel metal1 -3794 1646 -3674 1766 1 FreeSerif 160 0 0 0 A0
port 6 n
flabel metal2 -3228 -2190 -3108 -2070 1 FreeSerif 160 0 0 0 B2
port 7 n
flabel metal2 -3584 3886 -3464 4006 1 FreeSerif 160 0 0 0 B0
port 8 n
flabel metal2 -3220 -5452 -3100 -5332 1 FreeSerif 160 0 0 0 B3
port 9 n
flabel metal3 -2146 -202 -2026 -82 1 FreeSerif 160 0 0 0 A2
port 10 n
flabel metal2 -2952 -576 -2832 -456 1 FreeSerif 160 0 0 0 A1
port 11 n
flabel metal3 -3190 2678 -3070 2798 1 FreeSerif 160 0 0 0 A3
port 12 n
flabel metal2 12820 3054 12940 3174 1 FreeSerif 160 0 0 0 SO
port 13 n
flabel metal2 13166 -32 13262 54 1 FreeSerif 160 0 0 0 S1
port 14 n
flabel metal2 13182 -3394 13278 -3308 1 FreeSerif 160 0 0 0 S2
port 15 n
flabel metal2 6586 -6668 6682 -6582 1 FreeSerif 160 0 0 0 S5
port 16 n
flabel metal2 9878 -6670 9974 -6584 1 FreeSerif 160 0 0 0 S4
port 17 n
flabel metal2 13182 -6664 13278 -6578 1 FreeSerif 160 0 0 0 S3
port 18 n
flabel metal2 54 -6728 150 -6642 1 FreeSerif 160 0 0 0 S7
port 19 n
flabel metal2 3294 -6664 3390 -6578 1 FreeSerif 160 0 0 0 S6
port 20 n
<< end >>
