magic
tech sky130B
magscale 1 2
timestamp 1736704482
<< nwell >>
rect 1671 6310 4735 6311
rect 1671 5410 6439 6310
rect 4981 5409 6439 5410
rect 6903 5575 7933 5597
rect 6903 5165 8121 5575
rect 7641 5164 8121 5165
rect 7709 5089 8121 5164
rect -24166 3687 -22708 4587
rect -20875 3687 -19417 4587
rect -17584 3687 -16126 4587
rect -14293 3687 -12835 4587
rect -11002 3687 -9544 4587
rect -7712 3687 -6254 4587
rect -4421 3687 -2963 4587
rect -1130 3687 328 4587
rect 5557 3541 6850 4027
rect 7893 3373 10816 3374
rect 7893 3372 10870 3373
rect 7102 2835 11742 3372
rect -25114 1903 1213 2814
rect 7102 2797 11646 2835
rect 11737 2009 12827 2230
rect 11737 1653 13235 2009
rect 12823 1523 13235 1653
rect -25114 599 1213 1119
rect 7102 455 10816 456
rect 7102 417 11646 455
rect 7102 -120 11742 417
rect 5557 -987 6850 -501
rect 7893 -1155 10816 -1154
rect 7893 -1156 10870 -1155
rect 7102 -1693 11742 -1156
rect 7102 -1731 11646 -1693
rect -24483 -2203 -17802 -2161
rect -24483 -2689 -17776 -2203
rect 11737 -2519 12827 -2298
rect 11737 -2875 13235 -2519
rect 12823 -3005 13235 -2875
rect -24432 -4501 -23250 -3943
rect -22696 -4015 -21568 -3959
rect -22696 -4501 -21534 -4015
rect -21047 -4657 -7883 -3746
rect 7102 -4073 10816 -4072
rect 7102 -4111 11646 -4073
rect 7102 -4648 11742 -4111
rect -24432 -5307 -23304 -5251
rect -22696 -5307 -21568 -5251
rect -24432 -5793 -23274 -5307
rect -22696 -5793 -21540 -5307
rect 5557 -5415 6850 -4929
rect -21047 -5961 -7883 -5441
rect 7893 -5583 10816 -5582
rect 7893 -5584 10870 -5583
rect 7102 -6121 11742 -5584
rect 7102 -6159 11646 -6121
rect 11737 -6947 12827 -6726
rect -24432 -7280 -23304 -7224
rect -22695 -7280 -21567 -7224
rect -24432 -7766 -23272 -7280
rect -22695 -7766 -21538 -7280
rect -21047 -7922 -7883 -7011
rect 11737 -7303 13235 -6947
rect 12823 -7433 13235 -7303
rect 7102 -8501 10816 -8500
rect -24432 -8572 -23304 -8516
rect -22696 -8572 -21568 -8516
rect 7102 -8539 11646 -8501
rect -24432 -9058 -23271 -8572
rect -22696 -9058 -21534 -8572
rect -21047 -9226 -7883 -8706
rect 7102 -9076 11742 -8539
rect 5557 -10043 6850 -9557
rect 7893 -10211 10816 -10210
rect 7893 -10212 10870 -10211
rect -24432 -10544 -23304 -10488
rect -22695 -10544 -21567 -10488
rect -24432 -11030 -23271 -10544
rect -22695 -11030 -21538 -10544
rect -21047 -11186 -7883 -10275
rect 7102 -10749 11742 -10212
rect 7102 -10787 11646 -10749
rect 11737 -11575 12827 -11354
rect -24432 -11836 -23304 -11780
rect -22695 -11836 -21567 -11780
rect -24432 -12322 -23271 -11836
rect -22695 -12322 -21542 -11836
rect 11737 -11931 13235 -11575
rect -21047 -12490 -7883 -11970
rect 12823 -12061 13235 -11931
rect 7102 -13129 10816 -13128
rect 7102 -13167 11646 -13129
rect 7102 -13704 11742 -13167
rect -24605 -15384 -24173 -14880
rect -24605 -16065 -24172 -15384
rect -17898 -15553 -17321 -14463
rect -24604 -16569 -24172 -16065
rect -24604 -17278 -24167 -16569
rect -17898 -16953 -17321 -15863
rect -12543 -16873 -11643 -14057
rect -8339 -15748 -7797 -15248
rect -8339 -16160 -7796 -15748
rect -24599 -17782 -24167 -17278
rect -24599 -18397 -24152 -17782
rect -24584 -18901 -24152 -18397
rect -21778 -18436 -21236 -17936
rect -17898 -18353 -17321 -17263
rect -16187 -18307 -15645 -17807
rect -21778 -18848 -21235 -18436
rect -24584 -19591 -24150 -18901
rect -24582 -20095 -24150 -19591
rect -24582 -20791 -24119 -20095
rect -24551 -21295 -24119 -20791
rect -21778 -20768 -21236 -18848
rect -17898 -19753 -17321 -18663
rect -16187 -18719 -15644 -18307
rect -12543 -18331 -11641 -16873
rect -8339 -18080 -7797 -16160
rect -21778 -21171 -21250 -20768
rect -17898 -21153 -17321 -20063
rect -16187 -20639 -15645 -18719
rect -12543 -19830 -11643 -18331
rect -8339 -18483 -7811 -18080
rect -8339 -19020 -7809 -18483
rect -16187 -21042 -15659 -20639
rect -24551 -22072 -24118 -21295
rect -21778 -21708 -21248 -21171
rect -24551 -22094 -24120 -22072
rect -24552 -24109 -24120 -22094
rect -17898 -22553 -17321 -21463
rect -16187 -21579 -15657 -21042
rect -12543 -21288 -11641 -19830
rect -4932 -21067 -4446 -14103
rect -2216 -20684 -1730 -13720
rect 5557 -14571 6850 -14085
rect 7893 -14739 10816 -14738
rect 7893 -14740 10870 -14739
rect 7102 -15277 11742 -14740
rect 7102 -15315 11646 -15277
rect 11737 -16103 12827 -15882
rect 11737 -16459 13235 -16103
rect 12823 -16589 13235 -16459
rect 7102 -17657 10816 -17656
rect 7102 -17695 11646 -17657
rect 7102 -18232 11742 -17695
rect 15617 -18119 17009 -17611
rect 15617 -18120 17964 -18119
rect 15617 -18551 18408 -18120
rect 5557 -19099 6850 -18613
rect 7893 -19267 10816 -19266
rect 7893 -19268 10870 -19267
rect 7102 -19805 11742 -19268
rect 15617 -19561 17009 -18551
rect 17996 -18629 18408 -18551
rect 7102 -19843 11646 -19805
rect 11737 -20631 12827 -20410
rect 11737 -20987 13235 -20631
rect 12823 -21117 13235 -20987
rect -12543 -22409 -11643 -21288
rect 7102 -22185 10816 -22184
rect 7102 -22223 11646 -22185
rect -17898 -23953 -17321 -22863
rect -12543 -23867 -11641 -22409
rect 7102 -22760 11742 -22223
rect 5557 -23627 6850 -23141
rect 7893 -23795 10816 -23794
rect 7893 -23796 10870 -23795
rect -17898 -25353 -17321 -24263
rect -12543 -25177 -11643 -23867
rect 7102 -24333 11742 -23796
rect 7102 -24371 11646 -24333
rect 11737 -25159 12827 -24938
rect -12543 -26635 -11641 -25177
rect 11737 -25515 13235 -25159
rect 12823 -25645 13235 -25515
rect -12543 -27810 -11643 -26635
rect 7102 -26713 10816 -26712
rect 7102 -26751 11646 -26713
rect 7102 -27288 11742 -26751
rect -12543 -29268 -11641 -27810
rect 5557 -28155 6850 -27669
rect 7893 -28323 10816 -28322
rect 7893 -28324 10870 -28323
rect 7102 -28861 11742 -28324
rect 7102 -28899 11646 -28861
rect -12543 -30419 -11643 -29268
rect 11737 -29687 12827 -29466
rect 11737 -30043 13235 -29687
rect 12823 -30173 13235 -30043
rect -12543 -31877 -11641 -30419
rect 7102 -31241 10816 -31240
rect 7102 -31279 11646 -31241
rect 7102 -31816 11742 -31279
rect -12543 -34497 -11643 -31877
rect 5557 -32683 6850 -32197
rect 7893 -32851 10816 -32850
rect 7893 -32852 10870 -32851
rect 7102 -33389 11742 -32852
rect 7102 -33427 11646 -33389
rect 11737 -34215 12827 -33994
rect 11737 -34571 13235 -34215
rect 12823 -34701 13235 -34571
rect 7102 -35769 10816 -35768
rect 7102 -35807 11646 -35769
rect 7102 -36344 11742 -35807
rect 13088 -36406 13574 -35615
<< nmos >>
rect 1765 4914 1795 5044
rect 1857 4914 1887 5044
rect 1953 4914 1983 5044
rect 2049 4914 2079 5044
rect 2145 4914 2175 5044
rect 2241 4914 2271 5044
rect 2337 4914 2367 5044
rect 2433 4914 2463 5044
rect 2529 4914 2559 5044
rect 2625 4914 2655 5044
rect 2721 4914 2751 5044
rect 2817 4914 2847 5044
rect 2913 4914 2943 5044
rect 3005 4914 3035 5044
rect 3371 4914 3401 5044
rect 3463 4914 3493 5044
rect 3559 4914 3589 5044
rect 3655 4914 3685 5044
rect 3751 4914 3781 5044
rect 3847 4914 3877 5044
rect 3943 4914 3973 5044
rect 4039 4914 4069 5044
rect 4135 4914 4165 5044
rect 4231 4914 4261 5044
rect 4327 4914 4357 5044
rect 4423 4914 4453 5044
rect 4519 4914 4549 5044
rect 4611 4914 4641 5044
rect 5075 4912 5105 5042
rect 5167 4912 5197 5042
rect 5263 4912 5293 5042
rect 5359 4912 5389 5042
rect 5455 4912 5485 5042
rect 5551 4912 5581 5042
rect 5647 4912 5677 5042
rect 5743 4912 5773 5042
rect 5839 4912 5869 5042
rect 5935 4912 5965 5042
rect 6031 4912 6061 5042
rect 6127 4912 6157 5042
rect 6223 4912 6253 5042
rect 6315 4912 6345 5042
rect 7173 5005 7573 5035
rect 7173 4909 7573 4939
rect 7809 4933 8009 4963
rect 5658 3385 5858 3415
rect 6098 3385 6298 3415
rect 6538 3385 6738 3415
rect -24072 3190 -24042 3320
rect -23980 3190 -23950 3320
rect -23884 3190 -23854 3320
rect -23788 3190 -23758 3320
rect -23692 3190 -23662 3320
rect -23596 3190 -23566 3320
rect -23500 3190 -23470 3320
rect -23404 3190 -23374 3320
rect -23308 3190 -23278 3320
rect -23212 3190 -23182 3320
rect -23116 3190 -23086 3320
rect -23020 3190 -22990 3320
rect -22924 3190 -22894 3320
rect -22832 3190 -22802 3320
rect -20781 3190 -20751 3320
rect -20689 3190 -20659 3320
rect -20593 3190 -20563 3320
rect -20497 3190 -20467 3320
rect -20401 3190 -20371 3320
rect -20305 3190 -20275 3320
rect -20209 3190 -20179 3320
rect -20113 3190 -20083 3320
rect -20017 3190 -19987 3320
rect -19921 3190 -19891 3320
rect -19825 3190 -19795 3320
rect -19729 3190 -19699 3320
rect -19633 3190 -19603 3320
rect -19541 3190 -19511 3320
rect -17490 3190 -17460 3320
rect -17398 3190 -17368 3320
rect -17302 3190 -17272 3320
rect -17206 3190 -17176 3320
rect -17110 3190 -17080 3320
rect -17014 3190 -16984 3320
rect -16918 3190 -16888 3320
rect -16822 3190 -16792 3320
rect -16726 3190 -16696 3320
rect -16630 3190 -16600 3320
rect -16534 3190 -16504 3320
rect -16438 3190 -16408 3320
rect -16342 3190 -16312 3320
rect -16250 3190 -16220 3320
rect -14199 3190 -14169 3320
rect -14107 3190 -14077 3320
rect -14011 3190 -13981 3320
rect -13915 3190 -13885 3320
rect -13819 3190 -13789 3320
rect -13723 3190 -13693 3320
rect -13627 3190 -13597 3320
rect -13531 3190 -13501 3320
rect -13435 3190 -13405 3320
rect -13339 3190 -13309 3320
rect -13243 3190 -13213 3320
rect -13147 3190 -13117 3320
rect -13051 3190 -13021 3320
rect -12959 3190 -12929 3320
rect -10908 3190 -10878 3320
rect -10816 3190 -10786 3320
rect -10720 3190 -10690 3320
rect -10624 3190 -10594 3320
rect -10528 3190 -10498 3320
rect -10432 3190 -10402 3320
rect -10336 3190 -10306 3320
rect -10240 3190 -10210 3320
rect -10144 3190 -10114 3320
rect -10048 3190 -10018 3320
rect -9952 3190 -9922 3320
rect -9856 3190 -9826 3320
rect -9760 3190 -9730 3320
rect -9668 3190 -9638 3320
rect -7618 3190 -7588 3320
rect -7526 3190 -7496 3320
rect -7430 3190 -7400 3320
rect -7334 3190 -7304 3320
rect -7238 3190 -7208 3320
rect -7142 3190 -7112 3320
rect -7046 3190 -7016 3320
rect -6950 3190 -6920 3320
rect -6854 3190 -6824 3320
rect -6758 3190 -6728 3320
rect -6662 3190 -6632 3320
rect -6566 3190 -6536 3320
rect -6470 3190 -6440 3320
rect -6378 3190 -6348 3320
rect -4327 3190 -4297 3320
rect -4235 3190 -4205 3320
rect -4139 3190 -4109 3320
rect -4043 3190 -4013 3320
rect -3947 3190 -3917 3320
rect -3851 3190 -3821 3320
rect -3755 3190 -3725 3320
rect -3659 3190 -3629 3320
rect -3563 3190 -3533 3320
rect -3467 3190 -3437 3320
rect -3371 3190 -3341 3320
rect -3275 3190 -3245 3320
rect -3179 3190 -3149 3320
rect -3087 3190 -3057 3320
rect -1036 3190 -1006 3320
rect -944 3190 -914 3320
rect -848 3190 -818 3320
rect -752 3190 -722 3320
rect -656 3190 -626 3320
rect -560 3190 -530 3320
rect -464 3190 -434 3320
rect -368 3190 -338 3320
rect -272 3190 -242 3320
rect -176 3190 -146 3320
rect -80 3190 -50 3320
rect 16 3190 46 3320
rect 112 3190 142 3320
rect 204 3190 234 3320
rect 7422 1690 7452 2490
rect 7518 1690 7548 2490
rect 7614 1690 7644 2490
rect 7710 1690 7740 2490
rect 8370 1690 8400 2490
rect 8466 1690 8496 2490
rect 8562 1690 8592 2490
rect 8658 1690 8688 2490
rect 9306 1690 9336 2490
rect 9402 1690 9432 2490
rect 9498 1690 9528 2490
rect 9594 1690 9624 2490
rect 10237 1690 10267 2490
rect 10333 1690 10363 2490
rect 10429 1690 10459 2490
rect 10525 1690 10555 2490
rect 11164 1690 11194 2490
rect 11260 1690 11290 2490
rect 11356 1690 11386 2490
rect 11452 1690 11482 2490
rect -24746 1406 -24716 1536
rect -24654 1406 -24624 1536
rect -24558 1406 -24528 1536
rect -24462 1406 -24432 1536
rect -24366 1406 -24336 1536
rect -24270 1406 -24240 1536
rect -24174 1406 -24144 1536
rect -24078 1406 -24048 1536
rect -23982 1406 -23952 1536
rect -23886 1406 -23856 1536
rect -23790 1406 -23760 1536
rect -23694 1406 -23664 1536
rect -23598 1406 -23568 1536
rect -23506 1406 -23476 1536
rect -23187 1406 -23157 1536
rect -23095 1406 -23065 1536
rect -22999 1406 -22969 1536
rect -22903 1406 -22873 1536
rect -22807 1406 -22777 1536
rect -22711 1406 -22681 1536
rect -22615 1406 -22585 1536
rect -22519 1406 -22489 1536
rect -22423 1406 -22393 1536
rect -22327 1406 -22297 1536
rect -22231 1406 -22201 1536
rect -22135 1406 -22105 1536
rect -22039 1406 -22009 1536
rect -21947 1406 -21917 1536
rect -21455 1406 -21425 1536
rect -21363 1406 -21333 1536
rect -21267 1406 -21237 1536
rect -21171 1406 -21141 1536
rect -21075 1406 -21045 1536
rect -20979 1406 -20949 1536
rect -20883 1406 -20853 1536
rect -20787 1406 -20757 1536
rect -20691 1406 -20661 1536
rect -20595 1406 -20565 1536
rect -20499 1406 -20469 1536
rect -20403 1406 -20373 1536
rect -20307 1406 -20277 1536
rect -20215 1406 -20185 1536
rect -19896 1406 -19866 1536
rect -19804 1406 -19774 1536
rect -19708 1406 -19678 1536
rect -19612 1406 -19582 1536
rect -19516 1406 -19486 1536
rect -19420 1406 -19390 1536
rect -19324 1406 -19294 1536
rect -19228 1406 -19198 1536
rect -19132 1406 -19102 1536
rect -19036 1406 -19006 1536
rect -18940 1406 -18910 1536
rect -18844 1406 -18814 1536
rect -18748 1406 -18718 1536
rect -18656 1406 -18626 1536
rect -18164 1406 -18134 1536
rect -18072 1406 -18042 1536
rect -17976 1406 -17946 1536
rect -17880 1406 -17850 1536
rect -17784 1406 -17754 1536
rect -17688 1406 -17658 1536
rect -17592 1406 -17562 1536
rect -17496 1406 -17466 1536
rect -17400 1406 -17370 1536
rect -17304 1406 -17274 1536
rect -17208 1406 -17178 1536
rect -17112 1406 -17082 1536
rect -17016 1406 -16986 1536
rect -16924 1406 -16894 1536
rect -16605 1406 -16575 1536
rect -16513 1406 -16483 1536
rect -16417 1406 -16387 1536
rect -16321 1406 -16291 1536
rect -16225 1406 -16195 1536
rect -16129 1406 -16099 1536
rect -16033 1406 -16003 1536
rect -15937 1406 -15907 1536
rect -15841 1406 -15811 1536
rect -15745 1406 -15715 1536
rect -15649 1406 -15619 1536
rect -15553 1406 -15523 1536
rect -15457 1406 -15427 1536
rect -15365 1406 -15335 1536
rect -14873 1406 -14843 1536
rect -14781 1406 -14751 1536
rect -14685 1406 -14655 1536
rect -14589 1406 -14559 1536
rect -14493 1406 -14463 1536
rect -14397 1406 -14367 1536
rect -14301 1406 -14271 1536
rect -14205 1406 -14175 1536
rect -14109 1406 -14079 1536
rect -14013 1406 -13983 1536
rect -13917 1406 -13887 1536
rect -13821 1406 -13791 1536
rect -13725 1406 -13695 1536
rect -13633 1406 -13603 1536
rect -13314 1406 -13284 1536
rect -13222 1406 -13192 1536
rect -13126 1406 -13096 1536
rect -13030 1406 -13000 1536
rect -12934 1406 -12904 1536
rect -12838 1406 -12808 1536
rect -12742 1406 -12712 1536
rect -12646 1406 -12616 1536
rect -12550 1406 -12520 1536
rect -12454 1406 -12424 1536
rect -12358 1406 -12328 1536
rect -12262 1406 -12232 1536
rect -12166 1406 -12136 1536
rect -12074 1406 -12044 1536
rect -11582 1406 -11552 1536
rect -11490 1406 -11460 1536
rect -11394 1406 -11364 1536
rect -11298 1406 -11268 1536
rect -11202 1406 -11172 1536
rect -11106 1406 -11076 1536
rect -11010 1406 -10980 1536
rect -10914 1406 -10884 1536
rect -10818 1406 -10788 1536
rect -10722 1406 -10692 1536
rect -10626 1406 -10596 1536
rect -10530 1406 -10500 1536
rect -10434 1406 -10404 1536
rect -10342 1406 -10312 1536
rect -10023 1406 -9993 1536
rect -9931 1406 -9901 1536
rect -9835 1406 -9805 1536
rect -9739 1406 -9709 1536
rect -9643 1406 -9613 1536
rect -9547 1406 -9517 1536
rect -9451 1406 -9421 1536
rect -9355 1406 -9325 1536
rect -9259 1406 -9229 1536
rect -9163 1406 -9133 1536
rect -9067 1406 -9037 1536
rect -8971 1406 -8941 1536
rect -8875 1406 -8845 1536
rect -8783 1406 -8753 1536
rect -8292 1406 -8262 1536
rect -8200 1406 -8170 1536
rect -8104 1406 -8074 1536
rect -8008 1406 -7978 1536
rect -7912 1406 -7882 1536
rect -7816 1406 -7786 1536
rect -7720 1406 -7690 1536
rect -7624 1406 -7594 1536
rect -7528 1406 -7498 1536
rect -7432 1406 -7402 1536
rect -7336 1406 -7306 1536
rect -7240 1406 -7210 1536
rect -7144 1406 -7114 1536
rect -7052 1406 -7022 1536
rect -6733 1406 -6703 1536
rect -6641 1406 -6611 1536
rect -6545 1406 -6515 1536
rect -6449 1406 -6419 1536
rect -6353 1406 -6323 1536
rect -6257 1406 -6227 1536
rect -6161 1406 -6131 1536
rect -6065 1406 -6035 1536
rect -5969 1406 -5939 1536
rect -5873 1406 -5843 1536
rect -5777 1406 -5747 1536
rect -5681 1406 -5651 1536
rect -5585 1406 -5555 1536
rect -5493 1406 -5463 1536
rect -5001 1406 -4971 1536
rect -4909 1406 -4879 1536
rect -4813 1406 -4783 1536
rect -4717 1406 -4687 1536
rect -4621 1406 -4591 1536
rect -4525 1406 -4495 1536
rect -4429 1406 -4399 1536
rect -4333 1406 -4303 1536
rect -4237 1406 -4207 1536
rect -4141 1406 -4111 1536
rect -4045 1406 -4015 1536
rect -3949 1406 -3919 1536
rect -3853 1406 -3823 1536
rect -3761 1406 -3731 1536
rect -3442 1406 -3412 1536
rect -3350 1406 -3320 1536
rect -3254 1406 -3224 1536
rect -3158 1406 -3128 1536
rect -3062 1406 -3032 1536
rect -2966 1406 -2936 1536
rect -2870 1406 -2840 1536
rect -2774 1406 -2744 1536
rect -2678 1406 -2648 1536
rect -2582 1406 -2552 1536
rect -2486 1406 -2456 1536
rect -2390 1406 -2360 1536
rect -2294 1406 -2264 1536
rect -2202 1406 -2172 1536
rect -1710 1406 -1680 1536
rect -1618 1406 -1588 1536
rect -1522 1406 -1492 1536
rect -1426 1406 -1396 1536
rect -1330 1406 -1300 1536
rect -1234 1406 -1204 1536
rect -1138 1406 -1108 1536
rect -1042 1406 -1012 1536
rect -946 1406 -916 1536
rect -850 1406 -820 1536
rect -754 1406 -724 1536
rect -658 1406 -628 1536
rect -562 1406 -532 1536
rect -470 1406 -440 1536
rect -151 1406 -121 1536
rect -59 1406 -29 1536
rect 37 1406 67 1536
rect 133 1406 163 1536
rect 229 1406 259 1536
rect 325 1406 355 1536
rect 421 1406 451 1536
rect 517 1406 547 1536
rect 613 1406 643 1536
rect 709 1406 739 1536
rect 805 1406 835 1536
rect 901 1406 931 1536
rect 997 1406 1027 1536
rect 1089 1406 1119 1536
rect 7422 762 7452 1562
rect 7518 762 7548 1562
rect 7614 762 7644 1562
rect 7710 762 7740 1562
rect 8370 762 8400 1562
rect 8466 762 8496 1562
rect 8562 762 8592 1562
rect 8658 762 8688 1562
rect 9306 762 9336 1562
rect 9402 762 9432 1562
rect 9498 762 9528 1562
rect 9594 762 9624 1562
rect 10237 763 10267 1563
rect 10333 763 10363 1563
rect 10429 763 10459 1563
rect 10525 763 10555 1563
rect -24363 439 -23963 469
rect -23254 439 -22854 469
rect -22372 439 -21972 469
rect -21072 439 -20672 469
rect -19963 439 -19563 469
rect -19081 439 -18681 469
rect -17781 439 -17381 469
rect -16672 439 -16272 469
rect -15790 439 -15390 469
rect -14490 439 -14090 469
rect -13381 439 -12981 469
rect -12499 439 -12099 469
rect -11199 439 -10799 469
rect -10090 439 -9690 469
rect -9208 439 -8808 469
rect -7909 439 -7509 469
rect -6800 439 -6400 469
rect -5918 439 -5518 469
rect -4618 439 -4218 469
rect -3509 439 -3109 469
rect -2627 439 -2227 469
rect -1327 439 -927 469
rect -218 439 182 469
rect 664 439 1064 469
rect 11164 762 11194 1562
rect 11260 762 11290 1562
rect 11356 762 11386 1562
rect 11452 762 11482 1562
rect 12219 1320 12249 1520
rect 12315 1320 12345 1520
rect 12923 1367 13123 1397
rect -24363 343 -23963 373
rect -23254 343 -22854 373
rect -22372 343 -21972 373
rect -21072 343 -20672 373
rect -19963 343 -19563 373
rect -19081 343 -18681 373
rect -17781 343 -17381 373
rect -16672 343 -16272 373
rect -15790 343 -15390 373
rect -14490 343 -14090 373
rect -13381 343 -12981 373
rect -12499 343 -12099 373
rect -11199 343 -10799 373
rect -10090 343 -9690 373
rect -9208 343 -8808 373
rect -7909 343 -7509 373
rect -6800 343 -6400 373
rect -5918 343 -5518 373
rect -4618 343 -4218 373
rect -3509 343 -3109 373
rect -2627 343 -2227 373
rect -1327 343 -927 373
rect -218 343 182 373
rect 664 343 1064 373
rect 5658 -1143 5858 -1113
rect 6098 -1143 6298 -1113
rect 6538 -1143 6738 -1113
rect -24213 -2849 -23813 -2819
rect -23628 -2845 -23428 -2815
rect -22176 -2849 -21776 -2819
rect -21608 -2845 -21408 -2815
rect -20446 -2849 -20046 -2819
rect -19867 -2845 -19667 -2815
rect -18686 -2849 -18286 -2819
rect -18088 -2845 -17888 -2815
rect 7422 -2838 7452 -2038
rect 7518 -2838 7548 -2038
rect 7614 -2838 7644 -2038
rect 7710 -2838 7740 -2038
rect 8370 -2838 8400 -2038
rect 8466 -2838 8496 -2038
rect 8562 -2838 8592 -2038
rect 8658 -2838 8688 -2038
rect 9306 -2838 9336 -2038
rect 9402 -2838 9432 -2038
rect 9498 -2838 9528 -2038
rect 9594 -2838 9624 -2038
rect 10237 -2838 10267 -2038
rect 10333 -2838 10363 -2038
rect 10429 -2838 10459 -2038
rect 10525 -2838 10555 -2038
rect 11164 -2838 11194 -2038
rect 11260 -2838 11290 -2038
rect 11356 -2838 11386 -2038
rect 11452 -2838 11482 -2038
rect -24213 -2945 -23813 -2915
rect -22176 -2945 -21776 -2915
rect -20446 -2945 -20046 -2915
rect -18686 -2945 -18286 -2915
rect 7422 -3766 7452 -2966
rect 7518 -3766 7548 -2966
rect 7614 -3766 7644 -2966
rect 7710 -3766 7740 -2966
rect 8370 -3766 8400 -2966
rect 8466 -3766 8496 -2966
rect 8562 -3766 8592 -2966
rect 8658 -3766 8688 -2966
rect 9306 -3766 9336 -2966
rect 9402 -3766 9432 -2966
rect 9498 -3766 9528 -2966
rect 9594 -3766 9624 -2966
rect 10237 -3765 10267 -2965
rect 10333 -3765 10363 -2965
rect 10429 -3765 10459 -2965
rect 10525 -3765 10555 -2965
rect -24162 -4661 -23762 -4631
rect -23584 -4657 -23384 -4627
rect 11164 -3766 11194 -2966
rect 11260 -3766 11290 -2966
rect 11356 -3766 11386 -2966
rect 11452 -3766 11482 -2966
rect 12219 -3208 12249 -3008
rect 12315 -3208 12345 -3008
rect 12923 -3161 13123 -3131
rect -22426 -4661 -22026 -4631
rect -21846 -4657 -21646 -4627
rect -24162 -4757 -23762 -4727
rect -22426 -4757 -22026 -4727
rect -20679 -5154 -20649 -5024
rect -20587 -5154 -20557 -5024
rect -20491 -5154 -20461 -5024
rect -20395 -5154 -20365 -5024
rect -20299 -5154 -20269 -5024
rect -20203 -5154 -20173 -5024
rect -20107 -5154 -20077 -5024
rect -20011 -5154 -19981 -5024
rect -19915 -5154 -19885 -5024
rect -19819 -5154 -19789 -5024
rect -19723 -5154 -19693 -5024
rect -19627 -5154 -19597 -5024
rect -19531 -5154 -19501 -5024
rect -19439 -5154 -19409 -5024
rect -19120 -5154 -19090 -5024
rect -19028 -5154 -18998 -5024
rect -18932 -5154 -18902 -5024
rect -18836 -5154 -18806 -5024
rect -18740 -5154 -18710 -5024
rect -18644 -5154 -18614 -5024
rect -18548 -5154 -18518 -5024
rect -18452 -5154 -18422 -5024
rect -18356 -5154 -18326 -5024
rect -18260 -5154 -18230 -5024
rect -18164 -5154 -18134 -5024
rect -18068 -5154 -18038 -5024
rect -17972 -5154 -17942 -5024
rect -17880 -5154 -17850 -5024
rect -17388 -5154 -17358 -5024
rect -17296 -5154 -17266 -5024
rect -17200 -5154 -17170 -5024
rect -17104 -5154 -17074 -5024
rect -17008 -5154 -16978 -5024
rect -16912 -5154 -16882 -5024
rect -16816 -5154 -16786 -5024
rect -16720 -5154 -16690 -5024
rect -16624 -5154 -16594 -5024
rect -16528 -5154 -16498 -5024
rect -16432 -5154 -16402 -5024
rect -16336 -5154 -16306 -5024
rect -16240 -5154 -16210 -5024
rect -16148 -5154 -16118 -5024
rect -15829 -5154 -15799 -5024
rect -15737 -5154 -15707 -5024
rect -15641 -5154 -15611 -5024
rect -15545 -5154 -15515 -5024
rect -15449 -5154 -15419 -5024
rect -15353 -5154 -15323 -5024
rect -15257 -5154 -15227 -5024
rect -15161 -5154 -15131 -5024
rect -15065 -5154 -15035 -5024
rect -14969 -5154 -14939 -5024
rect -14873 -5154 -14843 -5024
rect -14777 -5154 -14747 -5024
rect -14681 -5154 -14651 -5024
rect -14589 -5154 -14559 -5024
rect -14097 -5154 -14067 -5024
rect -14005 -5154 -13975 -5024
rect -13909 -5154 -13879 -5024
rect -13813 -5154 -13783 -5024
rect -13717 -5154 -13687 -5024
rect -13621 -5154 -13591 -5024
rect -13525 -5154 -13495 -5024
rect -13429 -5154 -13399 -5024
rect -13333 -5154 -13303 -5024
rect -13237 -5154 -13207 -5024
rect -13141 -5154 -13111 -5024
rect -13045 -5154 -13015 -5024
rect -12949 -5154 -12919 -5024
rect -12857 -5154 -12827 -5024
rect -12538 -5154 -12508 -5024
rect -12446 -5154 -12416 -5024
rect -12350 -5154 -12320 -5024
rect -12254 -5154 -12224 -5024
rect -12158 -5154 -12128 -5024
rect -12062 -5154 -12032 -5024
rect -11966 -5154 -11936 -5024
rect -11870 -5154 -11840 -5024
rect -11774 -5154 -11744 -5024
rect -11678 -5154 -11648 -5024
rect -11582 -5154 -11552 -5024
rect -11486 -5154 -11456 -5024
rect -11390 -5154 -11360 -5024
rect -11298 -5154 -11268 -5024
rect -10806 -5154 -10776 -5024
rect -10714 -5154 -10684 -5024
rect -10618 -5154 -10588 -5024
rect -10522 -5154 -10492 -5024
rect -10426 -5154 -10396 -5024
rect -10330 -5154 -10300 -5024
rect -10234 -5154 -10204 -5024
rect -10138 -5154 -10108 -5024
rect -10042 -5154 -10012 -5024
rect -9946 -5154 -9916 -5024
rect -9850 -5154 -9820 -5024
rect -9754 -5154 -9724 -5024
rect -9658 -5154 -9628 -5024
rect -9566 -5154 -9536 -5024
rect -9247 -5154 -9217 -5024
rect -9155 -5154 -9125 -5024
rect -9059 -5154 -9029 -5024
rect -8963 -5154 -8933 -5024
rect -8867 -5154 -8837 -5024
rect -8771 -5154 -8741 -5024
rect -8675 -5154 -8645 -5024
rect -8579 -5154 -8549 -5024
rect -8483 -5154 -8453 -5024
rect -8387 -5154 -8357 -5024
rect -8291 -5154 -8261 -5024
rect -8195 -5154 -8165 -5024
rect -8099 -5154 -8069 -5024
rect -8007 -5154 -7977 -5024
rect 5658 -5571 5858 -5541
rect 6098 -5571 6298 -5541
rect 6538 -5571 6738 -5541
rect -24162 -5953 -23762 -5923
rect -23586 -5949 -23386 -5919
rect -22426 -5953 -22026 -5923
rect -21852 -5949 -21652 -5919
rect -24162 -6049 -23762 -6019
rect -22426 -6049 -22026 -6019
rect -20296 -6121 -19896 -6091
rect -19187 -6121 -18787 -6091
rect -18305 -6121 -17905 -6091
rect -17005 -6121 -16605 -6091
rect -15896 -6121 -15496 -6091
rect -15014 -6121 -14614 -6091
rect -13714 -6121 -13314 -6091
rect -12605 -6121 -12205 -6091
rect -11723 -6121 -11323 -6091
rect -10423 -6121 -10023 -6091
rect -9314 -6121 -8914 -6091
rect -8432 -6121 -8032 -6091
rect -20296 -6217 -19896 -6187
rect -19187 -6217 -18787 -6187
rect -18305 -6217 -17905 -6187
rect -17005 -6217 -16605 -6187
rect -15896 -6217 -15496 -6187
rect -15014 -6217 -14614 -6187
rect -13714 -6217 -13314 -6187
rect -12605 -6217 -12205 -6187
rect -11723 -6217 -11323 -6187
rect -10423 -6217 -10023 -6187
rect -9314 -6217 -8914 -6187
rect -8432 -6217 -8032 -6187
rect -24162 -7926 -23762 -7896
rect -23584 -7922 -23384 -7892
rect 7422 -7266 7452 -6466
rect 7518 -7266 7548 -6466
rect 7614 -7266 7644 -6466
rect 7710 -7266 7740 -6466
rect 8370 -7266 8400 -6466
rect 8466 -7266 8496 -6466
rect 8562 -7266 8592 -6466
rect 8658 -7266 8688 -6466
rect 9306 -7266 9336 -6466
rect 9402 -7266 9432 -6466
rect 9498 -7266 9528 -6466
rect 9594 -7266 9624 -6466
rect 10237 -7266 10267 -6466
rect 10333 -7266 10363 -6466
rect 10429 -7266 10459 -6466
rect 10525 -7266 10555 -6466
rect 11164 -7266 11194 -6466
rect 11260 -7266 11290 -6466
rect 11356 -7266 11386 -6466
rect 11452 -7266 11482 -6466
rect -22425 -7926 -22025 -7896
rect -21850 -7922 -21650 -7892
rect -24162 -8022 -23762 -7992
rect -22425 -8022 -22025 -7992
rect 7422 -8194 7452 -7394
rect 7518 -8194 7548 -7394
rect 7614 -8194 7644 -7394
rect 7710 -8194 7740 -7394
rect 8370 -8194 8400 -7394
rect 8466 -8194 8496 -7394
rect 8562 -8194 8592 -7394
rect 8658 -8194 8688 -7394
rect 9306 -8194 9336 -7394
rect 9402 -8194 9432 -7394
rect 9498 -8194 9528 -7394
rect 9594 -8194 9624 -7394
rect 10237 -8193 10267 -7393
rect 10333 -8193 10363 -7393
rect 10429 -8193 10459 -7393
rect 10525 -8193 10555 -7393
rect -20679 -8419 -20649 -8289
rect -20587 -8419 -20557 -8289
rect -20491 -8419 -20461 -8289
rect -20395 -8419 -20365 -8289
rect -20299 -8419 -20269 -8289
rect -20203 -8419 -20173 -8289
rect -20107 -8419 -20077 -8289
rect -20011 -8419 -19981 -8289
rect -19915 -8419 -19885 -8289
rect -19819 -8419 -19789 -8289
rect -19723 -8419 -19693 -8289
rect -19627 -8419 -19597 -8289
rect -19531 -8419 -19501 -8289
rect -19439 -8419 -19409 -8289
rect -19120 -8419 -19090 -8289
rect -19028 -8419 -18998 -8289
rect -18932 -8419 -18902 -8289
rect -18836 -8419 -18806 -8289
rect -18740 -8419 -18710 -8289
rect -18644 -8419 -18614 -8289
rect -18548 -8419 -18518 -8289
rect -18452 -8419 -18422 -8289
rect -18356 -8419 -18326 -8289
rect -18260 -8419 -18230 -8289
rect -18164 -8419 -18134 -8289
rect -18068 -8419 -18038 -8289
rect -17972 -8419 -17942 -8289
rect -17880 -8419 -17850 -8289
rect -17388 -8419 -17358 -8289
rect -17296 -8419 -17266 -8289
rect -17200 -8419 -17170 -8289
rect -17104 -8419 -17074 -8289
rect -17008 -8419 -16978 -8289
rect -16912 -8419 -16882 -8289
rect -16816 -8419 -16786 -8289
rect -16720 -8419 -16690 -8289
rect -16624 -8419 -16594 -8289
rect -16528 -8419 -16498 -8289
rect -16432 -8419 -16402 -8289
rect -16336 -8419 -16306 -8289
rect -16240 -8419 -16210 -8289
rect -16148 -8419 -16118 -8289
rect -15829 -8419 -15799 -8289
rect -15737 -8419 -15707 -8289
rect -15641 -8419 -15611 -8289
rect -15545 -8419 -15515 -8289
rect -15449 -8419 -15419 -8289
rect -15353 -8419 -15323 -8289
rect -15257 -8419 -15227 -8289
rect -15161 -8419 -15131 -8289
rect -15065 -8419 -15035 -8289
rect -14969 -8419 -14939 -8289
rect -14873 -8419 -14843 -8289
rect -14777 -8419 -14747 -8289
rect -14681 -8419 -14651 -8289
rect -14589 -8419 -14559 -8289
rect -14097 -8419 -14067 -8289
rect -14005 -8419 -13975 -8289
rect -13909 -8419 -13879 -8289
rect -13813 -8419 -13783 -8289
rect -13717 -8419 -13687 -8289
rect -13621 -8419 -13591 -8289
rect -13525 -8419 -13495 -8289
rect -13429 -8419 -13399 -8289
rect -13333 -8419 -13303 -8289
rect -13237 -8419 -13207 -8289
rect -13141 -8419 -13111 -8289
rect -13045 -8419 -13015 -8289
rect -12949 -8419 -12919 -8289
rect -12857 -8419 -12827 -8289
rect -12538 -8419 -12508 -8289
rect -12446 -8419 -12416 -8289
rect -12350 -8419 -12320 -8289
rect -12254 -8419 -12224 -8289
rect -12158 -8419 -12128 -8289
rect -12062 -8419 -12032 -8289
rect -11966 -8419 -11936 -8289
rect -11870 -8419 -11840 -8289
rect -11774 -8419 -11744 -8289
rect -11678 -8419 -11648 -8289
rect -11582 -8419 -11552 -8289
rect -11486 -8419 -11456 -8289
rect -11390 -8419 -11360 -8289
rect -11298 -8419 -11268 -8289
rect -10806 -8419 -10776 -8289
rect -10714 -8419 -10684 -8289
rect -10618 -8419 -10588 -8289
rect -10522 -8419 -10492 -8289
rect -10426 -8419 -10396 -8289
rect -10330 -8419 -10300 -8289
rect -10234 -8419 -10204 -8289
rect -10138 -8419 -10108 -8289
rect -10042 -8419 -10012 -8289
rect -9946 -8419 -9916 -8289
rect -9850 -8419 -9820 -8289
rect -9754 -8419 -9724 -8289
rect -9658 -8419 -9628 -8289
rect -9566 -8419 -9536 -8289
rect -9247 -8419 -9217 -8289
rect -9155 -8419 -9125 -8289
rect -9059 -8419 -9029 -8289
rect -8963 -8419 -8933 -8289
rect -8867 -8419 -8837 -8289
rect -8771 -8419 -8741 -8289
rect -8675 -8419 -8645 -8289
rect -8579 -8419 -8549 -8289
rect -8483 -8419 -8453 -8289
rect -8387 -8419 -8357 -8289
rect -8291 -8419 -8261 -8289
rect -8195 -8419 -8165 -8289
rect -8099 -8419 -8069 -8289
rect -8007 -8419 -7977 -8289
rect 11164 -8194 11194 -7394
rect 11260 -8194 11290 -7394
rect 11356 -8194 11386 -7394
rect 11452 -8194 11482 -7394
rect 12219 -7636 12249 -7436
rect 12315 -7636 12345 -7436
rect 12923 -7589 13123 -7559
rect -24162 -9218 -23762 -9188
rect -23583 -9214 -23383 -9184
rect -22426 -9218 -22026 -9188
rect -21846 -9214 -21646 -9184
rect -24162 -9314 -23762 -9284
rect -22426 -9314 -22026 -9284
rect -20296 -9386 -19896 -9356
rect -19187 -9386 -18787 -9356
rect -18305 -9386 -17905 -9356
rect -17005 -9386 -16605 -9356
rect -15896 -9386 -15496 -9356
rect -15014 -9386 -14614 -9356
rect -13714 -9386 -13314 -9356
rect -12605 -9386 -12205 -9356
rect -11723 -9386 -11323 -9356
rect -10423 -9386 -10023 -9356
rect -9314 -9386 -8914 -9356
rect -8432 -9386 -8032 -9356
rect -20296 -9482 -19896 -9452
rect -19187 -9482 -18787 -9452
rect -18305 -9482 -17905 -9452
rect -17005 -9482 -16605 -9452
rect -15896 -9482 -15496 -9452
rect -15014 -9482 -14614 -9452
rect -13714 -9482 -13314 -9452
rect -12605 -9482 -12205 -9452
rect -11723 -9482 -11323 -9452
rect -10423 -9482 -10023 -9452
rect -9314 -9482 -8914 -9452
rect -8432 -9482 -8032 -9452
rect 5658 -10199 5858 -10169
rect 6098 -10199 6298 -10169
rect 6538 -10199 6738 -10169
rect -24162 -11190 -23762 -11160
rect -23583 -11186 -23383 -11156
rect -22425 -11190 -22025 -11160
rect -21850 -11186 -21650 -11156
rect -24162 -11286 -23762 -11256
rect -22425 -11286 -22025 -11256
rect -20679 -11683 -20649 -11553
rect -20587 -11683 -20557 -11553
rect -20491 -11683 -20461 -11553
rect -20395 -11683 -20365 -11553
rect -20299 -11683 -20269 -11553
rect -20203 -11683 -20173 -11553
rect -20107 -11683 -20077 -11553
rect -20011 -11683 -19981 -11553
rect -19915 -11683 -19885 -11553
rect -19819 -11683 -19789 -11553
rect -19723 -11683 -19693 -11553
rect -19627 -11683 -19597 -11553
rect -19531 -11683 -19501 -11553
rect -19439 -11683 -19409 -11553
rect -19120 -11683 -19090 -11553
rect -19028 -11683 -18998 -11553
rect -18932 -11683 -18902 -11553
rect -18836 -11683 -18806 -11553
rect -18740 -11683 -18710 -11553
rect -18644 -11683 -18614 -11553
rect -18548 -11683 -18518 -11553
rect -18452 -11683 -18422 -11553
rect -18356 -11683 -18326 -11553
rect -18260 -11683 -18230 -11553
rect -18164 -11683 -18134 -11553
rect -18068 -11683 -18038 -11553
rect -17972 -11683 -17942 -11553
rect -17880 -11683 -17850 -11553
rect -17388 -11683 -17358 -11553
rect -17296 -11683 -17266 -11553
rect -17200 -11683 -17170 -11553
rect -17104 -11683 -17074 -11553
rect -17008 -11683 -16978 -11553
rect -16912 -11683 -16882 -11553
rect -16816 -11683 -16786 -11553
rect -16720 -11683 -16690 -11553
rect -16624 -11683 -16594 -11553
rect -16528 -11683 -16498 -11553
rect -16432 -11683 -16402 -11553
rect -16336 -11683 -16306 -11553
rect -16240 -11683 -16210 -11553
rect -16148 -11683 -16118 -11553
rect -15829 -11683 -15799 -11553
rect -15737 -11683 -15707 -11553
rect -15641 -11683 -15611 -11553
rect -15545 -11683 -15515 -11553
rect -15449 -11683 -15419 -11553
rect -15353 -11683 -15323 -11553
rect -15257 -11683 -15227 -11553
rect -15161 -11683 -15131 -11553
rect -15065 -11683 -15035 -11553
rect -14969 -11683 -14939 -11553
rect -14873 -11683 -14843 -11553
rect -14777 -11683 -14747 -11553
rect -14681 -11683 -14651 -11553
rect -14589 -11683 -14559 -11553
rect -14097 -11683 -14067 -11553
rect -14005 -11683 -13975 -11553
rect -13909 -11683 -13879 -11553
rect -13813 -11683 -13783 -11553
rect -13717 -11683 -13687 -11553
rect -13621 -11683 -13591 -11553
rect -13525 -11683 -13495 -11553
rect -13429 -11683 -13399 -11553
rect -13333 -11683 -13303 -11553
rect -13237 -11683 -13207 -11553
rect -13141 -11683 -13111 -11553
rect -13045 -11683 -13015 -11553
rect -12949 -11683 -12919 -11553
rect -12857 -11683 -12827 -11553
rect -12538 -11683 -12508 -11553
rect -12446 -11683 -12416 -11553
rect -12350 -11683 -12320 -11553
rect -12254 -11683 -12224 -11553
rect -12158 -11683 -12128 -11553
rect -12062 -11683 -12032 -11553
rect -11966 -11683 -11936 -11553
rect -11870 -11683 -11840 -11553
rect -11774 -11683 -11744 -11553
rect -11678 -11683 -11648 -11553
rect -11582 -11683 -11552 -11553
rect -11486 -11683 -11456 -11553
rect -11390 -11683 -11360 -11553
rect -11298 -11683 -11268 -11553
rect -10806 -11683 -10776 -11553
rect -10714 -11683 -10684 -11553
rect -10618 -11683 -10588 -11553
rect -10522 -11683 -10492 -11553
rect -10426 -11683 -10396 -11553
rect -10330 -11683 -10300 -11553
rect -10234 -11683 -10204 -11553
rect -10138 -11683 -10108 -11553
rect -10042 -11683 -10012 -11553
rect -9946 -11683 -9916 -11553
rect -9850 -11683 -9820 -11553
rect -9754 -11683 -9724 -11553
rect -9658 -11683 -9628 -11553
rect -9566 -11683 -9536 -11553
rect -9247 -11683 -9217 -11553
rect -9155 -11683 -9125 -11553
rect -9059 -11683 -9029 -11553
rect -8963 -11683 -8933 -11553
rect -8867 -11683 -8837 -11553
rect -8771 -11683 -8741 -11553
rect -8675 -11683 -8645 -11553
rect -8579 -11683 -8549 -11553
rect -8483 -11683 -8453 -11553
rect -8387 -11683 -8357 -11553
rect -8291 -11683 -8261 -11553
rect -8195 -11683 -8165 -11553
rect -8099 -11683 -8069 -11553
rect -8007 -11683 -7977 -11553
rect 7422 -11894 7452 -11094
rect 7518 -11894 7548 -11094
rect 7614 -11894 7644 -11094
rect 7710 -11894 7740 -11094
rect 8370 -11894 8400 -11094
rect 8466 -11894 8496 -11094
rect 8562 -11894 8592 -11094
rect 8658 -11894 8688 -11094
rect 9306 -11894 9336 -11094
rect 9402 -11894 9432 -11094
rect 9498 -11894 9528 -11094
rect 9594 -11894 9624 -11094
rect 10237 -11894 10267 -11094
rect 10333 -11894 10363 -11094
rect 10429 -11894 10459 -11094
rect 10525 -11894 10555 -11094
rect 11164 -11894 11194 -11094
rect 11260 -11894 11290 -11094
rect 11356 -11894 11386 -11094
rect 11452 -11894 11482 -11094
rect -24162 -12482 -23762 -12452
rect -23583 -12478 -23383 -12448
rect -22425 -12482 -22025 -12452
rect -21854 -12478 -21654 -12448
rect -24162 -12578 -23762 -12548
rect -22425 -12578 -22025 -12548
rect -20296 -12650 -19896 -12620
rect -19187 -12650 -18787 -12620
rect -18305 -12650 -17905 -12620
rect -17005 -12650 -16605 -12620
rect -15896 -12650 -15496 -12620
rect -15014 -12650 -14614 -12620
rect -13714 -12650 -13314 -12620
rect -12605 -12650 -12205 -12620
rect -11723 -12650 -11323 -12620
rect -10423 -12650 -10023 -12620
rect -9314 -12650 -8914 -12620
rect -8432 -12650 -8032 -12620
rect -20296 -12746 -19896 -12716
rect -19187 -12746 -18787 -12716
rect -18305 -12746 -17905 -12716
rect -17005 -12746 -16605 -12716
rect -15896 -12746 -15496 -12716
rect -15014 -12746 -14614 -12716
rect -13714 -12746 -13314 -12716
rect -12605 -12746 -12205 -12716
rect -11723 -12746 -11323 -12716
rect -10423 -12746 -10023 -12716
rect -9314 -12746 -8914 -12716
rect -8432 -12746 -8032 -12716
rect 7422 -12822 7452 -12022
rect 7518 -12822 7548 -12022
rect 7614 -12822 7644 -12022
rect 7710 -12822 7740 -12022
rect 8370 -12822 8400 -12022
rect 8466 -12822 8496 -12022
rect 8562 -12822 8592 -12022
rect 8658 -12822 8688 -12022
rect 9306 -12822 9336 -12022
rect 9402 -12822 9432 -12022
rect 9498 -12822 9528 -12022
rect 9594 -12822 9624 -12022
rect 10237 -12821 10267 -12021
rect 10333 -12821 10363 -12021
rect 10429 -12821 10459 -12021
rect 10525 -12821 10555 -12021
rect 11164 -12822 11194 -12022
rect 11260 -12822 11290 -12022
rect 11356 -12822 11386 -12022
rect 11452 -12822 11482 -12022
rect 12219 -12264 12249 -12064
rect 12315 -12264 12345 -12064
rect 12923 -12217 13123 -12187
rect -1604 -14032 -1574 -13832
rect -11276 -14181 -11146 -14151
rect -24043 -15316 -24013 -14916
rect -23947 -15316 -23917 -14916
rect -17188 -14975 -16988 -14945
rect -17188 -15071 -16988 -15041
rect -11276 -14273 -11146 -14243
rect -11276 -14369 -11146 -14339
rect -11276 -14465 -11146 -14435
rect -11276 -14561 -11146 -14531
rect -11276 -14657 -11146 -14627
rect -11276 -14753 -11146 -14723
rect -11276 -14849 -11146 -14819
rect -11276 -14945 -11146 -14915
rect -11276 -15041 -11146 -15011
rect -11276 -15137 -11146 -15107
rect -11276 -15233 -11146 -15203
rect -11276 -15329 -11146 -15299
rect -4320 -14403 -4290 -14203
rect -1604 -14411 -1574 -14211
rect -4320 -14843 -4290 -14643
rect -1604 -14851 -1574 -14651
rect 5658 -14727 5858 -14697
rect 6098 -14727 6298 -14697
rect 6538 -14727 6738 -14697
rect -4320 -15222 -4290 -15022
rect -1604 -15230 -1574 -15030
rect -11276 -15421 -11146 -15391
rect -7671 -15560 -7641 -15360
rect -4320 -15662 -4290 -15462
rect -1604 -15670 -1574 -15470
rect -7670 -16060 -7640 -15860
rect -4320 -16041 -4290 -15841
rect -24042 -16501 -24012 -16101
rect -23946 -16501 -23916 -16101
rect -1604 -16049 -1574 -15849
rect -17188 -16375 -16988 -16345
rect -17188 -16471 -16988 -16441
rect -7671 -16540 -7641 -16340
rect -4320 -16481 -4290 -16281
rect -1604 -16489 -1574 -16289
rect 7422 -16422 7452 -15622
rect 7518 -16422 7548 -15622
rect 7614 -16422 7644 -15622
rect 7710 -16422 7740 -15622
rect 8370 -16422 8400 -15622
rect 8466 -16422 8496 -15622
rect 8562 -16422 8592 -15622
rect 8658 -16422 8688 -15622
rect 9306 -16422 9336 -15622
rect 9402 -16422 9432 -15622
rect 9498 -16422 9528 -15622
rect 9594 -16422 9624 -15622
rect 10237 -16422 10267 -15622
rect 10333 -16422 10363 -15622
rect 10429 -16422 10459 -15622
rect 10525 -16422 10555 -15622
rect 11164 -16422 11194 -15622
rect 11260 -16422 11290 -15622
rect 11356 -16422 11386 -15622
rect 11452 -16422 11482 -15622
rect -11274 -16997 -11144 -16967
rect -24037 -17714 -24007 -17314
rect -23941 -17714 -23911 -17314
rect -17188 -17775 -16988 -17745
rect -17188 -17871 -16988 -17841
rect -21110 -18248 -21080 -18048
rect -15519 -18119 -15489 -17919
rect -11274 -17089 -11144 -17059
rect -11274 -17185 -11144 -17155
rect -11274 -17281 -11144 -17251
rect -11274 -17377 -11144 -17347
rect -11274 -17473 -11144 -17443
rect -11274 -17569 -11144 -17539
rect -11274 -17665 -11144 -17635
rect -11274 -17761 -11144 -17731
rect -11274 -17857 -11144 -17827
rect -11274 -17953 -11144 -17923
rect -11274 -18049 -11144 -18019
rect -11274 -18145 -11144 -18115
rect -7671 -17040 -7641 -16840
rect -4320 -16860 -4290 -16660
rect -1604 -16868 -1574 -16668
rect -4320 -17300 -4290 -17100
rect -7671 -17520 -7641 -17320
rect -1604 -17308 -1574 -17108
rect 7422 -17350 7452 -16550
rect 7518 -17350 7548 -16550
rect 7614 -17350 7644 -16550
rect 7710 -17350 7740 -16550
rect 8370 -17350 8400 -16550
rect 8466 -17350 8496 -16550
rect 8562 -17350 8592 -16550
rect 8658 -17350 8688 -16550
rect 9306 -17350 9336 -16550
rect 9402 -17350 9432 -16550
rect 9498 -17350 9528 -16550
rect 9594 -17350 9624 -16550
rect 10237 -17349 10267 -16549
rect 10333 -17349 10363 -16549
rect 10429 -17349 10459 -16549
rect 10525 -17349 10555 -16549
rect -4320 -17679 -4290 -17479
rect -1604 -17687 -1574 -17487
rect -7671 -17980 -7641 -17780
rect 11164 -17350 11194 -16550
rect 11260 -17350 11290 -16550
rect 11356 -17350 11386 -16550
rect 11452 -17350 11482 -16550
rect 12219 -16792 12249 -16592
rect 12315 -16792 12345 -16592
rect 12923 -16745 13123 -16715
rect 16209 -17249 16239 -17049
rect 16305 -17249 16335 -17049
rect 16401 -17249 16431 -17049
rect 16497 -17249 16527 -17049
rect -4320 -18119 -4290 -17919
rect -1604 -18127 -1574 -17927
rect -11274 -18237 -11144 -18207
rect -24022 -18833 -23992 -18433
rect -23926 -18833 -23896 -18433
rect -21109 -18748 -21079 -18548
rect -15518 -18619 -15488 -18419
rect -7685 -18440 -7655 -18240
rect -4320 -18498 -4290 -18298
rect -1604 -18506 -1574 -18306
rect -21110 -19228 -21080 -19028
rect -15519 -19099 -15489 -18899
rect -7683 -18920 -7653 -18720
rect -4320 -18938 -4290 -18738
rect -1604 -18946 -1574 -18746
rect -17188 -19175 -16988 -19145
rect -17188 -19271 -16988 -19241
rect -24020 -20027 -23990 -19627
rect -23924 -20027 -23894 -19627
rect -21110 -19728 -21080 -19528
rect -4320 -19317 -4290 -19117
rect -1604 -19325 -1574 -19125
rect 5658 -19255 5858 -19225
rect 6098 -19255 6298 -19225
rect 6538 -19255 6738 -19225
rect -15519 -19599 -15489 -19399
rect -4320 -19757 -4290 -19557
rect -1604 -19765 -1574 -19565
rect 17528 -18711 17928 -18681
rect 17528 -18807 17928 -18777
rect 18096 -18785 18296 -18755
rect -21110 -20208 -21080 -20008
rect -15519 -20079 -15489 -19879
rect -11274 -19954 -11144 -19924
rect -21110 -20668 -21080 -20468
rect -17188 -20575 -16988 -20545
rect -17188 -20671 -16988 -20641
rect -23989 -21227 -23959 -20827
rect -23893 -21227 -23863 -20827
rect -21124 -21128 -21094 -20928
rect -15519 -20539 -15489 -20339
rect -15533 -20999 -15503 -20799
rect -11274 -20046 -11144 -20016
rect -11274 -20142 -11144 -20112
rect -11274 -20238 -11144 -20208
rect -11274 -20334 -11144 -20304
rect -11274 -20430 -11144 -20400
rect -11274 -20526 -11144 -20496
rect -11274 -20622 -11144 -20592
rect -11274 -20718 -11144 -20688
rect -11274 -20814 -11144 -20784
rect -11274 -20910 -11144 -20880
rect -11274 -21006 -11144 -20976
rect -11274 -21102 -11144 -21072
rect -4320 -20136 -4290 -19936
rect -1604 -20144 -1574 -19944
rect 16209 -20123 16239 -19923
rect 16305 -20123 16335 -19923
rect 16401 -20123 16431 -19923
rect 16497 -20123 16527 -19923
rect -4320 -20576 -4290 -20376
rect -1604 -20584 -1574 -20384
rect -4320 -20955 -4290 -20755
rect 7422 -20950 7452 -20150
rect 7518 -20950 7548 -20150
rect 7614 -20950 7644 -20150
rect 7710 -20950 7740 -20150
rect 8370 -20950 8400 -20150
rect 8466 -20950 8496 -20150
rect 8562 -20950 8592 -20150
rect 8658 -20950 8688 -20150
rect 9306 -20950 9336 -20150
rect 9402 -20950 9432 -20150
rect 9498 -20950 9528 -20150
rect 9594 -20950 9624 -20150
rect 10237 -20950 10267 -20150
rect 10333 -20950 10363 -20150
rect 10429 -20950 10459 -20150
rect 10525 -20950 10555 -20150
rect 11164 -20950 11194 -20150
rect 11260 -20950 11290 -20150
rect 11356 -20950 11386 -20150
rect 11452 -20950 11482 -20150
rect -11274 -21194 -11144 -21164
rect -21122 -21608 -21092 -21408
rect -15531 -21479 -15501 -21279
rect 7422 -21878 7452 -21078
rect 7518 -21878 7548 -21078
rect 7614 -21878 7644 -21078
rect 7710 -21878 7740 -21078
rect 8370 -21878 8400 -21078
rect 8466 -21878 8496 -21078
rect 8562 -21878 8592 -21078
rect 8658 -21878 8688 -21078
rect 9306 -21878 9336 -21078
rect 9402 -21878 9432 -21078
rect 9498 -21878 9528 -21078
rect 9594 -21878 9624 -21078
rect 10237 -21877 10267 -21077
rect 10333 -21877 10363 -21077
rect 10429 -21877 10459 -21077
rect 10525 -21877 10555 -21077
rect -17188 -21975 -16988 -21945
rect -17188 -22071 -16988 -22041
rect -23990 -22530 -23960 -22130
rect -23894 -22530 -23864 -22130
rect 11164 -21878 11194 -21078
rect 11260 -21878 11290 -21078
rect 11356 -21878 11386 -21078
rect 11452 -21878 11482 -21078
rect 12219 -21320 12249 -21120
rect 12315 -21320 12345 -21120
rect 12923 -21273 13123 -21243
rect -11274 -22533 -11144 -22503
rect -17188 -23375 -16988 -23345
rect -23990 -23839 -23960 -23439
rect -23894 -23839 -23864 -23439
rect -17188 -23471 -16988 -23441
rect -11274 -22625 -11144 -22595
rect -11274 -22721 -11144 -22691
rect -11274 -22817 -11144 -22787
rect -11274 -22913 -11144 -22883
rect -11274 -23009 -11144 -22979
rect -11274 -23105 -11144 -23075
rect -11274 -23201 -11144 -23171
rect -11274 -23297 -11144 -23267
rect -11274 -23393 -11144 -23363
rect -11274 -23489 -11144 -23459
rect -11274 -23585 -11144 -23555
rect -11274 -23681 -11144 -23651
rect -11274 -23773 -11144 -23743
rect 5658 -23783 5858 -23753
rect 6098 -23783 6298 -23753
rect 6538 -23783 6738 -23753
rect -17188 -24775 -16988 -24745
rect -17188 -24871 -16988 -24841
rect -11274 -25301 -11144 -25271
rect -11274 -25393 -11144 -25363
rect -11274 -25489 -11144 -25459
rect -11274 -25585 -11144 -25555
rect -11274 -25681 -11144 -25651
rect -11274 -25777 -11144 -25747
rect -11274 -25873 -11144 -25843
rect -11274 -25969 -11144 -25939
rect -11274 -26065 -11144 -26035
rect -11274 -26161 -11144 -26131
rect -11274 -26257 -11144 -26227
rect -11274 -26353 -11144 -26323
rect -11274 -26449 -11144 -26419
rect 7422 -25478 7452 -24678
rect 7518 -25478 7548 -24678
rect 7614 -25478 7644 -24678
rect 7710 -25478 7740 -24678
rect 8370 -25478 8400 -24678
rect 8466 -25478 8496 -24678
rect 8562 -25478 8592 -24678
rect 8658 -25478 8688 -24678
rect 9306 -25478 9336 -24678
rect 9402 -25478 9432 -24678
rect 9498 -25478 9528 -24678
rect 9594 -25478 9624 -24678
rect 10237 -25478 10267 -24678
rect 10333 -25478 10363 -24678
rect 10429 -25478 10459 -24678
rect 10525 -25478 10555 -24678
rect 11164 -25478 11194 -24678
rect 11260 -25478 11290 -24678
rect 11356 -25478 11386 -24678
rect 11452 -25478 11482 -24678
rect 7422 -26406 7452 -25606
rect 7518 -26406 7548 -25606
rect 7614 -26406 7644 -25606
rect 7710 -26406 7740 -25606
rect 8370 -26406 8400 -25606
rect 8466 -26406 8496 -25606
rect 8562 -26406 8592 -25606
rect 8658 -26406 8688 -25606
rect 9306 -26406 9336 -25606
rect 9402 -26406 9432 -25606
rect 9498 -26406 9528 -25606
rect 9594 -26406 9624 -25606
rect 10237 -26405 10267 -25605
rect 10333 -26405 10363 -25605
rect 10429 -26405 10459 -25605
rect 10525 -26405 10555 -25605
rect -11274 -26541 -11144 -26511
rect 11164 -26406 11194 -25606
rect 11260 -26406 11290 -25606
rect 11356 -26406 11386 -25606
rect 11452 -26406 11482 -25606
rect 12219 -25848 12249 -25648
rect 12315 -25848 12345 -25648
rect 12923 -25801 13123 -25771
rect -11274 -27934 -11144 -27904
rect -11274 -28026 -11144 -27996
rect -11274 -28122 -11144 -28092
rect -11274 -28218 -11144 -28188
rect -11274 -28314 -11144 -28284
rect -11274 -28410 -11144 -28380
rect -11274 -28506 -11144 -28476
rect -11274 -28602 -11144 -28572
rect -11274 -28698 -11144 -28668
rect -11274 -28794 -11144 -28764
rect -11274 -28890 -11144 -28860
rect -11274 -28986 -11144 -28956
rect -11274 -29082 -11144 -29052
rect 5658 -28311 5858 -28281
rect 6098 -28311 6298 -28281
rect 6538 -28311 6738 -28281
rect -11274 -29174 -11144 -29144
rect 7422 -30006 7452 -29206
rect 7518 -30006 7548 -29206
rect 7614 -30006 7644 -29206
rect 7710 -30006 7740 -29206
rect 8370 -30006 8400 -29206
rect 8466 -30006 8496 -29206
rect 8562 -30006 8592 -29206
rect 8658 -30006 8688 -29206
rect 9306 -30006 9336 -29206
rect 9402 -30006 9432 -29206
rect 9498 -30006 9528 -29206
rect 9594 -30006 9624 -29206
rect 10237 -30006 10267 -29206
rect 10333 -30006 10363 -29206
rect 10429 -30006 10459 -29206
rect 10525 -30006 10555 -29206
rect 11164 -30006 11194 -29206
rect 11260 -30006 11290 -29206
rect 11356 -30006 11386 -29206
rect 11452 -30006 11482 -29206
rect -11274 -30543 -11144 -30513
rect -11274 -30635 -11144 -30605
rect -11274 -30731 -11144 -30701
rect -11274 -30827 -11144 -30797
rect -11274 -30923 -11144 -30893
rect -11274 -31019 -11144 -30989
rect -11274 -31115 -11144 -31085
rect -11274 -31211 -11144 -31181
rect -11274 -31307 -11144 -31277
rect -11274 -31403 -11144 -31373
rect -11274 -31499 -11144 -31469
rect -11274 -31595 -11144 -31565
rect -11274 -31691 -11144 -31661
rect 7422 -30934 7452 -30134
rect 7518 -30934 7548 -30134
rect 7614 -30934 7644 -30134
rect 7710 -30934 7740 -30134
rect 8370 -30934 8400 -30134
rect 8466 -30934 8496 -30134
rect 8562 -30934 8592 -30134
rect 8658 -30934 8688 -30134
rect 9306 -30934 9336 -30134
rect 9402 -30934 9432 -30134
rect 9498 -30934 9528 -30134
rect 9594 -30934 9624 -30134
rect 10237 -30933 10267 -30133
rect 10333 -30933 10363 -30133
rect 10429 -30933 10459 -30133
rect 10525 -30933 10555 -30133
rect 11164 -30934 11194 -30134
rect 11260 -30934 11290 -30134
rect 11356 -30934 11386 -30134
rect 11452 -30934 11482 -30134
rect 12219 -30376 12249 -30176
rect 12315 -30376 12345 -30176
rect 12923 -30329 13123 -30299
rect -11274 -31783 -11144 -31753
rect 5658 -32839 5858 -32809
rect 6098 -32839 6298 -32809
rect 6538 -32839 6738 -32809
rect -11276 -33163 -11146 -33133
rect -11276 -33255 -11146 -33225
rect -11276 -33351 -11146 -33321
rect -11276 -33447 -11146 -33417
rect -11276 -33543 -11146 -33513
rect -11276 -33639 -11146 -33609
rect -11276 -33735 -11146 -33705
rect -11276 -33831 -11146 -33801
rect -11276 -33927 -11146 -33897
rect -11276 -34023 -11146 -33993
rect -11276 -34119 -11146 -34089
rect -11276 -34215 -11146 -34185
rect -11276 -34311 -11146 -34281
rect -11276 -34403 -11146 -34373
rect 7422 -34534 7452 -33734
rect 7518 -34534 7548 -33734
rect 7614 -34534 7644 -33734
rect 7710 -34534 7740 -33734
rect 8370 -34534 8400 -33734
rect 8466 -34534 8496 -33734
rect 8562 -34534 8592 -33734
rect 8658 -34534 8688 -33734
rect 9306 -34534 9336 -33734
rect 9402 -34534 9432 -33734
rect 9498 -34534 9528 -33734
rect 9594 -34534 9624 -33734
rect 10237 -34534 10267 -33734
rect 10333 -34534 10363 -33734
rect 10429 -34534 10459 -33734
rect 10525 -34534 10555 -33734
rect 11164 -34534 11194 -33734
rect 11260 -34534 11290 -33734
rect 11356 -34534 11386 -33734
rect 11452 -34534 11482 -33734
rect 7422 -35462 7452 -34662
rect 7518 -35462 7548 -34662
rect 7614 -35462 7644 -34662
rect 7710 -35462 7740 -34662
rect 8370 -35462 8400 -34662
rect 8466 -35462 8496 -34662
rect 8562 -35462 8592 -34662
rect 8658 -35462 8688 -34662
rect 9306 -35462 9336 -34662
rect 9402 -35462 9432 -34662
rect 9498 -35462 9528 -34662
rect 9594 -35462 9624 -34662
rect 10237 -35461 10267 -34661
rect 10333 -35461 10363 -34661
rect 10429 -35461 10459 -34661
rect 10525 -35461 10555 -34661
rect 11164 -35462 11194 -34662
rect 11260 -35462 11290 -34662
rect 11356 -35462 11386 -34662
rect 11452 -35462 11482 -34662
rect 12219 -34904 12249 -34704
rect 12315 -34904 12345 -34704
rect 12923 -34857 13123 -34827
rect 12932 -35915 12962 -35715
rect 12932 -36294 12962 -36094
<< pmos >>
rect 1765 5534 1795 6084
rect 1857 5534 1887 6084
rect 1953 5534 1983 6084
rect 2049 5534 2079 6084
rect 2145 5534 2175 6084
rect 2241 5534 2271 6084
rect 2337 5534 2367 6084
rect 2433 5534 2463 6084
rect 2529 5534 2559 6084
rect 2625 5534 2655 6084
rect 2721 5534 2751 6084
rect 2817 5534 2847 6084
rect 2913 5534 2943 6084
rect 3005 5534 3035 6084
rect 3371 5534 3401 6084
rect 3463 5534 3493 6084
rect 3559 5534 3589 6084
rect 3655 5534 3685 6084
rect 3751 5534 3781 6084
rect 3847 5534 3877 6084
rect 3943 5534 3973 6084
rect 4039 5534 4069 6084
rect 4135 5534 4165 6084
rect 4231 5534 4261 6084
rect 4327 5534 4357 6084
rect 4423 5534 4453 6084
rect 4519 5534 4549 6084
rect 4611 5534 4641 6084
rect 5075 5532 5105 6082
rect 5167 5532 5197 6082
rect 5263 5532 5293 6082
rect 5359 5532 5389 6082
rect 5455 5532 5485 6082
rect 5551 5532 5581 6082
rect 5647 5532 5677 6082
rect 5743 5532 5773 6082
rect 5839 5532 5869 6082
rect 5935 5532 5965 6082
rect 6031 5532 6061 6082
rect 6127 5532 6157 6082
rect 6223 5532 6253 6082
rect 6315 5532 6345 6082
rect 7001 5227 7031 5441
rect 7097 5227 7127 5441
rect 7193 5227 7223 5441
rect 7289 5227 7319 5441
rect 7385 5227 7415 5441
rect 7481 5227 7511 5441
rect 7809 5379 8023 5409
rect 7809 5283 8023 5313
rect 7809 5187 8023 5217
rect -24072 3810 -24042 4360
rect -23980 3810 -23950 4360
rect -23884 3810 -23854 4360
rect -23788 3810 -23758 4360
rect -23692 3810 -23662 4360
rect -23596 3810 -23566 4360
rect -23500 3810 -23470 4360
rect -23404 3810 -23374 4360
rect -23308 3810 -23278 4360
rect -23212 3810 -23182 4360
rect -23116 3810 -23086 4360
rect -23020 3810 -22990 4360
rect -22924 3810 -22894 4360
rect -22832 3810 -22802 4360
rect -20781 3810 -20751 4360
rect -20689 3810 -20659 4360
rect -20593 3810 -20563 4360
rect -20497 3810 -20467 4360
rect -20401 3810 -20371 4360
rect -20305 3810 -20275 4360
rect -20209 3810 -20179 4360
rect -20113 3810 -20083 4360
rect -20017 3810 -19987 4360
rect -19921 3810 -19891 4360
rect -19825 3810 -19795 4360
rect -19729 3810 -19699 4360
rect -19633 3810 -19603 4360
rect -19541 3810 -19511 4360
rect -17490 3810 -17460 4360
rect -17398 3810 -17368 4360
rect -17302 3810 -17272 4360
rect -17206 3810 -17176 4360
rect -17110 3810 -17080 4360
rect -17014 3810 -16984 4360
rect -16918 3810 -16888 4360
rect -16822 3810 -16792 4360
rect -16726 3810 -16696 4360
rect -16630 3810 -16600 4360
rect -16534 3810 -16504 4360
rect -16438 3810 -16408 4360
rect -16342 3810 -16312 4360
rect -16250 3810 -16220 4360
rect -14199 3810 -14169 4360
rect -14107 3810 -14077 4360
rect -14011 3810 -13981 4360
rect -13915 3810 -13885 4360
rect -13819 3810 -13789 4360
rect -13723 3810 -13693 4360
rect -13627 3810 -13597 4360
rect -13531 3810 -13501 4360
rect -13435 3810 -13405 4360
rect -13339 3810 -13309 4360
rect -13243 3810 -13213 4360
rect -13147 3810 -13117 4360
rect -13051 3810 -13021 4360
rect -12959 3810 -12929 4360
rect -10908 3810 -10878 4360
rect -10816 3810 -10786 4360
rect -10720 3810 -10690 4360
rect -10624 3810 -10594 4360
rect -10528 3810 -10498 4360
rect -10432 3810 -10402 4360
rect -10336 3810 -10306 4360
rect -10240 3810 -10210 4360
rect -10144 3810 -10114 4360
rect -10048 3810 -10018 4360
rect -9952 3810 -9922 4360
rect -9856 3810 -9826 4360
rect -9760 3810 -9730 4360
rect -9668 3810 -9638 4360
rect -7618 3810 -7588 4360
rect -7526 3810 -7496 4360
rect -7430 3810 -7400 4360
rect -7334 3810 -7304 4360
rect -7238 3810 -7208 4360
rect -7142 3810 -7112 4360
rect -7046 3810 -7016 4360
rect -6950 3810 -6920 4360
rect -6854 3810 -6824 4360
rect -6758 3810 -6728 4360
rect -6662 3810 -6632 4360
rect -6566 3810 -6536 4360
rect -6470 3810 -6440 4360
rect -6378 3810 -6348 4360
rect -4327 3810 -4297 4360
rect -4235 3810 -4205 4360
rect -4139 3810 -4109 4360
rect -4043 3810 -4013 4360
rect -3947 3810 -3917 4360
rect -3851 3810 -3821 4360
rect -3755 3810 -3725 4360
rect -3659 3810 -3629 4360
rect -3563 3810 -3533 4360
rect -3467 3810 -3437 4360
rect -3371 3810 -3341 4360
rect -3275 3810 -3245 4360
rect -3179 3810 -3149 4360
rect -3087 3810 -3057 4360
rect -1036 3810 -1006 4360
rect -944 3810 -914 4360
rect -848 3810 -818 4360
rect -752 3810 -722 4360
rect -656 3810 -626 4360
rect -560 3810 -530 4360
rect -464 3810 -434 4360
rect -368 3810 -338 4360
rect -272 3810 -242 4360
rect -176 3810 -146 4360
rect -80 3810 -50 4360
rect 16 3810 46 4360
rect 112 3810 142 4360
rect 204 3810 234 4360
rect 5658 3831 5872 3861
rect 5658 3735 5872 3765
rect 5658 3639 5872 3669
rect 6098 3831 6312 3861
rect 6098 3735 6312 3765
rect 6098 3639 6312 3669
rect 6538 3831 6752 3861
rect 6538 3735 6752 3765
rect 6538 3639 6752 3669
rect 7200 2897 7230 3219
rect 7296 2897 7326 3219
rect 7392 2897 7422 3219
rect 7488 2897 7518 3219
rect 7584 2897 7614 3219
rect 7680 2897 7710 3219
rect 7776 2897 7806 3219
rect 7872 2897 7902 3219
rect 8148 2897 8178 3219
rect 8244 2897 8274 3219
rect 8340 2897 8370 3219
rect 8436 2897 8466 3219
rect 8532 2897 8562 3219
rect 8628 2897 8658 3219
rect 8724 2897 8754 3219
rect 8820 2897 8850 3219
rect 9084 2897 9114 3219
rect 9180 2897 9210 3219
rect 9276 2897 9306 3219
rect 9372 2897 9402 3219
rect 9468 2897 9498 3219
rect 9564 2897 9594 3219
rect 9660 2897 9690 3219
rect 9756 2897 9786 3219
rect 10015 2897 10045 3219
rect 10111 2897 10141 3219
rect 10207 2897 10237 3219
rect 10303 2897 10333 3219
rect 10399 2897 10429 3219
rect 10495 2897 10525 3219
rect 10591 2897 10621 3219
rect 10687 2897 10717 3219
rect 10942 2897 10972 3219
rect 11038 2897 11068 3219
rect 11134 2897 11164 3219
rect 11230 2897 11260 3219
rect 11326 2897 11356 3219
rect 11422 2897 11452 3219
rect 11518 2897 11548 3219
rect 11614 2897 11644 3219
rect -24746 2026 -24716 2576
rect -24654 2026 -24624 2576
rect -24558 2026 -24528 2576
rect -24462 2026 -24432 2576
rect -24366 2026 -24336 2576
rect -24270 2026 -24240 2576
rect -24174 2026 -24144 2576
rect -24078 2026 -24048 2576
rect -23982 2026 -23952 2576
rect -23886 2026 -23856 2576
rect -23790 2026 -23760 2576
rect -23694 2026 -23664 2576
rect -23598 2026 -23568 2576
rect -23506 2026 -23476 2576
rect -23187 2026 -23157 2576
rect -23095 2026 -23065 2576
rect -22999 2026 -22969 2576
rect -22903 2026 -22873 2576
rect -22807 2026 -22777 2576
rect -22711 2026 -22681 2576
rect -22615 2026 -22585 2576
rect -22519 2026 -22489 2576
rect -22423 2026 -22393 2576
rect -22327 2026 -22297 2576
rect -22231 2026 -22201 2576
rect -22135 2026 -22105 2576
rect -22039 2026 -22009 2576
rect -21947 2026 -21917 2576
rect -21455 2026 -21425 2576
rect -21363 2026 -21333 2576
rect -21267 2026 -21237 2576
rect -21171 2026 -21141 2576
rect -21075 2026 -21045 2576
rect -20979 2026 -20949 2576
rect -20883 2026 -20853 2576
rect -20787 2026 -20757 2576
rect -20691 2026 -20661 2576
rect -20595 2026 -20565 2576
rect -20499 2026 -20469 2576
rect -20403 2026 -20373 2576
rect -20307 2026 -20277 2576
rect -20215 2026 -20185 2576
rect -19896 2026 -19866 2576
rect -19804 2026 -19774 2576
rect -19708 2026 -19678 2576
rect -19612 2026 -19582 2576
rect -19516 2026 -19486 2576
rect -19420 2026 -19390 2576
rect -19324 2026 -19294 2576
rect -19228 2026 -19198 2576
rect -19132 2026 -19102 2576
rect -19036 2026 -19006 2576
rect -18940 2026 -18910 2576
rect -18844 2026 -18814 2576
rect -18748 2026 -18718 2576
rect -18656 2026 -18626 2576
rect -18164 2026 -18134 2576
rect -18072 2026 -18042 2576
rect -17976 2026 -17946 2576
rect -17880 2026 -17850 2576
rect -17784 2026 -17754 2576
rect -17688 2026 -17658 2576
rect -17592 2026 -17562 2576
rect -17496 2026 -17466 2576
rect -17400 2026 -17370 2576
rect -17304 2026 -17274 2576
rect -17208 2026 -17178 2576
rect -17112 2026 -17082 2576
rect -17016 2026 -16986 2576
rect -16924 2026 -16894 2576
rect -16605 2026 -16575 2576
rect -16513 2026 -16483 2576
rect -16417 2026 -16387 2576
rect -16321 2026 -16291 2576
rect -16225 2026 -16195 2576
rect -16129 2026 -16099 2576
rect -16033 2026 -16003 2576
rect -15937 2026 -15907 2576
rect -15841 2026 -15811 2576
rect -15745 2026 -15715 2576
rect -15649 2026 -15619 2576
rect -15553 2026 -15523 2576
rect -15457 2026 -15427 2576
rect -15365 2026 -15335 2576
rect -14873 2026 -14843 2576
rect -14781 2026 -14751 2576
rect -14685 2026 -14655 2576
rect -14589 2026 -14559 2576
rect -14493 2026 -14463 2576
rect -14397 2026 -14367 2576
rect -14301 2026 -14271 2576
rect -14205 2026 -14175 2576
rect -14109 2026 -14079 2576
rect -14013 2026 -13983 2576
rect -13917 2026 -13887 2576
rect -13821 2026 -13791 2576
rect -13725 2026 -13695 2576
rect -13633 2026 -13603 2576
rect -13314 2026 -13284 2576
rect -13222 2026 -13192 2576
rect -13126 2026 -13096 2576
rect -13030 2026 -13000 2576
rect -12934 2026 -12904 2576
rect -12838 2026 -12808 2576
rect -12742 2026 -12712 2576
rect -12646 2026 -12616 2576
rect -12550 2026 -12520 2576
rect -12454 2026 -12424 2576
rect -12358 2026 -12328 2576
rect -12262 2026 -12232 2576
rect -12166 2026 -12136 2576
rect -12074 2026 -12044 2576
rect -11582 2026 -11552 2576
rect -11490 2026 -11460 2576
rect -11394 2026 -11364 2576
rect -11298 2026 -11268 2576
rect -11202 2026 -11172 2576
rect -11106 2026 -11076 2576
rect -11010 2026 -10980 2576
rect -10914 2026 -10884 2576
rect -10818 2026 -10788 2576
rect -10722 2026 -10692 2576
rect -10626 2026 -10596 2576
rect -10530 2026 -10500 2576
rect -10434 2026 -10404 2576
rect -10342 2026 -10312 2576
rect -10023 2026 -9993 2576
rect -9931 2026 -9901 2576
rect -9835 2026 -9805 2576
rect -9739 2026 -9709 2576
rect -9643 2026 -9613 2576
rect -9547 2026 -9517 2576
rect -9451 2026 -9421 2576
rect -9355 2026 -9325 2576
rect -9259 2026 -9229 2576
rect -9163 2026 -9133 2576
rect -9067 2026 -9037 2576
rect -8971 2026 -8941 2576
rect -8875 2026 -8845 2576
rect -8783 2026 -8753 2576
rect -8292 2026 -8262 2576
rect -8200 2026 -8170 2576
rect -8104 2026 -8074 2576
rect -8008 2026 -7978 2576
rect -7912 2026 -7882 2576
rect -7816 2026 -7786 2576
rect -7720 2026 -7690 2576
rect -7624 2026 -7594 2576
rect -7528 2026 -7498 2576
rect -7432 2026 -7402 2576
rect -7336 2026 -7306 2576
rect -7240 2026 -7210 2576
rect -7144 2026 -7114 2576
rect -7052 2026 -7022 2576
rect -6733 2026 -6703 2576
rect -6641 2026 -6611 2576
rect -6545 2026 -6515 2576
rect -6449 2026 -6419 2576
rect -6353 2026 -6323 2576
rect -6257 2026 -6227 2576
rect -6161 2026 -6131 2576
rect -6065 2026 -6035 2576
rect -5969 2026 -5939 2576
rect -5873 2026 -5843 2576
rect -5777 2026 -5747 2576
rect -5681 2026 -5651 2576
rect -5585 2026 -5555 2576
rect -5493 2026 -5463 2576
rect -5001 2026 -4971 2576
rect -4909 2026 -4879 2576
rect -4813 2026 -4783 2576
rect -4717 2026 -4687 2576
rect -4621 2026 -4591 2576
rect -4525 2026 -4495 2576
rect -4429 2026 -4399 2576
rect -4333 2026 -4303 2576
rect -4237 2026 -4207 2576
rect -4141 2026 -4111 2576
rect -4045 2026 -4015 2576
rect -3949 2026 -3919 2576
rect -3853 2026 -3823 2576
rect -3761 2026 -3731 2576
rect -3442 2026 -3412 2576
rect -3350 2026 -3320 2576
rect -3254 2026 -3224 2576
rect -3158 2026 -3128 2576
rect -3062 2026 -3032 2576
rect -2966 2026 -2936 2576
rect -2870 2026 -2840 2576
rect -2774 2026 -2744 2576
rect -2678 2026 -2648 2576
rect -2582 2026 -2552 2576
rect -2486 2026 -2456 2576
rect -2390 2026 -2360 2576
rect -2294 2026 -2264 2576
rect -2202 2026 -2172 2576
rect -1710 2026 -1680 2576
rect -1618 2026 -1588 2576
rect -1522 2026 -1492 2576
rect -1426 2026 -1396 2576
rect -1330 2026 -1300 2576
rect -1234 2026 -1204 2576
rect -1138 2026 -1108 2576
rect -1042 2026 -1012 2576
rect -946 2026 -916 2576
rect -850 2026 -820 2576
rect -754 2026 -724 2576
rect -658 2026 -628 2576
rect -562 2026 -532 2576
rect -470 2026 -440 2576
rect -151 2026 -121 2576
rect -59 2026 -29 2576
rect 37 2026 67 2576
rect 133 2026 163 2576
rect 229 2026 259 2576
rect 325 2026 355 2576
rect 421 2026 451 2576
rect 517 2026 547 2576
rect 613 2026 643 2576
rect 709 2026 739 2576
rect 805 2026 835 2576
rect 901 2026 931 2576
rect 997 2026 1027 2576
rect 1089 2026 1119 2576
rect 11835 1753 11865 2009
rect 11931 1753 11961 2009
rect 12027 1753 12057 2009
rect 12123 1753 12153 2009
rect 12219 1753 12249 2009
rect 12315 1753 12345 2009
rect 12411 1753 12441 2009
rect 12507 1753 12537 2009
rect 12603 1753 12633 2009
rect 12699 1753 12729 2009
rect -24535 661 -24505 875
rect -24439 661 -24409 875
rect -24343 661 -24313 875
rect -24247 661 -24217 875
rect -24151 661 -24121 875
rect -24055 661 -24025 875
rect -23426 661 -23396 875
rect -23330 661 -23300 875
rect -23234 661 -23204 875
rect -23138 661 -23108 875
rect -23042 661 -23012 875
rect -22946 661 -22916 875
rect -22544 661 -22514 875
rect -22448 661 -22418 875
rect -22352 661 -22322 875
rect -22256 661 -22226 875
rect -22160 661 -22130 875
rect -22064 661 -22034 875
rect -21244 661 -21214 875
rect -21148 661 -21118 875
rect -21052 661 -21022 875
rect -20956 661 -20926 875
rect -20860 661 -20830 875
rect -20764 661 -20734 875
rect -20135 661 -20105 875
rect -20039 661 -20009 875
rect -19943 661 -19913 875
rect -19847 661 -19817 875
rect -19751 661 -19721 875
rect -19655 661 -19625 875
rect -19253 661 -19223 875
rect -19157 661 -19127 875
rect -19061 661 -19031 875
rect -18965 661 -18935 875
rect -18869 661 -18839 875
rect -18773 661 -18743 875
rect -17953 661 -17923 875
rect -17857 661 -17827 875
rect -17761 661 -17731 875
rect -17665 661 -17635 875
rect -17569 661 -17539 875
rect -17473 661 -17443 875
rect -16844 661 -16814 875
rect -16748 661 -16718 875
rect -16652 661 -16622 875
rect -16556 661 -16526 875
rect -16460 661 -16430 875
rect -16364 661 -16334 875
rect -15962 661 -15932 875
rect -15866 661 -15836 875
rect -15770 661 -15740 875
rect -15674 661 -15644 875
rect -15578 661 -15548 875
rect -15482 661 -15452 875
rect -14662 661 -14632 875
rect -14566 661 -14536 875
rect -14470 661 -14440 875
rect -14374 661 -14344 875
rect -14278 661 -14248 875
rect -14182 661 -14152 875
rect -13553 661 -13523 875
rect -13457 661 -13427 875
rect -13361 661 -13331 875
rect -13265 661 -13235 875
rect -13169 661 -13139 875
rect -13073 661 -13043 875
rect -12671 661 -12641 875
rect -12575 661 -12545 875
rect -12479 661 -12449 875
rect -12383 661 -12353 875
rect -12287 661 -12257 875
rect -12191 661 -12161 875
rect -11371 661 -11341 875
rect -11275 661 -11245 875
rect -11179 661 -11149 875
rect -11083 661 -11053 875
rect -10987 661 -10957 875
rect -10891 661 -10861 875
rect -10262 661 -10232 875
rect -10166 661 -10136 875
rect -10070 661 -10040 875
rect -9974 661 -9944 875
rect -9878 661 -9848 875
rect -9782 661 -9752 875
rect -9380 661 -9350 875
rect -9284 661 -9254 875
rect -9188 661 -9158 875
rect -9092 661 -9062 875
rect -8996 661 -8966 875
rect -8900 661 -8870 875
rect -8081 661 -8051 875
rect -7985 661 -7955 875
rect -7889 661 -7859 875
rect -7793 661 -7763 875
rect -7697 661 -7667 875
rect -7601 661 -7571 875
rect -6972 661 -6942 875
rect -6876 661 -6846 875
rect -6780 661 -6750 875
rect -6684 661 -6654 875
rect -6588 661 -6558 875
rect -6492 661 -6462 875
rect -6090 661 -6060 875
rect -5994 661 -5964 875
rect -5898 661 -5868 875
rect -5802 661 -5772 875
rect -5706 661 -5676 875
rect -5610 661 -5580 875
rect -4790 661 -4760 875
rect -4694 661 -4664 875
rect -4598 661 -4568 875
rect -4502 661 -4472 875
rect -4406 661 -4376 875
rect -4310 661 -4280 875
rect -3681 661 -3651 875
rect -3585 661 -3555 875
rect -3489 661 -3459 875
rect -3393 661 -3363 875
rect -3297 661 -3267 875
rect -3201 661 -3171 875
rect -2799 661 -2769 875
rect -2703 661 -2673 875
rect -2607 661 -2577 875
rect -2511 661 -2481 875
rect -2415 661 -2385 875
rect -2319 661 -2289 875
rect -1499 661 -1469 875
rect -1403 661 -1373 875
rect -1307 661 -1277 875
rect -1211 661 -1181 875
rect -1115 661 -1085 875
rect -1019 661 -989 875
rect -390 661 -360 875
rect -294 661 -264 875
rect -198 661 -168 875
rect -102 661 -72 875
rect -6 661 24 875
rect 90 661 120 875
rect 492 661 522 875
rect 588 661 618 875
rect 684 661 714 875
rect 780 661 810 875
rect 876 661 906 875
rect 972 661 1002 875
rect 12923 1813 13137 1843
rect 12923 1717 13137 1747
rect 12923 1621 13137 1651
rect 7200 33 7230 355
rect 7296 33 7326 355
rect 7392 33 7422 355
rect 7488 33 7518 355
rect 7584 33 7614 355
rect 7680 33 7710 355
rect 7776 33 7806 355
rect 7872 33 7902 355
rect 8148 33 8178 355
rect 8244 33 8274 355
rect 8340 33 8370 355
rect 8436 33 8466 355
rect 8532 33 8562 355
rect 8628 33 8658 355
rect 8724 33 8754 355
rect 8820 33 8850 355
rect 9084 33 9114 355
rect 9180 33 9210 355
rect 9276 33 9306 355
rect 9372 33 9402 355
rect 9468 33 9498 355
rect 9564 33 9594 355
rect 9660 33 9690 355
rect 9756 33 9786 355
rect 10015 34 10045 356
rect 10111 34 10141 356
rect 10207 34 10237 356
rect 10303 34 10333 356
rect 10399 34 10429 356
rect 10495 34 10525 356
rect 10591 34 10621 356
rect 10687 34 10717 356
rect 10942 33 10972 355
rect 11038 33 11068 355
rect 11134 33 11164 355
rect 11230 33 11260 355
rect 11326 33 11356 355
rect 11422 33 11452 355
rect 11518 33 11548 355
rect 11614 33 11644 355
rect 5658 -697 5872 -667
rect 5658 -793 5872 -763
rect 5658 -889 5872 -859
rect 6098 -697 6312 -667
rect 6098 -793 6312 -763
rect 6098 -889 6312 -859
rect 6538 -697 6752 -667
rect 6538 -793 6752 -763
rect 6538 -889 6752 -859
rect 7200 -1631 7230 -1309
rect 7296 -1631 7326 -1309
rect 7392 -1631 7422 -1309
rect 7488 -1631 7518 -1309
rect 7584 -1631 7614 -1309
rect 7680 -1631 7710 -1309
rect 7776 -1631 7806 -1309
rect 7872 -1631 7902 -1309
rect 8148 -1631 8178 -1309
rect 8244 -1631 8274 -1309
rect 8340 -1631 8370 -1309
rect 8436 -1631 8466 -1309
rect 8532 -1631 8562 -1309
rect 8628 -1631 8658 -1309
rect 8724 -1631 8754 -1309
rect 8820 -1631 8850 -1309
rect 9084 -1631 9114 -1309
rect 9180 -1631 9210 -1309
rect 9276 -1631 9306 -1309
rect 9372 -1631 9402 -1309
rect 9468 -1631 9498 -1309
rect 9564 -1631 9594 -1309
rect 9660 -1631 9690 -1309
rect 9756 -1631 9786 -1309
rect 10015 -1631 10045 -1309
rect 10111 -1631 10141 -1309
rect 10207 -1631 10237 -1309
rect 10303 -1631 10333 -1309
rect 10399 -1631 10429 -1309
rect 10495 -1631 10525 -1309
rect 10591 -1631 10621 -1309
rect 10687 -1631 10717 -1309
rect 10942 -1631 10972 -1309
rect 11038 -1631 11068 -1309
rect 11134 -1631 11164 -1309
rect 11230 -1631 11260 -1309
rect 11326 -1631 11356 -1309
rect 11422 -1631 11452 -1309
rect 11518 -1631 11548 -1309
rect 11614 -1631 11644 -1309
rect -24385 -2627 -24355 -2413
rect -24289 -2627 -24259 -2413
rect -24193 -2627 -24163 -2413
rect -24097 -2627 -24067 -2413
rect -24001 -2627 -23971 -2413
rect -23905 -2627 -23875 -2413
rect -23628 -2399 -23414 -2369
rect -23628 -2495 -23414 -2465
rect -23628 -2591 -23414 -2561
rect -22348 -2627 -22318 -2413
rect -22252 -2627 -22222 -2413
rect -22156 -2627 -22126 -2413
rect -22060 -2627 -22030 -2413
rect -21964 -2627 -21934 -2413
rect -21868 -2627 -21838 -2413
rect -21608 -2399 -21394 -2369
rect -21608 -2495 -21394 -2465
rect -21608 -2591 -21394 -2561
rect -20618 -2627 -20588 -2413
rect -20522 -2627 -20492 -2413
rect -20426 -2627 -20396 -2413
rect -20330 -2627 -20300 -2413
rect -20234 -2627 -20204 -2413
rect -20138 -2627 -20108 -2413
rect -19867 -2399 -19653 -2369
rect -19867 -2495 -19653 -2465
rect -19867 -2591 -19653 -2561
rect -18858 -2627 -18828 -2413
rect -18762 -2627 -18732 -2413
rect -18666 -2627 -18636 -2413
rect -18570 -2627 -18540 -2413
rect -18474 -2627 -18444 -2413
rect -18378 -2627 -18348 -2413
rect -18088 -2399 -17874 -2369
rect -18088 -2495 -17874 -2465
rect -18088 -2591 -17874 -2561
rect 11835 -2775 11865 -2519
rect 11931 -2775 11961 -2519
rect 12027 -2775 12057 -2519
rect 12123 -2775 12153 -2519
rect 12219 -2775 12249 -2519
rect 12315 -2775 12345 -2519
rect 12411 -2775 12441 -2519
rect 12507 -2775 12537 -2519
rect 12603 -2775 12633 -2519
rect 12699 -2775 12729 -2519
rect -24334 -4439 -24304 -4225
rect -24238 -4439 -24208 -4225
rect -24142 -4439 -24112 -4225
rect -24046 -4439 -24016 -4225
rect -23950 -4439 -23920 -4225
rect -23854 -4439 -23824 -4225
rect -23584 -4211 -23370 -4181
rect -23584 -4307 -23370 -4277
rect -23584 -4403 -23370 -4373
rect -22598 -4439 -22568 -4225
rect -22502 -4439 -22472 -4225
rect -22406 -4439 -22376 -4225
rect -22310 -4439 -22280 -4225
rect -22214 -4439 -22184 -4225
rect -22118 -4439 -22088 -4225
rect -21846 -4211 -21632 -4181
rect -21846 -4307 -21632 -4277
rect -21846 -4403 -21632 -4373
rect -20679 -4534 -20649 -3984
rect -20587 -4534 -20557 -3984
rect -20491 -4534 -20461 -3984
rect -20395 -4534 -20365 -3984
rect -20299 -4534 -20269 -3984
rect -20203 -4534 -20173 -3984
rect -20107 -4534 -20077 -3984
rect -20011 -4534 -19981 -3984
rect -19915 -4534 -19885 -3984
rect -19819 -4534 -19789 -3984
rect -19723 -4534 -19693 -3984
rect -19627 -4534 -19597 -3984
rect -19531 -4534 -19501 -3984
rect -19439 -4534 -19409 -3984
rect -19120 -4534 -19090 -3984
rect -19028 -4534 -18998 -3984
rect -18932 -4534 -18902 -3984
rect -18836 -4534 -18806 -3984
rect -18740 -4534 -18710 -3984
rect -18644 -4534 -18614 -3984
rect -18548 -4534 -18518 -3984
rect -18452 -4534 -18422 -3984
rect -18356 -4534 -18326 -3984
rect -18260 -4534 -18230 -3984
rect -18164 -4534 -18134 -3984
rect -18068 -4534 -18038 -3984
rect -17972 -4534 -17942 -3984
rect -17880 -4534 -17850 -3984
rect -17388 -4534 -17358 -3984
rect -17296 -4534 -17266 -3984
rect -17200 -4534 -17170 -3984
rect -17104 -4534 -17074 -3984
rect -17008 -4534 -16978 -3984
rect -16912 -4534 -16882 -3984
rect -16816 -4534 -16786 -3984
rect -16720 -4534 -16690 -3984
rect -16624 -4534 -16594 -3984
rect -16528 -4534 -16498 -3984
rect -16432 -4534 -16402 -3984
rect -16336 -4534 -16306 -3984
rect -16240 -4534 -16210 -3984
rect -16148 -4534 -16118 -3984
rect -15829 -4534 -15799 -3984
rect -15737 -4534 -15707 -3984
rect -15641 -4534 -15611 -3984
rect -15545 -4534 -15515 -3984
rect -15449 -4534 -15419 -3984
rect -15353 -4534 -15323 -3984
rect -15257 -4534 -15227 -3984
rect -15161 -4534 -15131 -3984
rect -15065 -4534 -15035 -3984
rect -14969 -4534 -14939 -3984
rect -14873 -4534 -14843 -3984
rect -14777 -4534 -14747 -3984
rect -14681 -4534 -14651 -3984
rect -14589 -4534 -14559 -3984
rect -14097 -4534 -14067 -3984
rect -14005 -4534 -13975 -3984
rect -13909 -4534 -13879 -3984
rect -13813 -4534 -13783 -3984
rect -13717 -4534 -13687 -3984
rect -13621 -4534 -13591 -3984
rect -13525 -4534 -13495 -3984
rect -13429 -4534 -13399 -3984
rect -13333 -4534 -13303 -3984
rect -13237 -4534 -13207 -3984
rect -13141 -4534 -13111 -3984
rect -13045 -4534 -13015 -3984
rect -12949 -4534 -12919 -3984
rect -12857 -4534 -12827 -3984
rect -12538 -4534 -12508 -3984
rect -12446 -4534 -12416 -3984
rect -12350 -4534 -12320 -3984
rect -12254 -4534 -12224 -3984
rect -12158 -4534 -12128 -3984
rect -12062 -4534 -12032 -3984
rect -11966 -4534 -11936 -3984
rect -11870 -4534 -11840 -3984
rect -11774 -4534 -11744 -3984
rect -11678 -4534 -11648 -3984
rect -11582 -4534 -11552 -3984
rect -11486 -4534 -11456 -3984
rect -11390 -4534 -11360 -3984
rect -11298 -4534 -11268 -3984
rect -10806 -4534 -10776 -3984
rect -10714 -4534 -10684 -3984
rect -10618 -4534 -10588 -3984
rect -10522 -4534 -10492 -3984
rect -10426 -4534 -10396 -3984
rect -10330 -4534 -10300 -3984
rect -10234 -4534 -10204 -3984
rect -10138 -4534 -10108 -3984
rect -10042 -4534 -10012 -3984
rect -9946 -4534 -9916 -3984
rect -9850 -4534 -9820 -3984
rect -9754 -4534 -9724 -3984
rect -9658 -4534 -9628 -3984
rect -9566 -4534 -9536 -3984
rect -9247 -4534 -9217 -3984
rect -9155 -4534 -9125 -3984
rect -9059 -4534 -9029 -3984
rect -8963 -4534 -8933 -3984
rect -8867 -4534 -8837 -3984
rect -8771 -4534 -8741 -3984
rect -8675 -4534 -8645 -3984
rect -8579 -4534 -8549 -3984
rect -8483 -4534 -8453 -3984
rect -8387 -4534 -8357 -3984
rect -8291 -4534 -8261 -3984
rect -8195 -4534 -8165 -3984
rect -8099 -4534 -8069 -3984
rect -8007 -4534 -7977 -3984
rect 12923 -2715 13137 -2685
rect 12923 -2811 13137 -2781
rect 12923 -2907 13137 -2877
rect 7200 -4495 7230 -4173
rect 7296 -4495 7326 -4173
rect 7392 -4495 7422 -4173
rect 7488 -4495 7518 -4173
rect 7584 -4495 7614 -4173
rect 7680 -4495 7710 -4173
rect 7776 -4495 7806 -4173
rect 7872 -4495 7902 -4173
rect 8148 -4495 8178 -4173
rect 8244 -4495 8274 -4173
rect 8340 -4495 8370 -4173
rect 8436 -4495 8466 -4173
rect 8532 -4495 8562 -4173
rect 8628 -4495 8658 -4173
rect 8724 -4495 8754 -4173
rect 8820 -4495 8850 -4173
rect 9084 -4495 9114 -4173
rect 9180 -4495 9210 -4173
rect 9276 -4495 9306 -4173
rect 9372 -4495 9402 -4173
rect 9468 -4495 9498 -4173
rect 9564 -4495 9594 -4173
rect 9660 -4495 9690 -4173
rect 9756 -4495 9786 -4173
rect 10015 -4494 10045 -4172
rect 10111 -4494 10141 -4172
rect 10207 -4494 10237 -4172
rect 10303 -4494 10333 -4172
rect 10399 -4494 10429 -4172
rect 10495 -4494 10525 -4172
rect 10591 -4494 10621 -4172
rect 10687 -4494 10717 -4172
rect 10942 -4495 10972 -4173
rect 11038 -4495 11068 -4173
rect 11134 -4495 11164 -4173
rect 11230 -4495 11260 -4173
rect 11326 -4495 11356 -4173
rect 11422 -4495 11452 -4173
rect 11518 -4495 11548 -4173
rect 11614 -4495 11644 -4173
rect 5658 -5125 5872 -5095
rect 5658 -5221 5872 -5191
rect 5658 -5317 5872 -5287
rect 6098 -5125 6312 -5095
rect 6098 -5221 6312 -5191
rect 6098 -5317 6312 -5287
rect 6538 -5125 6752 -5095
rect 6538 -5221 6752 -5191
rect 6538 -5317 6752 -5287
rect -24334 -5731 -24304 -5517
rect -24238 -5731 -24208 -5517
rect -24142 -5731 -24112 -5517
rect -24046 -5731 -24016 -5517
rect -23950 -5731 -23920 -5517
rect -23854 -5731 -23824 -5517
rect -23586 -5503 -23372 -5473
rect -23586 -5599 -23372 -5569
rect -23586 -5695 -23372 -5665
rect -22598 -5731 -22568 -5517
rect -22502 -5731 -22472 -5517
rect -22406 -5731 -22376 -5517
rect -22310 -5731 -22280 -5517
rect -22214 -5731 -22184 -5517
rect -22118 -5731 -22088 -5517
rect -21852 -5503 -21638 -5473
rect -21852 -5599 -21638 -5569
rect -21852 -5695 -21638 -5665
rect -20468 -5899 -20438 -5685
rect -20372 -5899 -20342 -5685
rect -20276 -5899 -20246 -5685
rect -20180 -5899 -20150 -5685
rect -20084 -5899 -20054 -5685
rect -19988 -5899 -19958 -5685
rect -19359 -5899 -19329 -5685
rect -19263 -5899 -19233 -5685
rect -19167 -5899 -19137 -5685
rect -19071 -5899 -19041 -5685
rect -18975 -5899 -18945 -5685
rect -18879 -5899 -18849 -5685
rect -18477 -5899 -18447 -5685
rect -18381 -5899 -18351 -5685
rect -18285 -5899 -18255 -5685
rect -18189 -5899 -18159 -5685
rect -18093 -5899 -18063 -5685
rect -17997 -5899 -17967 -5685
rect -17177 -5899 -17147 -5685
rect -17081 -5899 -17051 -5685
rect -16985 -5899 -16955 -5685
rect -16889 -5899 -16859 -5685
rect -16793 -5899 -16763 -5685
rect -16697 -5899 -16667 -5685
rect -16068 -5899 -16038 -5685
rect -15972 -5899 -15942 -5685
rect -15876 -5899 -15846 -5685
rect -15780 -5899 -15750 -5685
rect -15684 -5899 -15654 -5685
rect -15588 -5899 -15558 -5685
rect -15186 -5899 -15156 -5685
rect -15090 -5899 -15060 -5685
rect -14994 -5899 -14964 -5685
rect -14898 -5899 -14868 -5685
rect -14802 -5899 -14772 -5685
rect -14706 -5899 -14676 -5685
rect -13886 -5899 -13856 -5685
rect -13790 -5899 -13760 -5685
rect -13694 -5899 -13664 -5685
rect -13598 -5899 -13568 -5685
rect -13502 -5899 -13472 -5685
rect -13406 -5899 -13376 -5685
rect -12777 -5899 -12747 -5685
rect -12681 -5899 -12651 -5685
rect -12585 -5899 -12555 -5685
rect -12489 -5899 -12459 -5685
rect -12393 -5899 -12363 -5685
rect -12297 -5899 -12267 -5685
rect -11895 -5899 -11865 -5685
rect -11799 -5899 -11769 -5685
rect -11703 -5899 -11673 -5685
rect -11607 -5899 -11577 -5685
rect -11511 -5899 -11481 -5685
rect -11415 -5899 -11385 -5685
rect -10595 -5899 -10565 -5685
rect -10499 -5899 -10469 -5685
rect -10403 -5899 -10373 -5685
rect -10307 -5899 -10277 -5685
rect -10211 -5899 -10181 -5685
rect -10115 -5899 -10085 -5685
rect -9486 -5899 -9456 -5685
rect -9390 -5899 -9360 -5685
rect -9294 -5899 -9264 -5685
rect -9198 -5899 -9168 -5685
rect -9102 -5899 -9072 -5685
rect -9006 -5899 -8976 -5685
rect -8604 -5899 -8574 -5685
rect -8508 -5899 -8478 -5685
rect -8412 -5899 -8382 -5685
rect -8316 -5899 -8286 -5685
rect -8220 -5899 -8190 -5685
rect -8124 -5899 -8094 -5685
rect 7200 -6059 7230 -5737
rect 7296 -6059 7326 -5737
rect 7392 -6059 7422 -5737
rect 7488 -6059 7518 -5737
rect 7584 -6059 7614 -5737
rect 7680 -6059 7710 -5737
rect 7776 -6059 7806 -5737
rect 7872 -6059 7902 -5737
rect 8148 -6059 8178 -5737
rect 8244 -6059 8274 -5737
rect 8340 -6059 8370 -5737
rect 8436 -6059 8466 -5737
rect 8532 -6059 8562 -5737
rect 8628 -6059 8658 -5737
rect 8724 -6059 8754 -5737
rect 8820 -6059 8850 -5737
rect 9084 -6059 9114 -5737
rect 9180 -6059 9210 -5737
rect 9276 -6059 9306 -5737
rect 9372 -6059 9402 -5737
rect 9468 -6059 9498 -5737
rect 9564 -6059 9594 -5737
rect 9660 -6059 9690 -5737
rect 9756 -6059 9786 -5737
rect 10015 -6059 10045 -5737
rect 10111 -6059 10141 -5737
rect 10207 -6059 10237 -5737
rect 10303 -6059 10333 -5737
rect 10399 -6059 10429 -5737
rect 10495 -6059 10525 -5737
rect 10591 -6059 10621 -5737
rect 10687 -6059 10717 -5737
rect 10942 -6059 10972 -5737
rect 11038 -6059 11068 -5737
rect 11134 -6059 11164 -5737
rect 11230 -6059 11260 -5737
rect 11326 -6059 11356 -5737
rect 11422 -6059 11452 -5737
rect 11518 -6059 11548 -5737
rect 11614 -6059 11644 -5737
rect -24334 -7704 -24304 -7490
rect -24238 -7704 -24208 -7490
rect -24142 -7704 -24112 -7490
rect -24046 -7704 -24016 -7490
rect -23950 -7704 -23920 -7490
rect -23854 -7704 -23824 -7490
rect -23584 -7476 -23370 -7446
rect -23584 -7572 -23370 -7542
rect -23584 -7668 -23370 -7638
rect -22597 -7704 -22567 -7490
rect -22501 -7704 -22471 -7490
rect -22405 -7704 -22375 -7490
rect -22309 -7704 -22279 -7490
rect -22213 -7704 -22183 -7490
rect -22117 -7704 -22087 -7490
rect -21850 -7476 -21636 -7446
rect -21850 -7572 -21636 -7542
rect -21850 -7668 -21636 -7638
rect -20679 -7799 -20649 -7249
rect -20587 -7799 -20557 -7249
rect -20491 -7799 -20461 -7249
rect -20395 -7799 -20365 -7249
rect -20299 -7799 -20269 -7249
rect -20203 -7799 -20173 -7249
rect -20107 -7799 -20077 -7249
rect -20011 -7799 -19981 -7249
rect -19915 -7799 -19885 -7249
rect -19819 -7799 -19789 -7249
rect -19723 -7799 -19693 -7249
rect -19627 -7799 -19597 -7249
rect -19531 -7799 -19501 -7249
rect -19439 -7799 -19409 -7249
rect -19120 -7799 -19090 -7249
rect -19028 -7799 -18998 -7249
rect -18932 -7799 -18902 -7249
rect -18836 -7799 -18806 -7249
rect -18740 -7799 -18710 -7249
rect -18644 -7799 -18614 -7249
rect -18548 -7799 -18518 -7249
rect -18452 -7799 -18422 -7249
rect -18356 -7799 -18326 -7249
rect -18260 -7799 -18230 -7249
rect -18164 -7799 -18134 -7249
rect -18068 -7799 -18038 -7249
rect -17972 -7799 -17942 -7249
rect -17880 -7799 -17850 -7249
rect -17388 -7799 -17358 -7249
rect -17296 -7799 -17266 -7249
rect -17200 -7799 -17170 -7249
rect -17104 -7799 -17074 -7249
rect -17008 -7799 -16978 -7249
rect -16912 -7799 -16882 -7249
rect -16816 -7799 -16786 -7249
rect -16720 -7799 -16690 -7249
rect -16624 -7799 -16594 -7249
rect -16528 -7799 -16498 -7249
rect -16432 -7799 -16402 -7249
rect -16336 -7799 -16306 -7249
rect -16240 -7799 -16210 -7249
rect -16148 -7799 -16118 -7249
rect -15829 -7799 -15799 -7249
rect -15737 -7799 -15707 -7249
rect -15641 -7799 -15611 -7249
rect -15545 -7799 -15515 -7249
rect -15449 -7799 -15419 -7249
rect -15353 -7799 -15323 -7249
rect -15257 -7799 -15227 -7249
rect -15161 -7799 -15131 -7249
rect -15065 -7799 -15035 -7249
rect -14969 -7799 -14939 -7249
rect -14873 -7799 -14843 -7249
rect -14777 -7799 -14747 -7249
rect -14681 -7799 -14651 -7249
rect -14589 -7799 -14559 -7249
rect -14097 -7799 -14067 -7249
rect -14005 -7799 -13975 -7249
rect -13909 -7799 -13879 -7249
rect -13813 -7799 -13783 -7249
rect -13717 -7799 -13687 -7249
rect -13621 -7799 -13591 -7249
rect -13525 -7799 -13495 -7249
rect -13429 -7799 -13399 -7249
rect -13333 -7799 -13303 -7249
rect -13237 -7799 -13207 -7249
rect -13141 -7799 -13111 -7249
rect -13045 -7799 -13015 -7249
rect -12949 -7799 -12919 -7249
rect -12857 -7799 -12827 -7249
rect -12538 -7799 -12508 -7249
rect -12446 -7799 -12416 -7249
rect -12350 -7799 -12320 -7249
rect -12254 -7799 -12224 -7249
rect -12158 -7799 -12128 -7249
rect -12062 -7799 -12032 -7249
rect -11966 -7799 -11936 -7249
rect -11870 -7799 -11840 -7249
rect -11774 -7799 -11744 -7249
rect -11678 -7799 -11648 -7249
rect -11582 -7799 -11552 -7249
rect -11486 -7799 -11456 -7249
rect -11390 -7799 -11360 -7249
rect -11298 -7799 -11268 -7249
rect -10806 -7799 -10776 -7249
rect -10714 -7799 -10684 -7249
rect -10618 -7799 -10588 -7249
rect -10522 -7799 -10492 -7249
rect -10426 -7799 -10396 -7249
rect -10330 -7799 -10300 -7249
rect -10234 -7799 -10204 -7249
rect -10138 -7799 -10108 -7249
rect -10042 -7799 -10012 -7249
rect -9946 -7799 -9916 -7249
rect -9850 -7799 -9820 -7249
rect -9754 -7799 -9724 -7249
rect -9658 -7799 -9628 -7249
rect -9566 -7799 -9536 -7249
rect -9247 -7799 -9217 -7249
rect -9155 -7799 -9125 -7249
rect -9059 -7799 -9029 -7249
rect -8963 -7799 -8933 -7249
rect -8867 -7799 -8837 -7249
rect -8771 -7799 -8741 -7249
rect -8675 -7799 -8645 -7249
rect -8579 -7799 -8549 -7249
rect -8483 -7799 -8453 -7249
rect -8387 -7799 -8357 -7249
rect -8291 -7799 -8261 -7249
rect -8195 -7799 -8165 -7249
rect -8099 -7799 -8069 -7249
rect -8007 -7799 -7977 -7249
rect 11835 -7203 11865 -6947
rect 11931 -7203 11961 -6947
rect 12027 -7203 12057 -6947
rect 12123 -7203 12153 -6947
rect 12219 -7203 12249 -6947
rect 12315 -7203 12345 -6947
rect 12411 -7203 12441 -6947
rect 12507 -7203 12537 -6947
rect 12603 -7203 12633 -6947
rect 12699 -7203 12729 -6947
rect 12923 -7143 13137 -7113
rect 12923 -7239 13137 -7209
rect 12923 -7335 13137 -7305
rect -24334 -8996 -24304 -8782
rect -24238 -8996 -24208 -8782
rect -24142 -8996 -24112 -8782
rect -24046 -8996 -24016 -8782
rect -23950 -8996 -23920 -8782
rect -23854 -8996 -23824 -8782
rect -23583 -8768 -23369 -8738
rect -23583 -8864 -23369 -8834
rect -23583 -8960 -23369 -8930
rect -22598 -8996 -22568 -8782
rect -22502 -8996 -22472 -8782
rect -22406 -8996 -22376 -8782
rect -22310 -8996 -22280 -8782
rect -22214 -8996 -22184 -8782
rect -22118 -8996 -22088 -8782
rect -21846 -8768 -21632 -8738
rect -21846 -8864 -21632 -8834
rect -21846 -8960 -21632 -8930
rect 7200 -8923 7230 -8601
rect 7296 -8923 7326 -8601
rect 7392 -8923 7422 -8601
rect 7488 -8923 7518 -8601
rect 7584 -8923 7614 -8601
rect 7680 -8923 7710 -8601
rect 7776 -8923 7806 -8601
rect 7872 -8923 7902 -8601
rect 8148 -8923 8178 -8601
rect 8244 -8923 8274 -8601
rect 8340 -8923 8370 -8601
rect 8436 -8923 8466 -8601
rect 8532 -8923 8562 -8601
rect 8628 -8923 8658 -8601
rect 8724 -8923 8754 -8601
rect 8820 -8923 8850 -8601
rect 9084 -8923 9114 -8601
rect 9180 -8923 9210 -8601
rect 9276 -8923 9306 -8601
rect 9372 -8923 9402 -8601
rect 9468 -8923 9498 -8601
rect 9564 -8923 9594 -8601
rect 9660 -8923 9690 -8601
rect 9756 -8923 9786 -8601
rect 10015 -8922 10045 -8600
rect 10111 -8922 10141 -8600
rect 10207 -8922 10237 -8600
rect 10303 -8922 10333 -8600
rect 10399 -8922 10429 -8600
rect 10495 -8922 10525 -8600
rect 10591 -8922 10621 -8600
rect 10687 -8922 10717 -8600
rect 10942 -8923 10972 -8601
rect 11038 -8923 11068 -8601
rect 11134 -8923 11164 -8601
rect 11230 -8923 11260 -8601
rect 11326 -8923 11356 -8601
rect 11422 -8923 11452 -8601
rect 11518 -8923 11548 -8601
rect 11614 -8923 11644 -8601
rect -20468 -9164 -20438 -8950
rect -20372 -9164 -20342 -8950
rect -20276 -9164 -20246 -8950
rect -20180 -9164 -20150 -8950
rect -20084 -9164 -20054 -8950
rect -19988 -9164 -19958 -8950
rect -19359 -9164 -19329 -8950
rect -19263 -9164 -19233 -8950
rect -19167 -9164 -19137 -8950
rect -19071 -9164 -19041 -8950
rect -18975 -9164 -18945 -8950
rect -18879 -9164 -18849 -8950
rect -18477 -9164 -18447 -8950
rect -18381 -9164 -18351 -8950
rect -18285 -9164 -18255 -8950
rect -18189 -9164 -18159 -8950
rect -18093 -9164 -18063 -8950
rect -17997 -9164 -17967 -8950
rect -17177 -9164 -17147 -8950
rect -17081 -9164 -17051 -8950
rect -16985 -9164 -16955 -8950
rect -16889 -9164 -16859 -8950
rect -16793 -9164 -16763 -8950
rect -16697 -9164 -16667 -8950
rect -16068 -9164 -16038 -8950
rect -15972 -9164 -15942 -8950
rect -15876 -9164 -15846 -8950
rect -15780 -9164 -15750 -8950
rect -15684 -9164 -15654 -8950
rect -15588 -9164 -15558 -8950
rect -15186 -9164 -15156 -8950
rect -15090 -9164 -15060 -8950
rect -14994 -9164 -14964 -8950
rect -14898 -9164 -14868 -8950
rect -14802 -9164 -14772 -8950
rect -14706 -9164 -14676 -8950
rect -13886 -9164 -13856 -8950
rect -13790 -9164 -13760 -8950
rect -13694 -9164 -13664 -8950
rect -13598 -9164 -13568 -8950
rect -13502 -9164 -13472 -8950
rect -13406 -9164 -13376 -8950
rect -12777 -9164 -12747 -8950
rect -12681 -9164 -12651 -8950
rect -12585 -9164 -12555 -8950
rect -12489 -9164 -12459 -8950
rect -12393 -9164 -12363 -8950
rect -12297 -9164 -12267 -8950
rect -11895 -9164 -11865 -8950
rect -11799 -9164 -11769 -8950
rect -11703 -9164 -11673 -8950
rect -11607 -9164 -11577 -8950
rect -11511 -9164 -11481 -8950
rect -11415 -9164 -11385 -8950
rect -10595 -9164 -10565 -8950
rect -10499 -9164 -10469 -8950
rect -10403 -9164 -10373 -8950
rect -10307 -9164 -10277 -8950
rect -10211 -9164 -10181 -8950
rect -10115 -9164 -10085 -8950
rect -9486 -9164 -9456 -8950
rect -9390 -9164 -9360 -8950
rect -9294 -9164 -9264 -8950
rect -9198 -9164 -9168 -8950
rect -9102 -9164 -9072 -8950
rect -9006 -9164 -8976 -8950
rect -8604 -9164 -8574 -8950
rect -8508 -9164 -8478 -8950
rect -8412 -9164 -8382 -8950
rect -8316 -9164 -8286 -8950
rect -8220 -9164 -8190 -8950
rect -8124 -9164 -8094 -8950
rect 5658 -9753 5872 -9723
rect 5658 -9849 5872 -9819
rect 5658 -9945 5872 -9915
rect 6098 -9753 6312 -9723
rect 6098 -9849 6312 -9819
rect 6098 -9945 6312 -9915
rect 6538 -9753 6752 -9723
rect 6538 -9849 6752 -9819
rect 6538 -9945 6752 -9915
rect -24334 -10968 -24304 -10754
rect -24238 -10968 -24208 -10754
rect -24142 -10968 -24112 -10754
rect -24046 -10968 -24016 -10754
rect -23950 -10968 -23920 -10754
rect -23854 -10968 -23824 -10754
rect -23583 -10740 -23369 -10710
rect -23583 -10836 -23369 -10806
rect -23583 -10932 -23369 -10902
rect -22597 -10968 -22567 -10754
rect -22501 -10968 -22471 -10754
rect -22405 -10968 -22375 -10754
rect -22309 -10968 -22279 -10754
rect -22213 -10968 -22183 -10754
rect -22117 -10968 -22087 -10754
rect -21850 -10740 -21636 -10710
rect -21850 -10836 -21636 -10806
rect -21850 -10932 -21636 -10902
rect -20679 -11063 -20649 -10513
rect -20587 -11063 -20557 -10513
rect -20491 -11063 -20461 -10513
rect -20395 -11063 -20365 -10513
rect -20299 -11063 -20269 -10513
rect -20203 -11063 -20173 -10513
rect -20107 -11063 -20077 -10513
rect -20011 -11063 -19981 -10513
rect -19915 -11063 -19885 -10513
rect -19819 -11063 -19789 -10513
rect -19723 -11063 -19693 -10513
rect -19627 -11063 -19597 -10513
rect -19531 -11063 -19501 -10513
rect -19439 -11063 -19409 -10513
rect -19120 -11063 -19090 -10513
rect -19028 -11063 -18998 -10513
rect -18932 -11063 -18902 -10513
rect -18836 -11063 -18806 -10513
rect -18740 -11063 -18710 -10513
rect -18644 -11063 -18614 -10513
rect -18548 -11063 -18518 -10513
rect -18452 -11063 -18422 -10513
rect -18356 -11063 -18326 -10513
rect -18260 -11063 -18230 -10513
rect -18164 -11063 -18134 -10513
rect -18068 -11063 -18038 -10513
rect -17972 -11063 -17942 -10513
rect -17880 -11063 -17850 -10513
rect -17388 -11063 -17358 -10513
rect -17296 -11063 -17266 -10513
rect -17200 -11063 -17170 -10513
rect -17104 -11063 -17074 -10513
rect -17008 -11063 -16978 -10513
rect -16912 -11063 -16882 -10513
rect -16816 -11063 -16786 -10513
rect -16720 -11063 -16690 -10513
rect -16624 -11063 -16594 -10513
rect -16528 -11063 -16498 -10513
rect -16432 -11063 -16402 -10513
rect -16336 -11063 -16306 -10513
rect -16240 -11063 -16210 -10513
rect -16148 -11063 -16118 -10513
rect -15829 -11063 -15799 -10513
rect -15737 -11063 -15707 -10513
rect -15641 -11063 -15611 -10513
rect -15545 -11063 -15515 -10513
rect -15449 -11063 -15419 -10513
rect -15353 -11063 -15323 -10513
rect -15257 -11063 -15227 -10513
rect -15161 -11063 -15131 -10513
rect -15065 -11063 -15035 -10513
rect -14969 -11063 -14939 -10513
rect -14873 -11063 -14843 -10513
rect -14777 -11063 -14747 -10513
rect -14681 -11063 -14651 -10513
rect -14589 -11063 -14559 -10513
rect -14097 -11063 -14067 -10513
rect -14005 -11063 -13975 -10513
rect -13909 -11063 -13879 -10513
rect -13813 -11063 -13783 -10513
rect -13717 -11063 -13687 -10513
rect -13621 -11063 -13591 -10513
rect -13525 -11063 -13495 -10513
rect -13429 -11063 -13399 -10513
rect -13333 -11063 -13303 -10513
rect -13237 -11063 -13207 -10513
rect -13141 -11063 -13111 -10513
rect -13045 -11063 -13015 -10513
rect -12949 -11063 -12919 -10513
rect -12857 -11063 -12827 -10513
rect -12538 -11063 -12508 -10513
rect -12446 -11063 -12416 -10513
rect -12350 -11063 -12320 -10513
rect -12254 -11063 -12224 -10513
rect -12158 -11063 -12128 -10513
rect -12062 -11063 -12032 -10513
rect -11966 -11063 -11936 -10513
rect -11870 -11063 -11840 -10513
rect -11774 -11063 -11744 -10513
rect -11678 -11063 -11648 -10513
rect -11582 -11063 -11552 -10513
rect -11486 -11063 -11456 -10513
rect -11390 -11063 -11360 -10513
rect -11298 -11063 -11268 -10513
rect -10806 -11063 -10776 -10513
rect -10714 -11063 -10684 -10513
rect -10618 -11063 -10588 -10513
rect -10522 -11063 -10492 -10513
rect -10426 -11063 -10396 -10513
rect -10330 -11063 -10300 -10513
rect -10234 -11063 -10204 -10513
rect -10138 -11063 -10108 -10513
rect -10042 -11063 -10012 -10513
rect -9946 -11063 -9916 -10513
rect -9850 -11063 -9820 -10513
rect -9754 -11063 -9724 -10513
rect -9658 -11063 -9628 -10513
rect -9566 -11063 -9536 -10513
rect -9247 -11063 -9217 -10513
rect -9155 -11063 -9125 -10513
rect -9059 -11063 -9029 -10513
rect -8963 -11063 -8933 -10513
rect -8867 -11063 -8837 -10513
rect -8771 -11063 -8741 -10513
rect -8675 -11063 -8645 -10513
rect -8579 -11063 -8549 -10513
rect -8483 -11063 -8453 -10513
rect -8387 -11063 -8357 -10513
rect -8291 -11063 -8261 -10513
rect -8195 -11063 -8165 -10513
rect -8099 -11063 -8069 -10513
rect -8007 -11063 -7977 -10513
rect 7200 -10687 7230 -10365
rect 7296 -10687 7326 -10365
rect 7392 -10687 7422 -10365
rect 7488 -10687 7518 -10365
rect 7584 -10687 7614 -10365
rect 7680 -10687 7710 -10365
rect 7776 -10687 7806 -10365
rect 7872 -10687 7902 -10365
rect 8148 -10687 8178 -10365
rect 8244 -10687 8274 -10365
rect 8340 -10687 8370 -10365
rect 8436 -10687 8466 -10365
rect 8532 -10687 8562 -10365
rect 8628 -10687 8658 -10365
rect 8724 -10687 8754 -10365
rect 8820 -10687 8850 -10365
rect 9084 -10687 9114 -10365
rect 9180 -10687 9210 -10365
rect 9276 -10687 9306 -10365
rect 9372 -10687 9402 -10365
rect 9468 -10687 9498 -10365
rect 9564 -10687 9594 -10365
rect 9660 -10687 9690 -10365
rect 9756 -10687 9786 -10365
rect 10015 -10687 10045 -10365
rect 10111 -10687 10141 -10365
rect 10207 -10687 10237 -10365
rect 10303 -10687 10333 -10365
rect 10399 -10687 10429 -10365
rect 10495 -10687 10525 -10365
rect 10591 -10687 10621 -10365
rect 10687 -10687 10717 -10365
rect 10942 -10687 10972 -10365
rect 11038 -10687 11068 -10365
rect 11134 -10687 11164 -10365
rect 11230 -10687 11260 -10365
rect 11326 -10687 11356 -10365
rect 11422 -10687 11452 -10365
rect 11518 -10687 11548 -10365
rect 11614 -10687 11644 -10365
rect 11835 -11831 11865 -11575
rect 11931 -11831 11961 -11575
rect 12027 -11831 12057 -11575
rect 12123 -11831 12153 -11575
rect 12219 -11831 12249 -11575
rect 12315 -11831 12345 -11575
rect 12411 -11831 12441 -11575
rect 12507 -11831 12537 -11575
rect 12603 -11831 12633 -11575
rect 12699 -11831 12729 -11575
rect -24334 -12260 -24304 -12046
rect -24238 -12260 -24208 -12046
rect -24142 -12260 -24112 -12046
rect -24046 -12260 -24016 -12046
rect -23950 -12260 -23920 -12046
rect -23854 -12260 -23824 -12046
rect -23583 -12032 -23369 -12002
rect -23583 -12128 -23369 -12098
rect -23583 -12224 -23369 -12194
rect -22597 -12260 -22567 -12046
rect -22501 -12260 -22471 -12046
rect -22405 -12260 -22375 -12046
rect -22309 -12260 -22279 -12046
rect -22213 -12260 -22183 -12046
rect -22117 -12260 -22087 -12046
rect -21854 -12032 -21640 -12002
rect -21854 -12128 -21640 -12098
rect -21854 -12224 -21640 -12194
rect -20468 -12428 -20438 -12214
rect -20372 -12428 -20342 -12214
rect -20276 -12428 -20246 -12214
rect -20180 -12428 -20150 -12214
rect -20084 -12428 -20054 -12214
rect -19988 -12428 -19958 -12214
rect -19359 -12428 -19329 -12214
rect -19263 -12428 -19233 -12214
rect -19167 -12428 -19137 -12214
rect -19071 -12428 -19041 -12214
rect -18975 -12428 -18945 -12214
rect -18879 -12428 -18849 -12214
rect -18477 -12428 -18447 -12214
rect -18381 -12428 -18351 -12214
rect -18285 -12428 -18255 -12214
rect -18189 -12428 -18159 -12214
rect -18093 -12428 -18063 -12214
rect -17997 -12428 -17967 -12214
rect -17177 -12428 -17147 -12214
rect -17081 -12428 -17051 -12214
rect -16985 -12428 -16955 -12214
rect -16889 -12428 -16859 -12214
rect -16793 -12428 -16763 -12214
rect -16697 -12428 -16667 -12214
rect -16068 -12428 -16038 -12214
rect -15972 -12428 -15942 -12214
rect -15876 -12428 -15846 -12214
rect -15780 -12428 -15750 -12214
rect -15684 -12428 -15654 -12214
rect -15588 -12428 -15558 -12214
rect -15186 -12428 -15156 -12214
rect -15090 -12428 -15060 -12214
rect -14994 -12428 -14964 -12214
rect -14898 -12428 -14868 -12214
rect -14802 -12428 -14772 -12214
rect -14706 -12428 -14676 -12214
rect -13886 -12428 -13856 -12214
rect -13790 -12428 -13760 -12214
rect -13694 -12428 -13664 -12214
rect -13598 -12428 -13568 -12214
rect -13502 -12428 -13472 -12214
rect -13406 -12428 -13376 -12214
rect -12777 -12428 -12747 -12214
rect -12681 -12428 -12651 -12214
rect -12585 -12428 -12555 -12214
rect -12489 -12428 -12459 -12214
rect -12393 -12428 -12363 -12214
rect -12297 -12428 -12267 -12214
rect -11895 -12428 -11865 -12214
rect -11799 -12428 -11769 -12214
rect -11703 -12428 -11673 -12214
rect -11607 -12428 -11577 -12214
rect -11511 -12428 -11481 -12214
rect -11415 -12428 -11385 -12214
rect -10595 -12428 -10565 -12214
rect -10499 -12428 -10469 -12214
rect -10403 -12428 -10373 -12214
rect -10307 -12428 -10277 -12214
rect -10211 -12428 -10181 -12214
rect -10115 -12428 -10085 -12214
rect -9486 -12428 -9456 -12214
rect -9390 -12428 -9360 -12214
rect -9294 -12428 -9264 -12214
rect -9198 -12428 -9168 -12214
rect -9102 -12428 -9072 -12214
rect -9006 -12428 -8976 -12214
rect -8604 -12428 -8574 -12214
rect -8508 -12428 -8478 -12214
rect -8412 -12428 -8382 -12214
rect -8316 -12428 -8286 -12214
rect -8220 -12428 -8190 -12214
rect -8124 -12428 -8094 -12214
rect 12923 -11771 13137 -11741
rect 12923 -11867 13137 -11837
rect 12923 -11963 13137 -11933
rect 7200 -13551 7230 -13229
rect 7296 -13551 7326 -13229
rect 7392 -13551 7422 -13229
rect 7488 -13551 7518 -13229
rect 7584 -13551 7614 -13229
rect 7680 -13551 7710 -13229
rect 7776 -13551 7806 -13229
rect 7872 -13551 7902 -13229
rect 8148 -13551 8178 -13229
rect 8244 -13551 8274 -13229
rect 8340 -13551 8370 -13229
rect 8436 -13551 8466 -13229
rect 8532 -13551 8562 -13229
rect 8628 -13551 8658 -13229
rect 8724 -13551 8754 -13229
rect 8820 -13551 8850 -13229
rect 9084 -13551 9114 -13229
rect 9180 -13551 9210 -13229
rect 9276 -13551 9306 -13229
rect 9372 -13551 9402 -13229
rect 9468 -13551 9498 -13229
rect 9564 -13551 9594 -13229
rect 9660 -13551 9690 -13229
rect 9756 -13551 9786 -13229
rect 10015 -13550 10045 -13228
rect 10111 -13550 10141 -13228
rect 10207 -13550 10237 -13228
rect 10303 -13550 10333 -13228
rect 10399 -13550 10429 -13228
rect 10495 -13550 10525 -13228
rect 10591 -13550 10621 -13228
rect 10687 -13550 10717 -13228
rect 10942 -13551 10972 -13229
rect 11038 -13551 11068 -13229
rect 11134 -13551 11164 -13229
rect 11230 -13551 11260 -13229
rect 11326 -13551 11356 -13229
rect 11422 -13551 11452 -13229
rect 11518 -13551 11548 -13229
rect 11614 -13551 11644 -13229
rect -2050 -14032 -2020 -13818
rect -1954 -14032 -1924 -13818
rect -1858 -14032 -1828 -13818
rect -12316 -14181 -11766 -14151
rect -17677 -14591 -17421 -14561
rect -17677 -14687 -17421 -14657
rect -17677 -14783 -17421 -14753
rect -17677 -14879 -17421 -14849
rect -24449 -15008 -24235 -14978
rect -24449 -15104 -24235 -15074
rect -24449 -15200 -24235 -15170
rect -24449 -15296 -24235 -15266
rect -17677 -14975 -17421 -14945
rect -17677 -15071 -17421 -15041
rect -24449 -15392 -24235 -15362
rect -24449 -15488 -24235 -15458
rect -17677 -15167 -17421 -15137
rect -17677 -15263 -17421 -15233
rect -17677 -15359 -17421 -15329
rect -12316 -14273 -11766 -14243
rect -12316 -14369 -11766 -14339
rect -12316 -14465 -11766 -14435
rect -12316 -14561 -11766 -14531
rect -12316 -14657 -11766 -14627
rect -12316 -14753 -11766 -14723
rect -12316 -14849 -11766 -14819
rect -12316 -14945 -11766 -14915
rect -12316 -15041 -11766 -15011
rect -12316 -15137 -11766 -15107
rect -12316 -15233 -11766 -15203
rect -12316 -15329 -11766 -15299
rect -4766 -14417 -4736 -14203
rect -4670 -14417 -4640 -14203
rect -4574 -14417 -4544 -14203
rect -2050 -14411 -2020 -14197
rect -1954 -14411 -1924 -14197
rect -1858 -14411 -1828 -14197
rect 5658 -14281 5872 -14251
rect 5658 -14377 5872 -14347
rect 5658 -14473 5872 -14443
rect 6098 -14281 6312 -14251
rect 6098 -14377 6312 -14347
rect 6098 -14473 6312 -14443
rect 6538 -14281 6752 -14251
rect 6538 -14377 6752 -14347
rect 6538 -14473 6752 -14443
rect -4766 -14857 -4736 -14643
rect -4670 -14857 -4640 -14643
rect -4574 -14857 -4544 -14643
rect -2050 -14851 -2020 -14637
rect -1954 -14851 -1924 -14637
rect -1858 -14851 -1828 -14637
rect -4766 -15236 -4736 -15022
rect -4670 -15236 -4640 -15022
rect -4574 -15236 -4544 -15022
rect -2050 -15230 -2020 -15016
rect -1954 -15230 -1924 -15016
rect -1858 -15230 -1828 -15016
rect 7200 -15215 7230 -14893
rect 7296 -15215 7326 -14893
rect 7392 -15215 7422 -14893
rect 7488 -15215 7518 -14893
rect 7584 -15215 7614 -14893
rect 7680 -15215 7710 -14893
rect 7776 -15215 7806 -14893
rect 7872 -15215 7902 -14893
rect 8148 -15215 8178 -14893
rect 8244 -15215 8274 -14893
rect 8340 -15215 8370 -14893
rect 8436 -15215 8466 -14893
rect 8532 -15215 8562 -14893
rect 8628 -15215 8658 -14893
rect 8724 -15215 8754 -14893
rect 8820 -15215 8850 -14893
rect 9084 -15215 9114 -14893
rect 9180 -15215 9210 -14893
rect 9276 -15215 9306 -14893
rect 9372 -15215 9402 -14893
rect 9468 -15215 9498 -14893
rect 9564 -15215 9594 -14893
rect 9660 -15215 9690 -14893
rect 9756 -15215 9786 -14893
rect 10015 -15215 10045 -14893
rect 10111 -15215 10141 -14893
rect 10207 -15215 10237 -14893
rect 10303 -15215 10333 -14893
rect 10399 -15215 10429 -14893
rect 10495 -15215 10525 -14893
rect 10591 -15215 10621 -14893
rect 10687 -15215 10717 -14893
rect 10942 -15215 10972 -14893
rect 11038 -15215 11068 -14893
rect 11134 -15215 11164 -14893
rect 11230 -15215 11260 -14893
rect 11326 -15215 11356 -14893
rect 11422 -15215 11452 -14893
rect 11518 -15215 11548 -14893
rect 11614 -15215 11644 -14893
rect -12316 -15421 -11766 -15391
rect -17677 -15455 -17421 -15425
rect -8117 -15560 -8087 -15346
rect -8021 -15560 -7991 -15346
rect -7925 -15560 -7895 -15346
rect -4766 -15676 -4736 -15462
rect -4670 -15676 -4640 -15462
rect -4574 -15676 -4544 -15462
rect -2050 -15670 -2020 -15456
rect -1954 -15670 -1924 -15456
rect -1858 -15670 -1828 -15456
rect -17677 -15991 -17421 -15961
rect -17677 -16087 -17421 -16057
rect -8116 -16060 -8086 -15846
rect -8020 -16060 -7990 -15846
rect -7924 -16060 -7894 -15846
rect -4766 -16055 -4736 -15841
rect -4670 -16055 -4640 -15841
rect -4574 -16055 -4544 -15841
rect -24448 -16193 -24234 -16163
rect -24448 -16289 -24234 -16259
rect -24448 -16385 -24234 -16355
rect -24448 -16481 -24234 -16451
rect -2050 -16049 -2020 -15835
rect -1954 -16049 -1924 -15835
rect -1858 -16049 -1828 -15835
rect -17677 -16183 -17421 -16153
rect -17677 -16279 -17421 -16249
rect -17677 -16375 -17421 -16345
rect -17677 -16471 -17421 -16441
rect -24448 -16577 -24234 -16547
rect -24448 -16673 -24234 -16643
rect -17677 -16567 -17421 -16537
rect -8117 -16540 -8087 -16326
rect -8021 -16540 -7991 -16326
rect -7925 -16540 -7895 -16326
rect -4766 -16495 -4736 -16281
rect -4670 -16495 -4640 -16281
rect -4574 -16495 -4544 -16281
rect -2050 -16489 -2020 -16275
rect -1954 -16489 -1924 -16275
rect -1858 -16489 -1828 -16275
rect 11835 -16359 11865 -16103
rect 11931 -16359 11961 -16103
rect 12027 -16359 12057 -16103
rect 12123 -16359 12153 -16103
rect 12219 -16359 12249 -16103
rect 12315 -16359 12345 -16103
rect 12411 -16359 12441 -16103
rect 12507 -16359 12537 -16103
rect 12603 -16359 12633 -16103
rect 12699 -16359 12729 -16103
rect -17677 -16663 -17421 -16633
rect -17677 -16759 -17421 -16729
rect -17677 -16855 -17421 -16825
rect -12314 -16997 -11764 -16967
rect -24443 -17406 -24229 -17376
rect -24443 -17502 -24229 -17472
rect -24443 -17598 -24229 -17568
rect -24443 -17694 -24229 -17664
rect -17677 -17391 -17421 -17361
rect -17677 -17487 -17421 -17457
rect -17677 -17583 -17421 -17553
rect -17677 -17679 -17421 -17649
rect -24443 -17790 -24229 -17760
rect -17677 -17775 -17421 -17745
rect -24443 -17886 -24229 -17856
rect -17677 -17871 -17421 -17841
rect -21556 -18248 -21526 -18034
rect -21460 -18248 -21430 -18034
rect -21364 -18248 -21334 -18034
rect -17677 -17967 -17421 -17937
rect -17677 -18063 -17421 -18033
rect -15965 -18119 -15935 -17905
rect -15869 -18119 -15839 -17905
rect -15773 -18119 -15743 -17905
rect -17677 -18159 -17421 -18129
rect -12314 -17089 -11764 -17059
rect -12314 -17185 -11764 -17155
rect -12314 -17281 -11764 -17251
rect -12314 -17377 -11764 -17347
rect -12314 -17473 -11764 -17443
rect -12314 -17569 -11764 -17539
rect -12314 -17665 -11764 -17635
rect -12314 -17761 -11764 -17731
rect -12314 -17857 -11764 -17827
rect -12314 -17953 -11764 -17923
rect -12314 -18049 -11764 -18019
rect -12314 -18145 -11764 -18115
rect -8117 -17040 -8087 -16826
rect -8021 -17040 -7991 -16826
rect -7925 -17040 -7895 -16826
rect -4766 -16874 -4736 -16660
rect -4670 -16874 -4640 -16660
rect -4574 -16874 -4544 -16660
rect -2050 -16868 -2020 -16654
rect -1954 -16868 -1924 -16654
rect -1858 -16868 -1828 -16654
rect -8117 -17520 -8087 -17306
rect -8021 -17520 -7991 -17306
rect -7925 -17520 -7895 -17306
rect -4766 -17314 -4736 -17100
rect -4670 -17314 -4640 -17100
rect -4574 -17314 -4544 -17100
rect -2050 -17308 -2020 -17094
rect -1954 -17308 -1924 -17094
rect -1858 -17308 -1828 -17094
rect -4766 -17693 -4736 -17479
rect -4670 -17693 -4640 -17479
rect -4574 -17693 -4544 -17479
rect -2050 -17687 -2020 -17473
rect -1954 -17687 -1924 -17473
rect -1858 -17687 -1828 -17473
rect -8117 -17980 -8087 -17766
rect -8021 -17980 -7991 -17766
rect -7925 -17980 -7895 -17766
rect 12923 -16299 13137 -16269
rect 12923 -16395 13137 -16365
rect 12923 -16491 13137 -16461
rect -4766 -18133 -4736 -17919
rect -4670 -18133 -4640 -17919
rect -4574 -18133 -4544 -17919
rect -2050 -18127 -2020 -17913
rect -1954 -18127 -1924 -17913
rect -1858 -18127 -1828 -17913
rect 7200 -18079 7230 -17757
rect 7296 -18079 7326 -17757
rect 7392 -18079 7422 -17757
rect 7488 -18079 7518 -17757
rect 7584 -18079 7614 -17757
rect 7680 -18079 7710 -17757
rect 7776 -18079 7806 -17757
rect 7872 -18079 7902 -17757
rect 8148 -18079 8178 -17757
rect 8244 -18079 8274 -17757
rect 8340 -18079 8370 -17757
rect 8436 -18079 8466 -17757
rect 8532 -18079 8562 -17757
rect 8628 -18079 8658 -17757
rect 8724 -18079 8754 -17757
rect 8820 -18079 8850 -17757
rect 9084 -18079 9114 -17757
rect 9180 -18079 9210 -17757
rect 9276 -18079 9306 -17757
rect 9372 -18079 9402 -17757
rect 9468 -18079 9498 -17757
rect 9564 -18079 9594 -17757
rect 9660 -18079 9690 -17757
rect 9756 -18079 9786 -17757
rect 10015 -18078 10045 -17756
rect 10111 -18078 10141 -17756
rect 10207 -18078 10237 -17756
rect 10303 -18078 10333 -17756
rect 10399 -18078 10429 -17756
rect 10495 -18078 10525 -17756
rect 10591 -18078 10621 -17756
rect 10687 -18078 10717 -17756
rect 10942 -18079 10972 -17757
rect 11038 -18079 11068 -17757
rect 11134 -18079 11164 -17757
rect 11230 -18079 11260 -17757
rect 11326 -18079 11356 -17757
rect 11422 -18079 11452 -17757
rect 11518 -18079 11548 -17757
rect 11614 -18079 11644 -17757
rect -17677 -18255 -17421 -18225
rect -12314 -18237 -11764 -18207
rect -24428 -18525 -24214 -18495
rect -24428 -18621 -24214 -18591
rect -24428 -18717 -24214 -18687
rect -24428 -18813 -24214 -18783
rect -21555 -18748 -21525 -18534
rect -21459 -18748 -21429 -18534
rect -21363 -18748 -21333 -18534
rect -15964 -18619 -15934 -18405
rect -15868 -18619 -15838 -18405
rect -15772 -18619 -15742 -18405
rect -8131 -18440 -8101 -18226
rect -8035 -18440 -8005 -18226
rect -7939 -18440 -7909 -18226
rect -4766 -18512 -4736 -18298
rect -4670 -18512 -4640 -18298
rect -4574 -18512 -4544 -18298
rect -2050 -18506 -2020 -18292
rect -1954 -18506 -1924 -18292
rect -1858 -18506 -1828 -18292
rect 15825 -18523 15855 -17667
rect 15921 -18523 15951 -17667
rect 16017 -18523 16047 -17667
rect 16113 -18523 16143 -17667
rect 16209 -18523 16239 -17667
rect 16305 -18523 16335 -17667
rect 16401 -18523 16431 -17667
rect 16497 -18523 16527 -17667
rect 16593 -18523 16623 -17667
rect 16689 -18523 16719 -17667
rect 16785 -18523 16815 -17667
rect 16881 -18523 16911 -17667
rect 17356 -18489 17386 -18275
rect 17452 -18489 17482 -18275
rect 17548 -18489 17578 -18275
rect 17644 -18489 17674 -18275
rect 17740 -18489 17770 -18275
rect 17836 -18489 17866 -18275
rect -24428 -18909 -24214 -18879
rect -17677 -18791 -17421 -18761
rect -17677 -18887 -17421 -18857
rect -24428 -19005 -24214 -18975
rect -17677 -18983 -17421 -18953
rect -21556 -19228 -21526 -19014
rect -21460 -19228 -21430 -19014
rect -21364 -19228 -21334 -19014
rect -17677 -19079 -17421 -19049
rect -17677 -19175 -17421 -19145
rect -15965 -19099 -15935 -18885
rect -15869 -19099 -15839 -18885
rect -15773 -19099 -15743 -18885
rect -8129 -18920 -8099 -18706
rect -8033 -18920 -8003 -18706
rect -7937 -18920 -7907 -18706
rect 18096 -18339 18310 -18309
rect 18096 -18435 18310 -18405
rect 18096 -18531 18310 -18501
rect -4766 -18952 -4736 -18738
rect -4670 -18952 -4640 -18738
rect -4574 -18952 -4544 -18738
rect -2050 -18946 -2020 -18732
rect -1954 -18946 -1924 -18732
rect -1858 -18946 -1828 -18732
rect 5658 -18809 5872 -18779
rect 5658 -18905 5872 -18875
rect 5658 -19001 5872 -18971
rect 6098 -18809 6312 -18779
rect 6098 -18905 6312 -18875
rect 6098 -19001 6312 -18971
rect 6538 -18809 6752 -18779
rect 6538 -18905 6752 -18875
rect 6538 -19001 6752 -18971
rect -17677 -19271 -17421 -19241
rect -24426 -19719 -24212 -19689
rect -24426 -19815 -24212 -19785
rect -24426 -19911 -24212 -19881
rect -24426 -20007 -24212 -19977
rect -21556 -19728 -21526 -19514
rect -21460 -19728 -21430 -19514
rect -21364 -19728 -21334 -19514
rect -4766 -19331 -4736 -19117
rect -4670 -19331 -4640 -19117
rect -4574 -19331 -4544 -19117
rect -17677 -19367 -17421 -19337
rect -2050 -19325 -2020 -19111
rect -1954 -19325 -1924 -19111
rect -1858 -19325 -1828 -19111
rect -17677 -19463 -17421 -19433
rect -17677 -19559 -17421 -19529
rect -15965 -19599 -15935 -19385
rect -15869 -19599 -15839 -19385
rect -15773 -19599 -15743 -19385
rect -17677 -19655 -17421 -19625
rect -4766 -19771 -4736 -19557
rect -4670 -19771 -4640 -19557
rect -4574 -19771 -4544 -19557
rect -2050 -19765 -2020 -19551
rect -1954 -19765 -1924 -19551
rect -1858 -19765 -1828 -19551
rect 7200 -19743 7230 -19421
rect 7296 -19743 7326 -19421
rect 7392 -19743 7422 -19421
rect 7488 -19743 7518 -19421
rect 7584 -19743 7614 -19421
rect 7680 -19743 7710 -19421
rect 7776 -19743 7806 -19421
rect 7872 -19743 7902 -19421
rect 8148 -19743 8178 -19421
rect 8244 -19743 8274 -19421
rect 8340 -19743 8370 -19421
rect 8436 -19743 8466 -19421
rect 8532 -19743 8562 -19421
rect 8628 -19743 8658 -19421
rect 8724 -19743 8754 -19421
rect 8820 -19743 8850 -19421
rect 9084 -19743 9114 -19421
rect 9180 -19743 9210 -19421
rect 9276 -19743 9306 -19421
rect 9372 -19743 9402 -19421
rect 9468 -19743 9498 -19421
rect 9564 -19743 9594 -19421
rect 9660 -19743 9690 -19421
rect 9756 -19743 9786 -19421
rect 10015 -19743 10045 -19421
rect 10111 -19743 10141 -19421
rect 10207 -19743 10237 -19421
rect 10303 -19743 10333 -19421
rect 10399 -19743 10429 -19421
rect 10495 -19743 10525 -19421
rect 10591 -19743 10621 -19421
rect 10687 -19743 10717 -19421
rect 10942 -19743 10972 -19421
rect 11038 -19743 11068 -19421
rect 11134 -19743 11164 -19421
rect 11230 -19743 11260 -19421
rect 11326 -19743 11356 -19421
rect 11422 -19743 11452 -19421
rect 11518 -19743 11548 -19421
rect 11614 -19743 11644 -19421
rect 15825 -19505 15855 -18649
rect 15921 -19505 15951 -18649
rect 16017 -19505 16047 -18649
rect 16113 -19505 16143 -18649
rect 16209 -19505 16239 -18649
rect 16305 -19505 16335 -18649
rect 16401 -19505 16431 -18649
rect 16497 -19505 16527 -18649
rect 16593 -19505 16623 -18649
rect 16689 -19505 16719 -18649
rect 16785 -19505 16815 -18649
rect 16881 -19505 16911 -18649
rect -24426 -20103 -24212 -20073
rect -24426 -20199 -24212 -20169
rect -21556 -20208 -21526 -19994
rect -21460 -20208 -21430 -19994
rect -21364 -20208 -21334 -19994
rect -15965 -20079 -15935 -19865
rect -15869 -20079 -15839 -19865
rect -15773 -20079 -15743 -19865
rect -12314 -19954 -11764 -19924
rect -17677 -20191 -17421 -20161
rect -17677 -20287 -17421 -20257
rect -17677 -20383 -17421 -20353
rect -21556 -20668 -21526 -20454
rect -21460 -20668 -21430 -20454
rect -21364 -20668 -21334 -20454
rect -17677 -20479 -17421 -20449
rect -17677 -20575 -17421 -20545
rect -17677 -20671 -17421 -20641
rect -24395 -20919 -24181 -20889
rect -24395 -21015 -24181 -20985
rect -24395 -21111 -24181 -21081
rect -24395 -21207 -24181 -21177
rect -21570 -21128 -21540 -20914
rect -21474 -21128 -21444 -20914
rect -21378 -21128 -21348 -20914
rect -15965 -20539 -15935 -20325
rect -15869 -20539 -15839 -20325
rect -15773 -20539 -15743 -20325
rect -17677 -20767 -17421 -20737
rect -17677 -20863 -17421 -20833
rect -17677 -20959 -17421 -20929
rect -15979 -20999 -15949 -20785
rect -15883 -20999 -15853 -20785
rect -15787 -20999 -15757 -20785
rect -17677 -21055 -17421 -21025
rect -12314 -20046 -11764 -20016
rect -12314 -20142 -11764 -20112
rect -12314 -20238 -11764 -20208
rect -12314 -20334 -11764 -20304
rect -12314 -20430 -11764 -20400
rect -12314 -20526 -11764 -20496
rect -12314 -20622 -11764 -20592
rect -12314 -20718 -11764 -20688
rect -12314 -20814 -11764 -20784
rect -12314 -20910 -11764 -20880
rect -12314 -21006 -11764 -20976
rect -12314 -21102 -11764 -21072
rect -4766 -20150 -4736 -19936
rect -4670 -20150 -4640 -19936
rect -4574 -20150 -4544 -19936
rect -2050 -20144 -2020 -19930
rect -1954 -20144 -1924 -19930
rect -1858 -20144 -1828 -19930
rect -4766 -20590 -4736 -20376
rect -4670 -20590 -4640 -20376
rect -4574 -20590 -4544 -20376
rect -2050 -20584 -2020 -20370
rect -1954 -20584 -1924 -20370
rect -1858 -20584 -1828 -20370
rect -4766 -20969 -4736 -20755
rect -4670 -20969 -4640 -20755
rect -4574 -20969 -4544 -20755
rect 11835 -20887 11865 -20631
rect 11931 -20887 11961 -20631
rect 12027 -20887 12057 -20631
rect 12123 -20887 12153 -20631
rect 12219 -20887 12249 -20631
rect 12315 -20887 12345 -20631
rect 12411 -20887 12441 -20631
rect 12507 -20887 12537 -20631
rect 12603 -20887 12633 -20631
rect 12699 -20887 12729 -20631
rect -12314 -21194 -11764 -21164
rect -24395 -21303 -24181 -21273
rect -24395 -21399 -24181 -21369
rect -21568 -21608 -21538 -21394
rect -21472 -21608 -21442 -21394
rect -21376 -21608 -21346 -21394
rect -15977 -21479 -15947 -21265
rect -15881 -21479 -15851 -21265
rect -15785 -21479 -15755 -21265
rect -17677 -21591 -17421 -21561
rect -17677 -21687 -17421 -21657
rect -17677 -21783 -17421 -21753
rect -17677 -21879 -17421 -21849
rect -17677 -21975 -17421 -21945
rect -17677 -22071 -17421 -22041
rect -24396 -22222 -24182 -22192
rect -24396 -22318 -24182 -22288
rect -24396 -22414 -24182 -22384
rect -24396 -22510 -24182 -22480
rect -17677 -22167 -17421 -22137
rect -17677 -22263 -17421 -22233
rect 12923 -20827 13137 -20797
rect 12923 -20923 13137 -20893
rect 12923 -21019 13137 -20989
rect -17677 -22359 -17421 -22329
rect -17677 -22455 -17421 -22425
rect -24396 -22606 -24182 -22576
rect -12314 -22533 -11764 -22503
rect -24396 -22702 -24182 -22672
rect -17677 -22991 -17421 -22961
rect -17677 -23087 -17421 -23057
rect -17677 -23183 -17421 -23153
rect -17677 -23279 -17421 -23249
rect -17677 -23375 -17421 -23345
rect -24396 -23531 -24182 -23501
rect -24396 -23627 -24182 -23597
rect -24396 -23723 -24182 -23693
rect -24396 -23819 -24182 -23789
rect -17677 -23471 -17421 -23441
rect -24396 -23915 -24182 -23885
rect -17677 -23567 -17421 -23537
rect -17677 -23663 -17421 -23633
rect -17677 -23759 -17421 -23729
rect -12314 -22625 -11764 -22595
rect -12314 -22721 -11764 -22691
rect -12314 -22817 -11764 -22787
rect -12314 -22913 -11764 -22883
rect -12314 -23009 -11764 -22979
rect -12314 -23105 -11764 -23075
rect -12314 -23201 -11764 -23171
rect -12314 -23297 -11764 -23267
rect -12314 -23393 -11764 -23363
rect -12314 -23489 -11764 -23459
rect -12314 -23585 -11764 -23555
rect -12314 -23681 -11764 -23651
rect 7200 -22607 7230 -22285
rect 7296 -22607 7326 -22285
rect 7392 -22607 7422 -22285
rect 7488 -22607 7518 -22285
rect 7584 -22607 7614 -22285
rect 7680 -22607 7710 -22285
rect 7776 -22607 7806 -22285
rect 7872 -22607 7902 -22285
rect 8148 -22607 8178 -22285
rect 8244 -22607 8274 -22285
rect 8340 -22607 8370 -22285
rect 8436 -22607 8466 -22285
rect 8532 -22607 8562 -22285
rect 8628 -22607 8658 -22285
rect 8724 -22607 8754 -22285
rect 8820 -22607 8850 -22285
rect 9084 -22607 9114 -22285
rect 9180 -22607 9210 -22285
rect 9276 -22607 9306 -22285
rect 9372 -22607 9402 -22285
rect 9468 -22607 9498 -22285
rect 9564 -22607 9594 -22285
rect 9660 -22607 9690 -22285
rect 9756 -22607 9786 -22285
rect 10015 -22606 10045 -22284
rect 10111 -22606 10141 -22284
rect 10207 -22606 10237 -22284
rect 10303 -22606 10333 -22284
rect 10399 -22606 10429 -22284
rect 10495 -22606 10525 -22284
rect 10591 -22606 10621 -22284
rect 10687 -22606 10717 -22284
rect 10942 -22607 10972 -22285
rect 11038 -22607 11068 -22285
rect 11134 -22607 11164 -22285
rect 11230 -22607 11260 -22285
rect 11326 -22607 11356 -22285
rect 11422 -22607 11452 -22285
rect 11518 -22607 11548 -22285
rect 11614 -22607 11644 -22285
rect 5658 -23337 5872 -23307
rect 5658 -23433 5872 -23403
rect 5658 -23529 5872 -23499
rect 6098 -23337 6312 -23307
rect 6098 -23433 6312 -23403
rect 6098 -23529 6312 -23499
rect 6538 -23337 6752 -23307
rect 6538 -23433 6752 -23403
rect 6538 -23529 6752 -23499
rect -12314 -23773 -11764 -23743
rect -17677 -23855 -17421 -23825
rect -24396 -24011 -24182 -23981
rect 7200 -24271 7230 -23949
rect 7296 -24271 7326 -23949
rect 7392 -24271 7422 -23949
rect 7488 -24271 7518 -23949
rect 7584 -24271 7614 -23949
rect 7680 -24271 7710 -23949
rect 7776 -24271 7806 -23949
rect 7872 -24271 7902 -23949
rect 8148 -24271 8178 -23949
rect 8244 -24271 8274 -23949
rect 8340 -24271 8370 -23949
rect 8436 -24271 8466 -23949
rect 8532 -24271 8562 -23949
rect 8628 -24271 8658 -23949
rect 8724 -24271 8754 -23949
rect 8820 -24271 8850 -23949
rect 9084 -24271 9114 -23949
rect 9180 -24271 9210 -23949
rect 9276 -24271 9306 -23949
rect 9372 -24271 9402 -23949
rect 9468 -24271 9498 -23949
rect 9564 -24271 9594 -23949
rect 9660 -24271 9690 -23949
rect 9756 -24271 9786 -23949
rect 10015 -24271 10045 -23949
rect 10111 -24271 10141 -23949
rect 10207 -24271 10237 -23949
rect 10303 -24271 10333 -23949
rect 10399 -24271 10429 -23949
rect 10495 -24271 10525 -23949
rect 10591 -24271 10621 -23949
rect 10687 -24271 10717 -23949
rect 10942 -24271 10972 -23949
rect 11038 -24271 11068 -23949
rect 11134 -24271 11164 -23949
rect 11230 -24271 11260 -23949
rect 11326 -24271 11356 -23949
rect 11422 -24271 11452 -23949
rect 11518 -24271 11548 -23949
rect 11614 -24271 11644 -23949
rect -17677 -24391 -17421 -24361
rect -17677 -24487 -17421 -24457
rect -17677 -24583 -17421 -24553
rect -17677 -24679 -17421 -24649
rect -17677 -24775 -17421 -24745
rect -17677 -24871 -17421 -24841
rect -17677 -24967 -17421 -24937
rect -17677 -25063 -17421 -25033
rect -17677 -25159 -17421 -25129
rect -17677 -25255 -17421 -25225
rect -12314 -25301 -11764 -25271
rect -12314 -25393 -11764 -25363
rect -12314 -25489 -11764 -25459
rect -12314 -25585 -11764 -25555
rect -12314 -25681 -11764 -25651
rect -12314 -25777 -11764 -25747
rect -12314 -25873 -11764 -25843
rect -12314 -25969 -11764 -25939
rect -12314 -26065 -11764 -26035
rect -12314 -26161 -11764 -26131
rect -12314 -26257 -11764 -26227
rect -12314 -26353 -11764 -26323
rect -12314 -26449 -11764 -26419
rect 11835 -25415 11865 -25159
rect 11931 -25415 11961 -25159
rect 12027 -25415 12057 -25159
rect 12123 -25415 12153 -25159
rect 12219 -25415 12249 -25159
rect 12315 -25415 12345 -25159
rect 12411 -25415 12441 -25159
rect 12507 -25415 12537 -25159
rect 12603 -25415 12633 -25159
rect 12699 -25415 12729 -25159
rect -12314 -26541 -11764 -26511
rect 12923 -25355 13137 -25325
rect 12923 -25451 13137 -25421
rect 12923 -25547 13137 -25517
rect 7200 -27135 7230 -26813
rect 7296 -27135 7326 -26813
rect 7392 -27135 7422 -26813
rect 7488 -27135 7518 -26813
rect 7584 -27135 7614 -26813
rect 7680 -27135 7710 -26813
rect 7776 -27135 7806 -26813
rect 7872 -27135 7902 -26813
rect 8148 -27135 8178 -26813
rect 8244 -27135 8274 -26813
rect 8340 -27135 8370 -26813
rect 8436 -27135 8466 -26813
rect 8532 -27135 8562 -26813
rect 8628 -27135 8658 -26813
rect 8724 -27135 8754 -26813
rect 8820 -27135 8850 -26813
rect 9084 -27135 9114 -26813
rect 9180 -27135 9210 -26813
rect 9276 -27135 9306 -26813
rect 9372 -27135 9402 -26813
rect 9468 -27135 9498 -26813
rect 9564 -27135 9594 -26813
rect 9660 -27135 9690 -26813
rect 9756 -27135 9786 -26813
rect 10015 -27134 10045 -26812
rect 10111 -27134 10141 -26812
rect 10207 -27134 10237 -26812
rect 10303 -27134 10333 -26812
rect 10399 -27134 10429 -26812
rect 10495 -27134 10525 -26812
rect 10591 -27134 10621 -26812
rect 10687 -27134 10717 -26812
rect 10942 -27135 10972 -26813
rect 11038 -27135 11068 -26813
rect 11134 -27135 11164 -26813
rect 11230 -27135 11260 -26813
rect 11326 -27135 11356 -26813
rect 11422 -27135 11452 -26813
rect 11518 -27135 11548 -26813
rect 11614 -27135 11644 -26813
rect -12314 -27934 -11764 -27904
rect -12314 -28026 -11764 -27996
rect -12314 -28122 -11764 -28092
rect -12314 -28218 -11764 -28188
rect -12314 -28314 -11764 -28284
rect -12314 -28410 -11764 -28380
rect -12314 -28506 -11764 -28476
rect -12314 -28602 -11764 -28572
rect -12314 -28698 -11764 -28668
rect -12314 -28794 -11764 -28764
rect -12314 -28890 -11764 -28860
rect -12314 -28986 -11764 -28956
rect -12314 -29082 -11764 -29052
rect 5658 -27865 5872 -27835
rect 5658 -27961 5872 -27931
rect 5658 -28057 5872 -28027
rect 6098 -27865 6312 -27835
rect 6098 -27961 6312 -27931
rect 6098 -28057 6312 -28027
rect 6538 -27865 6752 -27835
rect 6538 -27961 6752 -27931
rect 6538 -28057 6752 -28027
rect 7200 -28799 7230 -28477
rect 7296 -28799 7326 -28477
rect 7392 -28799 7422 -28477
rect 7488 -28799 7518 -28477
rect 7584 -28799 7614 -28477
rect 7680 -28799 7710 -28477
rect 7776 -28799 7806 -28477
rect 7872 -28799 7902 -28477
rect 8148 -28799 8178 -28477
rect 8244 -28799 8274 -28477
rect 8340 -28799 8370 -28477
rect 8436 -28799 8466 -28477
rect 8532 -28799 8562 -28477
rect 8628 -28799 8658 -28477
rect 8724 -28799 8754 -28477
rect 8820 -28799 8850 -28477
rect 9084 -28799 9114 -28477
rect 9180 -28799 9210 -28477
rect 9276 -28799 9306 -28477
rect 9372 -28799 9402 -28477
rect 9468 -28799 9498 -28477
rect 9564 -28799 9594 -28477
rect 9660 -28799 9690 -28477
rect 9756 -28799 9786 -28477
rect 10015 -28799 10045 -28477
rect 10111 -28799 10141 -28477
rect 10207 -28799 10237 -28477
rect 10303 -28799 10333 -28477
rect 10399 -28799 10429 -28477
rect 10495 -28799 10525 -28477
rect 10591 -28799 10621 -28477
rect 10687 -28799 10717 -28477
rect 10942 -28799 10972 -28477
rect 11038 -28799 11068 -28477
rect 11134 -28799 11164 -28477
rect 11230 -28799 11260 -28477
rect 11326 -28799 11356 -28477
rect 11422 -28799 11452 -28477
rect 11518 -28799 11548 -28477
rect 11614 -28799 11644 -28477
rect -12314 -29174 -11764 -29144
rect 11835 -29943 11865 -29687
rect 11931 -29943 11961 -29687
rect 12027 -29943 12057 -29687
rect 12123 -29943 12153 -29687
rect 12219 -29943 12249 -29687
rect 12315 -29943 12345 -29687
rect 12411 -29943 12441 -29687
rect 12507 -29943 12537 -29687
rect 12603 -29943 12633 -29687
rect 12699 -29943 12729 -29687
rect -12314 -30543 -11764 -30513
rect -12314 -30635 -11764 -30605
rect -12314 -30731 -11764 -30701
rect -12314 -30827 -11764 -30797
rect -12314 -30923 -11764 -30893
rect -12314 -31019 -11764 -30989
rect -12314 -31115 -11764 -31085
rect -12314 -31211 -11764 -31181
rect -12314 -31307 -11764 -31277
rect -12314 -31403 -11764 -31373
rect -12314 -31499 -11764 -31469
rect -12314 -31595 -11764 -31565
rect -12314 -31691 -11764 -31661
rect 12923 -29883 13137 -29853
rect 12923 -29979 13137 -29949
rect 12923 -30075 13137 -30045
rect 7200 -31663 7230 -31341
rect 7296 -31663 7326 -31341
rect 7392 -31663 7422 -31341
rect 7488 -31663 7518 -31341
rect 7584 -31663 7614 -31341
rect 7680 -31663 7710 -31341
rect 7776 -31663 7806 -31341
rect 7872 -31663 7902 -31341
rect 8148 -31663 8178 -31341
rect 8244 -31663 8274 -31341
rect 8340 -31663 8370 -31341
rect 8436 -31663 8466 -31341
rect 8532 -31663 8562 -31341
rect 8628 -31663 8658 -31341
rect 8724 -31663 8754 -31341
rect 8820 -31663 8850 -31341
rect 9084 -31663 9114 -31341
rect 9180 -31663 9210 -31341
rect 9276 -31663 9306 -31341
rect 9372 -31663 9402 -31341
rect 9468 -31663 9498 -31341
rect 9564 -31663 9594 -31341
rect 9660 -31663 9690 -31341
rect 9756 -31663 9786 -31341
rect 10015 -31662 10045 -31340
rect 10111 -31662 10141 -31340
rect 10207 -31662 10237 -31340
rect 10303 -31662 10333 -31340
rect 10399 -31662 10429 -31340
rect 10495 -31662 10525 -31340
rect 10591 -31662 10621 -31340
rect 10687 -31662 10717 -31340
rect 10942 -31663 10972 -31341
rect 11038 -31663 11068 -31341
rect 11134 -31663 11164 -31341
rect 11230 -31663 11260 -31341
rect 11326 -31663 11356 -31341
rect 11422 -31663 11452 -31341
rect 11518 -31663 11548 -31341
rect 11614 -31663 11644 -31341
rect -12314 -31783 -11764 -31753
rect 5658 -32393 5872 -32363
rect 5658 -32489 5872 -32459
rect 5658 -32585 5872 -32555
rect 6098 -32393 6312 -32363
rect 6098 -32489 6312 -32459
rect 6098 -32585 6312 -32555
rect 6538 -32393 6752 -32363
rect 6538 -32489 6752 -32459
rect 6538 -32585 6752 -32555
rect -12316 -33163 -11766 -33133
rect -12316 -33255 -11766 -33225
rect -12316 -33351 -11766 -33321
rect -12316 -33447 -11766 -33417
rect -12316 -33543 -11766 -33513
rect -12316 -33639 -11766 -33609
rect -12316 -33735 -11766 -33705
rect -12316 -33831 -11766 -33801
rect -12316 -33927 -11766 -33897
rect -12316 -34023 -11766 -33993
rect -12316 -34119 -11766 -34089
rect -12316 -34215 -11766 -34185
rect -12316 -34311 -11766 -34281
rect 7200 -33327 7230 -33005
rect 7296 -33327 7326 -33005
rect 7392 -33327 7422 -33005
rect 7488 -33327 7518 -33005
rect 7584 -33327 7614 -33005
rect 7680 -33327 7710 -33005
rect 7776 -33327 7806 -33005
rect 7872 -33327 7902 -33005
rect 8148 -33327 8178 -33005
rect 8244 -33327 8274 -33005
rect 8340 -33327 8370 -33005
rect 8436 -33327 8466 -33005
rect 8532 -33327 8562 -33005
rect 8628 -33327 8658 -33005
rect 8724 -33327 8754 -33005
rect 8820 -33327 8850 -33005
rect 9084 -33327 9114 -33005
rect 9180 -33327 9210 -33005
rect 9276 -33327 9306 -33005
rect 9372 -33327 9402 -33005
rect 9468 -33327 9498 -33005
rect 9564 -33327 9594 -33005
rect 9660 -33327 9690 -33005
rect 9756 -33327 9786 -33005
rect 10015 -33327 10045 -33005
rect 10111 -33327 10141 -33005
rect 10207 -33327 10237 -33005
rect 10303 -33327 10333 -33005
rect 10399 -33327 10429 -33005
rect 10495 -33327 10525 -33005
rect 10591 -33327 10621 -33005
rect 10687 -33327 10717 -33005
rect 10942 -33327 10972 -33005
rect 11038 -33327 11068 -33005
rect 11134 -33327 11164 -33005
rect 11230 -33327 11260 -33005
rect 11326 -33327 11356 -33005
rect 11422 -33327 11452 -33005
rect 11518 -33327 11548 -33005
rect 11614 -33327 11644 -33005
rect -12316 -34403 -11766 -34373
rect 11835 -34471 11865 -34215
rect 11931 -34471 11961 -34215
rect 12027 -34471 12057 -34215
rect 12123 -34471 12153 -34215
rect 12219 -34471 12249 -34215
rect 12315 -34471 12345 -34215
rect 12411 -34471 12441 -34215
rect 12507 -34471 12537 -34215
rect 12603 -34471 12633 -34215
rect 12699 -34471 12729 -34215
rect 12923 -34411 13137 -34381
rect 12923 -34507 13137 -34477
rect 12923 -34603 13137 -34573
rect 7200 -36191 7230 -35869
rect 7296 -36191 7326 -35869
rect 7392 -36191 7422 -35869
rect 7488 -36191 7518 -35869
rect 7584 -36191 7614 -35869
rect 7680 -36191 7710 -35869
rect 7776 -36191 7806 -35869
rect 7872 -36191 7902 -35869
rect 8148 -36191 8178 -35869
rect 8244 -36191 8274 -35869
rect 8340 -36191 8370 -35869
rect 8436 -36191 8466 -35869
rect 8532 -36191 8562 -35869
rect 8628 -36191 8658 -35869
rect 8724 -36191 8754 -35869
rect 8820 -36191 8850 -35869
rect 9084 -36191 9114 -35869
rect 9180 -36191 9210 -35869
rect 9276 -36191 9306 -35869
rect 9372 -36191 9402 -35869
rect 9468 -36191 9498 -35869
rect 9564 -36191 9594 -35869
rect 9660 -36191 9690 -35869
rect 9756 -36191 9786 -35869
rect 10015 -36190 10045 -35868
rect 10111 -36190 10141 -35868
rect 10207 -36190 10237 -35868
rect 10303 -36190 10333 -35868
rect 10399 -36190 10429 -35868
rect 10495 -36190 10525 -35868
rect 10591 -36190 10621 -35868
rect 10687 -36190 10717 -35868
rect 10942 -36191 10972 -35869
rect 11038 -36191 11068 -35869
rect 11134 -36191 11164 -35869
rect 11230 -36191 11260 -35869
rect 11326 -36191 11356 -35869
rect 11422 -36191 11452 -35869
rect 11518 -36191 11548 -35869
rect 11614 -36191 11644 -35869
rect 13186 -35929 13216 -35715
rect 13282 -35929 13312 -35715
rect 13378 -35929 13408 -35715
rect 13186 -36308 13216 -36094
rect 13282 -36308 13312 -36094
rect 13378 -36308 13408 -36094
<< ndiff >>
rect 1707 5032 1765 5044
rect 1707 4926 1719 5032
rect 1753 4926 1765 5032
rect 1707 4914 1765 4926
rect 1795 5032 1857 5044
rect 1795 4926 1807 5032
rect 1841 4926 1857 5032
rect 1795 4914 1857 4926
rect 1887 5032 1953 5044
rect 1887 4926 1903 5032
rect 1937 4926 1953 5032
rect 1887 4914 1953 4926
rect 1983 5032 2049 5044
rect 1983 4926 1999 5032
rect 2033 4926 2049 5032
rect 1983 4914 2049 4926
rect 2079 5032 2145 5044
rect 2079 4926 2095 5032
rect 2129 4926 2145 5032
rect 2079 4914 2145 4926
rect 2175 5032 2241 5044
rect 2175 4926 2191 5032
rect 2225 4926 2241 5032
rect 2175 4914 2241 4926
rect 2271 5032 2337 5044
rect 2271 4926 2287 5032
rect 2321 4926 2337 5032
rect 2271 4914 2337 4926
rect 2367 5032 2433 5044
rect 2367 4926 2383 5032
rect 2417 4926 2433 5032
rect 2367 4914 2433 4926
rect 2463 5032 2529 5044
rect 2463 4926 2479 5032
rect 2513 4926 2529 5032
rect 2463 4914 2529 4926
rect 2559 5032 2625 5044
rect 2559 4926 2575 5032
rect 2609 4926 2625 5032
rect 2559 4914 2625 4926
rect 2655 5032 2721 5044
rect 2655 4926 2671 5032
rect 2705 4926 2721 5032
rect 2655 4914 2721 4926
rect 2751 5032 2817 5044
rect 2751 4926 2767 5032
rect 2801 4926 2817 5032
rect 2751 4914 2817 4926
rect 2847 5032 2913 5044
rect 2847 4926 2863 5032
rect 2897 4926 2913 5032
rect 2847 4914 2913 4926
rect 2943 5032 3005 5044
rect 2943 4926 2959 5032
rect 2993 4926 3005 5032
rect 2943 4914 3005 4926
rect 3035 5032 3093 5044
rect 3035 4926 3047 5032
rect 3081 4926 3093 5032
rect 3035 4914 3093 4926
rect 3313 5032 3371 5044
rect 3313 4926 3325 5032
rect 3359 4926 3371 5032
rect 3313 4914 3371 4926
rect 3401 5032 3463 5044
rect 3401 4926 3413 5032
rect 3447 4926 3463 5032
rect 3401 4914 3463 4926
rect 3493 5032 3559 5044
rect 3493 4926 3509 5032
rect 3543 4926 3559 5032
rect 3493 4914 3559 4926
rect 3589 5032 3655 5044
rect 3589 4926 3605 5032
rect 3639 4926 3655 5032
rect 3589 4914 3655 4926
rect 3685 5032 3751 5044
rect 3685 4926 3701 5032
rect 3735 4926 3751 5032
rect 3685 4914 3751 4926
rect 3781 5032 3847 5044
rect 3781 4926 3797 5032
rect 3831 4926 3847 5032
rect 3781 4914 3847 4926
rect 3877 5032 3943 5044
rect 3877 4926 3893 5032
rect 3927 4926 3943 5032
rect 3877 4914 3943 4926
rect 3973 5032 4039 5044
rect 3973 4926 3989 5032
rect 4023 4926 4039 5032
rect 3973 4914 4039 4926
rect 4069 5032 4135 5044
rect 4069 4926 4085 5032
rect 4119 4926 4135 5032
rect 4069 4914 4135 4926
rect 4165 5032 4231 5044
rect 4165 4926 4181 5032
rect 4215 4926 4231 5032
rect 4165 4914 4231 4926
rect 4261 5032 4327 5044
rect 4261 4926 4277 5032
rect 4311 4926 4327 5032
rect 4261 4914 4327 4926
rect 4357 5032 4423 5044
rect 4357 4926 4373 5032
rect 4407 4926 4423 5032
rect 4357 4914 4423 4926
rect 4453 5032 4519 5044
rect 4453 4926 4469 5032
rect 4503 4926 4519 5032
rect 4453 4914 4519 4926
rect 4549 5032 4611 5044
rect 4549 4926 4565 5032
rect 4599 4926 4611 5032
rect 4549 4914 4611 4926
rect 4641 5032 4699 5044
rect 4641 4926 4653 5032
rect 4687 4926 4699 5032
rect 4641 4914 4699 4926
rect 5017 5030 5075 5042
rect 5017 4924 5029 5030
rect 5063 4924 5075 5030
rect 5017 4912 5075 4924
rect 5105 5030 5167 5042
rect 5105 4924 5117 5030
rect 5151 4924 5167 5030
rect 5105 4912 5167 4924
rect 5197 5030 5263 5042
rect 5197 4924 5213 5030
rect 5247 4924 5263 5030
rect 5197 4912 5263 4924
rect 5293 5030 5359 5042
rect 5293 4924 5309 5030
rect 5343 4924 5359 5030
rect 5293 4912 5359 4924
rect 5389 5030 5455 5042
rect 5389 4924 5405 5030
rect 5439 4924 5455 5030
rect 5389 4912 5455 4924
rect 5485 5030 5551 5042
rect 5485 4924 5501 5030
rect 5535 4924 5551 5030
rect 5485 4912 5551 4924
rect 5581 5030 5647 5042
rect 5581 4924 5597 5030
rect 5631 4924 5647 5030
rect 5581 4912 5647 4924
rect 5677 5030 5743 5042
rect 5677 4924 5693 5030
rect 5727 4924 5743 5030
rect 5677 4912 5743 4924
rect 5773 5030 5839 5042
rect 5773 4924 5789 5030
rect 5823 4924 5839 5030
rect 5773 4912 5839 4924
rect 5869 5030 5935 5042
rect 5869 4924 5885 5030
rect 5919 4924 5935 5030
rect 5869 4912 5935 4924
rect 5965 5030 6031 5042
rect 5965 4924 5981 5030
rect 6015 4924 6031 5030
rect 5965 4912 6031 4924
rect 6061 5030 6127 5042
rect 6061 4924 6077 5030
rect 6111 4924 6127 5030
rect 6061 4912 6127 4924
rect 6157 5030 6223 5042
rect 6157 4924 6173 5030
rect 6207 4924 6223 5030
rect 6157 4912 6223 4924
rect 6253 5030 6315 5042
rect 6253 4924 6269 5030
rect 6303 4924 6315 5030
rect 6253 4912 6315 4924
rect 6345 5030 6403 5042
rect 6345 4924 6357 5030
rect 6391 4924 6403 5030
rect 6345 4912 6403 4924
rect 7173 5085 7573 5097
rect 7173 5051 7185 5085
rect 7561 5051 7573 5085
rect 7173 5035 7573 5051
rect 7809 5009 8009 5021
rect 7173 4939 7573 5005
rect 7809 4975 7821 5009
rect 7997 4975 8009 5009
rect 7809 4963 8009 4975
rect 7809 4921 8009 4933
rect 7173 4893 7573 4909
rect 7173 4859 7185 4893
rect 7561 4859 7573 4893
rect 7809 4887 7821 4921
rect 7997 4887 8009 4921
rect 7809 4875 8009 4887
rect 7173 4847 7573 4859
rect 5658 3461 5858 3473
rect 5658 3427 5670 3461
rect 5846 3427 5858 3461
rect 6098 3461 6298 3473
rect 5658 3415 5858 3427
rect 5658 3373 5858 3385
rect 5658 3339 5670 3373
rect 5846 3339 5858 3373
rect 6098 3427 6110 3461
rect 6286 3427 6298 3461
rect 6538 3461 6738 3473
rect 6098 3415 6298 3427
rect 6098 3373 6298 3385
rect 5658 3327 5858 3339
rect 6098 3339 6110 3373
rect 6286 3339 6298 3373
rect 6538 3427 6550 3461
rect 6726 3427 6738 3461
rect 6538 3415 6738 3427
rect 6538 3373 6738 3385
rect 6098 3327 6298 3339
rect 6538 3339 6550 3373
rect 6726 3339 6738 3373
rect 6538 3327 6738 3339
rect -24130 3308 -24072 3320
rect -24130 3202 -24118 3308
rect -24084 3202 -24072 3308
rect -24130 3190 -24072 3202
rect -24042 3308 -23980 3320
rect -24042 3202 -24030 3308
rect -23996 3202 -23980 3308
rect -24042 3190 -23980 3202
rect -23950 3308 -23884 3320
rect -23950 3202 -23934 3308
rect -23900 3202 -23884 3308
rect -23950 3190 -23884 3202
rect -23854 3308 -23788 3320
rect -23854 3202 -23838 3308
rect -23804 3202 -23788 3308
rect -23854 3190 -23788 3202
rect -23758 3308 -23692 3320
rect -23758 3202 -23742 3308
rect -23708 3202 -23692 3308
rect -23758 3190 -23692 3202
rect -23662 3308 -23596 3320
rect -23662 3202 -23646 3308
rect -23612 3202 -23596 3308
rect -23662 3190 -23596 3202
rect -23566 3308 -23500 3320
rect -23566 3202 -23550 3308
rect -23516 3202 -23500 3308
rect -23566 3190 -23500 3202
rect -23470 3308 -23404 3320
rect -23470 3202 -23454 3308
rect -23420 3202 -23404 3308
rect -23470 3190 -23404 3202
rect -23374 3308 -23308 3320
rect -23374 3202 -23358 3308
rect -23324 3202 -23308 3308
rect -23374 3190 -23308 3202
rect -23278 3308 -23212 3320
rect -23278 3202 -23262 3308
rect -23228 3202 -23212 3308
rect -23278 3190 -23212 3202
rect -23182 3308 -23116 3320
rect -23182 3202 -23166 3308
rect -23132 3202 -23116 3308
rect -23182 3190 -23116 3202
rect -23086 3308 -23020 3320
rect -23086 3202 -23070 3308
rect -23036 3202 -23020 3308
rect -23086 3190 -23020 3202
rect -22990 3308 -22924 3320
rect -22990 3202 -22974 3308
rect -22940 3202 -22924 3308
rect -22990 3190 -22924 3202
rect -22894 3308 -22832 3320
rect -22894 3202 -22878 3308
rect -22844 3202 -22832 3308
rect -22894 3190 -22832 3202
rect -22802 3308 -22744 3320
rect -22802 3202 -22790 3308
rect -22756 3202 -22744 3308
rect -22802 3190 -22744 3202
rect -20839 3308 -20781 3320
rect -20839 3202 -20827 3308
rect -20793 3202 -20781 3308
rect -20839 3190 -20781 3202
rect -20751 3308 -20689 3320
rect -20751 3202 -20739 3308
rect -20705 3202 -20689 3308
rect -20751 3190 -20689 3202
rect -20659 3308 -20593 3320
rect -20659 3202 -20643 3308
rect -20609 3202 -20593 3308
rect -20659 3190 -20593 3202
rect -20563 3308 -20497 3320
rect -20563 3202 -20547 3308
rect -20513 3202 -20497 3308
rect -20563 3190 -20497 3202
rect -20467 3308 -20401 3320
rect -20467 3202 -20451 3308
rect -20417 3202 -20401 3308
rect -20467 3190 -20401 3202
rect -20371 3308 -20305 3320
rect -20371 3202 -20355 3308
rect -20321 3202 -20305 3308
rect -20371 3190 -20305 3202
rect -20275 3308 -20209 3320
rect -20275 3202 -20259 3308
rect -20225 3202 -20209 3308
rect -20275 3190 -20209 3202
rect -20179 3308 -20113 3320
rect -20179 3202 -20163 3308
rect -20129 3202 -20113 3308
rect -20179 3190 -20113 3202
rect -20083 3308 -20017 3320
rect -20083 3202 -20067 3308
rect -20033 3202 -20017 3308
rect -20083 3190 -20017 3202
rect -19987 3308 -19921 3320
rect -19987 3202 -19971 3308
rect -19937 3202 -19921 3308
rect -19987 3190 -19921 3202
rect -19891 3308 -19825 3320
rect -19891 3202 -19875 3308
rect -19841 3202 -19825 3308
rect -19891 3190 -19825 3202
rect -19795 3308 -19729 3320
rect -19795 3202 -19779 3308
rect -19745 3202 -19729 3308
rect -19795 3190 -19729 3202
rect -19699 3308 -19633 3320
rect -19699 3202 -19683 3308
rect -19649 3202 -19633 3308
rect -19699 3190 -19633 3202
rect -19603 3308 -19541 3320
rect -19603 3202 -19587 3308
rect -19553 3202 -19541 3308
rect -19603 3190 -19541 3202
rect -19511 3308 -19453 3320
rect -19511 3202 -19499 3308
rect -19465 3202 -19453 3308
rect -19511 3190 -19453 3202
rect -17548 3308 -17490 3320
rect -17548 3202 -17536 3308
rect -17502 3202 -17490 3308
rect -17548 3190 -17490 3202
rect -17460 3308 -17398 3320
rect -17460 3202 -17448 3308
rect -17414 3202 -17398 3308
rect -17460 3190 -17398 3202
rect -17368 3308 -17302 3320
rect -17368 3202 -17352 3308
rect -17318 3202 -17302 3308
rect -17368 3190 -17302 3202
rect -17272 3308 -17206 3320
rect -17272 3202 -17256 3308
rect -17222 3202 -17206 3308
rect -17272 3190 -17206 3202
rect -17176 3308 -17110 3320
rect -17176 3202 -17160 3308
rect -17126 3202 -17110 3308
rect -17176 3190 -17110 3202
rect -17080 3308 -17014 3320
rect -17080 3202 -17064 3308
rect -17030 3202 -17014 3308
rect -17080 3190 -17014 3202
rect -16984 3308 -16918 3320
rect -16984 3202 -16968 3308
rect -16934 3202 -16918 3308
rect -16984 3190 -16918 3202
rect -16888 3308 -16822 3320
rect -16888 3202 -16872 3308
rect -16838 3202 -16822 3308
rect -16888 3190 -16822 3202
rect -16792 3308 -16726 3320
rect -16792 3202 -16776 3308
rect -16742 3202 -16726 3308
rect -16792 3190 -16726 3202
rect -16696 3308 -16630 3320
rect -16696 3202 -16680 3308
rect -16646 3202 -16630 3308
rect -16696 3190 -16630 3202
rect -16600 3308 -16534 3320
rect -16600 3202 -16584 3308
rect -16550 3202 -16534 3308
rect -16600 3190 -16534 3202
rect -16504 3308 -16438 3320
rect -16504 3202 -16488 3308
rect -16454 3202 -16438 3308
rect -16504 3190 -16438 3202
rect -16408 3308 -16342 3320
rect -16408 3202 -16392 3308
rect -16358 3202 -16342 3308
rect -16408 3190 -16342 3202
rect -16312 3308 -16250 3320
rect -16312 3202 -16296 3308
rect -16262 3202 -16250 3308
rect -16312 3190 -16250 3202
rect -16220 3308 -16162 3320
rect -16220 3202 -16208 3308
rect -16174 3202 -16162 3308
rect -16220 3190 -16162 3202
rect -14257 3308 -14199 3320
rect -14257 3202 -14245 3308
rect -14211 3202 -14199 3308
rect -14257 3190 -14199 3202
rect -14169 3308 -14107 3320
rect -14169 3202 -14157 3308
rect -14123 3202 -14107 3308
rect -14169 3190 -14107 3202
rect -14077 3308 -14011 3320
rect -14077 3202 -14061 3308
rect -14027 3202 -14011 3308
rect -14077 3190 -14011 3202
rect -13981 3308 -13915 3320
rect -13981 3202 -13965 3308
rect -13931 3202 -13915 3308
rect -13981 3190 -13915 3202
rect -13885 3308 -13819 3320
rect -13885 3202 -13869 3308
rect -13835 3202 -13819 3308
rect -13885 3190 -13819 3202
rect -13789 3308 -13723 3320
rect -13789 3202 -13773 3308
rect -13739 3202 -13723 3308
rect -13789 3190 -13723 3202
rect -13693 3308 -13627 3320
rect -13693 3202 -13677 3308
rect -13643 3202 -13627 3308
rect -13693 3190 -13627 3202
rect -13597 3308 -13531 3320
rect -13597 3202 -13581 3308
rect -13547 3202 -13531 3308
rect -13597 3190 -13531 3202
rect -13501 3308 -13435 3320
rect -13501 3202 -13485 3308
rect -13451 3202 -13435 3308
rect -13501 3190 -13435 3202
rect -13405 3308 -13339 3320
rect -13405 3202 -13389 3308
rect -13355 3202 -13339 3308
rect -13405 3190 -13339 3202
rect -13309 3308 -13243 3320
rect -13309 3202 -13293 3308
rect -13259 3202 -13243 3308
rect -13309 3190 -13243 3202
rect -13213 3308 -13147 3320
rect -13213 3202 -13197 3308
rect -13163 3202 -13147 3308
rect -13213 3190 -13147 3202
rect -13117 3308 -13051 3320
rect -13117 3202 -13101 3308
rect -13067 3202 -13051 3308
rect -13117 3190 -13051 3202
rect -13021 3308 -12959 3320
rect -13021 3202 -13005 3308
rect -12971 3202 -12959 3308
rect -13021 3190 -12959 3202
rect -12929 3308 -12871 3320
rect -12929 3202 -12917 3308
rect -12883 3202 -12871 3308
rect -12929 3190 -12871 3202
rect -10966 3308 -10908 3320
rect -10966 3202 -10954 3308
rect -10920 3202 -10908 3308
rect -10966 3190 -10908 3202
rect -10878 3308 -10816 3320
rect -10878 3202 -10866 3308
rect -10832 3202 -10816 3308
rect -10878 3190 -10816 3202
rect -10786 3308 -10720 3320
rect -10786 3202 -10770 3308
rect -10736 3202 -10720 3308
rect -10786 3190 -10720 3202
rect -10690 3308 -10624 3320
rect -10690 3202 -10674 3308
rect -10640 3202 -10624 3308
rect -10690 3190 -10624 3202
rect -10594 3308 -10528 3320
rect -10594 3202 -10578 3308
rect -10544 3202 -10528 3308
rect -10594 3190 -10528 3202
rect -10498 3308 -10432 3320
rect -10498 3202 -10482 3308
rect -10448 3202 -10432 3308
rect -10498 3190 -10432 3202
rect -10402 3308 -10336 3320
rect -10402 3202 -10386 3308
rect -10352 3202 -10336 3308
rect -10402 3190 -10336 3202
rect -10306 3308 -10240 3320
rect -10306 3202 -10290 3308
rect -10256 3202 -10240 3308
rect -10306 3190 -10240 3202
rect -10210 3308 -10144 3320
rect -10210 3202 -10194 3308
rect -10160 3202 -10144 3308
rect -10210 3190 -10144 3202
rect -10114 3308 -10048 3320
rect -10114 3202 -10098 3308
rect -10064 3202 -10048 3308
rect -10114 3190 -10048 3202
rect -10018 3308 -9952 3320
rect -10018 3202 -10002 3308
rect -9968 3202 -9952 3308
rect -10018 3190 -9952 3202
rect -9922 3308 -9856 3320
rect -9922 3202 -9906 3308
rect -9872 3202 -9856 3308
rect -9922 3190 -9856 3202
rect -9826 3308 -9760 3320
rect -9826 3202 -9810 3308
rect -9776 3202 -9760 3308
rect -9826 3190 -9760 3202
rect -9730 3308 -9668 3320
rect -9730 3202 -9714 3308
rect -9680 3202 -9668 3308
rect -9730 3190 -9668 3202
rect -9638 3308 -9580 3320
rect -9638 3202 -9626 3308
rect -9592 3202 -9580 3308
rect -9638 3190 -9580 3202
rect -7676 3308 -7618 3320
rect -7676 3202 -7664 3308
rect -7630 3202 -7618 3308
rect -7676 3190 -7618 3202
rect -7588 3308 -7526 3320
rect -7588 3202 -7576 3308
rect -7542 3202 -7526 3308
rect -7588 3190 -7526 3202
rect -7496 3308 -7430 3320
rect -7496 3202 -7480 3308
rect -7446 3202 -7430 3308
rect -7496 3190 -7430 3202
rect -7400 3308 -7334 3320
rect -7400 3202 -7384 3308
rect -7350 3202 -7334 3308
rect -7400 3190 -7334 3202
rect -7304 3308 -7238 3320
rect -7304 3202 -7288 3308
rect -7254 3202 -7238 3308
rect -7304 3190 -7238 3202
rect -7208 3308 -7142 3320
rect -7208 3202 -7192 3308
rect -7158 3202 -7142 3308
rect -7208 3190 -7142 3202
rect -7112 3308 -7046 3320
rect -7112 3202 -7096 3308
rect -7062 3202 -7046 3308
rect -7112 3190 -7046 3202
rect -7016 3308 -6950 3320
rect -7016 3202 -7000 3308
rect -6966 3202 -6950 3308
rect -7016 3190 -6950 3202
rect -6920 3308 -6854 3320
rect -6920 3202 -6904 3308
rect -6870 3202 -6854 3308
rect -6920 3190 -6854 3202
rect -6824 3308 -6758 3320
rect -6824 3202 -6808 3308
rect -6774 3202 -6758 3308
rect -6824 3190 -6758 3202
rect -6728 3308 -6662 3320
rect -6728 3202 -6712 3308
rect -6678 3202 -6662 3308
rect -6728 3190 -6662 3202
rect -6632 3308 -6566 3320
rect -6632 3202 -6616 3308
rect -6582 3202 -6566 3308
rect -6632 3190 -6566 3202
rect -6536 3308 -6470 3320
rect -6536 3202 -6520 3308
rect -6486 3202 -6470 3308
rect -6536 3190 -6470 3202
rect -6440 3308 -6378 3320
rect -6440 3202 -6424 3308
rect -6390 3202 -6378 3308
rect -6440 3190 -6378 3202
rect -6348 3308 -6290 3320
rect -6348 3202 -6336 3308
rect -6302 3202 -6290 3308
rect -6348 3190 -6290 3202
rect -4385 3308 -4327 3320
rect -4385 3202 -4373 3308
rect -4339 3202 -4327 3308
rect -4385 3190 -4327 3202
rect -4297 3308 -4235 3320
rect -4297 3202 -4285 3308
rect -4251 3202 -4235 3308
rect -4297 3190 -4235 3202
rect -4205 3308 -4139 3320
rect -4205 3202 -4189 3308
rect -4155 3202 -4139 3308
rect -4205 3190 -4139 3202
rect -4109 3308 -4043 3320
rect -4109 3202 -4093 3308
rect -4059 3202 -4043 3308
rect -4109 3190 -4043 3202
rect -4013 3308 -3947 3320
rect -4013 3202 -3997 3308
rect -3963 3202 -3947 3308
rect -4013 3190 -3947 3202
rect -3917 3308 -3851 3320
rect -3917 3202 -3901 3308
rect -3867 3202 -3851 3308
rect -3917 3190 -3851 3202
rect -3821 3308 -3755 3320
rect -3821 3202 -3805 3308
rect -3771 3202 -3755 3308
rect -3821 3190 -3755 3202
rect -3725 3308 -3659 3320
rect -3725 3202 -3709 3308
rect -3675 3202 -3659 3308
rect -3725 3190 -3659 3202
rect -3629 3308 -3563 3320
rect -3629 3202 -3613 3308
rect -3579 3202 -3563 3308
rect -3629 3190 -3563 3202
rect -3533 3308 -3467 3320
rect -3533 3202 -3517 3308
rect -3483 3202 -3467 3308
rect -3533 3190 -3467 3202
rect -3437 3308 -3371 3320
rect -3437 3202 -3421 3308
rect -3387 3202 -3371 3308
rect -3437 3190 -3371 3202
rect -3341 3308 -3275 3320
rect -3341 3202 -3325 3308
rect -3291 3202 -3275 3308
rect -3341 3190 -3275 3202
rect -3245 3308 -3179 3320
rect -3245 3202 -3229 3308
rect -3195 3202 -3179 3308
rect -3245 3190 -3179 3202
rect -3149 3308 -3087 3320
rect -3149 3202 -3133 3308
rect -3099 3202 -3087 3308
rect -3149 3190 -3087 3202
rect -3057 3308 -2999 3320
rect -3057 3202 -3045 3308
rect -3011 3202 -2999 3308
rect -3057 3190 -2999 3202
rect -1094 3308 -1036 3320
rect -1094 3202 -1082 3308
rect -1048 3202 -1036 3308
rect -1094 3190 -1036 3202
rect -1006 3308 -944 3320
rect -1006 3202 -994 3308
rect -960 3202 -944 3308
rect -1006 3190 -944 3202
rect -914 3308 -848 3320
rect -914 3202 -898 3308
rect -864 3202 -848 3308
rect -914 3190 -848 3202
rect -818 3308 -752 3320
rect -818 3202 -802 3308
rect -768 3202 -752 3308
rect -818 3190 -752 3202
rect -722 3308 -656 3320
rect -722 3202 -706 3308
rect -672 3202 -656 3308
rect -722 3190 -656 3202
rect -626 3308 -560 3320
rect -626 3202 -610 3308
rect -576 3202 -560 3308
rect -626 3190 -560 3202
rect -530 3308 -464 3320
rect -530 3202 -514 3308
rect -480 3202 -464 3308
rect -530 3190 -464 3202
rect -434 3308 -368 3320
rect -434 3202 -418 3308
rect -384 3202 -368 3308
rect -434 3190 -368 3202
rect -338 3308 -272 3320
rect -338 3202 -322 3308
rect -288 3202 -272 3308
rect -338 3190 -272 3202
rect -242 3308 -176 3320
rect -242 3202 -226 3308
rect -192 3202 -176 3308
rect -242 3190 -176 3202
rect -146 3308 -80 3320
rect -146 3202 -130 3308
rect -96 3202 -80 3308
rect -146 3190 -80 3202
rect -50 3308 16 3320
rect -50 3202 -34 3308
rect 0 3202 16 3308
rect -50 3190 16 3202
rect 46 3308 112 3320
rect 46 3202 62 3308
rect 96 3202 112 3308
rect 46 3190 112 3202
rect 142 3308 204 3320
rect 142 3202 158 3308
rect 192 3202 204 3308
rect 142 3190 204 3202
rect 234 3308 292 3320
rect 234 3202 246 3308
rect 280 3202 292 3308
rect 234 3190 292 3202
rect 7360 2478 7422 2490
rect 7360 1702 7372 2478
rect 7406 1702 7422 2478
rect 7360 1690 7422 1702
rect 7452 1690 7518 2490
rect 7548 1690 7614 2490
rect 7644 1690 7710 2490
rect 7740 2478 7802 2490
rect 7740 1702 7756 2478
rect 7790 1702 7802 2478
rect 7740 1690 7802 1702
rect 8308 2478 8370 2490
rect 8308 1702 8320 2478
rect 8354 1702 8370 2478
rect 8308 1690 8370 1702
rect 8400 1690 8466 2490
rect 8496 1690 8562 2490
rect 8592 1690 8658 2490
rect 8688 2478 8750 2490
rect 8688 1702 8704 2478
rect 8738 1702 8750 2478
rect 8688 1690 8750 1702
rect 9244 2478 9306 2490
rect 9244 1702 9256 2478
rect 9290 1702 9306 2478
rect 9244 1690 9306 1702
rect 9336 1690 9402 2490
rect 9432 1690 9498 2490
rect 9528 1690 9594 2490
rect 9624 2478 9686 2490
rect 9624 1702 9640 2478
rect 9674 1702 9686 2478
rect 9624 1690 9686 1702
rect 10175 2478 10237 2490
rect 10175 1702 10187 2478
rect 10221 1702 10237 2478
rect 10175 1690 10237 1702
rect 10267 1690 10333 2490
rect 10363 1690 10429 2490
rect 10459 1690 10525 2490
rect 10555 2478 10617 2490
rect 10555 1702 10571 2478
rect 10605 1702 10617 2478
rect 10555 1690 10617 1702
rect 11102 2478 11164 2490
rect 11102 1702 11114 2478
rect 11148 1702 11164 2478
rect 11102 1690 11164 1702
rect 11194 1690 11260 2490
rect 11290 1690 11356 2490
rect 11386 1690 11452 2490
rect 11482 2478 11544 2490
rect 11482 1702 11498 2478
rect 11532 1702 11544 2478
rect 11482 1690 11544 1702
rect 7360 1550 7422 1562
rect -24804 1524 -24746 1536
rect -24804 1418 -24792 1524
rect -24758 1418 -24746 1524
rect -24804 1406 -24746 1418
rect -24716 1524 -24654 1536
rect -24716 1418 -24704 1524
rect -24670 1418 -24654 1524
rect -24716 1406 -24654 1418
rect -24624 1524 -24558 1536
rect -24624 1418 -24608 1524
rect -24574 1418 -24558 1524
rect -24624 1406 -24558 1418
rect -24528 1524 -24462 1536
rect -24528 1418 -24512 1524
rect -24478 1418 -24462 1524
rect -24528 1406 -24462 1418
rect -24432 1524 -24366 1536
rect -24432 1418 -24416 1524
rect -24382 1418 -24366 1524
rect -24432 1406 -24366 1418
rect -24336 1524 -24270 1536
rect -24336 1418 -24320 1524
rect -24286 1418 -24270 1524
rect -24336 1406 -24270 1418
rect -24240 1524 -24174 1536
rect -24240 1418 -24224 1524
rect -24190 1418 -24174 1524
rect -24240 1406 -24174 1418
rect -24144 1524 -24078 1536
rect -24144 1418 -24128 1524
rect -24094 1418 -24078 1524
rect -24144 1406 -24078 1418
rect -24048 1524 -23982 1536
rect -24048 1418 -24032 1524
rect -23998 1418 -23982 1524
rect -24048 1406 -23982 1418
rect -23952 1524 -23886 1536
rect -23952 1418 -23936 1524
rect -23902 1418 -23886 1524
rect -23952 1406 -23886 1418
rect -23856 1524 -23790 1536
rect -23856 1418 -23840 1524
rect -23806 1418 -23790 1524
rect -23856 1406 -23790 1418
rect -23760 1524 -23694 1536
rect -23760 1418 -23744 1524
rect -23710 1418 -23694 1524
rect -23760 1406 -23694 1418
rect -23664 1524 -23598 1536
rect -23664 1418 -23648 1524
rect -23614 1418 -23598 1524
rect -23664 1406 -23598 1418
rect -23568 1524 -23506 1536
rect -23568 1418 -23552 1524
rect -23518 1418 -23506 1524
rect -23568 1406 -23506 1418
rect -23476 1524 -23418 1536
rect -23476 1418 -23464 1524
rect -23430 1418 -23418 1524
rect -23476 1406 -23418 1418
rect -23245 1524 -23187 1536
rect -23245 1418 -23233 1524
rect -23199 1418 -23187 1524
rect -23245 1406 -23187 1418
rect -23157 1524 -23095 1536
rect -23157 1418 -23145 1524
rect -23111 1418 -23095 1524
rect -23157 1406 -23095 1418
rect -23065 1524 -22999 1536
rect -23065 1418 -23049 1524
rect -23015 1418 -22999 1524
rect -23065 1406 -22999 1418
rect -22969 1524 -22903 1536
rect -22969 1418 -22953 1524
rect -22919 1418 -22903 1524
rect -22969 1406 -22903 1418
rect -22873 1524 -22807 1536
rect -22873 1418 -22857 1524
rect -22823 1418 -22807 1524
rect -22873 1406 -22807 1418
rect -22777 1524 -22711 1536
rect -22777 1418 -22761 1524
rect -22727 1418 -22711 1524
rect -22777 1406 -22711 1418
rect -22681 1524 -22615 1536
rect -22681 1418 -22665 1524
rect -22631 1418 -22615 1524
rect -22681 1406 -22615 1418
rect -22585 1524 -22519 1536
rect -22585 1418 -22569 1524
rect -22535 1418 -22519 1524
rect -22585 1406 -22519 1418
rect -22489 1524 -22423 1536
rect -22489 1418 -22473 1524
rect -22439 1418 -22423 1524
rect -22489 1406 -22423 1418
rect -22393 1524 -22327 1536
rect -22393 1418 -22377 1524
rect -22343 1418 -22327 1524
rect -22393 1406 -22327 1418
rect -22297 1524 -22231 1536
rect -22297 1418 -22281 1524
rect -22247 1418 -22231 1524
rect -22297 1406 -22231 1418
rect -22201 1524 -22135 1536
rect -22201 1418 -22185 1524
rect -22151 1418 -22135 1524
rect -22201 1406 -22135 1418
rect -22105 1524 -22039 1536
rect -22105 1418 -22089 1524
rect -22055 1418 -22039 1524
rect -22105 1406 -22039 1418
rect -22009 1524 -21947 1536
rect -22009 1418 -21993 1524
rect -21959 1418 -21947 1524
rect -22009 1406 -21947 1418
rect -21917 1524 -21859 1536
rect -21917 1418 -21905 1524
rect -21871 1418 -21859 1524
rect -21917 1406 -21859 1418
rect -21513 1524 -21455 1536
rect -21513 1418 -21501 1524
rect -21467 1418 -21455 1524
rect -21513 1406 -21455 1418
rect -21425 1524 -21363 1536
rect -21425 1418 -21413 1524
rect -21379 1418 -21363 1524
rect -21425 1406 -21363 1418
rect -21333 1524 -21267 1536
rect -21333 1418 -21317 1524
rect -21283 1418 -21267 1524
rect -21333 1406 -21267 1418
rect -21237 1524 -21171 1536
rect -21237 1418 -21221 1524
rect -21187 1418 -21171 1524
rect -21237 1406 -21171 1418
rect -21141 1524 -21075 1536
rect -21141 1418 -21125 1524
rect -21091 1418 -21075 1524
rect -21141 1406 -21075 1418
rect -21045 1524 -20979 1536
rect -21045 1418 -21029 1524
rect -20995 1418 -20979 1524
rect -21045 1406 -20979 1418
rect -20949 1524 -20883 1536
rect -20949 1418 -20933 1524
rect -20899 1418 -20883 1524
rect -20949 1406 -20883 1418
rect -20853 1524 -20787 1536
rect -20853 1418 -20837 1524
rect -20803 1418 -20787 1524
rect -20853 1406 -20787 1418
rect -20757 1524 -20691 1536
rect -20757 1418 -20741 1524
rect -20707 1418 -20691 1524
rect -20757 1406 -20691 1418
rect -20661 1524 -20595 1536
rect -20661 1418 -20645 1524
rect -20611 1418 -20595 1524
rect -20661 1406 -20595 1418
rect -20565 1524 -20499 1536
rect -20565 1418 -20549 1524
rect -20515 1418 -20499 1524
rect -20565 1406 -20499 1418
rect -20469 1524 -20403 1536
rect -20469 1418 -20453 1524
rect -20419 1418 -20403 1524
rect -20469 1406 -20403 1418
rect -20373 1524 -20307 1536
rect -20373 1418 -20357 1524
rect -20323 1418 -20307 1524
rect -20373 1406 -20307 1418
rect -20277 1524 -20215 1536
rect -20277 1418 -20261 1524
rect -20227 1418 -20215 1524
rect -20277 1406 -20215 1418
rect -20185 1524 -20127 1536
rect -20185 1418 -20173 1524
rect -20139 1418 -20127 1524
rect -20185 1406 -20127 1418
rect -19954 1524 -19896 1536
rect -19954 1418 -19942 1524
rect -19908 1418 -19896 1524
rect -19954 1406 -19896 1418
rect -19866 1524 -19804 1536
rect -19866 1418 -19854 1524
rect -19820 1418 -19804 1524
rect -19866 1406 -19804 1418
rect -19774 1524 -19708 1536
rect -19774 1418 -19758 1524
rect -19724 1418 -19708 1524
rect -19774 1406 -19708 1418
rect -19678 1524 -19612 1536
rect -19678 1418 -19662 1524
rect -19628 1418 -19612 1524
rect -19678 1406 -19612 1418
rect -19582 1524 -19516 1536
rect -19582 1418 -19566 1524
rect -19532 1418 -19516 1524
rect -19582 1406 -19516 1418
rect -19486 1524 -19420 1536
rect -19486 1418 -19470 1524
rect -19436 1418 -19420 1524
rect -19486 1406 -19420 1418
rect -19390 1524 -19324 1536
rect -19390 1418 -19374 1524
rect -19340 1418 -19324 1524
rect -19390 1406 -19324 1418
rect -19294 1524 -19228 1536
rect -19294 1418 -19278 1524
rect -19244 1418 -19228 1524
rect -19294 1406 -19228 1418
rect -19198 1524 -19132 1536
rect -19198 1418 -19182 1524
rect -19148 1418 -19132 1524
rect -19198 1406 -19132 1418
rect -19102 1524 -19036 1536
rect -19102 1418 -19086 1524
rect -19052 1418 -19036 1524
rect -19102 1406 -19036 1418
rect -19006 1524 -18940 1536
rect -19006 1418 -18990 1524
rect -18956 1418 -18940 1524
rect -19006 1406 -18940 1418
rect -18910 1524 -18844 1536
rect -18910 1418 -18894 1524
rect -18860 1418 -18844 1524
rect -18910 1406 -18844 1418
rect -18814 1524 -18748 1536
rect -18814 1418 -18798 1524
rect -18764 1418 -18748 1524
rect -18814 1406 -18748 1418
rect -18718 1524 -18656 1536
rect -18718 1418 -18702 1524
rect -18668 1418 -18656 1524
rect -18718 1406 -18656 1418
rect -18626 1524 -18568 1536
rect -18626 1418 -18614 1524
rect -18580 1418 -18568 1524
rect -18626 1406 -18568 1418
rect -18222 1524 -18164 1536
rect -18222 1418 -18210 1524
rect -18176 1418 -18164 1524
rect -18222 1406 -18164 1418
rect -18134 1524 -18072 1536
rect -18134 1418 -18122 1524
rect -18088 1418 -18072 1524
rect -18134 1406 -18072 1418
rect -18042 1524 -17976 1536
rect -18042 1418 -18026 1524
rect -17992 1418 -17976 1524
rect -18042 1406 -17976 1418
rect -17946 1524 -17880 1536
rect -17946 1418 -17930 1524
rect -17896 1418 -17880 1524
rect -17946 1406 -17880 1418
rect -17850 1524 -17784 1536
rect -17850 1418 -17834 1524
rect -17800 1418 -17784 1524
rect -17850 1406 -17784 1418
rect -17754 1524 -17688 1536
rect -17754 1418 -17738 1524
rect -17704 1418 -17688 1524
rect -17754 1406 -17688 1418
rect -17658 1524 -17592 1536
rect -17658 1418 -17642 1524
rect -17608 1418 -17592 1524
rect -17658 1406 -17592 1418
rect -17562 1524 -17496 1536
rect -17562 1418 -17546 1524
rect -17512 1418 -17496 1524
rect -17562 1406 -17496 1418
rect -17466 1524 -17400 1536
rect -17466 1418 -17450 1524
rect -17416 1418 -17400 1524
rect -17466 1406 -17400 1418
rect -17370 1524 -17304 1536
rect -17370 1418 -17354 1524
rect -17320 1418 -17304 1524
rect -17370 1406 -17304 1418
rect -17274 1524 -17208 1536
rect -17274 1418 -17258 1524
rect -17224 1418 -17208 1524
rect -17274 1406 -17208 1418
rect -17178 1524 -17112 1536
rect -17178 1418 -17162 1524
rect -17128 1418 -17112 1524
rect -17178 1406 -17112 1418
rect -17082 1524 -17016 1536
rect -17082 1418 -17066 1524
rect -17032 1418 -17016 1524
rect -17082 1406 -17016 1418
rect -16986 1524 -16924 1536
rect -16986 1418 -16970 1524
rect -16936 1418 -16924 1524
rect -16986 1406 -16924 1418
rect -16894 1524 -16836 1536
rect -16894 1418 -16882 1524
rect -16848 1418 -16836 1524
rect -16894 1406 -16836 1418
rect -16663 1524 -16605 1536
rect -16663 1418 -16651 1524
rect -16617 1418 -16605 1524
rect -16663 1406 -16605 1418
rect -16575 1524 -16513 1536
rect -16575 1418 -16563 1524
rect -16529 1418 -16513 1524
rect -16575 1406 -16513 1418
rect -16483 1524 -16417 1536
rect -16483 1418 -16467 1524
rect -16433 1418 -16417 1524
rect -16483 1406 -16417 1418
rect -16387 1524 -16321 1536
rect -16387 1418 -16371 1524
rect -16337 1418 -16321 1524
rect -16387 1406 -16321 1418
rect -16291 1524 -16225 1536
rect -16291 1418 -16275 1524
rect -16241 1418 -16225 1524
rect -16291 1406 -16225 1418
rect -16195 1524 -16129 1536
rect -16195 1418 -16179 1524
rect -16145 1418 -16129 1524
rect -16195 1406 -16129 1418
rect -16099 1524 -16033 1536
rect -16099 1418 -16083 1524
rect -16049 1418 -16033 1524
rect -16099 1406 -16033 1418
rect -16003 1524 -15937 1536
rect -16003 1418 -15987 1524
rect -15953 1418 -15937 1524
rect -16003 1406 -15937 1418
rect -15907 1524 -15841 1536
rect -15907 1418 -15891 1524
rect -15857 1418 -15841 1524
rect -15907 1406 -15841 1418
rect -15811 1524 -15745 1536
rect -15811 1418 -15795 1524
rect -15761 1418 -15745 1524
rect -15811 1406 -15745 1418
rect -15715 1524 -15649 1536
rect -15715 1418 -15699 1524
rect -15665 1418 -15649 1524
rect -15715 1406 -15649 1418
rect -15619 1524 -15553 1536
rect -15619 1418 -15603 1524
rect -15569 1418 -15553 1524
rect -15619 1406 -15553 1418
rect -15523 1524 -15457 1536
rect -15523 1418 -15507 1524
rect -15473 1418 -15457 1524
rect -15523 1406 -15457 1418
rect -15427 1524 -15365 1536
rect -15427 1418 -15411 1524
rect -15377 1418 -15365 1524
rect -15427 1406 -15365 1418
rect -15335 1524 -15277 1536
rect -15335 1418 -15323 1524
rect -15289 1418 -15277 1524
rect -15335 1406 -15277 1418
rect -14931 1524 -14873 1536
rect -14931 1418 -14919 1524
rect -14885 1418 -14873 1524
rect -14931 1406 -14873 1418
rect -14843 1524 -14781 1536
rect -14843 1418 -14831 1524
rect -14797 1418 -14781 1524
rect -14843 1406 -14781 1418
rect -14751 1524 -14685 1536
rect -14751 1418 -14735 1524
rect -14701 1418 -14685 1524
rect -14751 1406 -14685 1418
rect -14655 1524 -14589 1536
rect -14655 1418 -14639 1524
rect -14605 1418 -14589 1524
rect -14655 1406 -14589 1418
rect -14559 1524 -14493 1536
rect -14559 1418 -14543 1524
rect -14509 1418 -14493 1524
rect -14559 1406 -14493 1418
rect -14463 1524 -14397 1536
rect -14463 1418 -14447 1524
rect -14413 1418 -14397 1524
rect -14463 1406 -14397 1418
rect -14367 1524 -14301 1536
rect -14367 1418 -14351 1524
rect -14317 1418 -14301 1524
rect -14367 1406 -14301 1418
rect -14271 1524 -14205 1536
rect -14271 1418 -14255 1524
rect -14221 1418 -14205 1524
rect -14271 1406 -14205 1418
rect -14175 1524 -14109 1536
rect -14175 1418 -14159 1524
rect -14125 1418 -14109 1524
rect -14175 1406 -14109 1418
rect -14079 1524 -14013 1536
rect -14079 1418 -14063 1524
rect -14029 1418 -14013 1524
rect -14079 1406 -14013 1418
rect -13983 1524 -13917 1536
rect -13983 1418 -13967 1524
rect -13933 1418 -13917 1524
rect -13983 1406 -13917 1418
rect -13887 1524 -13821 1536
rect -13887 1418 -13871 1524
rect -13837 1418 -13821 1524
rect -13887 1406 -13821 1418
rect -13791 1524 -13725 1536
rect -13791 1418 -13775 1524
rect -13741 1418 -13725 1524
rect -13791 1406 -13725 1418
rect -13695 1524 -13633 1536
rect -13695 1418 -13679 1524
rect -13645 1418 -13633 1524
rect -13695 1406 -13633 1418
rect -13603 1524 -13545 1536
rect -13603 1418 -13591 1524
rect -13557 1418 -13545 1524
rect -13603 1406 -13545 1418
rect -13372 1524 -13314 1536
rect -13372 1418 -13360 1524
rect -13326 1418 -13314 1524
rect -13372 1406 -13314 1418
rect -13284 1524 -13222 1536
rect -13284 1418 -13272 1524
rect -13238 1418 -13222 1524
rect -13284 1406 -13222 1418
rect -13192 1524 -13126 1536
rect -13192 1418 -13176 1524
rect -13142 1418 -13126 1524
rect -13192 1406 -13126 1418
rect -13096 1524 -13030 1536
rect -13096 1418 -13080 1524
rect -13046 1418 -13030 1524
rect -13096 1406 -13030 1418
rect -13000 1524 -12934 1536
rect -13000 1418 -12984 1524
rect -12950 1418 -12934 1524
rect -13000 1406 -12934 1418
rect -12904 1524 -12838 1536
rect -12904 1418 -12888 1524
rect -12854 1418 -12838 1524
rect -12904 1406 -12838 1418
rect -12808 1524 -12742 1536
rect -12808 1418 -12792 1524
rect -12758 1418 -12742 1524
rect -12808 1406 -12742 1418
rect -12712 1524 -12646 1536
rect -12712 1418 -12696 1524
rect -12662 1418 -12646 1524
rect -12712 1406 -12646 1418
rect -12616 1524 -12550 1536
rect -12616 1418 -12600 1524
rect -12566 1418 -12550 1524
rect -12616 1406 -12550 1418
rect -12520 1524 -12454 1536
rect -12520 1418 -12504 1524
rect -12470 1418 -12454 1524
rect -12520 1406 -12454 1418
rect -12424 1524 -12358 1536
rect -12424 1418 -12408 1524
rect -12374 1418 -12358 1524
rect -12424 1406 -12358 1418
rect -12328 1524 -12262 1536
rect -12328 1418 -12312 1524
rect -12278 1418 -12262 1524
rect -12328 1406 -12262 1418
rect -12232 1524 -12166 1536
rect -12232 1418 -12216 1524
rect -12182 1418 -12166 1524
rect -12232 1406 -12166 1418
rect -12136 1524 -12074 1536
rect -12136 1418 -12120 1524
rect -12086 1418 -12074 1524
rect -12136 1406 -12074 1418
rect -12044 1524 -11986 1536
rect -12044 1418 -12032 1524
rect -11998 1418 -11986 1524
rect -12044 1406 -11986 1418
rect -11640 1524 -11582 1536
rect -11640 1418 -11628 1524
rect -11594 1418 -11582 1524
rect -11640 1406 -11582 1418
rect -11552 1524 -11490 1536
rect -11552 1418 -11540 1524
rect -11506 1418 -11490 1524
rect -11552 1406 -11490 1418
rect -11460 1524 -11394 1536
rect -11460 1418 -11444 1524
rect -11410 1418 -11394 1524
rect -11460 1406 -11394 1418
rect -11364 1524 -11298 1536
rect -11364 1418 -11348 1524
rect -11314 1418 -11298 1524
rect -11364 1406 -11298 1418
rect -11268 1524 -11202 1536
rect -11268 1418 -11252 1524
rect -11218 1418 -11202 1524
rect -11268 1406 -11202 1418
rect -11172 1524 -11106 1536
rect -11172 1418 -11156 1524
rect -11122 1418 -11106 1524
rect -11172 1406 -11106 1418
rect -11076 1524 -11010 1536
rect -11076 1418 -11060 1524
rect -11026 1418 -11010 1524
rect -11076 1406 -11010 1418
rect -10980 1524 -10914 1536
rect -10980 1418 -10964 1524
rect -10930 1418 -10914 1524
rect -10980 1406 -10914 1418
rect -10884 1524 -10818 1536
rect -10884 1418 -10868 1524
rect -10834 1418 -10818 1524
rect -10884 1406 -10818 1418
rect -10788 1524 -10722 1536
rect -10788 1418 -10772 1524
rect -10738 1418 -10722 1524
rect -10788 1406 -10722 1418
rect -10692 1524 -10626 1536
rect -10692 1418 -10676 1524
rect -10642 1418 -10626 1524
rect -10692 1406 -10626 1418
rect -10596 1524 -10530 1536
rect -10596 1418 -10580 1524
rect -10546 1418 -10530 1524
rect -10596 1406 -10530 1418
rect -10500 1524 -10434 1536
rect -10500 1418 -10484 1524
rect -10450 1418 -10434 1524
rect -10500 1406 -10434 1418
rect -10404 1524 -10342 1536
rect -10404 1418 -10388 1524
rect -10354 1418 -10342 1524
rect -10404 1406 -10342 1418
rect -10312 1524 -10254 1536
rect -10312 1418 -10300 1524
rect -10266 1418 -10254 1524
rect -10312 1406 -10254 1418
rect -10081 1524 -10023 1536
rect -10081 1418 -10069 1524
rect -10035 1418 -10023 1524
rect -10081 1406 -10023 1418
rect -9993 1524 -9931 1536
rect -9993 1418 -9981 1524
rect -9947 1418 -9931 1524
rect -9993 1406 -9931 1418
rect -9901 1524 -9835 1536
rect -9901 1418 -9885 1524
rect -9851 1418 -9835 1524
rect -9901 1406 -9835 1418
rect -9805 1524 -9739 1536
rect -9805 1418 -9789 1524
rect -9755 1418 -9739 1524
rect -9805 1406 -9739 1418
rect -9709 1524 -9643 1536
rect -9709 1418 -9693 1524
rect -9659 1418 -9643 1524
rect -9709 1406 -9643 1418
rect -9613 1524 -9547 1536
rect -9613 1418 -9597 1524
rect -9563 1418 -9547 1524
rect -9613 1406 -9547 1418
rect -9517 1524 -9451 1536
rect -9517 1418 -9501 1524
rect -9467 1418 -9451 1524
rect -9517 1406 -9451 1418
rect -9421 1524 -9355 1536
rect -9421 1418 -9405 1524
rect -9371 1418 -9355 1524
rect -9421 1406 -9355 1418
rect -9325 1524 -9259 1536
rect -9325 1418 -9309 1524
rect -9275 1418 -9259 1524
rect -9325 1406 -9259 1418
rect -9229 1524 -9163 1536
rect -9229 1418 -9213 1524
rect -9179 1418 -9163 1524
rect -9229 1406 -9163 1418
rect -9133 1524 -9067 1536
rect -9133 1418 -9117 1524
rect -9083 1418 -9067 1524
rect -9133 1406 -9067 1418
rect -9037 1524 -8971 1536
rect -9037 1418 -9021 1524
rect -8987 1418 -8971 1524
rect -9037 1406 -8971 1418
rect -8941 1524 -8875 1536
rect -8941 1418 -8925 1524
rect -8891 1418 -8875 1524
rect -8941 1406 -8875 1418
rect -8845 1524 -8783 1536
rect -8845 1418 -8829 1524
rect -8795 1418 -8783 1524
rect -8845 1406 -8783 1418
rect -8753 1524 -8695 1536
rect -8753 1418 -8741 1524
rect -8707 1418 -8695 1524
rect -8753 1406 -8695 1418
rect -8350 1524 -8292 1536
rect -8350 1418 -8338 1524
rect -8304 1418 -8292 1524
rect -8350 1406 -8292 1418
rect -8262 1524 -8200 1536
rect -8262 1418 -8250 1524
rect -8216 1418 -8200 1524
rect -8262 1406 -8200 1418
rect -8170 1524 -8104 1536
rect -8170 1418 -8154 1524
rect -8120 1418 -8104 1524
rect -8170 1406 -8104 1418
rect -8074 1524 -8008 1536
rect -8074 1418 -8058 1524
rect -8024 1418 -8008 1524
rect -8074 1406 -8008 1418
rect -7978 1524 -7912 1536
rect -7978 1418 -7962 1524
rect -7928 1418 -7912 1524
rect -7978 1406 -7912 1418
rect -7882 1524 -7816 1536
rect -7882 1418 -7866 1524
rect -7832 1418 -7816 1524
rect -7882 1406 -7816 1418
rect -7786 1524 -7720 1536
rect -7786 1418 -7770 1524
rect -7736 1418 -7720 1524
rect -7786 1406 -7720 1418
rect -7690 1524 -7624 1536
rect -7690 1418 -7674 1524
rect -7640 1418 -7624 1524
rect -7690 1406 -7624 1418
rect -7594 1524 -7528 1536
rect -7594 1418 -7578 1524
rect -7544 1418 -7528 1524
rect -7594 1406 -7528 1418
rect -7498 1524 -7432 1536
rect -7498 1418 -7482 1524
rect -7448 1418 -7432 1524
rect -7498 1406 -7432 1418
rect -7402 1524 -7336 1536
rect -7402 1418 -7386 1524
rect -7352 1418 -7336 1524
rect -7402 1406 -7336 1418
rect -7306 1524 -7240 1536
rect -7306 1418 -7290 1524
rect -7256 1418 -7240 1524
rect -7306 1406 -7240 1418
rect -7210 1524 -7144 1536
rect -7210 1418 -7194 1524
rect -7160 1418 -7144 1524
rect -7210 1406 -7144 1418
rect -7114 1524 -7052 1536
rect -7114 1418 -7098 1524
rect -7064 1418 -7052 1524
rect -7114 1406 -7052 1418
rect -7022 1524 -6964 1536
rect -7022 1418 -7010 1524
rect -6976 1418 -6964 1524
rect -7022 1406 -6964 1418
rect -6791 1524 -6733 1536
rect -6791 1418 -6779 1524
rect -6745 1418 -6733 1524
rect -6791 1406 -6733 1418
rect -6703 1524 -6641 1536
rect -6703 1418 -6691 1524
rect -6657 1418 -6641 1524
rect -6703 1406 -6641 1418
rect -6611 1524 -6545 1536
rect -6611 1418 -6595 1524
rect -6561 1418 -6545 1524
rect -6611 1406 -6545 1418
rect -6515 1524 -6449 1536
rect -6515 1418 -6499 1524
rect -6465 1418 -6449 1524
rect -6515 1406 -6449 1418
rect -6419 1524 -6353 1536
rect -6419 1418 -6403 1524
rect -6369 1418 -6353 1524
rect -6419 1406 -6353 1418
rect -6323 1524 -6257 1536
rect -6323 1418 -6307 1524
rect -6273 1418 -6257 1524
rect -6323 1406 -6257 1418
rect -6227 1524 -6161 1536
rect -6227 1418 -6211 1524
rect -6177 1418 -6161 1524
rect -6227 1406 -6161 1418
rect -6131 1524 -6065 1536
rect -6131 1418 -6115 1524
rect -6081 1418 -6065 1524
rect -6131 1406 -6065 1418
rect -6035 1524 -5969 1536
rect -6035 1418 -6019 1524
rect -5985 1418 -5969 1524
rect -6035 1406 -5969 1418
rect -5939 1524 -5873 1536
rect -5939 1418 -5923 1524
rect -5889 1418 -5873 1524
rect -5939 1406 -5873 1418
rect -5843 1524 -5777 1536
rect -5843 1418 -5827 1524
rect -5793 1418 -5777 1524
rect -5843 1406 -5777 1418
rect -5747 1524 -5681 1536
rect -5747 1418 -5731 1524
rect -5697 1418 -5681 1524
rect -5747 1406 -5681 1418
rect -5651 1524 -5585 1536
rect -5651 1418 -5635 1524
rect -5601 1418 -5585 1524
rect -5651 1406 -5585 1418
rect -5555 1524 -5493 1536
rect -5555 1418 -5539 1524
rect -5505 1418 -5493 1524
rect -5555 1406 -5493 1418
rect -5463 1524 -5405 1536
rect -5463 1418 -5451 1524
rect -5417 1418 -5405 1524
rect -5463 1406 -5405 1418
rect -5059 1524 -5001 1536
rect -5059 1418 -5047 1524
rect -5013 1418 -5001 1524
rect -5059 1406 -5001 1418
rect -4971 1524 -4909 1536
rect -4971 1418 -4959 1524
rect -4925 1418 -4909 1524
rect -4971 1406 -4909 1418
rect -4879 1524 -4813 1536
rect -4879 1418 -4863 1524
rect -4829 1418 -4813 1524
rect -4879 1406 -4813 1418
rect -4783 1524 -4717 1536
rect -4783 1418 -4767 1524
rect -4733 1418 -4717 1524
rect -4783 1406 -4717 1418
rect -4687 1524 -4621 1536
rect -4687 1418 -4671 1524
rect -4637 1418 -4621 1524
rect -4687 1406 -4621 1418
rect -4591 1524 -4525 1536
rect -4591 1418 -4575 1524
rect -4541 1418 -4525 1524
rect -4591 1406 -4525 1418
rect -4495 1524 -4429 1536
rect -4495 1418 -4479 1524
rect -4445 1418 -4429 1524
rect -4495 1406 -4429 1418
rect -4399 1524 -4333 1536
rect -4399 1418 -4383 1524
rect -4349 1418 -4333 1524
rect -4399 1406 -4333 1418
rect -4303 1524 -4237 1536
rect -4303 1418 -4287 1524
rect -4253 1418 -4237 1524
rect -4303 1406 -4237 1418
rect -4207 1524 -4141 1536
rect -4207 1418 -4191 1524
rect -4157 1418 -4141 1524
rect -4207 1406 -4141 1418
rect -4111 1524 -4045 1536
rect -4111 1418 -4095 1524
rect -4061 1418 -4045 1524
rect -4111 1406 -4045 1418
rect -4015 1524 -3949 1536
rect -4015 1418 -3999 1524
rect -3965 1418 -3949 1524
rect -4015 1406 -3949 1418
rect -3919 1524 -3853 1536
rect -3919 1418 -3903 1524
rect -3869 1418 -3853 1524
rect -3919 1406 -3853 1418
rect -3823 1524 -3761 1536
rect -3823 1418 -3807 1524
rect -3773 1418 -3761 1524
rect -3823 1406 -3761 1418
rect -3731 1524 -3673 1536
rect -3731 1418 -3719 1524
rect -3685 1418 -3673 1524
rect -3731 1406 -3673 1418
rect -3500 1524 -3442 1536
rect -3500 1418 -3488 1524
rect -3454 1418 -3442 1524
rect -3500 1406 -3442 1418
rect -3412 1524 -3350 1536
rect -3412 1418 -3400 1524
rect -3366 1418 -3350 1524
rect -3412 1406 -3350 1418
rect -3320 1524 -3254 1536
rect -3320 1418 -3304 1524
rect -3270 1418 -3254 1524
rect -3320 1406 -3254 1418
rect -3224 1524 -3158 1536
rect -3224 1418 -3208 1524
rect -3174 1418 -3158 1524
rect -3224 1406 -3158 1418
rect -3128 1524 -3062 1536
rect -3128 1418 -3112 1524
rect -3078 1418 -3062 1524
rect -3128 1406 -3062 1418
rect -3032 1524 -2966 1536
rect -3032 1418 -3016 1524
rect -2982 1418 -2966 1524
rect -3032 1406 -2966 1418
rect -2936 1524 -2870 1536
rect -2936 1418 -2920 1524
rect -2886 1418 -2870 1524
rect -2936 1406 -2870 1418
rect -2840 1524 -2774 1536
rect -2840 1418 -2824 1524
rect -2790 1418 -2774 1524
rect -2840 1406 -2774 1418
rect -2744 1524 -2678 1536
rect -2744 1418 -2728 1524
rect -2694 1418 -2678 1524
rect -2744 1406 -2678 1418
rect -2648 1524 -2582 1536
rect -2648 1418 -2632 1524
rect -2598 1418 -2582 1524
rect -2648 1406 -2582 1418
rect -2552 1524 -2486 1536
rect -2552 1418 -2536 1524
rect -2502 1418 -2486 1524
rect -2552 1406 -2486 1418
rect -2456 1524 -2390 1536
rect -2456 1418 -2440 1524
rect -2406 1418 -2390 1524
rect -2456 1406 -2390 1418
rect -2360 1524 -2294 1536
rect -2360 1418 -2344 1524
rect -2310 1418 -2294 1524
rect -2360 1406 -2294 1418
rect -2264 1524 -2202 1536
rect -2264 1418 -2248 1524
rect -2214 1418 -2202 1524
rect -2264 1406 -2202 1418
rect -2172 1524 -2114 1536
rect -2172 1418 -2160 1524
rect -2126 1418 -2114 1524
rect -2172 1406 -2114 1418
rect -1768 1524 -1710 1536
rect -1768 1418 -1756 1524
rect -1722 1418 -1710 1524
rect -1768 1406 -1710 1418
rect -1680 1524 -1618 1536
rect -1680 1418 -1668 1524
rect -1634 1418 -1618 1524
rect -1680 1406 -1618 1418
rect -1588 1524 -1522 1536
rect -1588 1418 -1572 1524
rect -1538 1418 -1522 1524
rect -1588 1406 -1522 1418
rect -1492 1524 -1426 1536
rect -1492 1418 -1476 1524
rect -1442 1418 -1426 1524
rect -1492 1406 -1426 1418
rect -1396 1524 -1330 1536
rect -1396 1418 -1380 1524
rect -1346 1418 -1330 1524
rect -1396 1406 -1330 1418
rect -1300 1524 -1234 1536
rect -1300 1418 -1284 1524
rect -1250 1418 -1234 1524
rect -1300 1406 -1234 1418
rect -1204 1524 -1138 1536
rect -1204 1418 -1188 1524
rect -1154 1418 -1138 1524
rect -1204 1406 -1138 1418
rect -1108 1524 -1042 1536
rect -1108 1418 -1092 1524
rect -1058 1418 -1042 1524
rect -1108 1406 -1042 1418
rect -1012 1524 -946 1536
rect -1012 1418 -996 1524
rect -962 1418 -946 1524
rect -1012 1406 -946 1418
rect -916 1524 -850 1536
rect -916 1418 -900 1524
rect -866 1418 -850 1524
rect -916 1406 -850 1418
rect -820 1524 -754 1536
rect -820 1418 -804 1524
rect -770 1418 -754 1524
rect -820 1406 -754 1418
rect -724 1524 -658 1536
rect -724 1418 -708 1524
rect -674 1418 -658 1524
rect -724 1406 -658 1418
rect -628 1524 -562 1536
rect -628 1418 -612 1524
rect -578 1418 -562 1524
rect -628 1406 -562 1418
rect -532 1524 -470 1536
rect -532 1418 -516 1524
rect -482 1418 -470 1524
rect -532 1406 -470 1418
rect -440 1524 -382 1536
rect -440 1418 -428 1524
rect -394 1418 -382 1524
rect -440 1406 -382 1418
rect -209 1524 -151 1536
rect -209 1418 -197 1524
rect -163 1418 -151 1524
rect -209 1406 -151 1418
rect -121 1524 -59 1536
rect -121 1418 -109 1524
rect -75 1418 -59 1524
rect -121 1406 -59 1418
rect -29 1524 37 1536
rect -29 1418 -13 1524
rect 21 1418 37 1524
rect -29 1406 37 1418
rect 67 1524 133 1536
rect 67 1418 83 1524
rect 117 1418 133 1524
rect 67 1406 133 1418
rect 163 1524 229 1536
rect 163 1418 179 1524
rect 213 1418 229 1524
rect 163 1406 229 1418
rect 259 1524 325 1536
rect 259 1418 275 1524
rect 309 1418 325 1524
rect 259 1406 325 1418
rect 355 1524 421 1536
rect 355 1418 371 1524
rect 405 1418 421 1524
rect 355 1406 421 1418
rect 451 1524 517 1536
rect 451 1418 467 1524
rect 501 1418 517 1524
rect 451 1406 517 1418
rect 547 1524 613 1536
rect 547 1418 563 1524
rect 597 1418 613 1524
rect 547 1406 613 1418
rect 643 1524 709 1536
rect 643 1418 659 1524
rect 693 1418 709 1524
rect 643 1406 709 1418
rect 739 1524 805 1536
rect 739 1418 755 1524
rect 789 1418 805 1524
rect 739 1406 805 1418
rect 835 1524 901 1536
rect 835 1418 851 1524
rect 885 1418 901 1524
rect 835 1406 901 1418
rect 931 1524 997 1536
rect 931 1418 947 1524
rect 981 1418 997 1524
rect 931 1406 997 1418
rect 1027 1524 1089 1536
rect 1027 1418 1043 1524
rect 1077 1418 1089 1524
rect 1027 1406 1089 1418
rect 1119 1524 1177 1536
rect 1119 1418 1131 1524
rect 1165 1418 1177 1524
rect 1119 1406 1177 1418
rect 7360 774 7372 1550
rect 7406 774 7422 1550
rect 7360 762 7422 774
rect 7452 762 7518 1562
rect 7548 762 7614 1562
rect 7644 762 7710 1562
rect 7740 1550 7802 1562
rect 7740 774 7756 1550
rect 7790 774 7802 1550
rect 7740 762 7802 774
rect 8308 1550 8370 1562
rect 8308 774 8320 1550
rect 8354 774 8370 1550
rect 8308 762 8370 774
rect 8400 762 8466 1562
rect 8496 762 8562 1562
rect 8592 762 8658 1562
rect 8688 1550 8750 1562
rect 8688 774 8704 1550
rect 8738 774 8750 1550
rect 8688 762 8750 774
rect 9244 1550 9306 1562
rect 9244 774 9256 1550
rect 9290 774 9306 1550
rect 9244 762 9306 774
rect 9336 762 9402 1562
rect 9432 762 9498 1562
rect 9528 762 9594 1562
rect 9624 1550 9686 1562
rect 9624 774 9640 1550
rect 9674 774 9686 1550
rect 9624 762 9686 774
rect 10175 1551 10237 1563
rect 10175 775 10187 1551
rect 10221 775 10237 1551
rect 10175 763 10237 775
rect 10267 763 10333 1563
rect 10363 763 10429 1563
rect 10459 763 10525 1563
rect 10555 1551 10617 1563
rect 10555 775 10571 1551
rect 10605 775 10617 1551
rect 10555 763 10617 775
rect 11102 1550 11164 1562
rect -24363 519 -23963 531
rect -24363 485 -24351 519
rect -23975 485 -23963 519
rect -24363 469 -23963 485
rect -24363 373 -23963 439
rect -23254 519 -22854 531
rect -23254 485 -23242 519
rect -22866 485 -22854 519
rect -23254 469 -22854 485
rect -23254 373 -22854 439
rect -22372 519 -21972 531
rect -22372 485 -22360 519
rect -21984 485 -21972 519
rect -22372 469 -21972 485
rect -22372 373 -21972 439
rect -21072 519 -20672 531
rect -21072 485 -21060 519
rect -20684 485 -20672 519
rect -21072 469 -20672 485
rect -21072 373 -20672 439
rect -19963 519 -19563 531
rect -19963 485 -19951 519
rect -19575 485 -19563 519
rect -19963 469 -19563 485
rect -19963 373 -19563 439
rect -19081 519 -18681 531
rect -19081 485 -19069 519
rect -18693 485 -18681 519
rect -19081 469 -18681 485
rect -19081 373 -18681 439
rect -17781 519 -17381 531
rect -17781 485 -17769 519
rect -17393 485 -17381 519
rect -17781 469 -17381 485
rect -17781 373 -17381 439
rect -16672 519 -16272 531
rect -16672 485 -16660 519
rect -16284 485 -16272 519
rect -16672 469 -16272 485
rect -16672 373 -16272 439
rect -15790 519 -15390 531
rect -15790 485 -15778 519
rect -15402 485 -15390 519
rect -15790 469 -15390 485
rect -15790 373 -15390 439
rect -14490 519 -14090 531
rect -14490 485 -14478 519
rect -14102 485 -14090 519
rect -14490 469 -14090 485
rect -14490 373 -14090 439
rect -13381 519 -12981 531
rect -13381 485 -13369 519
rect -12993 485 -12981 519
rect -13381 469 -12981 485
rect -13381 373 -12981 439
rect -12499 519 -12099 531
rect -12499 485 -12487 519
rect -12111 485 -12099 519
rect -12499 469 -12099 485
rect -12499 373 -12099 439
rect -11199 519 -10799 531
rect -11199 485 -11187 519
rect -10811 485 -10799 519
rect -11199 469 -10799 485
rect -11199 373 -10799 439
rect -10090 519 -9690 531
rect -10090 485 -10078 519
rect -9702 485 -9690 519
rect -10090 469 -9690 485
rect -10090 373 -9690 439
rect -9208 519 -8808 531
rect -9208 485 -9196 519
rect -8820 485 -8808 519
rect -9208 469 -8808 485
rect -9208 373 -8808 439
rect -7909 519 -7509 531
rect -7909 485 -7897 519
rect -7521 485 -7509 519
rect -7909 469 -7509 485
rect -7909 373 -7509 439
rect -6800 519 -6400 531
rect -6800 485 -6788 519
rect -6412 485 -6400 519
rect -6800 469 -6400 485
rect -6800 373 -6400 439
rect -5918 519 -5518 531
rect -5918 485 -5906 519
rect -5530 485 -5518 519
rect -5918 469 -5518 485
rect -5918 373 -5518 439
rect -4618 519 -4218 531
rect -4618 485 -4606 519
rect -4230 485 -4218 519
rect -4618 469 -4218 485
rect -4618 373 -4218 439
rect -3509 519 -3109 531
rect -3509 485 -3497 519
rect -3121 485 -3109 519
rect -3509 469 -3109 485
rect -3509 373 -3109 439
rect -2627 519 -2227 531
rect -2627 485 -2615 519
rect -2239 485 -2227 519
rect -2627 469 -2227 485
rect -2627 373 -2227 439
rect -1327 519 -927 531
rect -1327 485 -1315 519
rect -939 485 -927 519
rect -1327 469 -927 485
rect -1327 373 -927 439
rect -218 519 182 531
rect -218 485 -206 519
rect 170 485 182 519
rect -218 469 182 485
rect -218 373 182 439
rect 664 519 1064 531
rect 664 485 676 519
rect 1052 485 1064 519
rect 664 469 1064 485
rect 664 373 1064 439
rect 11102 774 11114 1550
rect 11148 774 11164 1550
rect 11102 762 11164 774
rect 11194 762 11260 1562
rect 11290 762 11356 1562
rect 11386 762 11452 1562
rect 11482 1550 11544 1562
rect 11482 774 11498 1550
rect 11532 774 11544 1550
rect 12157 1508 12219 1520
rect 12157 1332 12169 1508
rect 12203 1332 12219 1508
rect 12157 1320 12219 1332
rect 12249 1508 12315 1520
rect 12249 1332 12265 1508
rect 12299 1332 12315 1508
rect 12249 1320 12315 1332
rect 12345 1508 12407 1520
rect 12345 1332 12361 1508
rect 12395 1332 12407 1508
rect 12923 1443 13123 1455
rect 12923 1409 12935 1443
rect 13111 1409 13123 1443
rect 12923 1397 13123 1409
rect 12923 1355 13123 1367
rect 12345 1320 12407 1332
rect 12923 1321 12935 1355
rect 13111 1321 13123 1355
rect 12923 1309 13123 1321
rect 11482 762 11544 774
rect -24363 327 -23963 343
rect -24363 293 -24351 327
rect -23975 293 -23963 327
rect -23254 327 -22854 343
rect -24363 281 -23963 293
rect -23254 293 -23242 327
rect -22866 293 -22854 327
rect -22372 327 -21972 343
rect -23254 281 -22854 293
rect -22372 293 -22360 327
rect -21984 293 -21972 327
rect -21072 327 -20672 343
rect -22372 281 -21972 293
rect -21072 293 -21060 327
rect -20684 293 -20672 327
rect -19963 327 -19563 343
rect -21072 281 -20672 293
rect -19963 293 -19951 327
rect -19575 293 -19563 327
rect -19081 327 -18681 343
rect -19963 281 -19563 293
rect -19081 293 -19069 327
rect -18693 293 -18681 327
rect -17781 327 -17381 343
rect -19081 281 -18681 293
rect -17781 293 -17769 327
rect -17393 293 -17381 327
rect -16672 327 -16272 343
rect -17781 281 -17381 293
rect -16672 293 -16660 327
rect -16284 293 -16272 327
rect -15790 327 -15390 343
rect -16672 281 -16272 293
rect -15790 293 -15778 327
rect -15402 293 -15390 327
rect -14490 327 -14090 343
rect -15790 281 -15390 293
rect -14490 293 -14478 327
rect -14102 293 -14090 327
rect -13381 327 -12981 343
rect -14490 281 -14090 293
rect -13381 293 -13369 327
rect -12993 293 -12981 327
rect -12499 327 -12099 343
rect -13381 281 -12981 293
rect -12499 293 -12487 327
rect -12111 293 -12099 327
rect -11199 327 -10799 343
rect -12499 281 -12099 293
rect -11199 293 -11187 327
rect -10811 293 -10799 327
rect -10090 327 -9690 343
rect -11199 281 -10799 293
rect -10090 293 -10078 327
rect -9702 293 -9690 327
rect -9208 327 -8808 343
rect -10090 281 -9690 293
rect -9208 293 -9196 327
rect -8820 293 -8808 327
rect -7909 327 -7509 343
rect -9208 281 -8808 293
rect -7909 293 -7897 327
rect -7521 293 -7509 327
rect -6800 327 -6400 343
rect -7909 281 -7509 293
rect -6800 293 -6788 327
rect -6412 293 -6400 327
rect -5918 327 -5518 343
rect -6800 281 -6400 293
rect -5918 293 -5906 327
rect -5530 293 -5518 327
rect -4618 327 -4218 343
rect -5918 281 -5518 293
rect -4618 293 -4606 327
rect -4230 293 -4218 327
rect -3509 327 -3109 343
rect -4618 281 -4218 293
rect -3509 293 -3497 327
rect -3121 293 -3109 327
rect -2627 327 -2227 343
rect -3509 281 -3109 293
rect -2627 293 -2615 327
rect -2239 293 -2227 327
rect -1327 327 -927 343
rect -2627 281 -2227 293
rect -1327 293 -1315 327
rect -939 293 -927 327
rect -218 327 182 343
rect -1327 281 -927 293
rect -218 293 -206 327
rect 170 293 182 327
rect 664 327 1064 343
rect -218 281 182 293
rect 664 293 676 327
rect 1052 293 1064 327
rect 664 281 1064 293
rect 5658 -1067 5858 -1055
rect 5658 -1101 5670 -1067
rect 5846 -1101 5858 -1067
rect 6098 -1067 6298 -1055
rect 5658 -1113 5858 -1101
rect 5658 -1155 5858 -1143
rect 5658 -1189 5670 -1155
rect 5846 -1189 5858 -1155
rect 6098 -1101 6110 -1067
rect 6286 -1101 6298 -1067
rect 6538 -1067 6738 -1055
rect 6098 -1113 6298 -1101
rect 6098 -1155 6298 -1143
rect 5658 -1201 5858 -1189
rect 6098 -1189 6110 -1155
rect 6286 -1189 6298 -1155
rect 6538 -1101 6550 -1067
rect 6726 -1101 6738 -1067
rect 6538 -1113 6738 -1101
rect 6538 -1155 6738 -1143
rect 6098 -1201 6298 -1189
rect 6538 -1189 6550 -1155
rect 6726 -1189 6738 -1155
rect 6538 -1201 6738 -1189
rect 7360 -2050 7422 -2038
rect -24213 -2769 -23813 -2757
rect -24213 -2803 -24201 -2769
rect -23825 -2803 -23813 -2769
rect -23628 -2769 -23428 -2757
rect -24213 -2819 -23813 -2803
rect -23628 -2803 -23616 -2769
rect -23440 -2803 -23428 -2769
rect -23628 -2815 -23428 -2803
rect -24213 -2915 -23813 -2849
rect -23628 -2857 -23428 -2845
rect -23628 -2891 -23616 -2857
rect -23440 -2891 -23428 -2857
rect -23628 -2903 -23428 -2891
rect -22176 -2769 -21776 -2757
rect -22176 -2803 -22164 -2769
rect -21788 -2803 -21776 -2769
rect -21608 -2769 -21408 -2757
rect -22176 -2819 -21776 -2803
rect -21608 -2803 -21596 -2769
rect -21420 -2803 -21408 -2769
rect -21608 -2815 -21408 -2803
rect -22176 -2915 -21776 -2849
rect -21608 -2857 -21408 -2845
rect -21608 -2891 -21596 -2857
rect -21420 -2891 -21408 -2857
rect -21608 -2903 -21408 -2891
rect -20446 -2769 -20046 -2757
rect -20446 -2803 -20434 -2769
rect -20058 -2803 -20046 -2769
rect -19867 -2769 -19667 -2757
rect -20446 -2819 -20046 -2803
rect -19867 -2803 -19855 -2769
rect -19679 -2803 -19667 -2769
rect -19867 -2815 -19667 -2803
rect -20446 -2915 -20046 -2849
rect -19867 -2857 -19667 -2845
rect -19867 -2891 -19855 -2857
rect -19679 -2891 -19667 -2857
rect -19867 -2903 -19667 -2891
rect -18686 -2769 -18286 -2757
rect -18686 -2803 -18674 -2769
rect -18298 -2803 -18286 -2769
rect -18088 -2769 -17888 -2757
rect -18686 -2819 -18286 -2803
rect -18088 -2803 -18076 -2769
rect -17900 -2803 -17888 -2769
rect -18088 -2815 -17888 -2803
rect 7360 -2826 7372 -2050
rect 7406 -2826 7422 -2050
rect 7360 -2838 7422 -2826
rect 7452 -2838 7518 -2038
rect 7548 -2838 7614 -2038
rect 7644 -2838 7710 -2038
rect 7740 -2050 7802 -2038
rect 7740 -2826 7756 -2050
rect 7790 -2826 7802 -2050
rect 7740 -2838 7802 -2826
rect 8308 -2050 8370 -2038
rect 8308 -2826 8320 -2050
rect 8354 -2826 8370 -2050
rect 8308 -2838 8370 -2826
rect 8400 -2838 8466 -2038
rect 8496 -2838 8562 -2038
rect 8592 -2838 8658 -2038
rect 8688 -2050 8750 -2038
rect 8688 -2826 8704 -2050
rect 8738 -2826 8750 -2050
rect 8688 -2838 8750 -2826
rect 9244 -2050 9306 -2038
rect 9244 -2826 9256 -2050
rect 9290 -2826 9306 -2050
rect 9244 -2838 9306 -2826
rect 9336 -2838 9402 -2038
rect 9432 -2838 9498 -2038
rect 9528 -2838 9594 -2038
rect 9624 -2050 9686 -2038
rect 9624 -2826 9640 -2050
rect 9674 -2826 9686 -2050
rect 9624 -2838 9686 -2826
rect 10175 -2050 10237 -2038
rect 10175 -2826 10187 -2050
rect 10221 -2826 10237 -2050
rect 10175 -2838 10237 -2826
rect 10267 -2838 10333 -2038
rect 10363 -2838 10429 -2038
rect 10459 -2838 10525 -2038
rect 10555 -2050 10617 -2038
rect 10555 -2826 10571 -2050
rect 10605 -2826 10617 -2050
rect 10555 -2838 10617 -2826
rect 11102 -2050 11164 -2038
rect 11102 -2826 11114 -2050
rect 11148 -2826 11164 -2050
rect 11102 -2838 11164 -2826
rect 11194 -2838 11260 -2038
rect 11290 -2838 11356 -2038
rect 11386 -2838 11452 -2038
rect 11482 -2050 11544 -2038
rect 11482 -2826 11498 -2050
rect 11532 -2826 11544 -2050
rect 11482 -2838 11544 -2826
rect -18686 -2915 -18286 -2849
rect -18088 -2857 -17888 -2845
rect -18088 -2891 -18076 -2857
rect -17900 -2891 -17888 -2857
rect -18088 -2903 -17888 -2891
rect -24213 -2961 -23813 -2945
rect -24213 -2995 -24201 -2961
rect -23825 -2995 -23813 -2961
rect -24213 -3007 -23813 -2995
rect -22176 -2961 -21776 -2945
rect -22176 -2995 -22164 -2961
rect -21788 -2995 -21776 -2961
rect -22176 -3007 -21776 -2995
rect -20446 -2961 -20046 -2945
rect -20446 -2995 -20434 -2961
rect -20058 -2995 -20046 -2961
rect -20446 -3007 -20046 -2995
rect -18686 -2961 -18286 -2945
rect -18686 -2995 -18674 -2961
rect -18298 -2995 -18286 -2961
rect -18686 -3007 -18286 -2995
rect 7360 -2978 7422 -2966
rect 7360 -3754 7372 -2978
rect 7406 -3754 7422 -2978
rect 7360 -3766 7422 -3754
rect 7452 -3766 7518 -2966
rect 7548 -3766 7614 -2966
rect 7644 -3766 7710 -2966
rect 7740 -2978 7802 -2966
rect 7740 -3754 7756 -2978
rect 7790 -3754 7802 -2978
rect 7740 -3766 7802 -3754
rect 8308 -2978 8370 -2966
rect 8308 -3754 8320 -2978
rect 8354 -3754 8370 -2978
rect 8308 -3766 8370 -3754
rect 8400 -3766 8466 -2966
rect 8496 -3766 8562 -2966
rect 8592 -3766 8658 -2966
rect 8688 -2978 8750 -2966
rect 8688 -3754 8704 -2978
rect 8738 -3754 8750 -2978
rect 8688 -3766 8750 -3754
rect 9244 -2978 9306 -2966
rect 9244 -3754 9256 -2978
rect 9290 -3754 9306 -2978
rect 9244 -3766 9306 -3754
rect 9336 -3766 9402 -2966
rect 9432 -3766 9498 -2966
rect 9528 -3766 9594 -2966
rect 9624 -2978 9686 -2966
rect 9624 -3754 9640 -2978
rect 9674 -3754 9686 -2978
rect 9624 -3766 9686 -3754
rect 10175 -2977 10237 -2965
rect 10175 -3753 10187 -2977
rect 10221 -3753 10237 -2977
rect 10175 -3765 10237 -3753
rect 10267 -3765 10333 -2965
rect 10363 -3765 10429 -2965
rect 10459 -3765 10525 -2965
rect 10555 -2977 10617 -2965
rect 10555 -3753 10571 -2977
rect 10605 -3753 10617 -2977
rect 10555 -3765 10617 -3753
rect 11102 -2978 11164 -2966
rect -24162 -4581 -23762 -4569
rect -24162 -4615 -24150 -4581
rect -23774 -4615 -23762 -4581
rect -23584 -4581 -23384 -4569
rect -24162 -4631 -23762 -4615
rect -23584 -4615 -23572 -4581
rect -23396 -4615 -23384 -4581
rect -23584 -4627 -23384 -4615
rect -24162 -4727 -23762 -4661
rect -23584 -4669 -23384 -4657
rect -23584 -4703 -23572 -4669
rect -23396 -4703 -23384 -4669
rect -23584 -4715 -23384 -4703
rect 11102 -3754 11114 -2978
rect 11148 -3754 11164 -2978
rect 11102 -3766 11164 -3754
rect 11194 -3766 11260 -2966
rect 11290 -3766 11356 -2966
rect 11386 -3766 11452 -2966
rect 11482 -2978 11544 -2966
rect 11482 -3754 11498 -2978
rect 11532 -3754 11544 -2978
rect 12157 -3020 12219 -3008
rect 12157 -3196 12169 -3020
rect 12203 -3196 12219 -3020
rect 12157 -3208 12219 -3196
rect 12249 -3020 12315 -3008
rect 12249 -3196 12265 -3020
rect 12299 -3196 12315 -3020
rect 12249 -3208 12315 -3196
rect 12345 -3020 12407 -3008
rect 12345 -3196 12361 -3020
rect 12395 -3196 12407 -3020
rect 12923 -3085 13123 -3073
rect 12923 -3119 12935 -3085
rect 13111 -3119 13123 -3085
rect 12923 -3131 13123 -3119
rect 12923 -3173 13123 -3161
rect 12345 -3208 12407 -3196
rect 12923 -3207 12935 -3173
rect 13111 -3207 13123 -3173
rect 12923 -3219 13123 -3207
rect 11482 -3766 11544 -3754
rect -22426 -4581 -22026 -4569
rect -22426 -4615 -22414 -4581
rect -22038 -4615 -22026 -4581
rect -21846 -4581 -21646 -4569
rect -22426 -4631 -22026 -4615
rect -21846 -4615 -21834 -4581
rect -21658 -4615 -21646 -4581
rect -21846 -4627 -21646 -4615
rect -22426 -4727 -22026 -4661
rect -21846 -4669 -21646 -4657
rect -21846 -4703 -21834 -4669
rect -21658 -4703 -21646 -4669
rect -21846 -4715 -21646 -4703
rect -24162 -4773 -23762 -4757
rect -24162 -4807 -24150 -4773
rect -23774 -4807 -23762 -4773
rect -24162 -4819 -23762 -4807
rect -22426 -4773 -22026 -4757
rect -22426 -4807 -22414 -4773
rect -22038 -4807 -22026 -4773
rect -22426 -4819 -22026 -4807
rect -20737 -5036 -20679 -5024
rect -20737 -5142 -20725 -5036
rect -20691 -5142 -20679 -5036
rect -20737 -5154 -20679 -5142
rect -20649 -5036 -20587 -5024
rect -20649 -5142 -20637 -5036
rect -20603 -5142 -20587 -5036
rect -20649 -5154 -20587 -5142
rect -20557 -5036 -20491 -5024
rect -20557 -5142 -20541 -5036
rect -20507 -5142 -20491 -5036
rect -20557 -5154 -20491 -5142
rect -20461 -5036 -20395 -5024
rect -20461 -5142 -20445 -5036
rect -20411 -5142 -20395 -5036
rect -20461 -5154 -20395 -5142
rect -20365 -5036 -20299 -5024
rect -20365 -5142 -20349 -5036
rect -20315 -5142 -20299 -5036
rect -20365 -5154 -20299 -5142
rect -20269 -5036 -20203 -5024
rect -20269 -5142 -20253 -5036
rect -20219 -5142 -20203 -5036
rect -20269 -5154 -20203 -5142
rect -20173 -5036 -20107 -5024
rect -20173 -5142 -20157 -5036
rect -20123 -5142 -20107 -5036
rect -20173 -5154 -20107 -5142
rect -20077 -5036 -20011 -5024
rect -20077 -5142 -20061 -5036
rect -20027 -5142 -20011 -5036
rect -20077 -5154 -20011 -5142
rect -19981 -5036 -19915 -5024
rect -19981 -5142 -19965 -5036
rect -19931 -5142 -19915 -5036
rect -19981 -5154 -19915 -5142
rect -19885 -5036 -19819 -5024
rect -19885 -5142 -19869 -5036
rect -19835 -5142 -19819 -5036
rect -19885 -5154 -19819 -5142
rect -19789 -5036 -19723 -5024
rect -19789 -5142 -19773 -5036
rect -19739 -5142 -19723 -5036
rect -19789 -5154 -19723 -5142
rect -19693 -5036 -19627 -5024
rect -19693 -5142 -19677 -5036
rect -19643 -5142 -19627 -5036
rect -19693 -5154 -19627 -5142
rect -19597 -5036 -19531 -5024
rect -19597 -5142 -19581 -5036
rect -19547 -5142 -19531 -5036
rect -19597 -5154 -19531 -5142
rect -19501 -5036 -19439 -5024
rect -19501 -5142 -19485 -5036
rect -19451 -5142 -19439 -5036
rect -19501 -5154 -19439 -5142
rect -19409 -5036 -19351 -5024
rect -19409 -5142 -19397 -5036
rect -19363 -5142 -19351 -5036
rect -19409 -5154 -19351 -5142
rect -19178 -5036 -19120 -5024
rect -19178 -5142 -19166 -5036
rect -19132 -5142 -19120 -5036
rect -19178 -5154 -19120 -5142
rect -19090 -5036 -19028 -5024
rect -19090 -5142 -19078 -5036
rect -19044 -5142 -19028 -5036
rect -19090 -5154 -19028 -5142
rect -18998 -5036 -18932 -5024
rect -18998 -5142 -18982 -5036
rect -18948 -5142 -18932 -5036
rect -18998 -5154 -18932 -5142
rect -18902 -5036 -18836 -5024
rect -18902 -5142 -18886 -5036
rect -18852 -5142 -18836 -5036
rect -18902 -5154 -18836 -5142
rect -18806 -5036 -18740 -5024
rect -18806 -5142 -18790 -5036
rect -18756 -5142 -18740 -5036
rect -18806 -5154 -18740 -5142
rect -18710 -5036 -18644 -5024
rect -18710 -5142 -18694 -5036
rect -18660 -5142 -18644 -5036
rect -18710 -5154 -18644 -5142
rect -18614 -5036 -18548 -5024
rect -18614 -5142 -18598 -5036
rect -18564 -5142 -18548 -5036
rect -18614 -5154 -18548 -5142
rect -18518 -5036 -18452 -5024
rect -18518 -5142 -18502 -5036
rect -18468 -5142 -18452 -5036
rect -18518 -5154 -18452 -5142
rect -18422 -5036 -18356 -5024
rect -18422 -5142 -18406 -5036
rect -18372 -5142 -18356 -5036
rect -18422 -5154 -18356 -5142
rect -18326 -5036 -18260 -5024
rect -18326 -5142 -18310 -5036
rect -18276 -5142 -18260 -5036
rect -18326 -5154 -18260 -5142
rect -18230 -5036 -18164 -5024
rect -18230 -5142 -18214 -5036
rect -18180 -5142 -18164 -5036
rect -18230 -5154 -18164 -5142
rect -18134 -5036 -18068 -5024
rect -18134 -5142 -18118 -5036
rect -18084 -5142 -18068 -5036
rect -18134 -5154 -18068 -5142
rect -18038 -5036 -17972 -5024
rect -18038 -5142 -18022 -5036
rect -17988 -5142 -17972 -5036
rect -18038 -5154 -17972 -5142
rect -17942 -5036 -17880 -5024
rect -17942 -5142 -17926 -5036
rect -17892 -5142 -17880 -5036
rect -17942 -5154 -17880 -5142
rect -17850 -5036 -17792 -5024
rect -17850 -5142 -17838 -5036
rect -17804 -5142 -17792 -5036
rect -17850 -5154 -17792 -5142
rect -17446 -5036 -17388 -5024
rect -17446 -5142 -17434 -5036
rect -17400 -5142 -17388 -5036
rect -17446 -5154 -17388 -5142
rect -17358 -5036 -17296 -5024
rect -17358 -5142 -17346 -5036
rect -17312 -5142 -17296 -5036
rect -17358 -5154 -17296 -5142
rect -17266 -5036 -17200 -5024
rect -17266 -5142 -17250 -5036
rect -17216 -5142 -17200 -5036
rect -17266 -5154 -17200 -5142
rect -17170 -5036 -17104 -5024
rect -17170 -5142 -17154 -5036
rect -17120 -5142 -17104 -5036
rect -17170 -5154 -17104 -5142
rect -17074 -5036 -17008 -5024
rect -17074 -5142 -17058 -5036
rect -17024 -5142 -17008 -5036
rect -17074 -5154 -17008 -5142
rect -16978 -5036 -16912 -5024
rect -16978 -5142 -16962 -5036
rect -16928 -5142 -16912 -5036
rect -16978 -5154 -16912 -5142
rect -16882 -5036 -16816 -5024
rect -16882 -5142 -16866 -5036
rect -16832 -5142 -16816 -5036
rect -16882 -5154 -16816 -5142
rect -16786 -5036 -16720 -5024
rect -16786 -5142 -16770 -5036
rect -16736 -5142 -16720 -5036
rect -16786 -5154 -16720 -5142
rect -16690 -5036 -16624 -5024
rect -16690 -5142 -16674 -5036
rect -16640 -5142 -16624 -5036
rect -16690 -5154 -16624 -5142
rect -16594 -5036 -16528 -5024
rect -16594 -5142 -16578 -5036
rect -16544 -5142 -16528 -5036
rect -16594 -5154 -16528 -5142
rect -16498 -5036 -16432 -5024
rect -16498 -5142 -16482 -5036
rect -16448 -5142 -16432 -5036
rect -16498 -5154 -16432 -5142
rect -16402 -5036 -16336 -5024
rect -16402 -5142 -16386 -5036
rect -16352 -5142 -16336 -5036
rect -16402 -5154 -16336 -5142
rect -16306 -5036 -16240 -5024
rect -16306 -5142 -16290 -5036
rect -16256 -5142 -16240 -5036
rect -16306 -5154 -16240 -5142
rect -16210 -5036 -16148 -5024
rect -16210 -5142 -16194 -5036
rect -16160 -5142 -16148 -5036
rect -16210 -5154 -16148 -5142
rect -16118 -5036 -16060 -5024
rect -16118 -5142 -16106 -5036
rect -16072 -5142 -16060 -5036
rect -16118 -5154 -16060 -5142
rect -15887 -5036 -15829 -5024
rect -15887 -5142 -15875 -5036
rect -15841 -5142 -15829 -5036
rect -15887 -5154 -15829 -5142
rect -15799 -5036 -15737 -5024
rect -15799 -5142 -15787 -5036
rect -15753 -5142 -15737 -5036
rect -15799 -5154 -15737 -5142
rect -15707 -5036 -15641 -5024
rect -15707 -5142 -15691 -5036
rect -15657 -5142 -15641 -5036
rect -15707 -5154 -15641 -5142
rect -15611 -5036 -15545 -5024
rect -15611 -5142 -15595 -5036
rect -15561 -5142 -15545 -5036
rect -15611 -5154 -15545 -5142
rect -15515 -5036 -15449 -5024
rect -15515 -5142 -15499 -5036
rect -15465 -5142 -15449 -5036
rect -15515 -5154 -15449 -5142
rect -15419 -5036 -15353 -5024
rect -15419 -5142 -15403 -5036
rect -15369 -5142 -15353 -5036
rect -15419 -5154 -15353 -5142
rect -15323 -5036 -15257 -5024
rect -15323 -5142 -15307 -5036
rect -15273 -5142 -15257 -5036
rect -15323 -5154 -15257 -5142
rect -15227 -5036 -15161 -5024
rect -15227 -5142 -15211 -5036
rect -15177 -5142 -15161 -5036
rect -15227 -5154 -15161 -5142
rect -15131 -5036 -15065 -5024
rect -15131 -5142 -15115 -5036
rect -15081 -5142 -15065 -5036
rect -15131 -5154 -15065 -5142
rect -15035 -5036 -14969 -5024
rect -15035 -5142 -15019 -5036
rect -14985 -5142 -14969 -5036
rect -15035 -5154 -14969 -5142
rect -14939 -5036 -14873 -5024
rect -14939 -5142 -14923 -5036
rect -14889 -5142 -14873 -5036
rect -14939 -5154 -14873 -5142
rect -14843 -5036 -14777 -5024
rect -14843 -5142 -14827 -5036
rect -14793 -5142 -14777 -5036
rect -14843 -5154 -14777 -5142
rect -14747 -5036 -14681 -5024
rect -14747 -5142 -14731 -5036
rect -14697 -5142 -14681 -5036
rect -14747 -5154 -14681 -5142
rect -14651 -5036 -14589 -5024
rect -14651 -5142 -14635 -5036
rect -14601 -5142 -14589 -5036
rect -14651 -5154 -14589 -5142
rect -14559 -5036 -14501 -5024
rect -14559 -5142 -14547 -5036
rect -14513 -5142 -14501 -5036
rect -14559 -5154 -14501 -5142
rect -14155 -5036 -14097 -5024
rect -14155 -5142 -14143 -5036
rect -14109 -5142 -14097 -5036
rect -14155 -5154 -14097 -5142
rect -14067 -5036 -14005 -5024
rect -14067 -5142 -14055 -5036
rect -14021 -5142 -14005 -5036
rect -14067 -5154 -14005 -5142
rect -13975 -5036 -13909 -5024
rect -13975 -5142 -13959 -5036
rect -13925 -5142 -13909 -5036
rect -13975 -5154 -13909 -5142
rect -13879 -5036 -13813 -5024
rect -13879 -5142 -13863 -5036
rect -13829 -5142 -13813 -5036
rect -13879 -5154 -13813 -5142
rect -13783 -5036 -13717 -5024
rect -13783 -5142 -13767 -5036
rect -13733 -5142 -13717 -5036
rect -13783 -5154 -13717 -5142
rect -13687 -5036 -13621 -5024
rect -13687 -5142 -13671 -5036
rect -13637 -5142 -13621 -5036
rect -13687 -5154 -13621 -5142
rect -13591 -5036 -13525 -5024
rect -13591 -5142 -13575 -5036
rect -13541 -5142 -13525 -5036
rect -13591 -5154 -13525 -5142
rect -13495 -5036 -13429 -5024
rect -13495 -5142 -13479 -5036
rect -13445 -5142 -13429 -5036
rect -13495 -5154 -13429 -5142
rect -13399 -5036 -13333 -5024
rect -13399 -5142 -13383 -5036
rect -13349 -5142 -13333 -5036
rect -13399 -5154 -13333 -5142
rect -13303 -5036 -13237 -5024
rect -13303 -5142 -13287 -5036
rect -13253 -5142 -13237 -5036
rect -13303 -5154 -13237 -5142
rect -13207 -5036 -13141 -5024
rect -13207 -5142 -13191 -5036
rect -13157 -5142 -13141 -5036
rect -13207 -5154 -13141 -5142
rect -13111 -5036 -13045 -5024
rect -13111 -5142 -13095 -5036
rect -13061 -5142 -13045 -5036
rect -13111 -5154 -13045 -5142
rect -13015 -5036 -12949 -5024
rect -13015 -5142 -12999 -5036
rect -12965 -5142 -12949 -5036
rect -13015 -5154 -12949 -5142
rect -12919 -5036 -12857 -5024
rect -12919 -5142 -12903 -5036
rect -12869 -5142 -12857 -5036
rect -12919 -5154 -12857 -5142
rect -12827 -5036 -12769 -5024
rect -12827 -5142 -12815 -5036
rect -12781 -5142 -12769 -5036
rect -12827 -5154 -12769 -5142
rect -12596 -5036 -12538 -5024
rect -12596 -5142 -12584 -5036
rect -12550 -5142 -12538 -5036
rect -12596 -5154 -12538 -5142
rect -12508 -5036 -12446 -5024
rect -12508 -5142 -12496 -5036
rect -12462 -5142 -12446 -5036
rect -12508 -5154 -12446 -5142
rect -12416 -5036 -12350 -5024
rect -12416 -5142 -12400 -5036
rect -12366 -5142 -12350 -5036
rect -12416 -5154 -12350 -5142
rect -12320 -5036 -12254 -5024
rect -12320 -5142 -12304 -5036
rect -12270 -5142 -12254 -5036
rect -12320 -5154 -12254 -5142
rect -12224 -5036 -12158 -5024
rect -12224 -5142 -12208 -5036
rect -12174 -5142 -12158 -5036
rect -12224 -5154 -12158 -5142
rect -12128 -5036 -12062 -5024
rect -12128 -5142 -12112 -5036
rect -12078 -5142 -12062 -5036
rect -12128 -5154 -12062 -5142
rect -12032 -5036 -11966 -5024
rect -12032 -5142 -12016 -5036
rect -11982 -5142 -11966 -5036
rect -12032 -5154 -11966 -5142
rect -11936 -5036 -11870 -5024
rect -11936 -5142 -11920 -5036
rect -11886 -5142 -11870 -5036
rect -11936 -5154 -11870 -5142
rect -11840 -5036 -11774 -5024
rect -11840 -5142 -11824 -5036
rect -11790 -5142 -11774 -5036
rect -11840 -5154 -11774 -5142
rect -11744 -5036 -11678 -5024
rect -11744 -5142 -11728 -5036
rect -11694 -5142 -11678 -5036
rect -11744 -5154 -11678 -5142
rect -11648 -5036 -11582 -5024
rect -11648 -5142 -11632 -5036
rect -11598 -5142 -11582 -5036
rect -11648 -5154 -11582 -5142
rect -11552 -5036 -11486 -5024
rect -11552 -5142 -11536 -5036
rect -11502 -5142 -11486 -5036
rect -11552 -5154 -11486 -5142
rect -11456 -5036 -11390 -5024
rect -11456 -5142 -11440 -5036
rect -11406 -5142 -11390 -5036
rect -11456 -5154 -11390 -5142
rect -11360 -5036 -11298 -5024
rect -11360 -5142 -11344 -5036
rect -11310 -5142 -11298 -5036
rect -11360 -5154 -11298 -5142
rect -11268 -5036 -11210 -5024
rect -11268 -5142 -11256 -5036
rect -11222 -5142 -11210 -5036
rect -11268 -5154 -11210 -5142
rect -10864 -5036 -10806 -5024
rect -10864 -5142 -10852 -5036
rect -10818 -5142 -10806 -5036
rect -10864 -5154 -10806 -5142
rect -10776 -5036 -10714 -5024
rect -10776 -5142 -10764 -5036
rect -10730 -5142 -10714 -5036
rect -10776 -5154 -10714 -5142
rect -10684 -5036 -10618 -5024
rect -10684 -5142 -10668 -5036
rect -10634 -5142 -10618 -5036
rect -10684 -5154 -10618 -5142
rect -10588 -5036 -10522 -5024
rect -10588 -5142 -10572 -5036
rect -10538 -5142 -10522 -5036
rect -10588 -5154 -10522 -5142
rect -10492 -5036 -10426 -5024
rect -10492 -5142 -10476 -5036
rect -10442 -5142 -10426 -5036
rect -10492 -5154 -10426 -5142
rect -10396 -5036 -10330 -5024
rect -10396 -5142 -10380 -5036
rect -10346 -5142 -10330 -5036
rect -10396 -5154 -10330 -5142
rect -10300 -5036 -10234 -5024
rect -10300 -5142 -10284 -5036
rect -10250 -5142 -10234 -5036
rect -10300 -5154 -10234 -5142
rect -10204 -5036 -10138 -5024
rect -10204 -5142 -10188 -5036
rect -10154 -5142 -10138 -5036
rect -10204 -5154 -10138 -5142
rect -10108 -5036 -10042 -5024
rect -10108 -5142 -10092 -5036
rect -10058 -5142 -10042 -5036
rect -10108 -5154 -10042 -5142
rect -10012 -5036 -9946 -5024
rect -10012 -5142 -9996 -5036
rect -9962 -5142 -9946 -5036
rect -10012 -5154 -9946 -5142
rect -9916 -5036 -9850 -5024
rect -9916 -5142 -9900 -5036
rect -9866 -5142 -9850 -5036
rect -9916 -5154 -9850 -5142
rect -9820 -5036 -9754 -5024
rect -9820 -5142 -9804 -5036
rect -9770 -5142 -9754 -5036
rect -9820 -5154 -9754 -5142
rect -9724 -5036 -9658 -5024
rect -9724 -5142 -9708 -5036
rect -9674 -5142 -9658 -5036
rect -9724 -5154 -9658 -5142
rect -9628 -5036 -9566 -5024
rect -9628 -5142 -9612 -5036
rect -9578 -5142 -9566 -5036
rect -9628 -5154 -9566 -5142
rect -9536 -5036 -9478 -5024
rect -9536 -5142 -9524 -5036
rect -9490 -5142 -9478 -5036
rect -9536 -5154 -9478 -5142
rect -9305 -5036 -9247 -5024
rect -9305 -5142 -9293 -5036
rect -9259 -5142 -9247 -5036
rect -9305 -5154 -9247 -5142
rect -9217 -5036 -9155 -5024
rect -9217 -5142 -9205 -5036
rect -9171 -5142 -9155 -5036
rect -9217 -5154 -9155 -5142
rect -9125 -5036 -9059 -5024
rect -9125 -5142 -9109 -5036
rect -9075 -5142 -9059 -5036
rect -9125 -5154 -9059 -5142
rect -9029 -5036 -8963 -5024
rect -9029 -5142 -9013 -5036
rect -8979 -5142 -8963 -5036
rect -9029 -5154 -8963 -5142
rect -8933 -5036 -8867 -5024
rect -8933 -5142 -8917 -5036
rect -8883 -5142 -8867 -5036
rect -8933 -5154 -8867 -5142
rect -8837 -5036 -8771 -5024
rect -8837 -5142 -8821 -5036
rect -8787 -5142 -8771 -5036
rect -8837 -5154 -8771 -5142
rect -8741 -5036 -8675 -5024
rect -8741 -5142 -8725 -5036
rect -8691 -5142 -8675 -5036
rect -8741 -5154 -8675 -5142
rect -8645 -5036 -8579 -5024
rect -8645 -5142 -8629 -5036
rect -8595 -5142 -8579 -5036
rect -8645 -5154 -8579 -5142
rect -8549 -5036 -8483 -5024
rect -8549 -5142 -8533 -5036
rect -8499 -5142 -8483 -5036
rect -8549 -5154 -8483 -5142
rect -8453 -5036 -8387 -5024
rect -8453 -5142 -8437 -5036
rect -8403 -5142 -8387 -5036
rect -8453 -5154 -8387 -5142
rect -8357 -5036 -8291 -5024
rect -8357 -5142 -8341 -5036
rect -8307 -5142 -8291 -5036
rect -8357 -5154 -8291 -5142
rect -8261 -5036 -8195 -5024
rect -8261 -5142 -8245 -5036
rect -8211 -5142 -8195 -5036
rect -8261 -5154 -8195 -5142
rect -8165 -5036 -8099 -5024
rect -8165 -5142 -8149 -5036
rect -8115 -5142 -8099 -5036
rect -8165 -5154 -8099 -5142
rect -8069 -5036 -8007 -5024
rect -8069 -5142 -8053 -5036
rect -8019 -5142 -8007 -5036
rect -8069 -5154 -8007 -5142
rect -7977 -5036 -7919 -5024
rect -7977 -5142 -7965 -5036
rect -7931 -5142 -7919 -5036
rect -7977 -5154 -7919 -5142
rect 5658 -5495 5858 -5483
rect 5658 -5529 5670 -5495
rect 5846 -5529 5858 -5495
rect 6098 -5495 6298 -5483
rect 5658 -5541 5858 -5529
rect 5658 -5583 5858 -5571
rect 5658 -5617 5670 -5583
rect 5846 -5617 5858 -5583
rect 6098 -5529 6110 -5495
rect 6286 -5529 6298 -5495
rect 6538 -5495 6738 -5483
rect 6098 -5541 6298 -5529
rect 6098 -5583 6298 -5571
rect 5658 -5629 5858 -5617
rect 6098 -5617 6110 -5583
rect 6286 -5617 6298 -5583
rect 6538 -5529 6550 -5495
rect 6726 -5529 6738 -5495
rect 6538 -5541 6738 -5529
rect 6538 -5583 6738 -5571
rect 6098 -5629 6298 -5617
rect 6538 -5617 6550 -5583
rect 6726 -5617 6738 -5583
rect 6538 -5629 6738 -5617
rect -24162 -5873 -23762 -5861
rect -24162 -5907 -24150 -5873
rect -23774 -5907 -23762 -5873
rect -23586 -5873 -23386 -5861
rect -24162 -5923 -23762 -5907
rect -23586 -5907 -23574 -5873
rect -23398 -5907 -23386 -5873
rect -23586 -5919 -23386 -5907
rect -24162 -6019 -23762 -5953
rect -23586 -5961 -23386 -5949
rect -23586 -5995 -23574 -5961
rect -23398 -5995 -23386 -5961
rect -23586 -6007 -23386 -5995
rect -22426 -5873 -22026 -5861
rect -22426 -5907 -22414 -5873
rect -22038 -5907 -22026 -5873
rect -21852 -5873 -21652 -5861
rect -22426 -5923 -22026 -5907
rect -21852 -5907 -21840 -5873
rect -21664 -5907 -21652 -5873
rect -21852 -5919 -21652 -5907
rect -22426 -6019 -22026 -5953
rect -21852 -5961 -21652 -5949
rect -21852 -5995 -21840 -5961
rect -21664 -5995 -21652 -5961
rect -21852 -6007 -21652 -5995
rect -24162 -6065 -23762 -6049
rect -24162 -6099 -24150 -6065
rect -23774 -6099 -23762 -6065
rect -24162 -6111 -23762 -6099
rect -22426 -6065 -22026 -6049
rect -22426 -6099 -22414 -6065
rect -22038 -6099 -22026 -6065
rect -22426 -6111 -22026 -6099
rect -20296 -6041 -19896 -6029
rect -20296 -6075 -20284 -6041
rect -19908 -6075 -19896 -6041
rect -20296 -6091 -19896 -6075
rect -20296 -6187 -19896 -6121
rect -19187 -6041 -18787 -6029
rect -19187 -6075 -19175 -6041
rect -18799 -6075 -18787 -6041
rect -19187 -6091 -18787 -6075
rect -19187 -6187 -18787 -6121
rect -18305 -6041 -17905 -6029
rect -18305 -6075 -18293 -6041
rect -17917 -6075 -17905 -6041
rect -18305 -6091 -17905 -6075
rect -18305 -6187 -17905 -6121
rect -17005 -6041 -16605 -6029
rect -17005 -6075 -16993 -6041
rect -16617 -6075 -16605 -6041
rect -17005 -6091 -16605 -6075
rect -17005 -6187 -16605 -6121
rect -15896 -6041 -15496 -6029
rect -15896 -6075 -15884 -6041
rect -15508 -6075 -15496 -6041
rect -15896 -6091 -15496 -6075
rect -15896 -6187 -15496 -6121
rect -15014 -6041 -14614 -6029
rect -15014 -6075 -15002 -6041
rect -14626 -6075 -14614 -6041
rect -15014 -6091 -14614 -6075
rect -15014 -6187 -14614 -6121
rect -13714 -6041 -13314 -6029
rect -13714 -6075 -13702 -6041
rect -13326 -6075 -13314 -6041
rect -13714 -6091 -13314 -6075
rect -13714 -6187 -13314 -6121
rect -12605 -6041 -12205 -6029
rect -12605 -6075 -12593 -6041
rect -12217 -6075 -12205 -6041
rect -12605 -6091 -12205 -6075
rect -12605 -6187 -12205 -6121
rect -11723 -6041 -11323 -6029
rect -11723 -6075 -11711 -6041
rect -11335 -6075 -11323 -6041
rect -11723 -6091 -11323 -6075
rect -11723 -6187 -11323 -6121
rect -10423 -6041 -10023 -6029
rect -10423 -6075 -10411 -6041
rect -10035 -6075 -10023 -6041
rect -10423 -6091 -10023 -6075
rect -10423 -6187 -10023 -6121
rect -9314 -6041 -8914 -6029
rect -9314 -6075 -9302 -6041
rect -8926 -6075 -8914 -6041
rect -9314 -6091 -8914 -6075
rect -9314 -6187 -8914 -6121
rect -8432 -6041 -8032 -6029
rect -8432 -6075 -8420 -6041
rect -8044 -6075 -8032 -6041
rect -8432 -6091 -8032 -6075
rect -8432 -6187 -8032 -6121
rect -20296 -6233 -19896 -6217
rect -20296 -6267 -20284 -6233
rect -19908 -6267 -19896 -6233
rect -19187 -6233 -18787 -6217
rect -20296 -6279 -19896 -6267
rect -19187 -6267 -19175 -6233
rect -18799 -6267 -18787 -6233
rect -18305 -6233 -17905 -6217
rect -19187 -6279 -18787 -6267
rect -18305 -6267 -18293 -6233
rect -17917 -6267 -17905 -6233
rect -17005 -6233 -16605 -6217
rect -18305 -6279 -17905 -6267
rect -17005 -6267 -16993 -6233
rect -16617 -6267 -16605 -6233
rect -15896 -6233 -15496 -6217
rect -17005 -6279 -16605 -6267
rect -15896 -6267 -15884 -6233
rect -15508 -6267 -15496 -6233
rect -15014 -6233 -14614 -6217
rect -15896 -6279 -15496 -6267
rect -15014 -6267 -15002 -6233
rect -14626 -6267 -14614 -6233
rect -13714 -6233 -13314 -6217
rect -15014 -6279 -14614 -6267
rect -13714 -6267 -13702 -6233
rect -13326 -6267 -13314 -6233
rect -12605 -6233 -12205 -6217
rect -13714 -6279 -13314 -6267
rect -12605 -6267 -12593 -6233
rect -12217 -6267 -12205 -6233
rect -11723 -6233 -11323 -6217
rect -12605 -6279 -12205 -6267
rect -11723 -6267 -11711 -6233
rect -11335 -6267 -11323 -6233
rect -10423 -6233 -10023 -6217
rect -11723 -6279 -11323 -6267
rect -10423 -6267 -10411 -6233
rect -10035 -6267 -10023 -6233
rect -9314 -6233 -8914 -6217
rect -10423 -6279 -10023 -6267
rect -9314 -6267 -9302 -6233
rect -8926 -6267 -8914 -6233
rect -8432 -6233 -8032 -6217
rect -9314 -6279 -8914 -6267
rect -8432 -6267 -8420 -6233
rect -8044 -6267 -8032 -6233
rect -8432 -6279 -8032 -6267
rect 7360 -6478 7422 -6466
rect -24162 -7846 -23762 -7834
rect -24162 -7880 -24150 -7846
rect -23774 -7880 -23762 -7846
rect -23584 -7846 -23384 -7834
rect -24162 -7896 -23762 -7880
rect -23584 -7880 -23572 -7846
rect -23396 -7880 -23384 -7846
rect -23584 -7892 -23384 -7880
rect -24162 -7992 -23762 -7926
rect -23584 -7934 -23384 -7922
rect -23584 -7968 -23572 -7934
rect -23396 -7968 -23384 -7934
rect -23584 -7980 -23384 -7968
rect 7360 -7254 7372 -6478
rect 7406 -7254 7422 -6478
rect 7360 -7266 7422 -7254
rect 7452 -7266 7518 -6466
rect 7548 -7266 7614 -6466
rect 7644 -7266 7710 -6466
rect 7740 -6478 7802 -6466
rect 7740 -7254 7756 -6478
rect 7790 -7254 7802 -6478
rect 7740 -7266 7802 -7254
rect 8308 -6478 8370 -6466
rect 8308 -7254 8320 -6478
rect 8354 -7254 8370 -6478
rect 8308 -7266 8370 -7254
rect 8400 -7266 8466 -6466
rect 8496 -7266 8562 -6466
rect 8592 -7266 8658 -6466
rect 8688 -6478 8750 -6466
rect 8688 -7254 8704 -6478
rect 8738 -7254 8750 -6478
rect 8688 -7266 8750 -7254
rect 9244 -6478 9306 -6466
rect 9244 -7254 9256 -6478
rect 9290 -7254 9306 -6478
rect 9244 -7266 9306 -7254
rect 9336 -7266 9402 -6466
rect 9432 -7266 9498 -6466
rect 9528 -7266 9594 -6466
rect 9624 -6478 9686 -6466
rect 9624 -7254 9640 -6478
rect 9674 -7254 9686 -6478
rect 9624 -7266 9686 -7254
rect 10175 -6478 10237 -6466
rect 10175 -7254 10187 -6478
rect 10221 -7254 10237 -6478
rect 10175 -7266 10237 -7254
rect 10267 -7266 10333 -6466
rect 10363 -7266 10429 -6466
rect 10459 -7266 10525 -6466
rect 10555 -6478 10617 -6466
rect 10555 -7254 10571 -6478
rect 10605 -7254 10617 -6478
rect 10555 -7266 10617 -7254
rect 11102 -6478 11164 -6466
rect 11102 -7254 11114 -6478
rect 11148 -7254 11164 -6478
rect 11102 -7266 11164 -7254
rect 11194 -7266 11260 -6466
rect 11290 -7266 11356 -6466
rect 11386 -7266 11452 -6466
rect 11482 -6478 11544 -6466
rect 11482 -7254 11498 -6478
rect 11532 -7254 11544 -6478
rect 11482 -7266 11544 -7254
rect 7360 -7406 7422 -7394
rect -22425 -7846 -22025 -7834
rect -22425 -7880 -22413 -7846
rect -22037 -7880 -22025 -7846
rect -21850 -7846 -21650 -7834
rect -22425 -7896 -22025 -7880
rect -21850 -7880 -21838 -7846
rect -21662 -7880 -21650 -7846
rect -21850 -7892 -21650 -7880
rect -22425 -7992 -22025 -7926
rect -21850 -7934 -21650 -7922
rect -21850 -7968 -21838 -7934
rect -21662 -7968 -21650 -7934
rect -21850 -7980 -21650 -7968
rect -24162 -8038 -23762 -8022
rect -24162 -8072 -24150 -8038
rect -23774 -8072 -23762 -8038
rect -24162 -8084 -23762 -8072
rect -22425 -8038 -22025 -8022
rect -22425 -8072 -22413 -8038
rect -22037 -8072 -22025 -8038
rect -22425 -8084 -22025 -8072
rect 7360 -8182 7372 -7406
rect 7406 -8182 7422 -7406
rect 7360 -8194 7422 -8182
rect 7452 -8194 7518 -7394
rect 7548 -8194 7614 -7394
rect 7644 -8194 7710 -7394
rect 7740 -7406 7802 -7394
rect 7740 -8182 7756 -7406
rect 7790 -8182 7802 -7406
rect 7740 -8194 7802 -8182
rect 8308 -7406 8370 -7394
rect 8308 -8182 8320 -7406
rect 8354 -8182 8370 -7406
rect 8308 -8194 8370 -8182
rect 8400 -8194 8466 -7394
rect 8496 -8194 8562 -7394
rect 8592 -8194 8658 -7394
rect 8688 -7406 8750 -7394
rect 8688 -8182 8704 -7406
rect 8738 -8182 8750 -7406
rect 8688 -8194 8750 -8182
rect 9244 -7406 9306 -7394
rect 9244 -8182 9256 -7406
rect 9290 -8182 9306 -7406
rect 9244 -8194 9306 -8182
rect 9336 -8194 9402 -7394
rect 9432 -8194 9498 -7394
rect 9528 -8194 9594 -7394
rect 9624 -7406 9686 -7394
rect 9624 -8182 9640 -7406
rect 9674 -8182 9686 -7406
rect 9624 -8194 9686 -8182
rect 10175 -7405 10237 -7393
rect 10175 -8181 10187 -7405
rect 10221 -8181 10237 -7405
rect 10175 -8193 10237 -8181
rect 10267 -8193 10333 -7393
rect 10363 -8193 10429 -7393
rect 10459 -8193 10525 -7393
rect 10555 -7405 10617 -7393
rect 10555 -8181 10571 -7405
rect 10605 -8181 10617 -7405
rect 10555 -8193 10617 -8181
rect 11102 -7406 11164 -7394
rect -20737 -8301 -20679 -8289
rect -20737 -8407 -20725 -8301
rect -20691 -8407 -20679 -8301
rect -20737 -8419 -20679 -8407
rect -20649 -8301 -20587 -8289
rect -20649 -8407 -20637 -8301
rect -20603 -8407 -20587 -8301
rect -20649 -8419 -20587 -8407
rect -20557 -8301 -20491 -8289
rect -20557 -8407 -20541 -8301
rect -20507 -8407 -20491 -8301
rect -20557 -8419 -20491 -8407
rect -20461 -8301 -20395 -8289
rect -20461 -8407 -20445 -8301
rect -20411 -8407 -20395 -8301
rect -20461 -8419 -20395 -8407
rect -20365 -8301 -20299 -8289
rect -20365 -8407 -20349 -8301
rect -20315 -8407 -20299 -8301
rect -20365 -8419 -20299 -8407
rect -20269 -8301 -20203 -8289
rect -20269 -8407 -20253 -8301
rect -20219 -8407 -20203 -8301
rect -20269 -8419 -20203 -8407
rect -20173 -8301 -20107 -8289
rect -20173 -8407 -20157 -8301
rect -20123 -8407 -20107 -8301
rect -20173 -8419 -20107 -8407
rect -20077 -8301 -20011 -8289
rect -20077 -8407 -20061 -8301
rect -20027 -8407 -20011 -8301
rect -20077 -8419 -20011 -8407
rect -19981 -8301 -19915 -8289
rect -19981 -8407 -19965 -8301
rect -19931 -8407 -19915 -8301
rect -19981 -8419 -19915 -8407
rect -19885 -8301 -19819 -8289
rect -19885 -8407 -19869 -8301
rect -19835 -8407 -19819 -8301
rect -19885 -8419 -19819 -8407
rect -19789 -8301 -19723 -8289
rect -19789 -8407 -19773 -8301
rect -19739 -8407 -19723 -8301
rect -19789 -8419 -19723 -8407
rect -19693 -8301 -19627 -8289
rect -19693 -8407 -19677 -8301
rect -19643 -8407 -19627 -8301
rect -19693 -8419 -19627 -8407
rect -19597 -8301 -19531 -8289
rect -19597 -8407 -19581 -8301
rect -19547 -8407 -19531 -8301
rect -19597 -8419 -19531 -8407
rect -19501 -8301 -19439 -8289
rect -19501 -8407 -19485 -8301
rect -19451 -8407 -19439 -8301
rect -19501 -8419 -19439 -8407
rect -19409 -8301 -19351 -8289
rect -19409 -8407 -19397 -8301
rect -19363 -8407 -19351 -8301
rect -19409 -8419 -19351 -8407
rect -19178 -8301 -19120 -8289
rect -19178 -8407 -19166 -8301
rect -19132 -8407 -19120 -8301
rect -19178 -8419 -19120 -8407
rect -19090 -8301 -19028 -8289
rect -19090 -8407 -19078 -8301
rect -19044 -8407 -19028 -8301
rect -19090 -8419 -19028 -8407
rect -18998 -8301 -18932 -8289
rect -18998 -8407 -18982 -8301
rect -18948 -8407 -18932 -8301
rect -18998 -8419 -18932 -8407
rect -18902 -8301 -18836 -8289
rect -18902 -8407 -18886 -8301
rect -18852 -8407 -18836 -8301
rect -18902 -8419 -18836 -8407
rect -18806 -8301 -18740 -8289
rect -18806 -8407 -18790 -8301
rect -18756 -8407 -18740 -8301
rect -18806 -8419 -18740 -8407
rect -18710 -8301 -18644 -8289
rect -18710 -8407 -18694 -8301
rect -18660 -8407 -18644 -8301
rect -18710 -8419 -18644 -8407
rect -18614 -8301 -18548 -8289
rect -18614 -8407 -18598 -8301
rect -18564 -8407 -18548 -8301
rect -18614 -8419 -18548 -8407
rect -18518 -8301 -18452 -8289
rect -18518 -8407 -18502 -8301
rect -18468 -8407 -18452 -8301
rect -18518 -8419 -18452 -8407
rect -18422 -8301 -18356 -8289
rect -18422 -8407 -18406 -8301
rect -18372 -8407 -18356 -8301
rect -18422 -8419 -18356 -8407
rect -18326 -8301 -18260 -8289
rect -18326 -8407 -18310 -8301
rect -18276 -8407 -18260 -8301
rect -18326 -8419 -18260 -8407
rect -18230 -8301 -18164 -8289
rect -18230 -8407 -18214 -8301
rect -18180 -8407 -18164 -8301
rect -18230 -8419 -18164 -8407
rect -18134 -8301 -18068 -8289
rect -18134 -8407 -18118 -8301
rect -18084 -8407 -18068 -8301
rect -18134 -8419 -18068 -8407
rect -18038 -8301 -17972 -8289
rect -18038 -8407 -18022 -8301
rect -17988 -8407 -17972 -8301
rect -18038 -8419 -17972 -8407
rect -17942 -8301 -17880 -8289
rect -17942 -8407 -17926 -8301
rect -17892 -8407 -17880 -8301
rect -17942 -8419 -17880 -8407
rect -17850 -8301 -17792 -8289
rect -17850 -8407 -17838 -8301
rect -17804 -8407 -17792 -8301
rect -17850 -8419 -17792 -8407
rect -17446 -8301 -17388 -8289
rect -17446 -8407 -17434 -8301
rect -17400 -8407 -17388 -8301
rect -17446 -8419 -17388 -8407
rect -17358 -8301 -17296 -8289
rect -17358 -8407 -17346 -8301
rect -17312 -8407 -17296 -8301
rect -17358 -8419 -17296 -8407
rect -17266 -8301 -17200 -8289
rect -17266 -8407 -17250 -8301
rect -17216 -8407 -17200 -8301
rect -17266 -8419 -17200 -8407
rect -17170 -8301 -17104 -8289
rect -17170 -8407 -17154 -8301
rect -17120 -8407 -17104 -8301
rect -17170 -8419 -17104 -8407
rect -17074 -8301 -17008 -8289
rect -17074 -8407 -17058 -8301
rect -17024 -8407 -17008 -8301
rect -17074 -8419 -17008 -8407
rect -16978 -8301 -16912 -8289
rect -16978 -8407 -16962 -8301
rect -16928 -8407 -16912 -8301
rect -16978 -8419 -16912 -8407
rect -16882 -8301 -16816 -8289
rect -16882 -8407 -16866 -8301
rect -16832 -8407 -16816 -8301
rect -16882 -8419 -16816 -8407
rect -16786 -8301 -16720 -8289
rect -16786 -8407 -16770 -8301
rect -16736 -8407 -16720 -8301
rect -16786 -8419 -16720 -8407
rect -16690 -8301 -16624 -8289
rect -16690 -8407 -16674 -8301
rect -16640 -8407 -16624 -8301
rect -16690 -8419 -16624 -8407
rect -16594 -8301 -16528 -8289
rect -16594 -8407 -16578 -8301
rect -16544 -8407 -16528 -8301
rect -16594 -8419 -16528 -8407
rect -16498 -8301 -16432 -8289
rect -16498 -8407 -16482 -8301
rect -16448 -8407 -16432 -8301
rect -16498 -8419 -16432 -8407
rect -16402 -8301 -16336 -8289
rect -16402 -8407 -16386 -8301
rect -16352 -8407 -16336 -8301
rect -16402 -8419 -16336 -8407
rect -16306 -8301 -16240 -8289
rect -16306 -8407 -16290 -8301
rect -16256 -8407 -16240 -8301
rect -16306 -8419 -16240 -8407
rect -16210 -8301 -16148 -8289
rect -16210 -8407 -16194 -8301
rect -16160 -8407 -16148 -8301
rect -16210 -8419 -16148 -8407
rect -16118 -8301 -16060 -8289
rect -16118 -8407 -16106 -8301
rect -16072 -8407 -16060 -8301
rect -16118 -8419 -16060 -8407
rect -15887 -8301 -15829 -8289
rect -15887 -8407 -15875 -8301
rect -15841 -8407 -15829 -8301
rect -15887 -8419 -15829 -8407
rect -15799 -8301 -15737 -8289
rect -15799 -8407 -15787 -8301
rect -15753 -8407 -15737 -8301
rect -15799 -8419 -15737 -8407
rect -15707 -8301 -15641 -8289
rect -15707 -8407 -15691 -8301
rect -15657 -8407 -15641 -8301
rect -15707 -8419 -15641 -8407
rect -15611 -8301 -15545 -8289
rect -15611 -8407 -15595 -8301
rect -15561 -8407 -15545 -8301
rect -15611 -8419 -15545 -8407
rect -15515 -8301 -15449 -8289
rect -15515 -8407 -15499 -8301
rect -15465 -8407 -15449 -8301
rect -15515 -8419 -15449 -8407
rect -15419 -8301 -15353 -8289
rect -15419 -8407 -15403 -8301
rect -15369 -8407 -15353 -8301
rect -15419 -8419 -15353 -8407
rect -15323 -8301 -15257 -8289
rect -15323 -8407 -15307 -8301
rect -15273 -8407 -15257 -8301
rect -15323 -8419 -15257 -8407
rect -15227 -8301 -15161 -8289
rect -15227 -8407 -15211 -8301
rect -15177 -8407 -15161 -8301
rect -15227 -8419 -15161 -8407
rect -15131 -8301 -15065 -8289
rect -15131 -8407 -15115 -8301
rect -15081 -8407 -15065 -8301
rect -15131 -8419 -15065 -8407
rect -15035 -8301 -14969 -8289
rect -15035 -8407 -15019 -8301
rect -14985 -8407 -14969 -8301
rect -15035 -8419 -14969 -8407
rect -14939 -8301 -14873 -8289
rect -14939 -8407 -14923 -8301
rect -14889 -8407 -14873 -8301
rect -14939 -8419 -14873 -8407
rect -14843 -8301 -14777 -8289
rect -14843 -8407 -14827 -8301
rect -14793 -8407 -14777 -8301
rect -14843 -8419 -14777 -8407
rect -14747 -8301 -14681 -8289
rect -14747 -8407 -14731 -8301
rect -14697 -8407 -14681 -8301
rect -14747 -8419 -14681 -8407
rect -14651 -8301 -14589 -8289
rect -14651 -8407 -14635 -8301
rect -14601 -8407 -14589 -8301
rect -14651 -8419 -14589 -8407
rect -14559 -8301 -14501 -8289
rect -14559 -8407 -14547 -8301
rect -14513 -8407 -14501 -8301
rect -14559 -8419 -14501 -8407
rect -14155 -8301 -14097 -8289
rect -14155 -8407 -14143 -8301
rect -14109 -8407 -14097 -8301
rect -14155 -8419 -14097 -8407
rect -14067 -8301 -14005 -8289
rect -14067 -8407 -14055 -8301
rect -14021 -8407 -14005 -8301
rect -14067 -8419 -14005 -8407
rect -13975 -8301 -13909 -8289
rect -13975 -8407 -13959 -8301
rect -13925 -8407 -13909 -8301
rect -13975 -8419 -13909 -8407
rect -13879 -8301 -13813 -8289
rect -13879 -8407 -13863 -8301
rect -13829 -8407 -13813 -8301
rect -13879 -8419 -13813 -8407
rect -13783 -8301 -13717 -8289
rect -13783 -8407 -13767 -8301
rect -13733 -8407 -13717 -8301
rect -13783 -8419 -13717 -8407
rect -13687 -8301 -13621 -8289
rect -13687 -8407 -13671 -8301
rect -13637 -8407 -13621 -8301
rect -13687 -8419 -13621 -8407
rect -13591 -8301 -13525 -8289
rect -13591 -8407 -13575 -8301
rect -13541 -8407 -13525 -8301
rect -13591 -8419 -13525 -8407
rect -13495 -8301 -13429 -8289
rect -13495 -8407 -13479 -8301
rect -13445 -8407 -13429 -8301
rect -13495 -8419 -13429 -8407
rect -13399 -8301 -13333 -8289
rect -13399 -8407 -13383 -8301
rect -13349 -8407 -13333 -8301
rect -13399 -8419 -13333 -8407
rect -13303 -8301 -13237 -8289
rect -13303 -8407 -13287 -8301
rect -13253 -8407 -13237 -8301
rect -13303 -8419 -13237 -8407
rect -13207 -8301 -13141 -8289
rect -13207 -8407 -13191 -8301
rect -13157 -8407 -13141 -8301
rect -13207 -8419 -13141 -8407
rect -13111 -8301 -13045 -8289
rect -13111 -8407 -13095 -8301
rect -13061 -8407 -13045 -8301
rect -13111 -8419 -13045 -8407
rect -13015 -8301 -12949 -8289
rect -13015 -8407 -12999 -8301
rect -12965 -8407 -12949 -8301
rect -13015 -8419 -12949 -8407
rect -12919 -8301 -12857 -8289
rect -12919 -8407 -12903 -8301
rect -12869 -8407 -12857 -8301
rect -12919 -8419 -12857 -8407
rect -12827 -8301 -12769 -8289
rect -12827 -8407 -12815 -8301
rect -12781 -8407 -12769 -8301
rect -12827 -8419 -12769 -8407
rect -12596 -8301 -12538 -8289
rect -12596 -8407 -12584 -8301
rect -12550 -8407 -12538 -8301
rect -12596 -8419 -12538 -8407
rect -12508 -8301 -12446 -8289
rect -12508 -8407 -12496 -8301
rect -12462 -8407 -12446 -8301
rect -12508 -8419 -12446 -8407
rect -12416 -8301 -12350 -8289
rect -12416 -8407 -12400 -8301
rect -12366 -8407 -12350 -8301
rect -12416 -8419 -12350 -8407
rect -12320 -8301 -12254 -8289
rect -12320 -8407 -12304 -8301
rect -12270 -8407 -12254 -8301
rect -12320 -8419 -12254 -8407
rect -12224 -8301 -12158 -8289
rect -12224 -8407 -12208 -8301
rect -12174 -8407 -12158 -8301
rect -12224 -8419 -12158 -8407
rect -12128 -8301 -12062 -8289
rect -12128 -8407 -12112 -8301
rect -12078 -8407 -12062 -8301
rect -12128 -8419 -12062 -8407
rect -12032 -8301 -11966 -8289
rect -12032 -8407 -12016 -8301
rect -11982 -8407 -11966 -8301
rect -12032 -8419 -11966 -8407
rect -11936 -8301 -11870 -8289
rect -11936 -8407 -11920 -8301
rect -11886 -8407 -11870 -8301
rect -11936 -8419 -11870 -8407
rect -11840 -8301 -11774 -8289
rect -11840 -8407 -11824 -8301
rect -11790 -8407 -11774 -8301
rect -11840 -8419 -11774 -8407
rect -11744 -8301 -11678 -8289
rect -11744 -8407 -11728 -8301
rect -11694 -8407 -11678 -8301
rect -11744 -8419 -11678 -8407
rect -11648 -8301 -11582 -8289
rect -11648 -8407 -11632 -8301
rect -11598 -8407 -11582 -8301
rect -11648 -8419 -11582 -8407
rect -11552 -8301 -11486 -8289
rect -11552 -8407 -11536 -8301
rect -11502 -8407 -11486 -8301
rect -11552 -8419 -11486 -8407
rect -11456 -8301 -11390 -8289
rect -11456 -8407 -11440 -8301
rect -11406 -8407 -11390 -8301
rect -11456 -8419 -11390 -8407
rect -11360 -8301 -11298 -8289
rect -11360 -8407 -11344 -8301
rect -11310 -8407 -11298 -8301
rect -11360 -8419 -11298 -8407
rect -11268 -8301 -11210 -8289
rect -11268 -8407 -11256 -8301
rect -11222 -8407 -11210 -8301
rect -11268 -8419 -11210 -8407
rect -10864 -8301 -10806 -8289
rect -10864 -8407 -10852 -8301
rect -10818 -8407 -10806 -8301
rect -10864 -8419 -10806 -8407
rect -10776 -8301 -10714 -8289
rect -10776 -8407 -10764 -8301
rect -10730 -8407 -10714 -8301
rect -10776 -8419 -10714 -8407
rect -10684 -8301 -10618 -8289
rect -10684 -8407 -10668 -8301
rect -10634 -8407 -10618 -8301
rect -10684 -8419 -10618 -8407
rect -10588 -8301 -10522 -8289
rect -10588 -8407 -10572 -8301
rect -10538 -8407 -10522 -8301
rect -10588 -8419 -10522 -8407
rect -10492 -8301 -10426 -8289
rect -10492 -8407 -10476 -8301
rect -10442 -8407 -10426 -8301
rect -10492 -8419 -10426 -8407
rect -10396 -8301 -10330 -8289
rect -10396 -8407 -10380 -8301
rect -10346 -8407 -10330 -8301
rect -10396 -8419 -10330 -8407
rect -10300 -8301 -10234 -8289
rect -10300 -8407 -10284 -8301
rect -10250 -8407 -10234 -8301
rect -10300 -8419 -10234 -8407
rect -10204 -8301 -10138 -8289
rect -10204 -8407 -10188 -8301
rect -10154 -8407 -10138 -8301
rect -10204 -8419 -10138 -8407
rect -10108 -8301 -10042 -8289
rect -10108 -8407 -10092 -8301
rect -10058 -8407 -10042 -8301
rect -10108 -8419 -10042 -8407
rect -10012 -8301 -9946 -8289
rect -10012 -8407 -9996 -8301
rect -9962 -8407 -9946 -8301
rect -10012 -8419 -9946 -8407
rect -9916 -8301 -9850 -8289
rect -9916 -8407 -9900 -8301
rect -9866 -8407 -9850 -8301
rect -9916 -8419 -9850 -8407
rect -9820 -8301 -9754 -8289
rect -9820 -8407 -9804 -8301
rect -9770 -8407 -9754 -8301
rect -9820 -8419 -9754 -8407
rect -9724 -8301 -9658 -8289
rect -9724 -8407 -9708 -8301
rect -9674 -8407 -9658 -8301
rect -9724 -8419 -9658 -8407
rect -9628 -8301 -9566 -8289
rect -9628 -8407 -9612 -8301
rect -9578 -8407 -9566 -8301
rect -9628 -8419 -9566 -8407
rect -9536 -8301 -9478 -8289
rect -9536 -8407 -9524 -8301
rect -9490 -8407 -9478 -8301
rect -9536 -8419 -9478 -8407
rect -9305 -8301 -9247 -8289
rect -9305 -8407 -9293 -8301
rect -9259 -8407 -9247 -8301
rect -9305 -8419 -9247 -8407
rect -9217 -8301 -9155 -8289
rect -9217 -8407 -9205 -8301
rect -9171 -8407 -9155 -8301
rect -9217 -8419 -9155 -8407
rect -9125 -8301 -9059 -8289
rect -9125 -8407 -9109 -8301
rect -9075 -8407 -9059 -8301
rect -9125 -8419 -9059 -8407
rect -9029 -8301 -8963 -8289
rect -9029 -8407 -9013 -8301
rect -8979 -8407 -8963 -8301
rect -9029 -8419 -8963 -8407
rect -8933 -8301 -8867 -8289
rect -8933 -8407 -8917 -8301
rect -8883 -8407 -8867 -8301
rect -8933 -8419 -8867 -8407
rect -8837 -8301 -8771 -8289
rect -8837 -8407 -8821 -8301
rect -8787 -8407 -8771 -8301
rect -8837 -8419 -8771 -8407
rect -8741 -8301 -8675 -8289
rect -8741 -8407 -8725 -8301
rect -8691 -8407 -8675 -8301
rect -8741 -8419 -8675 -8407
rect -8645 -8301 -8579 -8289
rect -8645 -8407 -8629 -8301
rect -8595 -8407 -8579 -8301
rect -8645 -8419 -8579 -8407
rect -8549 -8301 -8483 -8289
rect -8549 -8407 -8533 -8301
rect -8499 -8407 -8483 -8301
rect -8549 -8419 -8483 -8407
rect -8453 -8301 -8387 -8289
rect -8453 -8407 -8437 -8301
rect -8403 -8407 -8387 -8301
rect -8453 -8419 -8387 -8407
rect -8357 -8301 -8291 -8289
rect -8357 -8407 -8341 -8301
rect -8307 -8407 -8291 -8301
rect -8357 -8419 -8291 -8407
rect -8261 -8301 -8195 -8289
rect -8261 -8407 -8245 -8301
rect -8211 -8407 -8195 -8301
rect -8261 -8419 -8195 -8407
rect -8165 -8301 -8099 -8289
rect -8165 -8407 -8149 -8301
rect -8115 -8407 -8099 -8301
rect -8165 -8419 -8099 -8407
rect -8069 -8301 -8007 -8289
rect -8069 -8407 -8053 -8301
rect -8019 -8407 -8007 -8301
rect -8069 -8419 -8007 -8407
rect -7977 -8301 -7919 -8289
rect -7977 -8407 -7965 -8301
rect -7931 -8407 -7919 -8301
rect -7977 -8419 -7919 -8407
rect 11102 -8182 11114 -7406
rect 11148 -8182 11164 -7406
rect 11102 -8194 11164 -8182
rect 11194 -8194 11260 -7394
rect 11290 -8194 11356 -7394
rect 11386 -8194 11452 -7394
rect 11482 -7406 11544 -7394
rect 11482 -8182 11498 -7406
rect 11532 -8182 11544 -7406
rect 12157 -7448 12219 -7436
rect 12157 -7624 12169 -7448
rect 12203 -7624 12219 -7448
rect 12157 -7636 12219 -7624
rect 12249 -7448 12315 -7436
rect 12249 -7624 12265 -7448
rect 12299 -7624 12315 -7448
rect 12249 -7636 12315 -7624
rect 12345 -7448 12407 -7436
rect 12345 -7624 12361 -7448
rect 12395 -7624 12407 -7448
rect 12923 -7513 13123 -7501
rect 12923 -7547 12935 -7513
rect 13111 -7547 13123 -7513
rect 12923 -7559 13123 -7547
rect 12923 -7601 13123 -7589
rect 12345 -7636 12407 -7624
rect 12923 -7635 12935 -7601
rect 13111 -7635 13123 -7601
rect 12923 -7647 13123 -7635
rect 11482 -8194 11544 -8182
rect -24162 -9138 -23762 -9126
rect -24162 -9172 -24150 -9138
rect -23774 -9172 -23762 -9138
rect -23583 -9138 -23383 -9126
rect -24162 -9188 -23762 -9172
rect -23583 -9172 -23571 -9138
rect -23395 -9172 -23383 -9138
rect -23583 -9184 -23383 -9172
rect -24162 -9284 -23762 -9218
rect -23583 -9226 -23383 -9214
rect -23583 -9260 -23571 -9226
rect -23395 -9260 -23383 -9226
rect -23583 -9272 -23383 -9260
rect -22426 -9138 -22026 -9126
rect -22426 -9172 -22414 -9138
rect -22038 -9172 -22026 -9138
rect -21846 -9138 -21646 -9126
rect -22426 -9188 -22026 -9172
rect -21846 -9172 -21834 -9138
rect -21658 -9172 -21646 -9138
rect -21846 -9184 -21646 -9172
rect -22426 -9284 -22026 -9218
rect -21846 -9226 -21646 -9214
rect -21846 -9260 -21834 -9226
rect -21658 -9260 -21646 -9226
rect -21846 -9272 -21646 -9260
rect -24162 -9330 -23762 -9314
rect -24162 -9364 -24150 -9330
rect -23774 -9364 -23762 -9330
rect -24162 -9376 -23762 -9364
rect -22426 -9330 -22026 -9314
rect -22426 -9364 -22414 -9330
rect -22038 -9364 -22026 -9330
rect -22426 -9376 -22026 -9364
rect -20296 -9306 -19896 -9294
rect -20296 -9340 -20284 -9306
rect -19908 -9340 -19896 -9306
rect -20296 -9356 -19896 -9340
rect -20296 -9452 -19896 -9386
rect -19187 -9306 -18787 -9294
rect -19187 -9340 -19175 -9306
rect -18799 -9340 -18787 -9306
rect -19187 -9356 -18787 -9340
rect -19187 -9452 -18787 -9386
rect -18305 -9306 -17905 -9294
rect -18305 -9340 -18293 -9306
rect -17917 -9340 -17905 -9306
rect -18305 -9356 -17905 -9340
rect -18305 -9452 -17905 -9386
rect -17005 -9306 -16605 -9294
rect -17005 -9340 -16993 -9306
rect -16617 -9340 -16605 -9306
rect -17005 -9356 -16605 -9340
rect -17005 -9452 -16605 -9386
rect -15896 -9306 -15496 -9294
rect -15896 -9340 -15884 -9306
rect -15508 -9340 -15496 -9306
rect -15896 -9356 -15496 -9340
rect -15896 -9452 -15496 -9386
rect -15014 -9306 -14614 -9294
rect -15014 -9340 -15002 -9306
rect -14626 -9340 -14614 -9306
rect -15014 -9356 -14614 -9340
rect -15014 -9452 -14614 -9386
rect -13714 -9306 -13314 -9294
rect -13714 -9340 -13702 -9306
rect -13326 -9340 -13314 -9306
rect -13714 -9356 -13314 -9340
rect -13714 -9452 -13314 -9386
rect -12605 -9306 -12205 -9294
rect -12605 -9340 -12593 -9306
rect -12217 -9340 -12205 -9306
rect -12605 -9356 -12205 -9340
rect -12605 -9452 -12205 -9386
rect -11723 -9306 -11323 -9294
rect -11723 -9340 -11711 -9306
rect -11335 -9340 -11323 -9306
rect -11723 -9356 -11323 -9340
rect -11723 -9452 -11323 -9386
rect -10423 -9306 -10023 -9294
rect -10423 -9340 -10411 -9306
rect -10035 -9340 -10023 -9306
rect -10423 -9356 -10023 -9340
rect -10423 -9452 -10023 -9386
rect -9314 -9306 -8914 -9294
rect -9314 -9340 -9302 -9306
rect -8926 -9340 -8914 -9306
rect -9314 -9356 -8914 -9340
rect -9314 -9452 -8914 -9386
rect -8432 -9306 -8032 -9294
rect -8432 -9340 -8420 -9306
rect -8044 -9340 -8032 -9306
rect -8432 -9356 -8032 -9340
rect -8432 -9452 -8032 -9386
rect -20296 -9498 -19896 -9482
rect -20296 -9532 -20284 -9498
rect -19908 -9532 -19896 -9498
rect -19187 -9498 -18787 -9482
rect -20296 -9544 -19896 -9532
rect -19187 -9532 -19175 -9498
rect -18799 -9532 -18787 -9498
rect -18305 -9498 -17905 -9482
rect -19187 -9544 -18787 -9532
rect -18305 -9532 -18293 -9498
rect -17917 -9532 -17905 -9498
rect -17005 -9498 -16605 -9482
rect -18305 -9544 -17905 -9532
rect -17005 -9532 -16993 -9498
rect -16617 -9532 -16605 -9498
rect -15896 -9498 -15496 -9482
rect -17005 -9544 -16605 -9532
rect -15896 -9532 -15884 -9498
rect -15508 -9532 -15496 -9498
rect -15014 -9498 -14614 -9482
rect -15896 -9544 -15496 -9532
rect -15014 -9532 -15002 -9498
rect -14626 -9532 -14614 -9498
rect -13714 -9498 -13314 -9482
rect -15014 -9544 -14614 -9532
rect -13714 -9532 -13702 -9498
rect -13326 -9532 -13314 -9498
rect -12605 -9498 -12205 -9482
rect -13714 -9544 -13314 -9532
rect -12605 -9532 -12593 -9498
rect -12217 -9532 -12205 -9498
rect -11723 -9498 -11323 -9482
rect -12605 -9544 -12205 -9532
rect -11723 -9532 -11711 -9498
rect -11335 -9532 -11323 -9498
rect -10423 -9498 -10023 -9482
rect -11723 -9544 -11323 -9532
rect -10423 -9532 -10411 -9498
rect -10035 -9532 -10023 -9498
rect -9314 -9498 -8914 -9482
rect -10423 -9544 -10023 -9532
rect -9314 -9532 -9302 -9498
rect -8926 -9532 -8914 -9498
rect -8432 -9498 -8032 -9482
rect -9314 -9544 -8914 -9532
rect -8432 -9532 -8420 -9498
rect -8044 -9532 -8032 -9498
rect -8432 -9544 -8032 -9532
rect 5658 -10123 5858 -10111
rect 5658 -10157 5670 -10123
rect 5846 -10157 5858 -10123
rect 6098 -10123 6298 -10111
rect 5658 -10169 5858 -10157
rect 5658 -10211 5858 -10199
rect 5658 -10245 5670 -10211
rect 5846 -10245 5858 -10211
rect 6098 -10157 6110 -10123
rect 6286 -10157 6298 -10123
rect 6538 -10123 6738 -10111
rect 6098 -10169 6298 -10157
rect 6098 -10211 6298 -10199
rect 5658 -10257 5858 -10245
rect 6098 -10245 6110 -10211
rect 6286 -10245 6298 -10211
rect 6538 -10157 6550 -10123
rect 6726 -10157 6738 -10123
rect 6538 -10169 6738 -10157
rect 6538 -10211 6738 -10199
rect 6098 -10257 6298 -10245
rect 6538 -10245 6550 -10211
rect 6726 -10245 6738 -10211
rect 6538 -10257 6738 -10245
rect -24162 -11110 -23762 -11098
rect -24162 -11144 -24150 -11110
rect -23774 -11144 -23762 -11110
rect -23583 -11110 -23383 -11098
rect -24162 -11160 -23762 -11144
rect -23583 -11144 -23571 -11110
rect -23395 -11144 -23383 -11110
rect -23583 -11156 -23383 -11144
rect -24162 -11256 -23762 -11190
rect -23583 -11198 -23383 -11186
rect -23583 -11232 -23571 -11198
rect -23395 -11232 -23383 -11198
rect -23583 -11244 -23383 -11232
rect -22425 -11110 -22025 -11098
rect -22425 -11144 -22413 -11110
rect -22037 -11144 -22025 -11110
rect -21850 -11110 -21650 -11098
rect -22425 -11160 -22025 -11144
rect -21850 -11144 -21838 -11110
rect -21662 -11144 -21650 -11110
rect -21850 -11156 -21650 -11144
rect -22425 -11256 -22025 -11190
rect -21850 -11198 -21650 -11186
rect -21850 -11232 -21838 -11198
rect -21662 -11232 -21650 -11198
rect -21850 -11244 -21650 -11232
rect -24162 -11302 -23762 -11286
rect -24162 -11336 -24150 -11302
rect -23774 -11336 -23762 -11302
rect -24162 -11348 -23762 -11336
rect -22425 -11302 -22025 -11286
rect -22425 -11336 -22413 -11302
rect -22037 -11336 -22025 -11302
rect -22425 -11348 -22025 -11336
rect 7360 -11106 7422 -11094
rect -20737 -11565 -20679 -11553
rect -20737 -11671 -20725 -11565
rect -20691 -11671 -20679 -11565
rect -20737 -11683 -20679 -11671
rect -20649 -11565 -20587 -11553
rect -20649 -11671 -20637 -11565
rect -20603 -11671 -20587 -11565
rect -20649 -11683 -20587 -11671
rect -20557 -11565 -20491 -11553
rect -20557 -11671 -20541 -11565
rect -20507 -11671 -20491 -11565
rect -20557 -11683 -20491 -11671
rect -20461 -11565 -20395 -11553
rect -20461 -11671 -20445 -11565
rect -20411 -11671 -20395 -11565
rect -20461 -11683 -20395 -11671
rect -20365 -11565 -20299 -11553
rect -20365 -11671 -20349 -11565
rect -20315 -11671 -20299 -11565
rect -20365 -11683 -20299 -11671
rect -20269 -11565 -20203 -11553
rect -20269 -11671 -20253 -11565
rect -20219 -11671 -20203 -11565
rect -20269 -11683 -20203 -11671
rect -20173 -11565 -20107 -11553
rect -20173 -11671 -20157 -11565
rect -20123 -11671 -20107 -11565
rect -20173 -11683 -20107 -11671
rect -20077 -11565 -20011 -11553
rect -20077 -11671 -20061 -11565
rect -20027 -11671 -20011 -11565
rect -20077 -11683 -20011 -11671
rect -19981 -11565 -19915 -11553
rect -19981 -11671 -19965 -11565
rect -19931 -11671 -19915 -11565
rect -19981 -11683 -19915 -11671
rect -19885 -11565 -19819 -11553
rect -19885 -11671 -19869 -11565
rect -19835 -11671 -19819 -11565
rect -19885 -11683 -19819 -11671
rect -19789 -11565 -19723 -11553
rect -19789 -11671 -19773 -11565
rect -19739 -11671 -19723 -11565
rect -19789 -11683 -19723 -11671
rect -19693 -11565 -19627 -11553
rect -19693 -11671 -19677 -11565
rect -19643 -11671 -19627 -11565
rect -19693 -11683 -19627 -11671
rect -19597 -11565 -19531 -11553
rect -19597 -11671 -19581 -11565
rect -19547 -11671 -19531 -11565
rect -19597 -11683 -19531 -11671
rect -19501 -11565 -19439 -11553
rect -19501 -11671 -19485 -11565
rect -19451 -11671 -19439 -11565
rect -19501 -11683 -19439 -11671
rect -19409 -11565 -19351 -11553
rect -19409 -11671 -19397 -11565
rect -19363 -11671 -19351 -11565
rect -19409 -11683 -19351 -11671
rect -19178 -11565 -19120 -11553
rect -19178 -11671 -19166 -11565
rect -19132 -11671 -19120 -11565
rect -19178 -11683 -19120 -11671
rect -19090 -11565 -19028 -11553
rect -19090 -11671 -19078 -11565
rect -19044 -11671 -19028 -11565
rect -19090 -11683 -19028 -11671
rect -18998 -11565 -18932 -11553
rect -18998 -11671 -18982 -11565
rect -18948 -11671 -18932 -11565
rect -18998 -11683 -18932 -11671
rect -18902 -11565 -18836 -11553
rect -18902 -11671 -18886 -11565
rect -18852 -11671 -18836 -11565
rect -18902 -11683 -18836 -11671
rect -18806 -11565 -18740 -11553
rect -18806 -11671 -18790 -11565
rect -18756 -11671 -18740 -11565
rect -18806 -11683 -18740 -11671
rect -18710 -11565 -18644 -11553
rect -18710 -11671 -18694 -11565
rect -18660 -11671 -18644 -11565
rect -18710 -11683 -18644 -11671
rect -18614 -11565 -18548 -11553
rect -18614 -11671 -18598 -11565
rect -18564 -11671 -18548 -11565
rect -18614 -11683 -18548 -11671
rect -18518 -11565 -18452 -11553
rect -18518 -11671 -18502 -11565
rect -18468 -11671 -18452 -11565
rect -18518 -11683 -18452 -11671
rect -18422 -11565 -18356 -11553
rect -18422 -11671 -18406 -11565
rect -18372 -11671 -18356 -11565
rect -18422 -11683 -18356 -11671
rect -18326 -11565 -18260 -11553
rect -18326 -11671 -18310 -11565
rect -18276 -11671 -18260 -11565
rect -18326 -11683 -18260 -11671
rect -18230 -11565 -18164 -11553
rect -18230 -11671 -18214 -11565
rect -18180 -11671 -18164 -11565
rect -18230 -11683 -18164 -11671
rect -18134 -11565 -18068 -11553
rect -18134 -11671 -18118 -11565
rect -18084 -11671 -18068 -11565
rect -18134 -11683 -18068 -11671
rect -18038 -11565 -17972 -11553
rect -18038 -11671 -18022 -11565
rect -17988 -11671 -17972 -11565
rect -18038 -11683 -17972 -11671
rect -17942 -11565 -17880 -11553
rect -17942 -11671 -17926 -11565
rect -17892 -11671 -17880 -11565
rect -17942 -11683 -17880 -11671
rect -17850 -11565 -17792 -11553
rect -17850 -11671 -17838 -11565
rect -17804 -11671 -17792 -11565
rect -17850 -11683 -17792 -11671
rect -17446 -11565 -17388 -11553
rect -17446 -11671 -17434 -11565
rect -17400 -11671 -17388 -11565
rect -17446 -11683 -17388 -11671
rect -17358 -11565 -17296 -11553
rect -17358 -11671 -17346 -11565
rect -17312 -11671 -17296 -11565
rect -17358 -11683 -17296 -11671
rect -17266 -11565 -17200 -11553
rect -17266 -11671 -17250 -11565
rect -17216 -11671 -17200 -11565
rect -17266 -11683 -17200 -11671
rect -17170 -11565 -17104 -11553
rect -17170 -11671 -17154 -11565
rect -17120 -11671 -17104 -11565
rect -17170 -11683 -17104 -11671
rect -17074 -11565 -17008 -11553
rect -17074 -11671 -17058 -11565
rect -17024 -11671 -17008 -11565
rect -17074 -11683 -17008 -11671
rect -16978 -11565 -16912 -11553
rect -16978 -11671 -16962 -11565
rect -16928 -11671 -16912 -11565
rect -16978 -11683 -16912 -11671
rect -16882 -11565 -16816 -11553
rect -16882 -11671 -16866 -11565
rect -16832 -11671 -16816 -11565
rect -16882 -11683 -16816 -11671
rect -16786 -11565 -16720 -11553
rect -16786 -11671 -16770 -11565
rect -16736 -11671 -16720 -11565
rect -16786 -11683 -16720 -11671
rect -16690 -11565 -16624 -11553
rect -16690 -11671 -16674 -11565
rect -16640 -11671 -16624 -11565
rect -16690 -11683 -16624 -11671
rect -16594 -11565 -16528 -11553
rect -16594 -11671 -16578 -11565
rect -16544 -11671 -16528 -11565
rect -16594 -11683 -16528 -11671
rect -16498 -11565 -16432 -11553
rect -16498 -11671 -16482 -11565
rect -16448 -11671 -16432 -11565
rect -16498 -11683 -16432 -11671
rect -16402 -11565 -16336 -11553
rect -16402 -11671 -16386 -11565
rect -16352 -11671 -16336 -11565
rect -16402 -11683 -16336 -11671
rect -16306 -11565 -16240 -11553
rect -16306 -11671 -16290 -11565
rect -16256 -11671 -16240 -11565
rect -16306 -11683 -16240 -11671
rect -16210 -11565 -16148 -11553
rect -16210 -11671 -16194 -11565
rect -16160 -11671 -16148 -11565
rect -16210 -11683 -16148 -11671
rect -16118 -11565 -16060 -11553
rect -16118 -11671 -16106 -11565
rect -16072 -11671 -16060 -11565
rect -16118 -11683 -16060 -11671
rect -15887 -11565 -15829 -11553
rect -15887 -11671 -15875 -11565
rect -15841 -11671 -15829 -11565
rect -15887 -11683 -15829 -11671
rect -15799 -11565 -15737 -11553
rect -15799 -11671 -15787 -11565
rect -15753 -11671 -15737 -11565
rect -15799 -11683 -15737 -11671
rect -15707 -11565 -15641 -11553
rect -15707 -11671 -15691 -11565
rect -15657 -11671 -15641 -11565
rect -15707 -11683 -15641 -11671
rect -15611 -11565 -15545 -11553
rect -15611 -11671 -15595 -11565
rect -15561 -11671 -15545 -11565
rect -15611 -11683 -15545 -11671
rect -15515 -11565 -15449 -11553
rect -15515 -11671 -15499 -11565
rect -15465 -11671 -15449 -11565
rect -15515 -11683 -15449 -11671
rect -15419 -11565 -15353 -11553
rect -15419 -11671 -15403 -11565
rect -15369 -11671 -15353 -11565
rect -15419 -11683 -15353 -11671
rect -15323 -11565 -15257 -11553
rect -15323 -11671 -15307 -11565
rect -15273 -11671 -15257 -11565
rect -15323 -11683 -15257 -11671
rect -15227 -11565 -15161 -11553
rect -15227 -11671 -15211 -11565
rect -15177 -11671 -15161 -11565
rect -15227 -11683 -15161 -11671
rect -15131 -11565 -15065 -11553
rect -15131 -11671 -15115 -11565
rect -15081 -11671 -15065 -11565
rect -15131 -11683 -15065 -11671
rect -15035 -11565 -14969 -11553
rect -15035 -11671 -15019 -11565
rect -14985 -11671 -14969 -11565
rect -15035 -11683 -14969 -11671
rect -14939 -11565 -14873 -11553
rect -14939 -11671 -14923 -11565
rect -14889 -11671 -14873 -11565
rect -14939 -11683 -14873 -11671
rect -14843 -11565 -14777 -11553
rect -14843 -11671 -14827 -11565
rect -14793 -11671 -14777 -11565
rect -14843 -11683 -14777 -11671
rect -14747 -11565 -14681 -11553
rect -14747 -11671 -14731 -11565
rect -14697 -11671 -14681 -11565
rect -14747 -11683 -14681 -11671
rect -14651 -11565 -14589 -11553
rect -14651 -11671 -14635 -11565
rect -14601 -11671 -14589 -11565
rect -14651 -11683 -14589 -11671
rect -14559 -11565 -14501 -11553
rect -14559 -11671 -14547 -11565
rect -14513 -11671 -14501 -11565
rect -14559 -11683 -14501 -11671
rect -14155 -11565 -14097 -11553
rect -14155 -11671 -14143 -11565
rect -14109 -11671 -14097 -11565
rect -14155 -11683 -14097 -11671
rect -14067 -11565 -14005 -11553
rect -14067 -11671 -14055 -11565
rect -14021 -11671 -14005 -11565
rect -14067 -11683 -14005 -11671
rect -13975 -11565 -13909 -11553
rect -13975 -11671 -13959 -11565
rect -13925 -11671 -13909 -11565
rect -13975 -11683 -13909 -11671
rect -13879 -11565 -13813 -11553
rect -13879 -11671 -13863 -11565
rect -13829 -11671 -13813 -11565
rect -13879 -11683 -13813 -11671
rect -13783 -11565 -13717 -11553
rect -13783 -11671 -13767 -11565
rect -13733 -11671 -13717 -11565
rect -13783 -11683 -13717 -11671
rect -13687 -11565 -13621 -11553
rect -13687 -11671 -13671 -11565
rect -13637 -11671 -13621 -11565
rect -13687 -11683 -13621 -11671
rect -13591 -11565 -13525 -11553
rect -13591 -11671 -13575 -11565
rect -13541 -11671 -13525 -11565
rect -13591 -11683 -13525 -11671
rect -13495 -11565 -13429 -11553
rect -13495 -11671 -13479 -11565
rect -13445 -11671 -13429 -11565
rect -13495 -11683 -13429 -11671
rect -13399 -11565 -13333 -11553
rect -13399 -11671 -13383 -11565
rect -13349 -11671 -13333 -11565
rect -13399 -11683 -13333 -11671
rect -13303 -11565 -13237 -11553
rect -13303 -11671 -13287 -11565
rect -13253 -11671 -13237 -11565
rect -13303 -11683 -13237 -11671
rect -13207 -11565 -13141 -11553
rect -13207 -11671 -13191 -11565
rect -13157 -11671 -13141 -11565
rect -13207 -11683 -13141 -11671
rect -13111 -11565 -13045 -11553
rect -13111 -11671 -13095 -11565
rect -13061 -11671 -13045 -11565
rect -13111 -11683 -13045 -11671
rect -13015 -11565 -12949 -11553
rect -13015 -11671 -12999 -11565
rect -12965 -11671 -12949 -11565
rect -13015 -11683 -12949 -11671
rect -12919 -11565 -12857 -11553
rect -12919 -11671 -12903 -11565
rect -12869 -11671 -12857 -11565
rect -12919 -11683 -12857 -11671
rect -12827 -11565 -12769 -11553
rect -12827 -11671 -12815 -11565
rect -12781 -11671 -12769 -11565
rect -12827 -11683 -12769 -11671
rect -12596 -11565 -12538 -11553
rect -12596 -11671 -12584 -11565
rect -12550 -11671 -12538 -11565
rect -12596 -11683 -12538 -11671
rect -12508 -11565 -12446 -11553
rect -12508 -11671 -12496 -11565
rect -12462 -11671 -12446 -11565
rect -12508 -11683 -12446 -11671
rect -12416 -11565 -12350 -11553
rect -12416 -11671 -12400 -11565
rect -12366 -11671 -12350 -11565
rect -12416 -11683 -12350 -11671
rect -12320 -11565 -12254 -11553
rect -12320 -11671 -12304 -11565
rect -12270 -11671 -12254 -11565
rect -12320 -11683 -12254 -11671
rect -12224 -11565 -12158 -11553
rect -12224 -11671 -12208 -11565
rect -12174 -11671 -12158 -11565
rect -12224 -11683 -12158 -11671
rect -12128 -11565 -12062 -11553
rect -12128 -11671 -12112 -11565
rect -12078 -11671 -12062 -11565
rect -12128 -11683 -12062 -11671
rect -12032 -11565 -11966 -11553
rect -12032 -11671 -12016 -11565
rect -11982 -11671 -11966 -11565
rect -12032 -11683 -11966 -11671
rect -11936 -11565 -11870 -11553
rect -11936 -11671 -11920 -11565
rect -11886 -11671 -11870 -11565
rect -11936 -11683 -11870 -11671
rect -11840 -11565 -11774 -11553
rect -11840 -11671 -11824 -11565
rect -11790 -11671 -11774 -11565
rect -11840 -11683 -11774 -11671
rect -11744 -11565 -11678 -11553
rect -11744 -11671 -11728 -11565
rect -11694 -11671 -11678 -11565
rect -11744 -11683 -11678 -11671
rect -11648 -11565 -11582 -11553
rect -11648 -11671 -11632 -11565
rect -11598 -11671 -11582 -11565
rect -11648 -11683 -11582 -11671
rect -11552 -11565 -11486 -11553
rect -11552 -11671 -11536 -11565
rect -11502 -11671 -11486 -11565
rect -11552 -11683 -11486 -11671
rect -11456 -11565 -11390 -11553
rect -11456 -11671 -11440 -11565
rect -11406 -11671 -11390 -11565
rect -11456 -11683 -11390 -11671
rect -11360 -11565 -11298 -11553
rect -11360 -11671 -11344 -11565
rect -11310 -11671 -11298 -11565
rect -11360 -11683 -11298 -11671
rect -11268 -11565 -11210 -11553
rect -11268 -11671 -11256 -11565
rect -11222 -11671 -11210 -11565
rect -11268 -11683 -11210 -11671
rect -10864 -11565 -10806 -11553
rect -10864 -11671 -10852 -11565
rect -10818 -11671 -10806 -11565
rect -10864 -11683 -10806 -11671
rect -10776 -11565 -10714 -11553
rect -10776 -11671 -10764 -11565
rect -10730 -11671 -10714 -11565
rect -10776 -11683 -10714 -11671
rect -10684 -11565 -10618 -11553
rect -10684 -11671 -10668 -11565
rect -10634 -11671 -10618 -11565
rect -10684 -11683 -10618 -11671
rect -10588 -11565 -10522 -11553
rect -10588 -11671 -10572 -11565
rect -10538 -11671 -10522 -11565
rect -10588 -11683 -10522 -11671
rect -10492 -11565 -10426 -11553
rect -10492 -11671 -10476 -11565
rect -10442 -11671 -10426 -11565
rect -10492 -11683 -10426 -11671
rect -10396 -11565 -10330 -11553
rect -10396 -11671 -10380 -11565
rect -10346 -11671 -10330 -11565
rect -10396 -11683 -10330 -11671
rect -10300 -11565 -10234 -11553
rect -10300 -11671 -10284 -11565
rect -10250 -11671 -10234 -11565
rect -10300 -11683 -10234 -11671
rect -10204 -11565 -10138 -11553
rect -10204 -11671 -10188 -11565
rect -10154 -11671 -10138 -11565
rect -10204 -11683 -10138 -11671
rect -10108 -11565 -10042 -11553
rect -10108 -11671 -10092 -11565
rect -10058 -11671 -10042 -11565
rect -10108 -11683 -10042 -11671
rect -10012 -11565 -9946 -11553
rect -10012 -11671 -9996 -11565
rect -9962 -11671 -9946 -11565
rect -10012 -11683 -9946 -11671
rect -9916 -11565 -9850 -11553
rect -9916 -11671 -9900 -11565
rect -9866 -11671 -9850 -11565
rect -9916 -11683 -9850 -11671
rect -9820 -11565 -9754 -11553
rect -9820 -11671 -9804 -11565
rect -9770 -11671 -9754 -11565
rect -9820 -11683 -9754 -11671
rect -9724 -11565 -9658 -11553
rect -9724 -11671 -9708 -11565
rect -9674 -11671 -9658 -11565
rect -9724 -11683 -9658 -11671
rect -9628 -11565 -9566 -11553
rect -9628 -11671 -9612 -11565
rect -9578 -11671 -9566 -11565
rect -9628 -11683 -9566 -11671
rect -9536 -11565 -9478 -11553
rect -9536 -11671 -9524 -11565
rect -9490 -11671 -9478 -11565
rect -9536 -11683 -9478 -11671
rect -9305 -11565 -9247 -11553
rect -9305 -11671 -9293 -11565
rect -9259 -11671 -9247 -11565
rect -9305 -11683 -9247 -11671
rect -9217 -11565 -9155 -11553
rect -9217 -11671 -9205 -11565
rect -9171 -11671 -9155 -11565
rect -9217 -11683 -9155 -11671
rect -9125 -11565 -9059 -11553
rect -9125 -11671 -9109 -11565
rect -9075 -11671 -9059 -11565
rect -9125 -11683 -9059 -11671
rect -9029 -11565 -8963 -11553
rect -9029 -11671 -9013 -11565
rect -8979 -11671 -8963 -11565
rect -9029 -11683 -8963 -11671
rect -8933 -11565 -8867 -11553
rect -8933 -11671 -8917 -11565
rect -8883 -11671 -8867 -11565
rect -8933 -11683 -8867 -11671
rect -8837 -11565 -8771 -11553
rect -8837 -11671 -8821 -11565
rect -8787 -11671 -8771 -11565
rect -8837 -11683 -8771 -11671
rect -8741 -11565 -8675 -11553
rect -8741 -11671 -8725 -11565
rect -8691 -11671 -8675 -11565
rect -8741 -11683 -8675 -11671
rect -8645 -11565 -8579 -11553
rect -8645 -11671 -8629 -11565
rect -8595 -11671 -8579 -11565
rect -8645 -11683 -8579 -11671
rect -8549 -11565 -8483 -11553
rect -8549 -11671 -8533 -11565
rect -8499 -11671 -8483 -11565
rect -8549 -11683 -8483 -11671
rect -8453 -11565 -8387 -11553
rect -8453 -11671 -8437 -11565
rect -8403 -11671 -8387 -11565
rect -8453 -11683 -8387 -11671
rect -8357 -11565 -8291 -11553
rect -8357 -11671 -8341 -11565
rect -8307 -11671 -8291 -11565
rect -8357 -11683 -8291 -11671
rect -8261 -11565 -8195 -11553
rect -8261 -11671 -8245 -11565
rect -8211 -11671 -8195 -11565
rect -8261 -11683 -8195 -11671
rect -8165 -11565 -8099 -11553
rect -8165 -11671 -8149 -11565
rect -8115 -11671 -8099 -11565
rect -8165 -11683 -8099 -11671
rect -8069 -11565 -8007 -11553
rect -8069 -11671 -8053 -11565
rect -8019 -11671 -8007 -11565
rect -8069 -11683 -8007 -11671
rect -7977 -11565 -7919 -11553
rect -7977 -11671 -7965 -11565
rect -7931 -11671 -7919 -11565
rect -7977 -11683 -7919 -11671
rect 7360 -11882 7372 -11106
rect 7406 -11882 7422 -11106
rect 7360 -11894 7422 -11882
rect 7452 -11894 7518 -11094
rect 7548 -11894 7614 -11094
rect 7644 -11894 7710 -11094
rect 7740 -11106 7802 -11094
rect 7740 -11882 7756 -11106
rect 7790 -11882 7802 -11106
rect 7740 -11894 7802 -11882
rect 8308 -11106 8370 -11094
rect 8308 -11882 8320 -11106
rect 8354 -11882 8370 -11106
rect 8308 -11894 8370 -11882
rect 8400 -11894 8466 -11094
rect 8496 -11894 8562 -11094
rect 8592 -11894 8658 -11094
rect 8688 -11106 8750 -11094
rect 8688 -11882 8704 -11106
rect 8738 -11882 8750 -11106
rect 8688 -11894 8750 -11882
rect 9244 -11106 9306 -11094
rect 9244 -11882 9256 -11106
rect 9290 -11882 9306 -11106
rect 9244 -11894 9306 -11882
rect 9336 -11894 9402 -11094
rect 9432 -11894 9498 -11094
rect 9528 -11894 9594 -11094
rect 9624 -11106 9686 -11094
rect 9624 -11882 9640 -11106
rect 9674 -11882 9686 -11106
rect 9624 -11894 9686 -11882
rect 10175 -11106 10237 -11094
rect 10175 -11882 10187 -11106
rect 10221 -11882 10237 -11106
rect 10175 -11894 10237 -11882
rect 10267 -11894 10333 -11094
rect 10363 -11894 10429 -11094
rect 10459 -11894 10525 -11094
rect 10555 -11106 10617 -11094
rect 10555 -11882 10571 -11106
rect 10605 -11882 10617 -11106
rect 10555 -11894 10617 -11882
rect 11102 -11106 11164 -11094
rect 11102 -11882 11114 -11106
rect 11148 -11882 11164 -11106
rect 11102 -11894 11164 -11882
rect 11194 -11894 11260 -11094
rect 11290 -11894 11356 -11094
rect 11386 -11894 11452 -11094
rect 11482 -11106 11544 -11094
rect 11482 -11882 11498 -11106
rect 11532 -11882 11544 -11106
rect 11482 -11894 11544 -11882
rect 7360 -12034 7422 -12022
rect -24162 -12402 -23762 -12390
rect -24162 -12436 -24150 -12402
rect -23774 -12436 -23762 -12402
rect -23583 -12402 -23383 -12390
rect -24162 -12452 -23762 -12436
rect -23583 -12436 -23571 -12402
rect -23395 -12436 -23383 -12402
rect -23583 -12448 -23383 -12436
rect -24162 -12548 -23762 -12482
rect -23583 -12490 -23383 -12478
rect -23583 -12524 -23571 -12490
rect -23395 -12524 -23383 -12490
rect -23583 -12536 -23383 -12524
rect -22425 -12402 -22025 -12390
rect -22425 -12436 -22413 -12402
rect -22037 -12436 -22025 -12402
rect -21854 -12402 -21654 -12390
rect -22425 -12452 -22025 -12436
rect -21854 -12436 -21842 -12402
rect -21666 -12436 -21654 -12402
rect -21854 -12448 -21654 -12436
rect -22425 -12548 -22025 -12482
rect -21854 -12490 -21654 -12478
rect -21854 -12524 -21842 -12490
rect -21666 -12524 -21654 -12490
rect -21854 -12536 -21654 -12524
rect -24162 -12594 -23762 -12578
rect -24162 -12628 -24150 -12594
rect -23774 -12628 -23762 -12594
rect -24162 -12640 -23762 -12628
rect -22425 -12594 -22025 -12578
rect -22425 -12628 -22413 -12594
rect -22037 -12628 -22025 -12594
rect -22425 -12640 -22025 -12628
rect -20296 -12570 -19896 -12558
rect -20296 -12604 -20284 -12570
rect -19908 -12604 -19896 -12570
rect -20296 -12620 -19896 -12604
rect -20296 -12716 -19896 -12650
rect -19187 -12570 -18787 -12558
rect -19187 -12604 -19175 -12570
rect -18799 -12604 -18787 -12570
rect -19187 -12620 -18787 -12604
rect -19187 -12716 -18787 -12650
rect -18305 -12570 -17905 -12558
rect -18305 -12604 -18293 -12570
rect -17917 -12604 -17905 -12570
rect -18305 -12620 -17905 -12604
rect -18305 -12716 -17905 -12650
rect -17005 -12570 -16605 -12558
rect -17005 -12604 -16993 -12570
rect -16617 -12604 -16605 -12570
rect -17005 -12620 -16605 -12604
rect -17005 -12716 -16605 -12650
rect -15896 -12570 -15496 -12558
rect -15896 -12604 -15884 -12570
rect -15508 -12604 -15496 -12570
rect -15896 -12620 -15496 -12604
rect -15896 -12716 -15496 -12650
rect -15014 -12570 -14614 -12558
rect -15014 -12604 -15002 -12570
rect -14626 -12604 -14614 -12570
rect -15014 -12620 -14614 -12604
rect -15014 -12716 -14614 -12650
rect -13714 -12570 -13314 -12558
rect -13714 -12604 -13702 -12570
rect -13326 -12604 -13314 -12570
rect -13714 -12620 -13314 -12604
rect -13714 -12716 -13314 -12650
rect -12605 -12570 -12205 -12558
rect -12605 -12604 -12593 -12570
rect -12217 -12604 -12205 -12570
rect -12605 -12620 -12205 -12604
rect -12605 -12716 -12205 -12650
rect -11723 -12570 -11323 -12558
rect -11723 -12604 -11711 -12570
rect -11335 -12604 -11323 -12570
rect -11723 -12620 -11323 -12604
rect -11723 -12716 -11323 -12650
rect -10423 -12570 -10023 -12558
rect -10423 -12604 -10411 -12570
rect -10035 -12604 -10023 -12570
rect -10423 -12620 -10023 -12604
rect -10423 -12716 -10023 -12650
rect -9314 -12570 -8914 -12558
rect -9314 -12604 -9302 -12570
rect -8926 -12604 -8914 -12570
rect -9314 -12620 -8914 -12604
rect -9314 -12716 -8914 -12650
rect -8432 -12570 -8032 -12558
rect -8432 -12604 -8420 -12570
rect -8044 -12604 -8032 -12570
rect -8432 -12620 -8032 -12604
rect -8432 -12716 -8032 -12650
rect -20296 -12762 -19896 -12746
rect -20296 -12796 -20284 -12762
rect -19908 -12796 -19896 -12762
rect -19187 -12762 -18787 -12746
rect -20296 -12808 -19896 -12796
rect -19187 -12796 -19175 -12762
rect -18799 -12796 -18787 -12762
rect -18305 -12762 -17905 -12746
rect -19187 -12808 -18787 -12796
rect -18305 -12796 -18293 -12762
rect -17917 -12796 -17905 -12762
rect -17005 -12762 -16605 -12746
rect -18305 -12808 -17905 -12796
rect -17005 -12796 -16993 -12762
rect -16617 -12796 -16605 -12762
rect -15896 -12762 -15496 -12746
rect -17005 -12808 -16605 -12796
rect -15896 -12796 -15884 -12762
rect -15508 -12796 -15496 -12762
rect -15014 -12762 -14614 -12746
rect -15896 -12808 -15496 -12796
rect -15014 -12796 -15002 -12762
rect -14626 -12796 -14614 -12762
rect -13714 -12762 -13314 -12746
rect -15014 -12808 -14614 -12796
rect -13714 -12796 -13702 -12762
rect -13326 -12796 -13314 -12762
rect -12605 -12762 -12205 -12746
rect -13714 -12808 -13314 -12796
rect -12605 -12796 -12593 -12762
rect -12217 -12796 -12205 -12762
rect -11723 -12762 -11323 -12746
rect -12605 -12808 -12205 -12796
rect -11723 -12796 -11711 -12762
rect -11335 -12796 -11323 -12762
rect -10423 -12762 -10023 -12746
rect -11723 -12808 -11323 -12796
rect -10423 -12796 -10411 -12762
rect -10035 -12796 -10023 -12762
rect -9314 -12762 -8914 -12746
rect -10423 -12808 -10023 -12796
rect -9314 -12796 -9302 -12762
rect -8926 -12796 -8914 -12762
rect -8432 -12762 -8032 -12746
rect -9314 -12808 -8914 -12796
rect -8432 -12796 -8420 -12762
rect -8044 -12796 -8032 -12762
rect -8432 -12808 -8032 -12796
rect 7360 -12810 7372 -12034
rect 7406 -12810 7422 -12034
rect 7360 -12822 7422 -12810
rect 7452 -12822 7518 -12022
rect 7548 -12822 7614 -12022
rect 7644 -12822 7710 -12022
rect 7740 -12034 7802 -12022
rect 7740 -12810 7756 -12034
rect 7790 -12810 7802 -12034
rect 7740 -12822 7802 -12810
rect 8308 -12034 8370 -12022
rect 8308 -12810 8320 -12034
rect 8354 -12810 8370 -12034
rect 8308 -12822 8370 -12810
rect 8400 -12822 8466 -12022
rect 8496 -12822 8562 -12022
rect 8592 -12822 8658 -12022
rect 8688 -12034 8750 -12022
rect 8688 -12810 8704 -12034
rect 8738 -12810 8750 -12034
rect 8688 -12822 8750 -12810
rect 9244 -12034 9306 -12022
rect 9244 -12810 9256 -12034
rect 9290 -12810 9306 -12034
rect 9244 -12822 9306 -12810
rect 9336 -12822 9402 -12022
rect 9432 -12822 9498 -12022
rect 9528 -12822 9594 -12022
rect 9624 -12034 9686 -12022
rect 9624 -12810 9640 -12034
rect 9674 -12810 9686 -12034
rect 9624 -12822 9686 -12810
rect 10175 -12033 10237 -12021
rect 10175 -12809 10187 -12033
rect 10221 -12809 10237 -12033
rect 10175 -12821 10237 -12809
rect 10267 -12821 10333 -12021
rect 10363 -12821 10429 -12021
rect 10459 -12821 10525 -12021
rect 10555 -12033 10617 -12021
rect 10555 -12809 10571 -12033
rect 10605 -12809 10617 -12033
rect 10555 -12821 10617 -12809
rect 11102 -12034 11164 -12022
rect 11102 -12810 11114 -12034
rect 11148 -12810 11164 -12034
rect 11102 -12822 11164 -12810
rect 11194 -12822 11260 -12022
rect 11290 -12822 11356 -12022
rect 11386 -12822 11452 -12022
rect 11482 -12034 11544 -12022
rect 11482 -12810 11498 -12034
rect 11532 -12810 11544 -12034
rect 12157 -12076 12219 -12064
rect 12157 -12252 12169 -12076
rect 12203 -12252 12219 -12076
rect 12157 -12264 12219 -12252
rect 12249 -12076 12315 -12064
rect 12249 -12252 12265 -12076
rect 12299 -12252 12315 -12076
rect 12249 -12264 12315 -12252
rect 12345 -12076 12407 -12064
rect 12345 -12252 12361 -12076
rect 12395 -12252 12407 -12076
rect 12923 -12141 13123 -12129
rect 12923 -12175 12935 -12141
rect 13111 -12175 13123 -12141
rect 12923 -12187 13123 -12175
rect 12923 -12229 13123 -12217
rect 12345 -12264 12407 -12252
rect 12923 -12263 12935 -12229
rect 13111 -12263 13123 -12229
rect 12923 -12275 13123 -12263
rect 11482 -12822 11544 -12810
rect -1662 -13844 -1604 -13832
rect -1662 -14020 -1650 -13844
rect -1616 -14020 -1604 -13844
rect -1662 -14032 -1604 -14020
rect -1574 -13844 -1516 -13832
rect -1574 -14020 -1562 -13844
rect -1528 -14020 -1516 -13844
rect -1574 -14032 -1516 -14020
rect -11276 -14105 -11146 -14093
rect -11276 -14139 -11264 -14105
rect -11158 -14139 -11146 -14105
rect -11276 -14151 -11146 -14139
rect -24105 -14928 -24043 -14916
rect -24105 -15304 -24093 -14928
rect -24059 -15304 -24043 -14928
rect -24105 -15316 -24043 -15304
rect -24013 -15316 -23947 -14916
rect -23917 -14928 -23855 -14916
rect -23917 -15304 -23901 -14928
rect -23867 -15304 -23855 -14928
rect -17188 -14895 -16988 -14883
rect -17188 -14929 -17176 -14895
rect -17000 -14929 -16988 -14895
rect -17188 -14945 -16988 -14929
rect -17188 -14991 -16988 -14975
rect -17188 -15025 -17176 -14991
rect -17000 -15025 -16988 -14991
rect -17188 -15041 -16988 -15025
rect -23917 -15316 -23855 -15304
rect -17188 -15087 -16988 -15071
rect -17188 -15121 -17176 -15087
rect -17000 -15121 -16988 -15087
rect -17188 -15133 -16988 -15121
rect -11276 -14193 -11146 -14181
rect -11276 -14227 -11264 -14193
rect -11158 -14227 -11146 -14193
rect -11276 -14243 -11146 -14227
rect -11276 -14289 -11146 -14273
rect -11276 -14323 -11264 -14289
rect -11158 -14323 -11146 -14289
rect -11276 -14339 -11146 -14323
rect -11276 -14385 -11146 -14369
rect -11276 -14419 -11264 -14385
rect -11158 -14419 -11146 -14385
rect -11276 -14435 -11146 -14419
rect -11276 -14481 -11146 -14465
rect -11276 -14515 -11264 -14481
rect -11158 -14515 -11146 -14481
rect -11276 -14531 -11146 -14515
rect -11276 -14577 -11146 -14561
rect -11276 -14611 -11264 -14577
rect -11158 -14611 -11146 -14577
rect -11276 -14627 -11146 -14611
rect -11276 -14673 -11146 -14657
rect -11276 -14707 -11264 -14673
rect -11158 -14707 -11146 -14673
rect -11276 -14723 -11146 -14707
rect -11276 -14769 -11146 -14753
rect -11276 -14803 -11264 -14769
rect -11158 -14803 -11146 -14769
rect -11276 -14819 -11146 -14803
rect -11276 -14865 -11146 -14849
rect -11276 -14899 -11264 -14865
rect -11158 -14899 -11146 -14865
rect -11276 -14915 -11146 -14899
rect -11276 -14961 -11146 -14945
rect -11276 -14995 -11264 -14961
rect -11158 -14995 -11146 -14961
rect -11276 -15011 -11146 -14995
rect -11276 -15057 -11146 -15041
rect -11276 -15091 -11264 -15057
rect -11158 -15091 -11146 -15057
rect -11276 -15107 -11146 -15091
rect -11276 -15153 -11146 -15137
rect -11276 -15187 -11264 -15153
rect -11158 -15187 -11146 -15153
rect -11276 -15203 -11146 -15187
rect -11276 -15249 -11146 -15233
rect -11276 -15283 -11264 -15249
rect -11158 -15283 -11146 -15249
rect -11276 -15299 -11146 -15283
rect -11276 -15345 -11146 -15329
rect -11276 -15379 -11264 -15345
rect -11158 -15379 -11146 -15345
rect -11276 -15391 -11146 -15379
rect -4378 -14215 -4320 -14203
rect -4378 -14391 -4366 -14215
rect -4332 -14391 -4320 -14215
rect -4378 -14403 -4320 -14391
rect -4290 -14215 -4232 -14203
rect -4290 -14391 -4278 -14215
rect -4244 -14391 -4232 -14215
rect -4290 -14403 -4232 -14391
rect -1662 -14223 -1604 -14211
rect -1662 -14399 -1650 -14223
rect -1616 -14399 -1604 -14223
rect -1662 -14411 -1604 -14399
rect -1574 -14223 -1516 -14211
rect -1574 -14399 -1562 -14223
rect -1528 -14399 -1516 -14223
rect -1574 -14411 -1516 -14399
rect -4378 -14655 -4320 -14643
rect -4378 -14831 -4366 -14655
rect -4332 -14831 -4320 -14655
rect -4378 -14843 -4320 -14831
rect -4290 -14655 -4232 -14643
rect -4290 -14831 -4278 -14655
rect -4244 -14831 -4232 -14655
rect -4290 -14843 -4232 -14831
rect 5658 -14651 5858 -14639
rect -1662 -14663 -1604 -14651
rect -1662 -14839 -1650 -14663
rect -1616 -14839 -1604 -14663
rect -1662 -14851 -1604 -14839
rect -1574 -14663 -1516 -14651
rect -1574 -14839 -1562 -14663
rect -1528 -14839 -1516 -14663
rect -1574 -14851 -1516 -14839
rect 5658 -14685 5670 -14651
rect 5846 -14685 5858 -14651
rect 6098 -14651 6298 -14639
rect 5658 -14697 5858 -14685
rect 5658 -14739 5858 -14727
rect 5658 -14773 5670 -14739
rect 5846 -14773 5858 -14739
rect 6098 -14685 6110 -14651
rect 6286 -14685 6298 -14651
rect 6538 -14651 6738 -14639
rect 6098 -14697 6298 -14685
rect 6098 -14739 6298 -14727
rect 5658 -14785 5858 -14773
rect 6098 -14773 6110 -14739
rect 6286 -14773 6298 -14739
rect 6538 -14685 6550 -14651
rect 6726 -14685 6738 -14651
rect 6538 -14697 6738 -14685
rect 6538 -14739 6738 -14727
rect 6098 -14785 6298 -14773
rect 6538 -14773 6550 -14739
rect 6726 -14773 6738 -14739
rect 6538 -14785 6738 -14773
rect -4378 -15034 -4320 -15022
rect -4378 -15210 -4366 -15034
rect -4332 -15210 -4320 -15034
rect -4378 -15222 -4320 -15210
rect -4290 -15034 -4232 -15022
rect -4290 -15210 -4278 -15034
rect -4244 -15210 -4232 -15034
rect -4290 -15222 -4232 -15210
rect -1662 -15042 -1604 -15030
rect -1662 -15218 -1650 -15042
rect -1616 -15218 -1604 -15042
rect -1662 -15230 -1604 -15218
rect -1574 -15042 -1516 -15030
rect -1574 -15218 -1562 -15042
rect -1528 -15218 -1516 -15042
rect -1574 -15230 -1516 -15218
rect -11276 -15433 -11146 -15421
rect -11276 -15467 -11264 -15433
rect -11158 -15467 -11146 -15433
rect -11276 -15479 -11146 -15467
rect -7729 -15372 -7671 -15360
rect -7729 -15548 -7717 -15372
rect -7683 -15548 -7671 -15372
rect -7729 -15560 -7671 -15548
rect -7641 -15372 -7583 -15360
rect -7641 -15548 -7629 -15372
rect -7595 -15548 -7583 -15372
rect -7641 -15560 -7583 -15548
rect -4378 -15474 -4320 -15462
rect -4378 -15650 -4366 -15474
rect -4332 -15650 -4320 -15474
rect -4378 -15662 -4320 -15650
rect -4290 -15474 -4232 -15462
rect -4290 -15650 -4278 -15474
rect -4244 -15650 -4232 -15474
rect -4290 -15662 -4232 -15650
rect -1662 -15482 -1604 -15470
rect -1662 -15658 -1650 -15482
rect -1616 -15658 -1604 -15482
rect -1662 -15670 -1604 -15658
rect -1574 -15482 -1516 -15470
rect -1574 -15658 -1562 -15482
rect -1528 -15658 -1516 -15482
rect -1574 -15670 -1516 -15658
rect 7360 -15634 7422 -15622
rect -7728 -15872 -7670 -15860
rect -7728 -16048 -7716 -15872
rect -7682 -16048 -7670 -15872
rect -7728 -16060 -7670 -16048
rect -7640 -15872 -7582 -15860
rect -7640 -16048 -7628 -15872
rect -7594 -16048 -7582 -15872
rect -7640 -16060 -7582 -16048
rect -4378 -15853 -4320 -15841
rect -4378 -16029 -4366 -15853
rect -4332 -16029 -4320 -15853
rect -4378 -16041 -4320 -16029
rect -4290 -15853 -4232 -15841
rect -4290 -16029 -4278 -15853
rect -4244 -16029 -4232 -15853
rect -4290 -16041 -4232 -16029
rect -24104 -16113 -24042 -16101
rect -24104 -16489 -24092 -16113
rect -24058 -16489 -24042 -16113
rect -24104 -16501 -24042 -16489
rect -24012 -16501 -23946 -16101
rect -23916 -16113 -23854 -16101
rect -23916 -16489 -23900 -16113
rect -23866 -16489 -23854 -16113
rect -1662 -15861 -1604 -15849
rect -1662 -16037 -1650 -15861
rect -1616 -16037 -1604 -15861
rect -1662 -16049 -1604 -16037
rect -1574 -15861 -1516 -15849
rect -1574 -16037 -1562 -15861
rect -1528 -16037 -1516 -15861
rect -1574 -16049 -1516 -16037
rect -17188 -16295 -16988 -16283
rect -17188 -16329 -17176 -16295
rect -17000 -16329 -16988 -16295
rect -17188 -16345 -16988 -16329
rect -17188 -16391 -16988 -16375
rect -17188 -16425 -17176 -16391
rect -17000 -16425 -16988 -16391
rect -17188 -16441 -16988 -16425
rect -23916 -16501 -23854 -16489
rect -17188 -16487 -16988 -16471
rect -17188 -16521 -17176 -16487
rect -17000 -16521 -16988 -16487
rect -17188 -16533 -16988 -16521
rect -7729 -16352 -7671 -16340
rect -7729 -16528 -7717 -16352
rect -7683 -16528 -7671 -16352
rect -7729 -16540 -7671 -16528
rect -7641 -16352 -7583 -16340
rect -7641 -16528 -7629 -16352
rect -7595 -16528 -7583 -16352
rect -7641 -16540 -7583 -16528
rect -4378 -16293 -4320 -16281
rect -4378 -16469 -4366 -16293
rect -4332 -16469 -4320 -16293
rect -4378 -16481 -4320 -16469
rect -4290 -16293 -4232 -16281
rect -4290 -16469 -4278 -16293
rect -4244 -16469 -4232 -16293
rect -4290 -16481 -4232 -16469
rect -1662 -16301 -1604 -16289
rect -1662 -16477 -1650 -16301
rect -1616 -16477 -1604 -16301
rect -1662 -16489 -1604 -16477
rect -1574 -16301 -1516 -16289
rect -1574 -16477 -1562 -16301
rect -1528 -16477 -1516 -16301
rect -1574 -16489 -1516 -16477
rect 7360 -16410 7372 -15634
rect 7406 -16410 7422 -15634
rect 7360 -16422 7422 -16410
rect 7452 -16422 7518 -15622
rect 7548 -16422 7614 -15622
rect 7644 -16422 7710 -15622
rect 7740 -15634 7802 -15622
rect 7740 -16410 7756 -15634
rect 7790 -16410 7802 -15634
rect 7740 -16422 7802 -16410
rect 8308 -15634 8370 -15622
rect 8308 -16410 8320 -15634
rect 8354 -16410 8370 -15634
rect 8308 -16422 8370 -16410
rect 8400 -16422 8466 -15622
rect 8496 -16422 8562 -15622
rect 8592 -16422 8658 -15622
rect 8688 -15634 8750 -15622
rect 8688 -16410 8704 -15634
rect 8738 -16410 8750 -15634
rect 8688 -16422 8750 -16410
rect 9244 -15634 9306 -15622
rect 9244 -16410 9256 -15634
rect 9290 -16410 9306 -15634
rect 9244 -16422 9306 -16410
rect 9336 -16422 9402 -15622
rect 9432 -16422 9498 -15622
rect 9528 -16422 9594 -15622
rect 9624 -15634 9686 -15622
rect 9624 -16410 9640 -15634
rect 9674 -16410 9686 -15634
rect 9624 -16422 9686 -16410
rect 10175 -15634 10237 -15622
rect 10175 -16410 10187 -15634
rect 10221 -16410 10237 -15634
rect 10175 -16422 10237 -16410
rect 10267 -16422 10333 -15622
rect 10363 -16422 10429 -15622
rect 10459 -16422 10525 -15622
rect 10555 -15634 10617 -15622
rect 10555 -16410 10571 -15634
rect 10605 -16410 10617 -15634
rect 10555 -16422 10617 -16410
rect 11102 -15634 11164 -15622
rect 11102 -16410 11114 -15634
rect 11148 -16410 11164 -15634
rect 11102 -16422 11164 -16410
rect 11194 -16422 11260 -15622
rect 11290 -16422 11356 -15622
rect 11386 -16422 11452 -15622
rect 11482 -15634 11544 -15622
rect 11482 -16410 11498 -15634
rect 11532 -16410 11544 -15634
rect 11482 -16422 11544 -16410
rect 7360 -16562 7422 -16550
rect -11274 -16921 -11144 -16909
rect -11274 -16955 -11262 -16921
rect -11156 -16955 -11144 -16921
rect -11274 -16967 -11144 -16955
rect -24099 -17326 -24037 -17314
rect -24099 -17702 -24087 -17326
rect -24053 -17702 -24037 -17326
rect -24099 -17714 -24037 -17702
rect -24007 -17714 -23941 -17314
rect -23911 -17326 -23849 -17314
rect -23911 -17702 -23895 -17326
rect -23861 -17702 -23849 -17326
rect -23911 -17714 -23849 -17702
rect -17188 -17695 -16988 -17683
rect -17188 -17729 -17176 -17695
rect -17000 -17729 -16988 -17695
rect -17188 -17745 -16988 -17729
rect -17188 -17791 -16988 -17775
rect -17188 -17825 -17176 -17791
rect -17000 -17825 -16988 -17791
rect -17188 -17841 -16988 -17825
rect -21168 -18060 -21110 -18048
rect -21168 -18236 -21156 -18060
rect -21122 -18236 -21110 -18060
rect -21168 -18248 -21110 -18236
rect -21080 -18060 -21022 -18048
rect -21080 -18236 -21068 -18060
rect -21034 -18236 -21022 -18060
rect -21080 -18248 -21022 -18236
rect -17188 -17887 -16988 -17871
rect -17188 -17921 -17176 -17887
rect -17000 -17921 -16988 -17887
rect -17188 -17933 -16988 -17921
rect -15577 -17931 -15519 -17919
rect -15577 -18107 -15565 -17931
rect -15531 -18107 -15519 -17931
rect -15577 -18119 -15519 -18107
rect -15489 -17931 -15431 -17919
rect -15489 -18107 -15477 -17931
rect -15443 -18107 -15431 -17931
rect -15489 -18119 -15431 -18107
rect -11274 -17009 -11144 -16997
rect -11274 -17043 -11262 -17009
rect -11156 -17043 -11144 -17009
rect -11274 -17059 -11144 -17043
rect -11274 -17105 -11144 -17089
rect -11274 -17139 -11262 -17105
rect -11156 -17139 -11144 -17105
rect -11274 -17155 -11144 -17139
rect -11274 -17201 -11144 -17185
rect -11274 -17235 -11262 -17201
rect -11156 -17235 -11144 -17201
rect -11274 -17251 -11144 -17235
rect -11274 -17297 -11144 -17281
rect -11274 -17331 -11262 -17297
rect -11156 -17331 -11144 -17297
rect -11274 -17347 -11144 -17331
rect -11274 -17393 -11144 -17377
rect -11274 -17427 -11262 -17393
rect -11156 -17427 -11144 -17393
rect -11274 -17443 -11144 -17427
rect -11274 -17489 -11144 -17473
rect -11274 -17523 -11262 -17489
rect -11156 -17523 -11144 -17489
rect -11274 -17539 -11144 -17523
rect -11274 -17585 -11144 -17569
rect -11274 -17619 -11262 -17585
rect -11156 -17619 -11144 -17585
rect -11274 -17635 -11144 -17619
rect -11274 -17681 -11144 -17665
rect -11274 -17715 -11262 -17681
rect -11156 -17715 -11144 -17681
rect -11274 -17731 -11144 -17715
rect -11274 -17777 -11144 -17761
rect -11274 -17811 -11262 -17777
rect -11156 -17811 -11144 -17777
rect -11274 -17827 -11144 -17811
rect -11274 -17873 -11144 -17857
rect -11274 -17907 -11262 -17873
rect -11156 -17907 -11144 -17873
rect -11274 -17923 -11144 -17907
rect -11274 -17969 -11144 -17953
rect -11274 -18003 -11262 -17969
rect -11156 -18003 -11144 -17969
rect -11274 -18019 -11144 -18003
rect -11274 -18065 -11144 -18049
rect -11274 -18099 -11262 -18065
rect -11156 -18099 -11144 -18065
rect -11274 -18115 -11144 -18099
rect -11274 -18161 -11144 -18145
rect -11274 -18195 -11262 -18161
rect -11156 -18195 -11144 -18161
rect -11274 -18207 -11144 -18195
rect -7729 -16852 -7671 -16840
rect -7729 -17028 -7717 -16852
rect -7683 -17028 -7671 -16852
rect -7729 -17040 -7671 -17028
rect -7641 -16852 -7583 -16840
rect -7641 -17028 -7629 -16852
rect -7595 -17028 -7583 -16852
rect -7641 -17040 -7583 -17028
rect -4378 -16672 -4320 -16660
rect -4378 -16848 -4366 -16672
rect -4332 -16848 -4320 -16672
rect -4378 -16860 -4320 -16848
rect -4290 -16672 -4232 -16660
rect -4290 -16848 -4278 -16672
rect -4244 -16848 -4232 -16672
rect -4290 -16860 -4232 -16848
rect -1662 -16680 -1604 -16668
rect -1662 -16856 -1650 -16680
rect -1616 -16856 -1604 -16680
rect -1662 -16868 -1604 -16856
rect -1574 -16680 -1516 -16668
rect -1574 -16856 -1562 -16680
rect -1528 -16856 -1516 -16680
rect -1574 -16868 -1516 -16856
rect -4378 -17112 -4320 -17100
rect -4378 -17288 -4366 -17112
rect -4332 -17288 -4320 -17112
rect -4378 -17300 -4320 -17288
rect -4290 -17112 -4232 -17100
rect -4290 -17288 -4278 -17112
rect -4244 -17288 -4232 -17112
rect -4290 -17300 -4232 -17288
rect -7729 -17332 -7671 -17320
rect -7729 -17508 -7717 -17332
rect -7683 -17508 -7671 -17332
rect -7729 -17520 -7671 -17508
rect -7641 -17332 -7583 -17320
rect -7641 -17508 -7629 -17332
rect -7595 -17508 -7583 -17332
rect -7641 -17520 -7583 -17508
rect -1662 -17120 -1604 -17108
rect -1662 -17296 -1650 -17120
rect -1616 -17296 -1604 -17120
rect -1662 -17308 -1604 -17296
rect -1574 -17120 -1516 -17108
rect -1574 -17296 -1562 -17120
rect -1528 -17296 -1516 -17120
rect -1574 -17308 -1516 -17296
rect 7360 -17338 7372 -16562
rect 7406 -17338 7422 -16562
rect 7360 -17350 7422 -17338
rect 7452 -17350 7518 -16550
rect 7548 -17350 7614 -16550
rect 7644 -17350 7710 -16550
rect 7740 -16562 7802 -16550
rect 7740 -17338 7756 -16562
rect 7790 -17338 7802 -16562
rect 7740 -17350 7802 -17338
rect 8308 -16562 8370 -16550
rect 8308 -17338 8320 -16562
rect 8354 -17338 8370 -16562
rect 8308 -17350 8370 -17338
rect 8400 -17350 8466 -16550
rect 8496 -17350 8562 -16550
rect 8592 -17350 8658 -16550
rect 8688 -16562 8750 -16550
rect 8688 -17338 8704 -16562
rect 8738 -17338 8750 -16562
rect 8688 -17350 8750 -17338
rect 9244 -16562 9306 -16550
rect 9244 -17338 9256 -16562
rect 9290 -17338 9306 -16562
rect 9244 -17350 9306 -17338
rect 9336 -17350 9402 -16550
rect 9432 -17350 9498 -16550
rect 9528 -17350 9594 -16550
rect 9624 -16562 9686 -16550
rect 9624 -17338 9640 -16562
rect 9674 -17338 9686 -16562
rect 9624 -17350 9686 -17338
rect 10175 -16561 10237 -16549
rect 10175 -17337 10187 -16561
rect 10221 -17337 10237 -16561
rect 10175 -17349 10237 -17337
rect 10267 -17349 10333 -16549
rect 10363 -17349 10429 -16549
rect 10459 -17349 10525 -16549
rect 10555 -16561 10617 -16549
rect 10555 -17337 10571 -16561
rect 10605 -17337 10617 -16561
rect 10555 -17349 10617 -17337
rect 11102 -16562 11164 -16550
rect -4378 -17491 -4320 -17479
rect -4378 -17667 -4366 -17491
rect -4332 -17667 -4320 -17491
rect -4378 -17679 -4320 -17667
rect -4290 -17491 -4232 -17479
rect -4290 -17667 -4278 -17491
rect -4244 -17667 -4232 -17491
rect -4290 -17679 -4232 -17667
rect -1662 -17499 -1604 -17487
rect -1662 -17675 -1650 -17499
rect -1616 -17675 -1604 -17499
rect -1662 -17687 -1604 -17675
rect -1574 -17499 -1516 -17487
rect -1574 -17675 -1562 -17499
rect -1528 -17675 -1516 -17499
rect -1574 -17687 -1516 -17675
rect -7729 -17792 -7671 -17780
rect -7729 -17968 -7717 -17792
rect -7683 -17968 -7671 -17792
rect -7729 -17980 -7671 -17968
rect -7641 -17792 -7583 -17780
rect -7641 -17968 -7629 -17792
rect -7595 -17968 -7583 -17792
rect -7641 -17980 -7583 -17968
rect 11102 -17338 11114 -16562
rect 11148 -17338 11164 -16562
rect 11102 -17350 11164 -17338
rect 11194 -17350 11260 -16550
rect 11290 -17350 11356 -16550
rect 11386 -17350 11452 -16550
rect 11482 -16562 11544 -16550
rect 11482 -17338 11498 -16562
rect 11532 -17338 11544 -16562
rect 12157 -16604 12219 -16592
rect 12157 -16780 12169 -16604
rect 12203 -16780 12219 -16604
rect 12157 -16792 12219 -16780
rect 12249 -16604 12315 -16592
rect 12249 -16780 12265 -16604
rect 12299 -16780 12315 -16604
rect 12249 -16792 12315 -16780
rect 12345 -16604 12407 -16592
rect 12345 -16780 12361 -16604
rect 12395 -16780 12407 -16604
rect 12923 -16669 13123 -16657
rect 12923 -16703 12935 -16669
rect 13111 -16703 13123 -16669
rect 12923 -16715 13123 -16703
rect 12923 -16757 13123 -16745
rect 12345 -16792 12407 -16780
rect 12923 -16791 12935 -16757
rect 13111 -16791 13123 -16757
rect 12923 -16803 13123 -16791
rect 16147 -17061 16209 -17049
rect 16147 -17237 16159 -17061
rect 16193 -17237 16209 -17061
rect 16147 -17249 16209 -17237
rect 16239 -17061 16305 -17049
rect 16239 -17237 16255 -17061
rect 16289 -17237 16305 -17061
rect 16239 -17249 16305 -17237
rect 16335 -17061 16401 -17049
rect 16335 -17237 16351 -17061
rect 16385 -17237 16401 -17061
rect 16335 -17249 16401 -17237
rect 16431 -17061 16497 -17049
rect 16431 -17237 16447 -17061
rect 16481 -17237 16497 -17061
rect 16431 -17249 16497 -17237
rect 16527 -17061 16589 -17049
rect 16527 -17237 16543 -17061
rect 16577 -17237 16589 -17061
rect 16527 -17249 16589 -17237
rect 11482 -17350 11544 -17338
rect -4378 -17931 -4320 -17919
rect -4378 -18107 -4366 -17931
rect -4332 -18107 -4320 -17931
rect -4378 -18119 -4320 -18107
rect -4290 -17931 -4232 -17919
rect -4290 -18107 -4278 -17931
rect -4244 -18107 -4232 -17931
rect -4290 -18119 -4232 -18107
rect -1662 -17939 -1604 -17927
rect -1662 -18115 -1650 -17939
rect -1616 -18115 -1604 -17939
rect -1662 -18127 -1604 -18115
rect -1574 -17939 -1516 -17927
rect -1574 -18115 -1562 -17939
rect -1528 -18115 -1516 -17939
rect -1574 -18127 -1516 -18115
rect -11274 -18249 -11144 -18237
rect -11274 -18283 -11262 -18249
rect -11156 -18283 -11144 -18249
rect -11274 -18295 -11144 -18283
rect -24084 -18445 -24022 -18433
rect -24084 -18821 -24072 -18445
rect -24038 -18821 -24022 -18445
rect -24084 -18833 -24022 -18821
rect -23992 -18833 -23926 -18433
rect -23896 -18445 -23834 -18433
rect -23896 -18821 -23880 -18445
rect -23846 -18821 -23834 -18445
rect -21167 -18560 -21109 -18548
rect -21167 -18736 -21155 -18560
rect -21121 -18736 -21109 -18560
rect -21167 -18748 -21109 -18736
rect -21079 -18560 -21021 -18548
rect -21079 -18736 -21067 -18560
rect -21033 -18736 -21021 -18560
rect -21079 -18748 -21021 -18736
rect -15576 -18431 -15518 -18419
rect -15576 -18607 -15564 -18431
rect -15530 -18607 -15518 -18431
rect -15576 -18619 -15518 -18607
rect -15488 -18431 -15430 -18419
rect -15488 -18607 -15476 -18431
rect -15442 -18607 -15430 -18431
rect -15488 -18619 -15430 -18607
rect -7743 -18252 -7685 -18240
rect -7743 -18428 -7731 -18252
rect -7697 -18428 -7685 -18252
rect -7743 -18440 -7685 -18428
rect -7655 -18252 -7597 -18240
rect -7655 -18428 -7643 -18252
rect -7609 -18428 -7597 -18252
rect -7655 -18440 -7597 -18428
rect -4378 -18310 -4320 -18298
rect -4378 -18486 -4366 -18310
rect -4332 -18486 -4320 -18310
rect -4378 -18498 -4320 -18486
rect -4290 -18310 -4232 -18298
rect -4290 -18486 -4278 -18310
rect -4244 -18486 -4232 -18310
rect -4290 -18498 -4232 -18486
rect -1662 -18318 -1604 -18306
rect -1662 -18494 -1650 -18318
rect -1616 -18494 -1604 -18318
rect -1662 -18506 -1604 -18494
rect -1574 -18318 -1516 -18306
rect -1574 -18494 -1562 -18318
rect -1528 -18494 -1516 -18318
rect -1574 -18506 -1516 -18494
rect -23896 -18833 -23834 -18821
rect -21168 -19040 -21110 -19028
rect -21168 -19216 -21156 -19040
rect -21122 -19216 -21110 -19040
rect -21168 -19228 -21110 -19216
rect -21080 -19040 -21022 -19028
rect -21080 -19216 -21068 -19040
rect -21034 -19216 -21022 -19040
rect -21080 -19228 -21022 -19216
rect -17188 -19095 -16988 -19083
rect -17188 -19129 -17176 -19095
rect -17000 -19129 -16988 -19095
rect -17188 -19145 -16988 -19129
rect -15577 -18911 -15519 -18899
rect -15577 -19087 -15565 -18911
rect -15531 -19087 -15519 -18911
rect -15577 -19099 -15519 -19087
rect -15489 -18911 -15431 -18899
rect -15489 -19087 -15477 -18911
rect -15443 -19087 -15431 -18911
rect -15489 -19099 -15431 -19087
rect -7741 -18732 -7683 -18720
rect -7741 -18908 -7729 -18732
rect -7695 -18908 -7683 -18732
rect -7741 -18920 -7683 -18908
rect -7653 -18732 -7595 -18720
rect -7653 -18908 -7641 -18732
rect -7607 -18908 -7595 -18732
rect -7653 -18920 -7595 -18908
rect -4378 -18750 -4320 -18738
rect -4378 -18926 -4366 -18750
rect -4332 -18926 -4320 -18750
rect -4378 -18938 -4320 -18926
rect -4290 -18750 -4232 -18738
rect -4290 -18926 -4278 -18750
rect -4244 -18926 -4232 -18750
rect -4290 -18938 -4232 -18926
rect -1662 -18758 -1604 -18746
rect -1662 -18934 -1650 -18758
rect -1616 -18934 -1604 -18758
rect -1662 -18946 -1604 -18934
rect -1574 -18758 -1516 -18746
rect -1574 -18934 -1562 -18758
rect -1528 -18934 -1516 -18758
rect -1574 -18946 -1516 -18934
rect -17188 -19191 -16988 -19175
rect -17188 -19225 -17176 -19191
rect -17000 -19225 -16988 -19191
rect -17188 -19241 -16988 -19225
rect -24082 -19639 -24020 -19627
rect -24082 -20015 -24070 -19639
rect -24036 -20015 -24020 -19639
rect -24082 -20027 -24020 -20015
rect -23990 -20027 -23924 -19627
rect -23894 -19639 -23832 -19627
rect -23894 -20015 -23878 -19639
rect -23844 -20015 -23832 -19639
rect -21168 -19540 -21110 -19528
rect -21168 -19716 -21156 -19540
rect -21122 -19716 -21110 -19540
rect -21168 -19728 -21110 -19716
rect -21080 -19540 -21022 -19528
rect -21080 -19716 -21068 -19540
rect -21034 -19716 -21022 -19540
rect -21080 -19728 -21022 -19716
rect -17188 -19287 -16988 -19271
rect -17188 -19321 -17176 -19287
rect -17000 -19321 -16988 -19287
rect -17188 -19333 -16988 -19321
rect -4378 -19129 -4320 -19117
rect -4378 -19305 -4366 -19129
rect -4332 -19305 -4320 -19129
rect -4378 -19317 -4320 -19305
rect -4290 -19129 -4232 -19117
rect -4290 -19305 -4278 -19129
rect -4244 -19305 -4232 -19129
rect -4290 -19317 -4232 -19305
rect -1662 -19137 -1604 -19125
rect -1662 -19313 -1650 -19137
rect -1616 -19313 -1604 -19137
rect -1662 -19325 -1604 -19313
rect -1574 -19137 -1516 -19125
rect -1574 -19313 -1562 -19137
rect -1528 -19313 -1516 -19137
rect -1574 -19325 -1516 -19313
rect 5658 -19179 5858 -19167
rect 5658 -19213 5670 -19179
rect 5846 -19213 5858 -19179
rect 6098 -19179 6298 -19167
rect 5658 -19225 5858 -19213
rect 5658 -19267 5858 -19255
rect 5658 -19301 5670 -19267
rect 5846 -19301 5858 -19267
rect 6098 -19213 6110 -19179
rect 6286 -19213 6298 -19179
rect 6538 -19179 6738 -19167
rect 6098 -19225 6298 -19213
rect 6098 -19267 6298 -19255
rect 5658 -19313 5858 -19301
rect 6098 -19301 6110 -19267
rect 6286 -19301 6298 -19267
rect 6538 -19213 6550 -19179
rect 6726 -19213 6738 -19179
rect 6538 -19225 6738 -19213
rect 6538 -19267 6738 -19255
rect 6098 -19313 6298 -19301
rect 6538 -19301 6550 -19267
rect 6726 -19301 6738 -19267
rect 6538 -19313 6738 -19301
rect -15577 -19411 -15519 -19399
rect -15577 -19587 -15565 -19411
rect -15531 -19587 -15519 -19411
rect -15577 -19599 -15519 -19587
rect -15489 -19411 -15431 -19399
rect -15489 -19587 -15477 -19411
rect -15443 -19587 -15431 -19411
rect -15489 -19599 -15431 -19587
rect -4378 -19569 -4320 -19557
rect -4378 -19745 -4366 -19569
rect -4332 -19745 -4320 -19569
rect -4378 -19757 -4320 -19745
rect -4290 -19569 -4232 -19557
rect -4290 -19745 -4278 -19569
rect -4244 -19745 -4232 -19569
rect -4290 -19757 -4232 -19745
rect -1662 -19577 -1604 -19565
rect -1662 -19753 -1650 -19577
rect -1616 -19753 -1604 -19577
rect -1662 -19765 -1604 -19753
rect -1574 -19577 -1516 -19565
rect -1574 -19753 -1562 -19577
rect -1528 -19753 -1516 -19577
rect -1574 -19765 -1516 -19753
rect 17528 -18631 17928 -18619
rect 17528 -18665 17540 -18631
rect 17916 -18665 17928 -18631
rect 17528 -18681 17928 -18665
rect 18096 -18709 18296 -18697
rect 17528 -18777 17928 -18711
rect 18096 -18743 18108 -18709
rect 18284 -18743 18296 -18709
rect 18096 -18755 18296 -18743
rect 18096 -18797 18296 -18785
rect 17528 -18823 17928 -18807
rect 17528 -18857 17540 -18823
rect 17916 -18857 17928 -18823
rect 18096 -18831 18108 -18797
rect 18284 -18831 18296 -18797
rect 18096 -18843 18296 -18831
rect 17528 -18869 17928 -18857
rect -23894 -20027 -23832 -20015
rect -21168 -20020 -21110 -20008
rect -21168 -20196 -21156 -20020
rect -21122 -20196 -21110 -20020
rect -21168 -20208 -21110 -20196
rect -21080 -20020 -21022 -20008
rect -21080 -20196 -21068 -20020
rect -21034 -20196 -21022 -20020
rect -21080 -20208 -21022 -20196
rect -15577 -19891 -15519 -19879
rect -15577 -20067 -15565 -19891
rect -15531 -20067 -15519 -19891
rect -15577 -20079 -15519 -20067
rect -15489 -19891 -15431 -19879
rect -15489 -20067 -15477 -19891
rect -15443 -20067 -15431 -19891
rect -15489 -20079 -15431 -20067
rect -11274 -19878 -11144 -19866
rect -11274 -19912 -11262 -19878
rect -11156 -19912 -11144 -19878
rect -11274 -19924 -11144 -19912
rect -21168 -20480 -21110 -20468
rect -21168 -20656 -21156 -20480
rect -21122 -20656 -21110 -20480
rect -21168 -20668 -21110 -20656
rect -21080 -20480 -21022 -20468
rect -21080 -20656 -21068 -20480
rect -21034 -20656 -21022 -20480
rect -21080 -20668 -21022 -20656
rect -17188 -20495 -16988 -20483
rect -17188 -20529 -17176 -20495
rect -17000 -20529 -16988 -20495
rect -17188 -20545 -16988 -20529
rect -17188 -20591 -16988 -20575
rect -17188 -20625 -17176 -20591
rect -17000 -20625 -16988 -20591
rect -17188 -20641 -16988 -20625
rect -24051 -20839 -23989 -20827
rect -24051 -21215 -24039 -20839
rect -24005 -21215 -23989 -20839
rect -24051 -21227 -23989 -21215
rect -23959 -21227 -23893 -20827
rect -23863 -20839 -23801 -20827
rect -23863 -21215 -23847 -20839
rect -23813 -21215 -23801 -20839
rect -21182 -20940 -21124 -20928
rect -21182 -21116 -21170 -20940
rect -21136 -21116 -21124 -20940
rect -21182 -21128 -21124 -21116
rect -21094 -20940 -21036 -20928
rect -21094 -21116 -21082 -20940
rect -21048 -21116 -21036 -20940
rect -21094 -21128 -21036 -21116
rect -17188 -20687 -16988 -20671
rect -17188 -20721 -17176 -20687
rect -17000 -20721 -16988 -20687
rect -17188 -20733 -16988 -20721
rect -15577 -20351 -15519 -20339
rect -15577 -20527 -15565 -20351
rect -15531 -20527 -15519 -20351
rect -15577 -20539 -15519 -20527
rect -15489 -20351 -15431 -20339
rect -15489 -20527 -15477 -20351
rect -15443 -20527 -15431 -20351
rect -15489 -20539 -15431 -20527
rect -15591 -20811 -15533 -20799
rect -15591 -20987 -15579 -20811
rect -15545 -20987 -15533 -20811
rect -15591 -20999 -15533 -20987
rect -15503 -20811 -15445 -20799
rect -15503 -20987 -15491 -20811
rect -15457 -20987 -15445 -20811
rect -15503 -20999 -15445 -20987
rect -11274 -19966 -11144 -19954
rect -11274 -20000 -11262 -19966
rect -11156 -20000 -11144 -19966
rect -11274 -20016 -11144 -20000
rect -11274 -20062 -11144 -20046
rect -11274 -20096 -11262 -20062
rect -11156 -20096 -11144 -20062
rect -11274 -20112 -11144 -20096
rect -11274 -20158 -11144 -20142
rect -11274 -20192 -11262 -20158
rect -11156 -20192 -11144 -20158
rect -11274 -20208 -11144 -20192
rect -11274 -20254 -11144 -20238
rect -11274 -20288 -11262 -20254
rect -11156 -20288 -11144 -20254
rect -11274 -20304 -11144 -20288
rect -11274 -20350 -11144 -20334
rect -11274 -20384 -11262 -20350
rect -11156 -20384 -11144 -20350
rect -11274 -20400 -11144 -20384
rect -11274 -20446 -11144 -20430
rect -11274 -20480 -11262 -20446
rect -11156 -20480 -11144 -20446
rect -11274 -20496 -11144 -20480
rect -11274 -20542 -11144 -20526
rect -11274 -20576 -11262 -20542
rect -11156 -20576 -11144 -20542
rect -11274 -20592 -11144 -20576
rect -11274 -20638 -11144 -20622
rect -11274 -20672 -11262 -20638
rect -11156 -20672 -11144 -20638
rect -11274 -20688 -11144 -20672
rect -11274 -20734 -11144 -20718
rect -11274 -20768 -11262 -20734
rect -11156 -20768 -11144 -20734
rect -11274 -20784 -11144 -20768
rect -11274 -20830 -11144 -20814
rect -11274 -20864 -11262 -20830
rect -11156 -20864 -11144 -20830
rect -11274 -20880 -11144 -20864
rect -11274 -20926 -11144 -20910
rect -11274 -20960 -11262 -20926
rect -11156 -20960 -11144 -20926
rect -11274 -20976 -11144 -20960
rect -11274 -21022 -11144 -21006
rect -11274 -21056 -11262 -21022
rect -11156 -21056 -11144 -21022
rect -11274 -21072 -11144 -21056
rect -23863 -21227 -23801 -21215
rect -11274 -21118 -11144 -21102
rect -11274 -21152 -11262 -21118
rect -11156 -21152 -11144 -21118
rect -11274 -21164 -11144 -21152
rect -4378 -19948 -4320 -19936
rect -4378 -20124 -4366 -19948
rect -4332 -20124 -4320 -19948
rect -4378 -20136 -4320 -20124
rect -4290 -19948 -4232 -19936
rect -4290 -20124 -4278 -19948
rect -4244 -20124 -4232 -19948
rect -4290 -20136 -4232 -20124
rect -1662 -19956 -1604 -19944
rect -1662 -20132 -1650 -19956
rect -1616 -20132 -1604 -19956
rect -1662 -20144 -1604 -20132
rect -1574 -19956 -1516 -19944
rect -1574 -20132 -1562 -19956
rect -1528 -20132 -1516 -19956
rect -1574 -20144 -1516 -20132
rect 16147 -19935 16209 -19923
rect 16147 -20111 16159 -19935
rect 16193 -20111 16209 -19935
rect 16147 -20123 16209 -20111
rect 16239 -19935 16305 -19923
rect 16239 -20111 16255 -19935
rect 16289 -20111 16305 -19935
rect 16239 -20123 16305 -20111
rect 16335 -19935 16401 -19923
rect 16335 -20111 16351 -19935
rect 16385 -20111 16401 -19935
rect 16335 -20123 16401 -20111
rect 16431 -19935 16497 -19923
rect 16431 -20111 16447 -19935
rect 16481 -20111 16497 -19935
rect 16431 -20123 16497 -20111
rect 16527 -19935 16589 -19923
rect 16527 -20111 16543 -19935
rect 16577 -20111 16589 -19935
rect 16527 -20123 16589 -20111
rect 7360 -20162 7422 -20150
rect -4378 -20388 -4320 -20376
rect -4378 -20564 -4366 -20388
rect -4332 -20564 -4320 -20388
rect -4378 -20576 -4320 -20564
rect -4290 -20388 -4232 -20376
rect -4290 -20564 -4278 -20388
rect -4244 -20564 -4232 -20388
rect -4290 -20576 -4232 -20564
rect -1662 -20396 -1604 -20384
rect -1662 -20572 -1650 -20396
rect -1616 -20572 -1604 -20396
rect -1662 -20584 -1604 -20572
rect -1574 -20396 -1516 -20384
rect -1574 -20572 -1562 -20396
rect -1528 -20572 -1516 -20396
rect -1574 -20584 -1516 -20572
rect -4378 -20767 -4320 -20755
rect -4378 -20943 -4366 -20767
rect -4332 -20943 -4320 -20767
rect -4378 -20955 -4320 -20943
rect -4290 -20767 -4232 -20755
rect -4290 -20943 -4278 -20767
rect -4244 -20943 -4232 -20767
rect -4290 -20955 -4232 -20943
rect 7360 -20938 7372 -20162
rect 7406 -20938 7422 -20162
rect 7360 -20950 7422 -20938
rect 7452 -20950 7518 -20150
rect 7548 -20950 7614 -20150
rect 7644 -20950 7710 -20150
rect 7740 -20162 7802 -20150
rect 7740 -20938 7756 -20162
rect 7790 -20938 7802 -20162
rect 7740 -20950 7802 -20938
rect 8308 -20162 8370 -20150
rect 8308 -20938 8320 -20162
rect 8354 -20938 8370 -20162
rect 8308 -20950 8370 -20938
rect 8400 -20950 8466 -20150
rect 8496 -20950 8562 -20150
rect 8592 -20950 8658 -20150
rect 8688 -20162 8750 -20150
rect 8688 -20938 8704 -20162
rect 8738 -20938 8750 -20162
rect 8688 -20950 8750 -20938
rect 9244 -20162 9306 -20150
rect 9244 -20938 9256 -20162
rect 9290 -20938 9306 -20162
rect 9244 -20950 9306 -20938
rect 9336 -20950 9402 -20150
rect 9432 -20950 9498 -20150
rect 9528 -20950 9594 -20150
rect 9624 -20162 9686 -20150
rect 9624 -20938 9640 -20162
rect 9674 -20938 9686 -20162
rect 9624 -20950 9686 -20938
rect 10175 -20162 10237 -20150
rect 10175 -20938 10187 -20162
rect 10221 -20938 10237 -20162
rect 10175 -20950 10237 -20938
rect 10267 -20950 10333 -20150
rect 10363 -20950 10429 -20150
rect 10459 -20950 10525 -20150
rect 10555 -20162 10617 -20150
rect 10555 -20938 10571 -20162
rect 10605 -20938 10617 -20162
rect 10555 -20950 10617 -20938
rect 11102 -20162 11164 -20150
rect 11102 -20938 11114 -20162
rect 11148 -20938 11164 -20162
rect 11102 -20950 11164 -20938
rect 11194 -20950 11260 -20150
rect 11290 -20950 11356 -20150
rect 11386 -20950 11452 -20150
rect 11482 -20162 11544 -20150
rect 11482 -20938 11498 -20162
rect 11532 -20938 11544 -20162
rect 11482 -20950 11544 -20938
rect 7360 -21090 7422 -21078
rect -11274 -21206 -11144 -21194
rect -21180 -21420 -21122 -21408
rect -21180 -21596 -21168 -21420
rect -21134 -21596 -21122 -21420
rect -21180 -21608 -21122 -21596
rect -21092 -21420 -21034 -21408
rect -21092 -21596 -21080 -21420
rect -21046 -21596 -21034 -21420
rect -21092 -21608 -21034 -21596
rect -15589 -21291 -15531 -21279
rect -15589 -21467 -15577 -21291
rect -15543 -21467 -15531 -21291
rect -15589 -21479 -15531 -21467
rect -15501 -21291 -15443 -21279
rect -15501 -21467 -15489 -21291
rect -15455 -21467 -15443 -21291
rect -15501 -21479 -15443 -21467
rect -11274 -21240 -11262 -21206
rect -11156 -21240 -11144 -21206
rect -11274 -21252 -11144 -21240
rect 7360 -21866 7372 -21090
rect 7406 -21866 7422 -21090
rect 7360 -21878 7422 -21866
rect 7452 -21878 7518 -21078
rect 7548 -21878 7614 -21078
rect 7644 -21878 7710 -21078
rect 7740 -21090 7802 -21078
rect 7740 -21866 7756 -21090
rect 7790 -21866 7802 -21090
rect 7740 -21878 7802 -21866
rect 8308 -21090 8370 -21078
rect 8308 -21866 8320 -21090
rect 8354 -21866 8370 -21090
rect 8308 -21878 8370 -21866
rect 8400 -21878 8466 -21078
rect 8496 -21878 8562 -21078
rect 8592 -21878 8658 -21078
rect 8688 -21090 8750 -21078
rect 8688 -21866 8704 -21090
rect 8738 -21866 8750 -21090
rect 8688 -21878 8750 -21866
rect 9244 -21090 9306 -21078
rect 9244 -21866 9256 -21090
rect 9290 -21866 9306 -21090
rect 9244 -21878 9306 -21866
rect 9336 -21878 9402 -21078
rect 9432 -21878 9498 -21078
rect 9528 -21878 9594 -21078
rect 9624 -21090 9686 -21078
rect 9624 -21866 9640 -21090
rect 9674 -21866 9686 -21090
rect 9624 -21878 9686 -21866
rect 10175 -21089 10237 -21077
rect 10175 -21865 10187 -21089
rect 10221 -21865 10237 -21089
rect 10175 -21877 10237 -21865
rect 10267 -21877 10333 -21077
rect 10363 -21877 10429 -21077
rect 10459 -21877 10525 -21077
rect 10555 -21089 10617 -21077
rect 10555 -21865 10571 -21089
rect 10605 -21865 10617 -21089
rect 10555 -21877 10617 -21865
rect 11102 -21090 11164 -21078
rect -17188 -21895 -16988 -21883
rect -17188 -21929 -17176 -21895
rect -17000 -21929 -16988 -21895
rect -17188 -21945 -16988 -21929
rect -17188 -21991 -16988 -21975
rect -17188 -22025 -17176 -21991
rect -17000 -22025 -16988 -21991
rect -17188 -22041 -16988 -22025
rect -24052 -22142 -23990 -22130
rect -24052 -22518 -24040 -22142
rect -24006 -22518 -23990 -22142
rect -24052 -22530 -23990 -22518
rect -23960 -22530 -23894 -22130
rect -23864 -22142 -23802 -22130
rect -23864 -22518 -23848 -22142
rect -23814 -22518 -23802 -22142
rect -23864 -22530 -23802 -22518
rect -17188 -22087 -16988 -22071
rect -17188 -22121 -17176 -22087
rect -17000 -22121 -16988 -22087
rect -17188 -22133 -16988 -22121
rect 11102 -21866 11114 -21090
rect 11148 -21866 11164 -21090
rect 11102 -21878 11164 -21866
rect 11194 -21878 11260 -21078
rect 11290 -21878 11356 -21078
rect 11386 -21878 11452 -21078
rect 11482 -21090 11544 -21078
rect 11482 -21866 11498 -21090
rect 11532 -21866 11544 -21090
rect 12157 -21132 12219 -21120
rect 12157 -21308 12169 -21132
rect 12203 -21308 12219 -21132
rect 12157 -21320 12219 -21308
rect 12249 -21132 12315 -21120
rect 12249 -21308 12265 -21132
rect 12299 -21308 12315 -21132
rect 12249 -21320 12315 -21308
rect 12345 -21132 12407 -21120
rect 12345 -21308 12361 -21132
rect 12395 -21308 12407 -21132
rect 12923 -21197 13123 -21185
rect 12923 -21231 12935 -21197
rect 13111 -21231 13123 -21197
rect 12923 -21243 13123 -21231
rect 12923 -21285 13123 -21273
rect 12345 -21320 12407 -21308
rect 12923 -21319 12935 -21285
rect 13111 -21319 13123 -21285
rect 12923 -21331 13123 -21319
rect 11482 -21878 11544 -21866
rect -11274 -22457 -11144 -22445
rect -11274 -22491 -11262 -22457
rect -11156 -22491 -11144 -22457
rect -11274 -22503 -11144 -22491
rect -17188 -23295 -16988 -23283
rect -17188 -23329 -17176 -23295
rect -17000 -23329 -16988 -23295
rect -17188 -23345 -16988 -23329
rect -17188 -23391 -16988 -23375
rect -24052 -23451 -23990 -23439
rect -24052 -23827 -24040 -23451
rect -24006 -23827 -23990 -23451
rect -24052 -23839 -23990 -23827
rect -23960 -23839 -23894 -23439
rect -23864 -23451 -23802 -23439
rect -23864 -23827 -23848 -23451
rect -23814 -23827 -23802 -23451
rect -17188 -23425 -17176 -23391
rect -17000 -23425 -16988 -23391
rect -17188 -23441 -16988 -23425
rect -23864 -23839 -23802 -23827
rect -17188 -23487 -16988 -23471
rect -17188 -23521 -17176 -23487
rect -17000 -23521 -16988 -23487
rect -17188 -23533 -16988 -23521
rect -11274 -22545 -11144 -22533
rect -11274 -22579 -11262 -22545
rect -11156 -22579 -11144 -22545
rect -11274 -22595 -11144 -22579
rect -11274 -22641 -11144 -22625
rect -11274 -22675 -11262 -22641
rect -11156 -22675 -11144 -22641
rect -11274 -22691 -11144 -22675
rect -11274 -22737 -11144 -22721
rect -11274 -22771 -11262 -22737
rect -11156 -22771 -11144 -22737
rect -11274 -22787 -11144 -22771
rect -11274 -22833 -11144 -22817
rect -11274 -22867 -11262 -22833
rect -11156 -22867 -11144 -22833
rect -11274 -22883 -11144 -22867
rect -11274 -22929 -11144 -22913
rect -11274 -22963 -11262 -22929
rect -11156 -22963 -11144 -22929
rect -11274 -22979 -11144 -22963
rect -11274 -23025 -11144 -23009
rect -11274 -23059 -11262 -23025
rect -11156 -23059 -11144 -23025
rect -11274 -23075 -11144 -23059
rect -11274 -23121 -11144 -23105
rect -11274 -23155 -11262 -23121
rect -11156 -23155 -11144 -23121
rect -11274 -23171 -11144 -23155
rect -11274 -23217 -11144 -23201
rect -11274 -23251 -11262 -23217
rect -11156 -23251 -11144 -23217
rect -11274 -23267 -11144 -23251
rect -11274 -23313 -11144 -23297
rect -11274 -23347 -11262 -23313
rect -11156 -23347 -11144 -23313
rect -11274 -23363 -11144 -23347
rect -11274 -23409 -11144 -23393
rect -11274 -23443 -11262 -23409
rect -11156 -23443 -11144 -23409
rect -11274 -23459 -11144 -23443
rect -11274 -23505 -11144 -23489
rect -11274 -23539 -11262 -23505
rect -11156 -23539 -11144 -23505
rect -11274 -23555 -11144 -23539
rect -11274 -23601 -11144 -23585
rect -11274 -23635 -11262 -23601
rect -11156 -23635 -11144 -23601
rect -11274 -23651 -11144 -23635
rect -11274 -23697 -11144 -23681
rect -11274 -23731 -11262 -23697
rect -11156 -23731 -11144 -23697
rect -11274 -23743 -11144 -23731
rect 5658 -23707 5858 -23695
rect -11274 -23785 -11144 -23773
rect -11274 -23819 -11262 -23785
rect -11156 -23819 -11144 -23785
rect 5658 -23741 5670 -23707
rect 5846 -23741 5858 -23707
rect 6098 -23707 6298 -23695
rect 5658 -23753 5858 -23741
rect 5658 -23795 5858 -23783
rect -11274 -23831 -11144 -23819
rect 5658 -23829 5670 -23795
rect 5846 -23829 5858 -23795
rect 6098 -23741 6110 -23707
rect 6286 -23741 6298 -23707
rect 6538 -23707 6738 -23695
rect 6098 -23753 6298 -23741
rect 6098 -23795 6298 -23783
rect 5658 -23841 5858 -23829
rect 6098 -23829 6110 -23795
rect 6286 -23829 6298 -23795
rect 6538 -23741 6550 -23707
rect 6726 -23741 6738 -23707
rect 6538 -23753 6738 -23741
rect 6538 -23795 6738 -23783
rect 6098 -23841 6298 -23829
rect 6538 -23829 6550 -23795
rect 6726 -23829 6738 -23795
rect 6538 -23841 6738 -23829
rect -17188 -24695 -16988 -24683
rect -17188 -24729 -17176 -24695
rect -17000 -24729 -16988 -24695
rect -17188 -24745 -16988 -24729
rect -17188 -24791 -16988 -24775
rect -17188 -24825 -17176 -24791
rect -17000 -24825 -16988 -24791
rect -17188 -24841 -16988 -24825
rect -17188 -24887 -16988 -24871
rect -17188 -24921 -17176 -24887
rect -17000 -24921 -16988 -24887
rect -17188 -24933 -16988 -24921
rect 7360 -24690 7422 -24678
rect -11274 -25225 -11144 -25213
rect -11274 -25259 -11262 -25225
rect -11156 -25259 -11144 -25225
rect -11274 -25271 -11144 -25259
rect -11274 -25313 -11144 -25301
rect -11274 -25347 -11262 -25313
rect -11156 -25347 -11144 -25313
rect -11274 -25363 -11144 -25347
rect -11274 -25409 -11144 -25393
rect -11274 -25443 -11262 -25409
rect -11156 -25443 -11144 -25409
rect -11274 -25459 -11144 -25443
rect -11274 -25505 -11144 -25489
rect -11274 -25539 -11262 -25505
rect -11156 -25539 -11144 -25505
rect -11274 -25555 -11144 -25539
rect -11274 -25601 -11144 -25585
rect -11274 -25635 -11262 -25601
rect -11156 -25635 -11144 -25601
rect -11274 -25651 -11144 -25635
rect -11274 -25697 -11144 -25681
rect -11274 -25731 -11262 -25697
rect -11156 -25731 -11144 -25697
rect -11274 -25747 -11144 -25731
rect -11274 -25793 -11144 -25777
rect -11274 -25827 -11262 -25793
rect -11156 -25827 -11144 -25793
rect -11274 -25843 -11144 -25827
rect -11274 -25889 -11144 -25873
rect -11274 -25923 -11262 -25889
rect -11156 -25923 -11144 -25889
rect -11274 -25939 -11144 -25923
rect -11274 -25985 -11144 -25969
rect -11274 -26019 -11262 -25985
rect -11156 -26019 -11144 -25985
rect -11274 -26035 -11144 -26019
rect -11274 -26081 -11144 -26065
rect -11274 -26115 -11262 -26081
rect -11156 -26115 -11144 -26081
rect -11274 -26131 -11144 -26115
rect -11274 -26177 -11144 -26161
rect -11274 -26211 -11262 -26177
rect -11156 -26211 -11144 -26177
rect -11274 -26227 -11144 -26211
rect -11274 -26273 -11144 -26257
rect -11274 -26307 -11262 -26273
rect -11156 -26307 -11144 -26273
rect -11274 -26323 -11144 -26307
rect -11274 -26369 -11144 -26353
rect -11274 -26403 -11262 -26369
rect -11156 -26403 -11144 -26369
rect -11274 -26419 -11144 -26403
rect -11274 -26465 -11144 -26449
rect -11274 -26499 -11262 -26465
rect -11156 -26499 -11144 -26465
rect -11274 -26511 -11144 -26499
rect 7360 -25466 7372 -24690
rect 7406 -25466 7422 -24690
rect 7360 -25478 7422 -25466
rect 7452 -25478 7518 -24678
rect 7548 -25478 7614 -24678
rect 7644 -25478 7710 -24678
rect 7740 -24690 7802 -24678
rect 7740 -25466 7756 -24690
rect 7790 -25466 7802 -24690
rect 7740 -25478 7802 -25466
rect 8308 -24690 8370 -24678
rect 8308 -25466 8320 -24690
rect 8354 -25466 8370 -24690
rect 8308 -25478 8370 -25466
rect 8400 -25478 8466 -24678
rect 8496 -25478 8562 -24678
rect 8592 -25478 8658 -24678
rect 8688 -24690 8750 -24678
rect 8688 -25466 8704 -24690
rect 8738 -25466 8750 -24690
rect 8688 -25478 8750 -25466
rect 9244 -24690 9306 -24678
rect 9244 -25466 9256 -24690
rect 9290 -25466 9306 -24690
rect 9244 -25478 9306 -25466
rect 9336 -25478 9402 -24678
rect 9432 -25478 9498 -24678
rect 9528 -25478 9594 -24678
rect 9624 -24690 9686 -24678
rect 9624 -25466 9640 -24690
rect 9674 -25466 9686 -24690
rect 9624 -25478 9686 -25466
rect 10175 -24690 10237 -24678
rect 10175 -25466 10187 -24690
rect 10221 -25466 10237 -24690
rect 10175 -25478 10237 -25466
rect 10267 -25478 10333 -24678
rect 10363 -25478 10429 -24678
rect 10459 -25478 10525 -24678
rect 10555 -24690 10617 -24678
rect 10555 -25466 10571 -24690
rect 10605 -25466 10617 -24690
rect 10555 -25478 10617 -25466
rect 11102 -24690 11164 -24678
rect 11102 -25466 11114 -24690
rect 11148 -25466 11164 -24690
rect 11102 -25478 11164 -25466
rect 11194 -25478 11260 -24678
rect 11290 -25478 11356 -24678
rect 11386 -25478 11452 -24678
rect 11482 -24690 11544 -24678
rect 11482 -25466 11498 -24690
rect 11532 -25466 11544 -24690
rect 11482 -25478 11544 -25466
rect 7360 -25618 7422 -25606
rect 7360 -26394 7372 -25618
rect 7406 -26394 7422 -25618
rect 7360 -26406 7422 -26394
rect 7452 -26406 7518 -25606
rect 7548 -26406 7614 -25606
rect 7644 -26406 7710 -25606
rect 7740 -25618 7802 -25606
rect 7740 -26394 7756 -25618
rect 7790 -26394 7802 -25618
rect 7740 -26406 7802 -26394
rect 8308 -25618 8370 -25606
rect 8308 -26394 8320 -25618
rect 8354 -26394 8370 -25618
rect 8308 -26406 8370 -26394
rect 8400 -26406 8466 -25606
rect 8496 -26406 8562 -25606
rect 8592 -26406 8658 -25606
rect 8688 -25618 8750 -25606
rect 8688 -26394 8704 -25618
rect 8738 -26394 8750 -25618
rect 8688 -26406 8750 -26394
rect 9244 -25618 9306 -25606
rect 9244 -26394 9256 -25618
rect 9290 -26394 9306 -25618
rect 9244 -26406 9306 -26394
rect 9336 -26406 9402 -25606
rect 9432 -26406 9498 -25606
rect 9528 -26406 9594 -25606
rect 9624 -25618 9686 -25606
rect 9624 -26394 9640 -25618
rect 9674 -26394 9686 -25618
rect 9624 -26406 9686 -26394
rect 10175 -25617 10237 -25605
rect 10175 -26393 10187 -25617
rect 10221 -26393 10237 -25617
rect 10175 -26405 10237 -26393
rect 10267 -26405 10333 -25605
rect 10363 -26405 10429 -25605
rect 10459 -26405 10525 -25605
rect 10555 -25617 10617 -25605
rect 10555 -26393 10571 -25617
rect 10605 -26393 10617 -25617
rect 10555 -26405 10617 -26393
rect 11102 -25618 11164 -25606
rect -11274 -26553 -11144 -26541
rect -11274 -26587 -11262 -26553
rect -11156 -26587 -11144 -26553
rect -11274 -26599 -11144 -26587
rect 11102 -26394 11114 -25618
rect 11148 -26394 11164 -25618
rect 11102 -26406 11164 -26394
rect 11194 -26406 11260 -25606
rect 11290 -26406 11356 -25606
rect 11386 -26406 11452 -25606
rect 11482 -25618 11544 -25606
rect 11482 -26394 11498 -25618
rect 11532 -26394 11544 -25618
rect 12157 -25660 12219 -25648
rect 12157 -25836 12169 -25660
rect 12203 -25836 12219 -25660
rect 12157 -25848 12219 -25836
rect 12249 -25660 12315 -25648
rect 12249 -25836 12265 -25660
rect 12299 -25836 12315 -25660
rect 12249 -25848 12315 -25836
rect 12345 -25660 12407 -25648
rect 12345 -25836 12361 -25660
rect 12395 -25836 12407 -25660
rect 12923 -25725 13123 -25713
rect 12923 -25759 12935 -25725
rect 13111 -25759 13123 -25725
rect 12923 -25771 13123 -25759
rect 12923 -25813 13123 -25801
rect 12345 -25848 12407 -25836
rect 12923 -25847 12935 -25813
rect 13111 -25847 13123 -25813
rect 12923 -25859 13123 -25847
rect 11482 -26406 11544 -26394
rect -11274 -27858 -11144 -27846
rect -11274 -27892 -11262 -27858
rect -11156 -27892 -11144 -27858
rect -11274 -27904 -11144 -27892
rect -11274 -27946 -11144 -27934
rect -11274 -27980 -11262 -27946
rect -11156 -27980 -11144 -27946
rect -11274 -27996 -11144 -27980
rect -11274 -28042 -11144 -28026
rect -11274 -28076 -11262 -28042
rect -11156 -28076 -11144 -28042
rect -11274 -28092 -11144 -28076
rect -11274 -28138 -11144 -28122
rect -11274 -28172 -11262 -28138
rect -11156 -28172 -11144 -28138
rect -11274 -28188 -11144 -28172
rect -11274 -28234 -11144 -28218
rect -11274 -28268 -11262 -28234
rect -11156 -28268 -11144 -28234
rect -11274 -28284 -11144 -28268
rect -11274 -28330 -11144 -28314
rect -11274 -28364 -11262 -28330
rect -11156 -28364 -11144 -28330
rect -11274 -28380 -11144 -28364
rect -11274 -28426 -11144 -28410
rect -11274 -28460 -11262 -28426
rect -11156 -28460 -11144 -28426
rect -11274 -28476 -11144 -28460
rect -11274 -28522 -11144 -28506
rect -11274 -28556 -11262 -28522
rect -11156 -28556 -11144 -28522
rect -11274 -28572 -11144 -28556
rect -11274 -28618 -11144 -28602
rect -11274 -28652 -11262 -28618
rect -11156 -28652 -11144 -28618
rect -11274 -28668 -11144 -28652
rect -11274 -28714 -11144 -28698
rect -11274 -28748 -11262 -28714
rect -11156 -28748 -11144 -28714
rect -11274 -28764 -11144 -28748
rect -11274 -28810 -11144 -28794
rect -11274 -28844 -11262 -28810
rect -11156 -28844 -11144 -28810
rect -11274 -28860 -11144 -28844
rect -11274 -28906 -11144 -28890
rect -11274 -28940 -11262 -28906
rect -11156 -28940 -11144 -28906
rect -11274 -28956 -11144 -28940
rect -11274 -29002 -11144 -28986
rect -11274 -29036 -11262 -29002
rect -11156 -29036 -11144 -29002
rect -11274 -29052 -11144 -29036
rect -11274 -29098 -11144 -29082
rect -11274 -29132 -11262 -29098
rect -11156 -29132 -11144 -29098
rect -11274 -29144 -11144 -29132
rect 5658 -28235 5858 -28223
rect 5658 -28269 5670 -28235
rect 5846 -28269 5858 -28235
rect 6098 -28235 6298 -28223
rect 5658 -28281 5858 -28269
rect 5658 -28323 5858 -28311
rect 5658 -28357 5670 -28323
rect 5846 -28357 5858 -28323
rect 6098 -28269 6110 -28235
rect 6286 -28269 6298 -28235
rect 6538 -28235 6738 -28223
rect 6098 -28281 6298 -28269
rect 6098 -28323 6298 -28311
rect 5658 -28369 5858 -28357
rect 6098 -28357 6110 -28323
rect 6286 -28357 6298 -28323
rect 6538 -28269 6550 -28235
rect 6726 -28269 6738 -28235
rect 6538 -28281 6738 -28269
rect 6538 -28323 6738 -28311
rect 6098 -28369 6298 -28357
rect 6538 -28357 6550 -28323
rect 6726 -28357 6738 -28323
rect 6538 -28369 6738 -28357
rect -11274 -29186 -11144 -29174
rect -11274 -29220 -11262 -29186
rect -11156 -29220 -11144 -29186
rect -11274 -29232 -11144 -29220
rect 7360 -29218 7422 -29206
rect 7360 -29994 7372 -29218
rect 7406 -29994 7422 -29218
rect 7360 -30006 7422 -29994
rect 7452 -30006 7518 -29206
rect 7548 -30006 7614 -29206
rect 7644 -30006 7710 -29206
rect 7740 -29218 7802 -29206
rect 7740 -29994 7756 -29218
rect 7790 -29994 7802 -29218
rect 7740 -30006 7802 -29994
rect 8308 -29218 8370 -29206
rect 8308 -29994 8320 -29218
rect 8354 -29994 8370 -29218
rect 8308 -30006 8370 -29994
rect 8400 -30006 8466 -29206
rect 8496 -30006 8562 -29206
rect 8592 -30006 8658 -29206
rect 8688 -29218 8750 -29206
rect 8688 -29994 8704 -29218
rect 8738 -29994 8750 -29218
rect 8688 -30006 8750 -29994
rect 9244 -29218 9306 -29206
rect 9244 -29994 9256 -29218
rect 9290 -29994 9306 -29218
rect 9244 -30006 9306 -29994
rect 9336 -30006 9402 -29206
rect 9432 -30006 9498 -29206
rect 9528 -30006 9594 -29206
rect 9624 -29218 9686 -29206
rect 9624 -29994 9640 -29218
rect 9674 -29994 9686 -29218
rect 9624 -30006 9686 -29994
rect 10175 -29218 10237 -29206
rect 10175 -29994 10187 -29218
rect 10221 -29994 10237 -29218
rect 10175 -30006 10237 -29994
rect 10267 -30006 10333 -29206
rect 10363 -30006 10429 -29206
rect 10459 -30006 10525 -29206
rect 10555 -29218 10617 -29206
rect 10555 -29994 10571 -29218
rect 10605 -29994 10617 -29218
rect 10555 -30006 10617 -29994
rect 11102 -29218 11164 -29206
rect 11102 -29994 11114 -29218
rect 11148 -29994 11164 -29218
rect 11102 -30006 11164 -29994
rect 11194 -30006 11260 -29206
rect 11290 -30006 11356 -29206
rect 11386 -30006 11452 -29206
rect 11482 -29218 11544 -29206
rect 11482 -29994 11498 -29218
rect 11532 -29994 11544 -29218
rect 11482 -30006 11544 -29994
rect 7360 -30146 7422 -30134
rect -11274 -30467 -11144 -30455
rect -11274 -30501 -11262 -30467
rect -11156 -30501 -11144 -30467
rect -11274 -30513 -11144 -30501
rect -11274 -30555 -11144 -30543
rect -11274 -30589 -11262 -30555
rect -11156 -30589 -11144 -30555
rect -11274 -30605 -11144 -30589
rect -11274 -30651 -11144 -30635
rect -11274 -30685 -11262 -30651
rect -11156 -30685 -11144 -30651
rect -11274 -30701 -11144 -30685
rect -11274 -30747 -11144 -30731
rect -11274 -30781 -11262 -30747
rect -11156 -30781 -11144 -30747
rect -11274 -30797 -11144 -30781
rect -11274 -30843 -11144 -30827
rect -11274 -30877 -11262 -30843
rect -11156 -30877 -11144 -30843
rect -11274 -30893 -11144 -30877
rect -11274 -30939 -11144 -30923
rect -11274 -30973 -11262 -30939
rect -11156 -30973 -11144 -30939
rect -11274 -30989 -11144 -30973
rect -11274 -31035 -11144 -31019
rect -11274 -31069 -11262 -31035
rect -11156 -31069 -11144 -31035
rect -11274 -31085 -11144 -31069
rect -11274 -31131 -11144 -31115
rect -11274 -31165 -11262 -31131
rect -11156 -31165 -11144 -31131
rect -11274 -31181 -11144 -31165
rect -11274 -31227 -11144 -31211
rect -11274 -31261 -11262 -31227
rect -11156 -31261 -11144 -31227
rect -11274 -31277 -11144 -31261
rect -11274 -31323 -11144 -31307
rect -11274 -31357 -11262 -31323
rect -11156 -31357 -11144 -31323
rect -11274 -31373 -11144 -31357
rect -11274 -31419 -11144 -31403
rect -11274 -31453 -11262 -31419
rect -11156 -31453 -11144 -31419
rect -11274 -31469 -11144 -31453
rect -11274 -31515 -11144 -31499
rect -11274 -31549 -11262 -31515
rect -11156 -31549 -11144 -31515
rect -11274 -31565 -11144 -31549
rect -11274 -31611 -11144 -31595
rect -11274 -31645 -11262 -31611
rect -11156 -31645 -11144 -31611
rect -11274 -31661 -11144 -31645
rect -11274 -31707 -11144 -31691
rect -11274 -31741 -11262 -31707
rect -11156 -31741 -11144 -31707
rect -11274 -31753 -11144 -31741
rect 7360 -30922 7372 -30146
rect 7406 -30922 7422 -30146
rect 7360 -30934 7422 -30922
rect 7452 -30934 7518 -30134
rect 7548 -30934 7614 -30134
rect 7644 -30934 7710 -30134
rect 7740 -30146 7802 -30134
rect 7740 -30922 7756 -30146
rect 7790 -30922 7802 -30146
rect 7740 -30934 7802 -30922
rect 8308 -30146 8370 -30134
rect 8308 -30922 8320 -30146
rect 8354 -30922 8370 -30146
rect 8308 -30934 8370 -30922
rect 8400 -30934 8466 -30134
rect 8496 -30934 8562 -30134
rect 8592 -30934 8658 -30134
rect 8688 -30146 8750 -30134
rect 8688 -30922 8704 -30146
rect 8738 -30922 8750 -30146
rect 8688 -30934 8750 -30922
rect 9244 -30146 9306 -30134
rect 9244 -30922 9256 -30146
rect 9290 -30922 9306 -30146
rect 9244 -30934 9306 -30922
rect 9336 -30934 9402 -30134
rect 9432 -30934 9498 -30134
rect 9528 -30934 9594 -30134
rect 9624 -30146 9686 -30134
rect 9624 -30922 9640 -30146
rect 9674 -30922 9686 -30146
rect 9624 -30934 9686 -30922
rect 10175 -30145 10237 -30133
rect 10175 -30921 10187 -30145
rect 10221 -30921 10237 -30145
rect 10175 -30933 10237 -30921
rect 10267 -30933 10333 -30133
rect 10363 -30933 10429 -30133
rect 10459 -30933 10525 -30133
rect 10555 -30145 10617 -30133
rect 10555 -30921 10571 -30145
rect 10605 -30921 10617 -30145
rect 10555 -30933 10617 -30921
rect 11102 -30146 11164 -30134
rect 11102 -30922 11114 -30146
rect 11148 -30922 11164 -30146
rect 11102 -30934 11164 -30922
rect 11194 -30934 11260 -30134
rect 11290 -30934 11356 -30134
rect 11386 -30934 11452 -30134
rect 11482 -30146 11544 -30134
rect 11482 -30922 11498 -30146
rect 11532 -30922 11544 -30146
rect 12157 -30188 12219 -30176
rect 12157 -30364 12169 -30188
rect 12203 -30364 12219 -30188
rect 12157 -30376 12219 -30364
rect 12249 -30188 12315 -30176
rect 12249 -30364 12265 -30188
rect 12299 -30364 12315 -30188
rect 12249 -30376 12315 -30364
rect 12345 -30188 12407 -30176
rect 12345 -30364 12361 -30188
rect 12395 -30364 12407 -30188
rect 12923 -30253 13123 -30241
rect 12923 -30287 12935 -30253
rect 13111 -30287 13123 -30253
rect 12923 -30299 13123 -30287
rect 12923 -30341 13123 -30329
rect 12345 -30376 12407 -30364
rect 12923 -30375 12935 -30341
rect 13111 -30375 13123 -30341
rect 12923 -30387 13123 -30375
rect 11482 -30934 11544 -30922
rect -11274 -31795 -11144 -31783
rect -11274 -31829 -11262 -31795
rect -11156 -31829 -11144 -31795
rect -11274 -31841 -11144 -31829
rect 5658 -32763 5858 -32751
rect 5658 -32797 5670 -32763
rect 5846 -32797 5858 -32763
rect 6098 -32763 6298 -32751
rect 5658 -32809 5858 -32797
rect 5658 -32851 5858 -32839
rect 5658 -32885 5670 -32851
rect 5846 -32885 5858 -32851
rect 6098 -32797 6110 -32763
rect 6286 -32797 6298 -32763
rect 6538 -32763 6738 -32751
rect 6098 -32809 6298 -32797
rect 6098 -32851 6298 -32839
rect 5658 -32897 5858 -32885
rect 6098 -32885 6110 -32851
rect 6286 -32885 6298 -32851
rect 6538 -32797 6550 -32763
rect 6726 -32797 6738 -32763
rect 6538 -32809 6738 -32797
rect 6538 -32851 6738 -32839
rect 6098 -32897 6298 -32885
rect 6538 -32885 6550 -32851
rect 6726 -32885 6738 -32851
rect 6538 -32897 6738 -32885
rect -11276 -33087 -11146 -33075
rect -11276 -33121 -11264 -33087
rect -11158 -33121 -11146 -33087
rect -11276 -33133 -11146 -33121
rect -11276 -33175 -11146 -33163
rect -11276 -33209 -11264 -33175
rect -11158 -33209 -11146 -33175
rect -11276 -33225 -11146 -33209
rect -11276 -33271 -11146 -33255
rect -11276 -33305 -11264 -33271
rect -11158 -33305 -11146 -33271
rect -11276 -33321 -11146 -33305
rect -11276 -33367 -11146 -33351
rect -11276 -33401 -11264 -33367
rect -11158 -33401 -11146 -33367
rect -11276 -33417 -11146 -33401
rect -11276 -33463 -11146 -33447
rect -11276 -33497 -11264 -33463
rect -11158 -33497 -11146 -33463
rect -11276 -33513 -11146 -33497
rect -11276 -33559 -11146 -33543
rect -11276 -33593 -11264 -33559
rect -11158 -33593 -11146 -33559
rect -11276 -33609 -11146 -33593
rect -11276 -33655 -11146 -33639
rect -11276 -33689 -11264 -33655
rect -11158 -33689 -11146 -33655
rect -11276 -33705 -11146 -33689
rect -11276 -33751 -11146 -33735
rect -11276 -33785 -11264 -33751
rect -11158 -33785 -11146 -33751
rect -11276 -33801 -11146 -33785
rect -11276 -33847 -11146 -33831
rect -11276 -33881 -11264 -33847
rect -11158 -33881 -11146 -33847
rect -11276 -33897 -11146 -33881
rect -11276 -33943 -11146 -33927
rect -11276 -33977 -11264 -33943
rect -11158 -33977 -11146 -33943
rect -11276 -33993 -11146 -33977
rect -11276 -34039 -11146 -34023
rect -11276 -34073 -11264 -34039
rect -11158 -34073 -11146 -34039
rect -11276 -34089 -11146 -34073
rect -11276 -34135 -11146 -34119
rect -11276 -34169 -11264 -34135
rect -11158 -34169 -11146 -34135
rect -11276 -34185 -11146 -34169
rect -11276 -34231 -11146 -34215
rect -11276 -34265 -11264 -34231
rect -11158 -34265 -11146 -34231
rect -11276 -34281 -11146 -34265
rect -11276 -34327 -11146 -34311
rect -11276 -34361 -11264 -34327
rect -11158 -34361 -11146 -34327
rect -11276 -34373 -11146 -34361
rect 7360 -33746 7422 -33734
rect -11276 -34415 -11146 -34403
rect -11276 -34449 -11264 -34415
rect -11158 -34449 -11146 -34415
rect -11276 -34461 -11146 -34449
rect 7360 -34522 7372 -33746
rect 7406 -34522 7422 -33746
rect 7360 -34534 7422 -34522
rect 7452 -34534 7518 -33734
rect 7548 -34534 7614 -33734
rect 7644 -34534 7710 -33734
rect 7740 -33746 7802 -33734
rect 7740 -34522 7756 -33746
rect 7790 -34522 7802 -33746
rect 7740 -34534 7802 -34522
rect 8308 -33746 8370 -33734
rect 8308 -34522 8320 -33746
rect 8354 -34522 8370 -33746
rect 8308 -34534 8370 -34522
rect 8400 -34534 8466 -33734
rect 8496 -34534 8562 -33734
rect 8592 -34534 8658 -33734
rect 8688 -33746 8750 -33734
rect 8688 -34522 8704 -33746
rect 8738 -34522 8750 -33746
rect 8688 -34534 8750 -34522
rect 9244 -33746 9306 -33734
rect 9244 -34522 9256 -33746
rect 9290 -34522 9306 -33746
rect 9244 -34534 9306 -34522
rect 9336 -34534 9402 -33734
rect 9432 -34534 9498 -33734
rect 9528 -34534 9594 -33734
rect 9624 -33746 9686 -33734
rect 9624 -34522 9640 -33746
rect 9674 -34522 9686 -33746
rect 9624 -34534 9686 -34522
rect 10175 -33746 10237 -33734
rect 10175 -34522 10187 -33746
rect 10221 -34522 10237 -33746
rect 10175 -34534 10237 -34522
rect 10267 -34534 10333 -33734
rect 10363 -34534 10429 -33734
rect 10459 -34534 10525 -33734
rect 10555 -33746 10617 -33734
rect 10555 -34522 10571 -33746
rect 10605 -34522 10617 -33746
rect 10555 -34534 10617 -34522
rect 11102 -33746 11164 -33734
rect 11102 -34522 11114 -33746
rect 11148 -34522 11164 -33746
rect 11102 -34534 11164 -34522
rect 11194 -34534 11260 -33734
rect 11290 -34534 11356 -33734
rect 11386 -34534 11452 -33734
rect 11482 -33746 11544 -33734
rect 11482 -34522 11498 -33746
rect 11532 -34522 11544 -33746
rect 11482 -34534 11544 -34522
rect 7360 -34674 7422 -34662
rect 7360 -35450 7372 -34674
rect 7406 -35450 7422 -34674
rect 7360 -35462 7422 -35450
rect 7452 -35462 7518 -34662
rect 7548 -35462 7614 -34662
rect 7644 -35462 7710 -34662
rect 7740 -34674 7802 -34662
rect 7740 -35450 7756 -34674
rect 7790 -35450 7802 -34674
rect 7740 -35462 7802 -35450
rect 8308 -34674 8370 -34662
rect 8308 -35450 8320 -34674
rect 8354 -35450 8370 -34674
rect 8308 -35462 8370 -35450
rect 8400 -35462 8466 -34662
rect 8496 -35462 8562 -34662
rect 8592 -35462 8658 -34662
rect 8688 -34674 8750 -34662
rect 8688 -35450 8704 -34674
rect 8738 -35450 8750 -34674
rect 8688 -35462 8750 -35450
rect 9244 -34674 9306 -34662
rect 9244 -35450 9256 -34674
rect 9290 -35450 9306 -34674
rect 9244 -35462 9306 -35450
rect 9336 -35462 9402 -34662
rect 9432 -35462 9498 -34662
rect 9528 -35462 9594 -34662
rect 9624 -34674 9686 -34662
rect 9624 -35450 9640 -34674
rect 9674 -35450 9686 -34674
rect 9624 -35462 9686 -35450
rect 10175 -34673 10237 -34661
rect 10175 -35449 10187 -34673
rect 10221 -35449 10237 -34673
rect 10175 -35461 10237 -35449
rect 10267 -35461 10333 -34661
rect 10363 -35461 10429 -34661
rect 10459 -35461 10525 -34661
rect 10555 -34673 10617 -34661
rect 10555 -35449 10571 -34673
rect 10605 -35449 10617 -34673
rect 10555 -35461 10617 -35449
rect 11102 -34674 11164 -34662
rect 11102 -35450 11114 -34674
rect 11148 -35450 11164 -34674
rect 11102 -35462 11164 -35450
rect 11194 -35462 11260 -34662
rect 11290 -35462 11356 -34662
rect 11386 -35462 11452 -34662
rect 11482 -34674 11544 -34662
rect 11482 -35450 11498 -34674
rect 11532 -35450 11544 -34674
rect 12157 -34716 12219 -34704
rect 12157 -34892 12169 -34716
rect 12203 -34892 12219 -34716
rect 12157 -34904 12219 -34892
rect 12249 -34716 12315 -34704
rect 12249 -34892 12265 -34716
rect 12299 -34892 12315 -34716
rect 12249 -34904 12315 -34892
rect 12345 -34716 12407 -34704
rect 12345 -34892 12361 -34716
rect 12395 -34892 12407 -34716
rect 12923 -34781 13123 -34769
rect 12923 -34815 12935 -34781
rect 13111 -34815 13123 -34781
rect 12923 -34827 13123 -34815
rect 12923 -34869 13123 -34857
rect 12345 -34904 12407 -34892
rect 12923 -34903 12935 -34869
rect 13111 -34903 13123 -34869
rect 12923 -34915 13123 -34903
rect 11482 -35462 11544 -35450
rect 12874 -35727 12932 -35715
rect 12874 -35903 12886 -35727
rect 12920 -35903 12932 -35727
rect 12874 -35915 12932 -35903
rect 12962 -35727 13020 -35715
rect 12962 -35903 12974 -35727
rect 13008 -35903 13020 -35727
rect 12962 -35915 13020 -35903
rect 12874 -36106 12932 -36094
rect 12874 -36282 12886 -36106
rect 12920 -36282 12932 -36106
rect 12874 -36294 12932 -36282
rect 12962 -36106 13020 -36094
rect 12962 -36282 12974 -36106
rect 13008 -36282 13020 -36106
rect 12962 -36294 13020 -36282
<< pdiff >>
rect 1707 6072 1765 6084
rect 1707 5546 1719 6072
rect 1753 5546 1765 6072
rect 1707 5534 1765 5546
rect 1795 6072 1857 6084
rect 1795 5546 1807 6072
rect 1841 5546 1857 6072
rect 1795 5534 1857 5546
rect 1887 6072 1953 6084
rect 1887 5546 1903 6072
rect 1937 5546 1953 6072
rect 1887 5534 1953 5546
rect 1983 6072 2049 6084
rect 1983 5546 1999 6072
rect 2033 5546 2049 6072
rect 1983 5534 2049 5546
rect 2079 6072 2145 6084
rect 2079 5546 2095 6072
rect 2129 5546 2145 6072
rect 2079 5534 2145 5546
rect 2175 6072 2241 6084
rect 2175 5546 2191 6072
rect 2225 5546 2241 6072
rect 2175 5534 2241 5546
rect 2271 6072 2337 6084
rect 2271 5546 2287 6072
rect 2321 5546 2337 6072
rect 2271 5534 2337 5546
rect 2367 6072 2433 6084
rect 2367 5546 2383 6072
rect 2417 5546 2433 6072
rect 2367 5534 2433 5546
rect 2463 6072 2529 6084
rect 2463 5546 2479 6072
rect 2513 5546 2529 6072
rect 2463 5534 2529 5546
rect 2559 6072 2625 6084
rect 2559 5546 2575 6072
rect 2609 5546 2625 6072
rect 2559 5534 2625 5546
rect 2655 6072 2721 6084
rect 2655 5546 2671 6072
rect 2705 5546 2721 6072
rect 2655 5534 2721 5546
rect 2751 6072 2817 6084
rect 2751 5546 2767 6072
rect 2801 5546 2817 6072
rect 2751 5534 2817 5546
rect 2847 6072 2913 6084
rect 2847 5546 2863 6072
rect 2897 5546 2913 6072
rect 2847 5534 2913 5546
rect 2943 6072 3005 6084
rect 2943 5546 2959 6072
rect 2993 5546 3005 6072
rect 2943 5534 3005 5546
rect 3035 6072 3093 6084
rect 3035 5546 3047 6072
rect 3081 5546 3093 6072
rect 3035 5534 3093 5546
rect 3313 6072 3371 6084
rect 3313 5546 3325 6072
rect 3359 5546 3371 6072
rect 3313 5534 3371 5546
rect 3401 6072 3463 6084
rect 3401 5546 3413 6072
rect 3447 5546 3463 6072
rect 3401 5534 3463 5546
rect 3493 6072 3559 6084
rect 3493 5546 3509 6072
rect 3543 5546 3559 6072
rect 3493 5534 3559 5546
rect 3589 6072 3655 6084
rect 3589 5546 3605 6072
rect 3639 5546 3655 6072
rect 3589 5534 3655 5546
rect 3685 6072 3751 6084
rect 3685 5546 3701 6072
rect 3735 5546 3751 6072
rect 3685 5534 3751 5546
rect 3781 6072 3847 6084
rect 3781 5546 3797 6072
rect 3831 5546 3847 6072
rect 3781 5534 3847 5546
rect 3877 6072 3943 6084
rect 3877 5546 3893 6072
rect 3927 5546 3943 6072
rect 3877 5534 3943 5546
rect 3973 6072 4039 6084
rect 3973 5546 3989 6072
rect 4023 5546 4039 6072
rect 3973 5534 4039 5546
rect 4069 6072 4135 6084
rect 4069 5546 4085 6072
rect 4119 5546 4135 6072
rect 4069 5534 4135 5546
rect 4165 6072 4231 6084
rect 4165 5546 4181 6072
rect 4215 5546 4231 6072
rect 4165 5534 4231 5546
rect 4261 6072 4327 6084
rect 4261 5546 4277 6072
rect 4311 5546 4327 6072
rect 4261 5534 4327 5546
rect 4357 6072 4423 6084
rect 4357 5546 4373 6072
rect 4407 5546 4423 6072
rect 4357 5534 4423 5546
rect 4453 6072 4519 6084
rect 4453 5546 4469 6072
rect 4503 5546 4519 6072
rect 4453 5534 4519 5546
rect 4549 6072 4611 6084
rect 4549 5546 4565 6072
rect 4599 5546 4611 6072
rect 4549 5534 4611 5546
rect 4641 6072 4699 6084
rect 4641 5546 4653 6072
rect 4687 5546 4699 6072
rect 4641 5534 4699 5546
rect 5017 6070 5075 6082
rect 5017 5544 5029 6070
rect 5063 5544 5075 6070
rect 5017 5532 5075 5544
rect 5105 6070 5167 6082
rect 5105 5544 5117 6070
rect 5151 5544 5167 6070
rect 5105 5532 5167 5544
rect 5197 6070 5263 6082
rect 5197 5544 5213 6070
rect 5247 5544 5263 6070
rect 5197 5532 5263 5544
rect 5293 6070 5359 6082
rect 5293 5544 5309 6070
rect 5343 5544 5359 6070
rect 5293 5532 5359 5544
rect 5389 6070 5455 6082
rect 5389 5544 5405 6070
rect 5439 5544 5455 6070
rect 5389 5532 5455 5544
rect 5485 6070 5551 6082
rect 5485 5544 5501 6070
rect 5535 5544 5551 6070
rect 5485 5532 5551 5544
rect 5581 6070 5647 6082
rect 5581 5544 5597 6070
rect 5631 5544 5647 6070
rect 5581 5532 5647 5544
rect 5677 6070 5743 6082
rect 5677 5544 5693 6070
rect 5727 5544 5743 6070
rect 5677 5532 5743 5544
rect 5773 6070 5839 6082
rect 5773 5544 5789 6070
rect 5823 5544 5839 6070
rect 5773 5532 5839 5544
rect 5869 6070 5935 6082
rect 5869 5544 5885 6070
rect 5919 5544 5935 6070
rect 5869 5532 5935 5544
rect 5965 6070 6031 6082
rect 5965 5544 5981 6070
rect 6015 5544 6031 6070
rect 5965 5532 6031 5544
rect 6061 6070 6127 6082
rect 6061 5544 6077 6070
rect 6111 5544 6127 6070
rect 6061 5532 6127 5544
rect 6157 6070 6223 6082
rect 6157 5544 6173 6070
rect 6207 5544 6223 6070
rect 6157 5532 6223 5544
rect 6253 6070 6315 6082
rect 6253 5544 6269 6070
rect 6303 5544 6315 6070
rect 6253 5532 6315 5544
rect 6345 6070 6403 6082
rect 6345 5544 6357 6070
rect 6391 5544 6403 6070
rect 6345 5532 6403 5544
rect 7809 5459 8023 5471
rect 6939 5429 7001 5441
rect 6939 5239 6951 5429
rect 6985 5239 7001 5429
rect 6939 5227 7001 5239
rect 7031 5429 7097 5441
rect 7031 5239 7047 5429
rect 7081 5239 7097 5429
rect 7031 5227 7097 5239
rect 7127 5429 7193 5441
rect 7127 5239 7143 5429
rect 7177 5239 7193 5429
rect 7127 5227 7193 5239
rect 7223 5429 7289 5441
rect 7223 5239 7239 5429
rect 7273 5239 7289 5429
rect 7223 5227 7289 5239
rect 7319 5429 7385 5441
rect 7319 5239 7335 5429
rect 7369 5239 7385 5429
rect 7319 5227 7385 5239
rect 7415 5429 7481 5441
rect 7415 5239 7431 5429
rect 7465 5239 7481 5429
rect 7415 5227 7481 5239
rect 7511 5429 7573 5441
rect 7511 5239 7527 5429
rect 7561 5239 7573 5429
rect 7511 5227 7573 5239
rect 7809 5425 7821 5459
rect 8011 5425 8023 5459
rect 7809 5409 8023 5425
rect 7809 5363 8023 5379
rect 7809 5329 7821 5363
rect 8015 5329 8023 5363
rect 7809 5313 8023 5329
rect 7809 5267 8023 5283
rect 7809 5233 7821 5267
rect 8011 5233 8023 5267
rect 7809 5217 8023 5233
rect 7809 5171 8023 5187
rect 7809 5137 7821 5171
rect 8015 5137 8023 5171
rect 7809 5125 8023 5137
rect -24130 4348 -24072 4360
rect -24130 3822 -24118 4348
rect -24084 3822 -24072 4348
rect -24130 3810 -24072 3822
rect -24042 4348 -23980 4360
rect -24042 3822 -24030 4348
rect -23996 3822 -23980 4348
rect -24042 3810 -23980 3822
rect -23950 4348 -23884 4360
rect -23950 3822 -23934 4348
rect -23900 3822 -23884 4348
rect -23950 3810 -23884 3822
rect -23854 4348 -23788 4360
rect -23854 3822 -23838 4348
rect -23804 3822 -23788 4348
rect -23854 3810 -23788 3822
rect -23758 4348 -23692 4360
rect -23758 3822 -23742 4348
rect -23708 3822 -23692 4348
rect -23758 3810 -23692 3822
rect -23662 4348 -23596 4360
rect -23662 3822 -23646 4348
rect -23612 3822 -23596 4348
rect -23662 3810 -23596 3822
rect -23566 4348 -23500 4360
rect -23566 3822 -23550 4348
rect -23516 3822 -23500 4348
rect -23566 3810 -23500 3822
rect -23470 4348 -23404 4360
rect -23470 3822 -23454 4348
rect -23420 3822 -23404 4348
rect -23470 3810 -23404 3822
rect -23374 4348 -23308 4360
rect -23374 3822 -23358 4348
rect -23324 3822 -23308 4348
rect -23374 3810 -23308 3822
rect -23278 4348 -23212 4360
rect -23278 3822 -23262 4348
rect -23228 3822 -23212 4348
rect -23278 3810 -23212 3822
rect -23182 4348 -23116 4360
rect -23182 3822 -23166 4348
rect -23132 3822 -23116 4348
rect -23182 3810 -23116 3822
rect -23086 4348 -23020 4360
rect -23086 3822 -23070 4348
rect -23036 3822 -23020 4348
rect -23086 3810 -23020 3822
rect -22990 4348 -22924 4360
rect -22990 3822 -22974 4348
rect -22940 3822 -22924 4348
rect -22990 3810 -22924 3822
rect -22894 4348 -22832 4360
rect -22894 3822 -22878 4348
rect -22844 3822 -22832 4348
rect -22894 3810 -22832 3822
rect -22802 4348 -22744 4360
rect -22802 3822 -22790 4348
rect -22756 3822 -22744 4348
rect -22802 3810 -22744 3822
rect -20839 4348 -20781 4360
rect -20839 3822 -20827 4348
rect -20793 3822 -20781 4348
rect -20839 3810 -20781 3822
rect -20751 4348 -20689 4360
rect -20751 3822 -20739 4348
rect -20705 3822 -20689 4348
rect -20751 3810 -20689 3822
rect -20659 4348 -20593 4360
rect -20659 3822 -20643 4348
rect -20609 3822 -20593 4348
rect -20659 3810 -20593 3822
rect -20563 4348 -20497 4360
rect -20563 3822 -20547 4348
rect -20513 3822 -20497 4348
rect -20563 3810 -20497 3822
rect -20467 4348 -20401 4360
rect -20467 3822 -20451 4348
rect -20417 3822 -20401 4348
rect -20467 3810 -20401 3822
rect -20371 4348 -20305 4360
rect -20371 3822 -20355 4348
rect -20321 3822 -20305 4348
rect -20371 3810 -20305 3822
rect -20275 4348 -20209 4360
rect -20275 3822 -20259 4348
rect -20225 3822 -20209 4348
rect -20275 3810 -20209 3822
rect -20179 4348 -20113 4360
rect -20179 3822 -20163 4348
rect -20129 3822 -20113 4348
rect -20179 3810 -20113 3822
rect -20083 4348 -20017 4360
rect -20083 3822 -20067 4348
rect -20033 3822 -20017 4348
rect -20083 3810 -20017 3822
rect -19987 4348 -19921 4360
rect -19987 3822 -19971 4348
rect -19937 3822 -19921 4348
rect -19987 3810 -19921 3822
rect -19891 4348 -19825 4360
rect -19891 3822 -19875 4348
rect -19841 3822 -19825 4348
rect -19891 3810 -19825 3822
rect -19795 4348 -19729 4360
rect -19795 3822 -19779 4348
rect -19745 3822 -19729 4348
rect -19795 3810 -19729 3822
rect -19699 4348 -19633 4360
rect -19699 3822 -19683 4348
rect -19649 3822 -19633 4348
rect -19699 3810 -19633 3822
rect -19603 4348 -19541 4360
rect -19603 3822 -19587 4348
rect -19553 3822 -19541 4348
rect -19603 3810 -19541 3822
rect -19511 4348 -19453 4360
rect -19511 3822 -19499 4348
rect -19465 3822 -19453 4348
rect -19511 3810 -19453 3822
rect -17548 4348 -17490 4360
rect -17548 3822 -17536 4348
rect -17502 3822 -17490 4348
rect -17548 3810 -17490 3822
rect -17460 4348 -17398 4360
rect -17460 3822 -17448 4348
rect -17414 3822 -17398 4348
rect -17460 3810 -17398 3822
rect -17368 4348 -17302 4360
rect -17368 3822 -17352 4348
rect -17318 3822 -17302 4348
rect -17368 3810 -17302 3822
rect -17272 4348 -17206 4360
rect -17272 3822 -17256 4348
rect -17222 3822 -17206 4348
rect -17272 3810 -17206 3822
rect -17176 4348 -17110 4360
rect -17176 3822 -17160 4348
rect -17126 3822 -17110 4348
rect -17176 3810 -17110 3822
rect -17080 4348 -17014 4360
rect -17080 3822 -17064 4348
rect -17030 3822 -17014 4348
rect -17080 3810 -17014 3822
rect -16984 4348 -16918 4360
rect -16984 3822 -16968 4348
rect -16934 3822 -16918 4348
rect -16984 3810 -16918 3822
rect -16888 4348 -16822 4360
rect -16888 3822 -16872 4348
rect -16838 3822 -16822 4348
rect -16888 3810 -16822 3822
rect -16792 4348 -16726 4360
rect -16792 3822 -16776 4348
rect -16742 3822 -16726 4348
rect -16792 3810 -16726 3822
rect -16696 4348 -16630 4360
rect -16696 3822 -16680 4348
rect -16646 3822 -16630 4348
rect -16696 3810 -16630 3822
rect -16600 4348 -16534 4360
rect -16600 3822 -16584 4348
rect -16550 3822 -16534 4348
rect -16600 3810 -16534 3822
rect -16504 4348 -16438 4360
rect -16504 3822 -16488 4348
rect -16454 3822 -16438 4348
rect -16504 3810 -16438 3822
rect -16408 4348 -16342 4360
rect -16408 3822 -16392 4348
rect -16358 3822 -16342 4348
rect -16408 3810 -16342 3822
rect -16312 4348 -16250 4360
rect -16312 3822 -16296 4348
rect -16262 3822 -16250 4348
rect -16312 3810 -16250 3822
rect -16220 4348 -16162 4360
rect -16220 3822 -16208 4348
rect -16174 3822 -16162 4348
rect -16220 3810 -16162 3822
rect -14257 4348 -14199 4360
rect -14257 3822 -14245 4348
rect -14211 3822 -14199 4348
rect -14257 3810 -14199 3822
rect -14169 4348 -14107 4360
rect -14169 3822 -14157 4348
rect -14123 3822 -14107 4348
rect -14169 3810 -14107 3822
rect -14077 4348 -14011 4360
rect -14077 3822 -14061 4348
rect -14027 3822 -14011 4348
rect -14077 3810 -14011 3822
rect -13981 4348 -13915 4360
rect -13981 3822 -13965 4348
rect -13931 3822 -13915 4348
rect -13981 3810 -13915 3822
rect -13885 4348 -13819 4360
rect -13885 3822 -13869 4348
rect -13835 3822 -13819 4348
rect -13885 3810 -13819 3822
rect -13789 4348 -13723 4360
rect -13789 3822 -13773 4348
rect -13739 3822 -13723 4348
rect -13789 3810 -13723 3822
rect -13693 4348 -13627 4360
rect -13693 3822 -13677 4348
rect -13643 3822 -13627 4348
rect -13693 3810 -13627 3822
rect -13597 4348 -13531 4360
rect -13597 3822 -13581 4348
rect -13547 3822 -13531 4348
rect -13597 3810 -13531 3822
rect -13501 4348 -13435 4360
rect -13501 3822 -13485 4348
rect -13451 3822 -13435 4348
rect -13501 3810 -13435 3822
rect -13405 4348 -13339 4360
rect -13405 3822 -13389 4348
rect -13355 3822 -13339 4348
rect -13405 3810 -13339 3822
rect -13309 4348 -13243 4360
rect -13309 3822 -13293 4348
rect -13259 3822 -13243 4348
rect -13309 3810 -13243 3822
rect -13213 4348 -13147 4360
rect -13213 3822 -13197 4348
rect -13163 3822 -13147 4348
rect -13213 3810 -13147 3822
rect -13117 4348 -13051 4360
rect -13117 3822 -13101 4348
rect -13067 3822 -13051 4348
rect -13117 3810 -13051 3822
rect -13021 4348 -12959 4360
rect -13021 3822 -13005 4348
rect -12971 3822 -12959 4348
rect -13021 3810 -12959 3822
rect -12929 4348 -12871 4360
rect -12929 3822 -12917 4348
rect -12883 3822 -12871 4348
rect -12929 3810 -12871 3822
rect -10966 4348 -10908 4360
rect -10966 3822 -10954 4348
rect -10920 3822 -10908 4348
rect -10966 3810 -10908 3822
rect -10878 4348 -10816 4360
rect -10878 3822 -10866 4348
rect -10832 3822 -10816 4348
rect -10878 3810 -10816 3822
rect -10786 4348 -10720 4360
rect -10786 3822 -10770 4348
rect -10736 3822 -10720 4348
rect -10786 3810 -10720 3822
rect -10690 4348 -10624 4360
rect -10690 3822 -10674 4348
rect -10640 3822 -10624 4348
rect -10690 3810 -10624 3822
rect -10594 4348 -10528 4360
rect -10594 3822 -10578 4348
rect -10544 3822 -10528 4348
rect -10594 3810 -10528 3822
rect -10498 4348 -10432 4360
rect -10498 3822 -10482 4348
rect -10448 3822 -10432 4348
rect -10498 3810 -10432 3822
rect -10402 4348 -10336 4360
rect -10402 3822 -10386 4348
rect -10352 3822 -10336 4348
rect -10402 3810 -10336 3822
rect -10306 4348 -10240 4360
rect -10306 3822 -10290 4348
rect -10256 3822 -10240 4348
rect -10306 3810 -10240 3822
rect -10210 4348 -10144 4360
rect -10210 3822 -10194 4348
rect -10160 3822 -10144 4348
rect -10210 3810 -10144 3822
rect -10114 4348 -10048 4360
rect -10114 3822 -10098 4348
rect -10064 3822 -10048 4348
rect -10114 3810 -10048 3822
rect -10018 4348 -9952 4360
rect -10018 3822 -10002 4348
rect -9968 3822 -9952 4348
rect -10018 3810 -9952 3822
rect -9922 4348 -9856 4360
rect -9922 3822 -9906 4348
rect -9872 3822 -9856 4348
rect -9922 3810 -9856 3822
rect -9826 4348 -9760 4360
rect -9826 3822 -9810 4348
rect -9776 3822 -9760 4348
rect -9826 3810 -9760 3822
rect -9730 4348 -9668 4360
rect -9730 3822 -9714 4348
rect -9680 3822 -9668 4348
rect -9730 3810 -9668 3822
rect -9638 4348 -9580 4360
rect -9638 3822 -9626 4348
rect -9592 3822 -9580 4348
rect -9638 3810 -9580 3822
rect -7676 4348 -7618 4360
rect -7676 3822 -7664 4348
rect -7630 3822 -7618 4348
rect -7676 3810 -7618 3822
rect -7588 4348 -7526 4360
rect -7588 3822 -7576 4348
rect -7542 3822 -7526 4348
rect -7588 3810 -7526 3822
rect -7496 4348 -7430 4360
rect -7496 3822 -7480 4348
rect -7446 3822 -7430 4348
rect -7496 3810 -7430 3822
rect -7400 4348 -7334 4360
rect -7400 3822 -7384 4348
rect -7350 3822 -7334 4348
rect -7400 3810 -7334 3822
rect -7304 4348 -7238 4360
rect -7304 3822 -7288 4348
rect -7254 3822 -7238 4348
rect -7304 3810 -7238 3822
rect -7208 4348 -7142 4360
rect -7208 3822 -7192 4348
rect -7158 3822 -7142 4348
rect -7208 3810 -7142 3822
rect -7112 4348 -7046 4360
rect -7112 3822 -7096 4348
rect -7062 3822 -7046 4348
rect -7112 3810 -7046 3822
rect -7016 4348 -6950 4360
rect -7016 3822 -7000 4348
rect -6966 3822 -6950 4348
rect -7016 3810 -6950 3822
rect -6920 4348 -6854 4360
rect -6920 3822 -6904 4348
rect -6870 3822 -6854 4348
rect -6920 3810 -6854 3822
rect -6824 4348 -6758 4360
rect -6824 3822 -6808 4348
rect -6774 3822 -6758 4348
rect -6824 3810 -6758 3822
rect -6728 4348 -6662 4360
rect -6728 3822 -6712 4348
rect -6678 3822 -6662 4348
rect -6728 3810 -6662 3822
rect -6632 4348 -6566 4360
rect -6632 3822 -6616 4348
rect -6582 3822 -6566 4348
rect -6632 3810 -6566 3822
rect -6536 4348 -6470 4360
rect -6536 3822 -6520 4348
rect -6486 3822 -6470 4348
rect -6536 3810 -6470 3822
rect -6440 4348 -6378 4360
rect -6440 3822 -6424 4348
rect -6390 3822 -6378 4348
rect -6440 3810 -6378 3822
rect -6348 4348 -6290 4360
rect -6348 3822 -6336 4348
rect -6302 3822 -6290 4348
rect -6348 3810 -6290 3822
rect -4385 4348 -4327 4360
rect -4385 3822 -4373 4348
rect -4339 3822 -4327 4348
rect -4385 3810 -4327 3822
rect -4297 4348 -4235 4360
rect -4297 3822 -4285 4348
rect -4251 3822 -4235 4348
rect -4297 3810 -4235 3822
rect -4205 4348 -4139 4360
rect -4205 3822 -4189 4348
rect -4155 3822 -4139 4348
rect -4205 3810 -4139 3822
rect -4109 4348 -4043 4360
rect -4109 3822 -4093 4348
rect -4059 3822 -4043 4348
rect -4109 3810 -4043 3822
rect -4013 4348 -3947 4360
rect -4013 3822 -3997 4348
rect -3963 3822 -3947 4348
rect -4013 3810 -3947 3822
rect -3917 4348 -3851 4360
rect -3917 3822 -3901 4348
rect -3867 3822 -3851 4348
rect -3917 3810 -3851 3822
rect -3821 4348 -3755 4360
rect -3821 3822 -3805 4348
rect -3771 3822 -3755 4348
rect -3821 3810 -3755 3822
rect -3725 4348 -3659 4360
rect -3725 3822 -3709 4348
rect -3675 3822 -3659 4348
rect -3725 3810 -3659 3822
rect -3629 4348 -3563 4360
rect -3629 3822 -3613 4348
rect -3579 3822 -3563 4348
rect -3629 3810 -3563 3822
rect -3533 4348 -3467 4360
rect -3533 3822 -3517 4348
rect -3483 3822 -3467 4348
rect -3533 3810 -3467 3822
rect -3437 4348 -3371 4360
rect -3437 3822 -3421 4348
rect -3387 3822 -3371 4348
rect -3437 3810 -3371 3822
rect -3341 4348 -3275 4360
rect -3341 3822 -3325 4348
rect -3291 3822 -3275 4348
rect -3341 3810 -3275 3822
rect -3245 4348 -3179 4360
rect -3245 3822 -3229 4348
rect -3195 3822 -3179 4348
rect -3245 3810 -3179 3822
rect -3149 4348 -3087 4360
rect -3149 3822 -3133 4348
rect -3099 3822 -3087 4348
rect -3149 3810 -3087 3822
rect -3057 4348 -2999 4360
rect -3057 3822 -3045 4348
rect -3011 3822 -2999 4348
rect -3057 3810 -2999 3822
rect -1094 4348 -1036 4360
rect -1094 3822 -1082 4348
rect -1048 3822 -1036 4348
rect -1094 3810 -1036 3822
rect -1006 4348 -944 4360
rect -1006 3822 -994 4348
rect -960 3822 -944 4348
rect -1006 3810 -944 3822
rect -914 4348 -848 4360
rect -914 3822 -898 4348
rect -864 3822 -848 4348
rect -914 3810 -848 3822
rect -818 4348 -752 4360
rect -818 3822 -802 4348
rect -768 3822 -752 4348
rect -818 3810 -752 3822
rect -722 4348 -656 4360
rect -722 3822 -706 4348
rect -672 3822 -656 4348
rect -722 3810 -656 3822
rect -626 4348 -560 4360
rect -626 3822 -610 4348
rect -576 3822 -560 4348
rect -626 3810 -560 3822
rect -530 4348 -464 4360
rect -530 3822 -514 4348
rect -480 3822 -464 4348
rect -530 3810 -464 3822
rect -434 4348 -368 4360
rect -434 3822 -418 4348
rect -384 3822 -368 4348
rect -434 3810 -368 3822
rect -338 4348 -272 4360
rect -338 3822 -322 4348
rect -288 3822 -272 4348
rect -338 3810 -272 3822
rect -242 4348 -176 4360
rect -242 3822 -226 4348
rect -192 3822 -176 4348
rect -242 3810 -176 3822
rect -146 4348 -80 4360
rect -146 3822 -130 4348
rect -96 3822 -80 4348
rect -146 3810 -80 3822
rect -50 4348 16 4360
rect -50 3822 -34 4348
rect 0 3822 16 4348
rect -50 3810 16 3822
rect 46 4348 112 4360
rect 46 3822 62 4348
rect 96 3822 112 4348
rect 46 3810 112 3822
rect 142 4348 204 4360
rect 142 3822 158 4348
rect 192 3822 204 4348
rect 142 3810 204 3822
rect 234 4348 292 4360
rect 234 3822 246 4348
rect 280 3822 292 4348
rect 5658 3911 5872 3923
rect 234 3810 292 3822
rect 5658 3877 5670 3911
rect 5860 3877 5872 3911
rect 6098 3911 6312 3923
rect 5658 3861 5872 3877
rect 5658 3815 5872 3831
rect 5658 3781 5670 3815
rect 5864 3781 5872 3815
rect 5658 3765 5872 3781
rect 5658 3719 5872 3735
rect 5658 3685 5670 3719
rect 5860 3685 5872 3719
rect 5658 3669 5872 3685
rect 5658 3623 5872 3639
rect 5658 3589 5670 3623
rect 5864 3589 5872 3623
rect 6098 3877 6110 3911
rect 6300 3877 6312 3911
rect 6538 3911 6752 3923
rect 6098 3861 6312 3877
rect 6098 3815 6312 3831
rect 6098 3781 6110 3815
rect 6304 3781 6312 3815
rect 6098 3765 6312 3781
rect 6098 3719 6312 3735
rect 6098 3685 6110 3719
rect 6300 3685 6312 3719
rect 6098 3669 6312 3685
rect 6098 3623 6312 3639
rect 5658 3577 5872 3589
rect 6098 3589 6110 3623
rect 6304 3589 6312 3623
rect 6538 3877 6550 3911
rect 6740 3877 6752 3911
rect 6538 3861 6752 3877
rect 6538 3815 6752 3831
rect 6538 3781 6550 3815
rect 6744 3781 6752 3815
rect 6538 3765 6752 3781
rect 6538 3719 6752 3735
rect 6538 3685 6550 3719
rect 6740 3685 6752 3719
rect 6538 3669 6752 3685
rect 6538 3623 6752 3639
rect 6098 3577 6312 3589
rect 6538 3589 6550 3623
rect 6744 3589 6752 3623
rect 6538 3577 6752 3589
rect 7138 3207 7200 3219
rect 7138 2909 7150 3207
rect 7184 2909 7200 3207
rect 7138 2897 7200 2909
rect 7230 3207 7296 3219
rect 7230 2909 7246 3207
rect 7280 2909 7296 3207
rect 7230 2897 7296 2909
rect 7326 3207 7392 3219
rect 7326 2909 7342 3207
rect 7376 2909 7392 3207
rect 7326 2897 7392 2909
rect 7422 3207 7488 3219
rect 7422 2909 7438 3207
rect 7472 2909 7488 3207
rect 7422 2897 7488 2909
rect 7518 3207 7584 3219
rect 7518 2909 7534 3207
rect 7568 2909 7584 3207
rect 7518 2897 7584 2909
rect 7614 3207 7680 3219
rect 7614 2909 7630 3207
rect 7664 2909 7680 3207
rect 7614 2897 7680 2909
rect 7710 3207 7776 3219
rect 7710 2909 7726 3207
rect 7760 2909 7776 3207
rect 7710 2897 7776 2909
rect 7806 3207 7872 3219
rect 7806 2909 7822 3207
rect 7856 2909 7872 3207
rect 7806 2897 7872 2909
rect 7902 3207 7964 3219
rect 7902 2909 7918 3207
rect 7952 2909 7964 3207
rect 7902 2897 7964 2909
rect 8086 3207 8148 3219
rect 8086 2909 8098 3207
rect 8132 2909 8148 3207
rect 8086 2897 8148 2909
rect 8178 3207 8244 3219
rect 8178 2909 8194 3207
rect 8228 2909 8244 3207
rect 8178 2897 8244 2909
rect 8274 3207 8340 3219
rect 8274 2909 8290 3207
rect 8324 2909 8340 3207
rect 8274 2897 8340 2909
rect 8370 3207 8436 3219
rect 8370 2909 8386 3207
rect 8420 2909 8436 3207
rect 8370 2897 8436 2909
rect 8466 3207 8532 3219
rect 8466 2909 8482 3207
rect 8516 2909 8532 3207
rect 8466 2897 8532 2909
rect 8562 3207 8628 3219
rect 8562 2909 8578 3207
rect 8612 2909 8628 3207
rect 8562 2897 8628 2909
rect 8658 3207 8724 3219
rect 8658 2909 8674 3207
rect 8708 2909 8724 3207
rect 8658 2897 8724 2909
rect 8754 3207 8820 3219
rect 8754 2909 8770 3207
rect 8804 2909 8820 3207
rect 8754 2897 8820 2909
rect 8850 3207 8912 3219
rect 8850 2909 8866 3207
rect 8900 2909 8912 3207
rect 8850 2897 8912 2909
rect 9022 3207 9084 3219
rect 9022 2909 9034 3207
rect 9068 2909 9084 3207
rect 9022 2897 9084 2909
rect 9114 3207 9180 3219
rect 9114 2909 9130 3207
rect 9164 2909 9180 3207
rect 9114 2897 9180 2909
rect 9210 3207 9276 3219
rect 9210 2909 9226 3207
rect 9260 2909 9276 3207
rect 9210 2897 9276 2909
rect 9306 3207 9372 3219
rect 9306 2909 9322 3207
rect 9356 2909 9372 3207
rect 9306 2897 9372 2909
rect 9402 3207 9468 3219
rect 9402 2909 9418 3207
rect 9452 2909 9468 3207
rect 9402 2897 9468 2909
rect 9498 3207 9564 3219
rect 9498 2909 9514 3207
rect 9548 2909 9564 3207
rect 9498 2897 9564 2909
rect 9594 3207 9660 3219
rect 9594 2909 9610 3207
rect 9644 2909 9660 3207
rect 9594 2897 9660 2909
rect 9690 3207 9756 3219
rect 9690 2909 9706 3207
rect 9740 2909 9756 3207
rect 9690 2897 9756 2909
rect 9786 3207 9848 3219
rect 9786 2909 9802 3207
rect 9836 2909 9848 3207
rect 9786 2897 9848 2909
rect 9953 3207 10015 3219
rect 9953 2909 9965 3207
rect 9999 2909 10015 3207
rect 9953 2897 10015 2909
rect 10045 3207 10111 3219
rect 10045 2909 10061 3207
rect 10095 2909 10111 3207
rect 10045 2897 10111 2909
rect 10141 3207 10207 3219
rect 10141 2909 10157 3207
rect 10191 2909 10207 3207
rect 10141 2897 10207 2909
rect 10237 3207 10303 3219
rect 10237 2909 10253 3207
rect 10287 2909 10303 3207
rect 10237 2897 10303 2909
rect 10333 3207 10399 3219
rect 10333 2909 10349 3207
rect 10383 2909 10399 3207
rect 10333 2897 10399 2909
rect 10429 3207 10495 3219
rect 10429 2909 10445 3207
rect 10479 2909 10495 3207
rect 10429 2897 10495 2909
rect 10525 3207 10591 3219
rect 10525 2909 10541 3207
rect 10575 2909 10591 3207
rect 10525 2897 10591 2909
rect 10621 3207 10687 3219
rect 10621 2909 10637 3207
rect 10671 2909 10687 3207
rect 10621 2897 10687 2909
rect 10717 3207 10779 3219
rect 10717 2909 10733 3207
rect 10767 2909 10779 3207
rect 10717 2897 10779 2909
rect 10880 3207 10942 3219
rect 10880 2909 10892 3207
rect 10926 2909 10942 3207
rect 10880 2897 10942 2909
rect 10972 3207 11038 3219
rect 10972 2909 10988 3207
rect 11022 2909 11038 3207
rect 10972 2897 11038 2909
rect 11068 3207 11134 3219
rect 11068 2909 11084 3207
rect 11118 2909 11134 3207
rect 11068 2897 11134 2909
rect 11164 3207 11230 3219
rect 11164 2909 11180 3207
rect 11214 2909 11230 3207
rect 11164 2897 11230 2909
rect 11260 3207 11326 3219
rect 11260 2909 11276 3207
rect 11310 2909 11326 3207
rect 11260 2897 11326 2909
rect 11356 3207 11422 3219
rect 11356 2909 11372 3207
rect 11406 2909 11422 3207
rect 11356 2897 11422 2909
rect 11452 3207 11518 3219
rect 11452 2909 11468 3207
rect 11502 2909 11518 3207
rect 11452 2897 11518 2909
rect 11548 3207 11614 3219
rect 11548 2909 11564 3207
rect 11598 2909 11614 3207
rect 11548 2897 11614 2909
rect 11644 3207 11706 3219
rect 11644 2909 11660 3207
rect 11694 2909 11706 3207
rect 11644 2897 11706 2909
rect -24804 2564 -24746 2576
rect -24804 2038 -24792 2564
rect -24758 2038 -24746 2564
rect -24804 2026 -24746 2038
rect -24716 2564 -24654 2576
rect -24716 2038 -24704 2564
rect -24670 2038 -24654 2564
rect -24716 2026 -24654 2038
rect -24624 2564 -24558 2576
rect -24624 2038 -24608 2564
rect -24574 2038 -24558 2564
rect -24624 2026 -24558 2038
rect -24528 2564 -24462 2576
rect -24528 2038 -24512 2564
rect -24478 2038 -24462 2564
rect -24528 2026 -24462 2038
rect -24432 2564 -24366 2576
rect -24432 2038 -24416 2564
rect -24382 2038 -24366 2564
rect -24432 2026 -24366 2038
rect -24336 2564 -24270 2576
rect -24336 2038 -24320 2564
rect -24286 2038 -24270 2564
rect -24336 2026 -24270 2038
rect -24240 2564 -24174 2576
rect -24240 2038 -24224 2564
rect -24190 2038 -24174 2564
rect -24240 2026 -24174 2038
rect -24144 2564 -24078 2576
rect -24144 2038 -24128 2564
rect -24094 2038 -24078 2564
rect -24144 2026 -24078 2038
rect -24048 2564 -23982 2576
rect -24048 2038 -24032 2564
rect -23998 2038 -23982 2564
rect -24048 2026 -23982 2038
rect -23952 2564 -23886 2576
rect -23952 2038 -23936 2564
rect -23902 2038 -23886 2564
rect -23952 2026 -23886 2038
rect -23856 2564 -23790 2576
rect -23856 2038 -23840 2564
rect -23806 2038 -23790 2564
rect -23856 2026 -23790 2038
rect -23760 2564 -23694 2576
rect -23760 2038 -23744 2564
rect -23710 2038 -23694 2564
rect -23760 2026 -23694 2038
rect -23664 2564 -23598 2576
rect -23664 2038 -23648 2564
rect -23614 2038 -23598 2564
rect -23664 2026 -23598 2038
rect -23568 2564 -23506 2576
rect -23568 2038 -23552 2564
rect -23518 2038 -23506 2564
rect -23568 2026 -23506 2038
rect -23476 2564 -23418 2576
rect -23476 2038 -23464 2564
rect -23430 2038 -23418 2564
rect -23476 2026 -23418 2038
rect -23245 2564 -23187 2576
rect -23245 2038 -23233 2564
rect -23199 2038 -23187 2564
rect -23245 2026 -23187 2038
rect -23157 2564 -23095 2576
rect -23157 2038 -23145 2564
rect -23111 2038 -23095 2564
rect -23157 2026 -23095 2038
rect -23065 2564 -22999 2576
rect -23065 2038 -23049 2564
rect -23015 2038 -22999 2564
rect -23065 2026 -22999 2038
rect -22969 2564 -22903 2576
rect -22969 2038 -22953 2564
rect -22919 2038 -22903 2564
rect -22969 2026 -22903 2038
rect -22873 2564 -22807 2576
rect -22873 2038 -22857 2564
rect -22823 2038 -22807 2564
rect -22873 2026 -22807 2038
rect -22777 2564 -22711 2576
rect -22777 2038 -22761 2564
rect -22727 2038 -22711 2564
rect -22777 2026 -22711 2038
rect -22681 2564 -22615 2576
rect -22681 2038 -22665 2564
rect -22631 2038 -22615 2564
rect -22681 2026 -22615 2038
rect -22585 2564 -22519 2576
rect -22585 2038 -22569 2564
rect -22535 2038 -22519 2564
rect -22585 2026 -22519 2038
rect -22489 2564 -22423 2576
rect -22489 2038 -22473 2564
rect -22439 2038 -22423 2564
rect -22489 2026 -22423 2038
rect -22393 2564 -22327 2576
rect -22393 2038 -22377 2564
rect -22343 2038 -22327 2564
rect -22393 2026 -22327 2038
rect -22297 2564 -22231 2576
rect -22297 2038 -22281 2564
rect -22247 2038 -22231 2564
rect -22297 2026 -22231 2038
rect -22201 2564 -22135 2576
rect -22201 2038 -22185 2564
rect -22151 2038 -22135 2564
rect -22201 2026 -22135 2038
rect -22105 2564 -22039 2576
rect -22105 2038 -22089 2564
rect -22055 2038 -22039 2564
rect -22105 2026 -22039 2038
rect -22009 2564 -21947 2576
rect -22009 2038 -21993 2564
rect -21959 2038 -21947 2564
rect -22009 2026 -21947 2038
rect -21917 2564 -21859 2576
rect -21917 2038 -21905 2564
rect -21871 2038 -21859 2564
rect -21917 2026 -21859 2038
rect -21513 2564 -21455 2576
rect -21513 2038 -21501 2564
rect -21467 2038 -21455 2564
rect -21513 2026 -21455 2038
rect -21425 2564 -21363 2576
rect -21425 2038 -21413 2564
rect -21379 2038 -21363 2564
rect -21425 2026 -21363 2038
rect -21333 2564 -21267 2576
rect -21333 2038 -21317 2564
rect -21283 2038 -21267 2564
rect -21333 2026 -21267 2038
rect -21237 2564 -21171 2576
rect -21237 2038 -21221 2564
rect -21187 2038 -21171 2564
rect -21237 2026 -21171 2038
rect -21141 2564 -21075 2576
rect -21141 2038 -21125 2564
rect -21091 2038 -21075 2564
rect -21141 2026 -21075 2038
rect -21045 2564 -20979 2576
rect -21045 2038 -21029 2564
rect -20995 2038 -20979 2564
rect -21045 2026 -20979 2038
rect -20949 2564 -20883 2576
rect -20949 2038 -20933 2564
rect -20899 2038 -20883 2564
rect -20949 2026 -20883 2038
rect -20853 2564 -20787 2576
rect -20853 2038 -20837 2564
rect -20803 2038 -20787 2564
rect -20853 2026 -20787 2038
rect -20757 2564 -20691 2576
rect -20757 2038 -20741 2564
rect -20707 2038 -20691 2564
rect -20757 2026 -20691 2038
rect -20661 2564 -20595 2576
rect -20661 2038 -20645 2564
rect -20611 2038 -20595 2564
rect -20661 2026 -20595 2038
rect -20565 2564 -20499 2576
rect -20565 2038 -20549 2564
rect -20515 2038 -20499 2564
rect -20565 2026 -20499 2038
rect -20469 2564 -20403 2576
rect -20469 2038 -20453 2564
rect -20419 2038 -20403 2564
rect -20469 2026 -20403 2038
rect -20373 2564 -20307 2576
rect -20373 2038 -20357 2564
rect -20323 2038 -20307 2564
rect -20373 2026 -20307 2038
rect -20277 2564 -20215 2576
rect -20277 2038 -20261 2564
rect -20227 2038 -20215 2564
rect -20277 2026 -20215 2038
rect -20185 2564 -20127 2576
rect -20185 2038 -20173 2564
rect -20139 2038 -20127 2564
rect -20185 2026 -20127 2038
rect -19954 2564 -19896 2576
rect -19954 2038 -19942 2564
rect -19908 2038 -19896 2564
rect -19954 2026 -19896 2038
rect -19866 2564 -19804 2576
rect -19866 2038 -19854 2564
rect -19820 2038 -19804 2564
rect -19866 2026 -19804 2038
rect -19774 2564 -19708 2576
rect -19774 2038 -19758 2564
rect -19724 2038 -19708 2564
rect -19774 2026 -19708 2038
rect -19678 2564 -19612 2576
rect -19678 2038 -19662 2564
rect -19628 2038 -19612 2564
rect -19678 2026 -19612 2038
rect -19582 2564 -19516 2576
rect -19582 2038 -19566 2564
rect -19532 2038 -19516 2564
rect -19582 2026 -19516 2038
rect -19486 2564 -19420 2576
rect -19486 2038 -19470 2564
rect -19436 2038 -19420 2564
rect -19486 2026 -19420 2038
rect -19390 2564 -19324 2576
rect -19390 2038 -19374 2564
rect -19340 2038 -19324 2564
rect -19390 2026 -19324 2038
rect -19294 2564 -19228 2576
rect -19294 2038 -19278 2564
rect -19244 2038 -19228 2564
rect -19294 2026 -19228 2038
rect -19198 2564 -19132 2576
rect -19198 2038 -19182 2564
rect -19148 2038 -19132 2564
rect -19198 2026 -19132 2038
rect -19102 2564 -19036 2576
rect -19102 2038 -19086 2564
rect -19052 2038 -19036 2564
rect -19102 2026 -19036 2038
rect -19006 2564 -18940 2576
rect -19006 2038 -18990 2564
rect -18956 2038 -18940 2564
rect -19006 2026 -18940 2038
rect -18910 2564 -18844 2576
rect -18910 2038 -18894 2564
rect -18860 2038 -18844 2564
rect -18910 2026 -18844 2038
rect -18814 2564 -18748 2576
rect -18814 2038 -18798 2564
rect -18764 2038 -18748 2564
rect -18814 2026 -18748 2038
rect -18718 2564 -18656 2576
rect -18718 2038 -18702 2564
rect -18668 2038 -18656 2564
rect -18718 2026 -18656 2038
rect -18626 2564 -18568 2576
rect -18626 2038 -18614 2564
rect -18580 2038 -18568 2564
rect -18626 2026 -18568 2038
rect -18222 2564 -18164 2576
rect -18222 2038 -18210 2564
rect -18176 2038 -18164 2564
rect -18222 2026 -18164 2038
rect -18134 2564 -18072 2576
rect -18134 2038 -18122 2564
rect -18088 2038 -18072 2564
rect -18134 2026 -18072 2038
rect -18042 2564 -17976 2576
rect -18042 2038 -18026 2564
rect -17992 2038 -17976 2564
rect -18042 2026 -17976 2038
rect -17946 2564 -17880 2576
rect -17946 2038 -17930 2564
rect -17896 2038 -17880 2564
rect -17946 2026 -17880 2038
rect -17850 2564 -17784 2576
rect -17850 2038 -17834 2564
rect -17800 2038 -17784 2564
rect -17850 2026 -17784 2038
rect -17754 2564 -17688 2576
rect -17754 2038 -17738 2564
rect -17704 2038 -17688 2564
rect -17754 2026 -17688 2038
rect -17658 2564 -17592 2576
rect -17658 2038 -17642 2564
rect -17608 2038 -17592 2564
rect -17658 2026 -17592 2038
rect -17562 2564 -17496 2576
rect -17562 2038 -17546 2564
rect -17512 2038 -17496 2564
rect -17562 2026 -17496 2038
rect -17466 2564 -17400 2576
rect -17466 2038 -17450 2564
rect -17416 2038 -17400 2564
rect -17466 2026 -17400 2038
rect -17370 2564 -17304 2576
rect -17370 2038 -17354 2564
rect -17320 2038 -17304 2564
rect -17370 2026 -17304 2038
rect -17274 2564 -17208 2576
rect -17274 2038 -17258 2564
rect -17224 2038 -17208 2564
rect -17274 2026 -17208 2038
rect -17178 2564 -17112 2576
rect -17178 2038 -17162 2564
rect -17128 2038 -17112 2564
rect -17178 2026 -17112 2038
rect -17082 2564 -17016 2576
rect -17082 2038 -17066 2564
rect -17032 2038 -17016 2564
rect -17082 2026 -17016 2038
rect -16986 2564 -16924 2576
rect -16986 2038 -16970 2564
rect -16936 2038 -16924 2564
rect -16986 2026 -16924 2038
rect -16894 2564 -16836 2576
rect -16894 2038 -16882 2564
rect -16848 2038 -16836 2564
rect -16894 2026 -16836 2038
rect -16663 2564 -16605 2576
rect -16663 2038 -16651 2564
rect -16617 2038 -16605 2564
rect -16663 2026 -16605 2038
rect -16575 2564 -16513 2576
rect -16575 2038 -16563 2564
rect -16529 2038 -16513 2564
rect -16575 2026 -16513 2038
rect -16483 2564 -16417 2576
rect -16483 2038 -16467 2564
rect -16433 2038 -16417 2564
rect -16483 2026 -16417 2038
rect -16387 2564 -16321 2576
rect -16387 2038 -16371 2564
rect -16337 2038 -16321 2564
rect -16387 2026 -16321 2038
rect -16291 2564 -16225 2576
rect -16291 2038 -16275 2564
rect -16241 2038 -16225 2564
rect -16291 2026 -16225 2038
rect -16195 2564 -16129 2576
rect -16195 2038 -16179 2564
rect -16145 2038 -16129 2564
rect -16195 2026 -16129 2038
rect -16099 2564 -16033 2576
rect -16099 2038 -16083 2564
rect -16049 2038 -16033 2564
rect -16099 2026 -16033 2038
rect -16003 2564 -15937 2576
rect -16003 2038 -15987 2564
rect -15953 2038 -15937 2564
rect -16003 2026 -15937 2038
rect -15907 2564 -15841 2576
rect -15907 2038 -15891 2564
rect -15857 2038 -15841 2564
rect -15907 2026 -15841 2038
rect -15811 2564 -15745 2576
rect -15811 2038 -15795 2564
rect -15761 2038 -15745 2564
rect -15811 2026 -15745 2038
rect -15715 2564 -15649 2576
rect -15715 2038 -15699 2564
rect -15665 2038 -15649 2564
rect -15715 2026 -15649 2038
rect -15619 2564 -15553 2576
rect -15619 2038 -15603 2564
rect -15569 2038 -15553 2564
rect -15619 2026 -15553 2038
rect -15523 2564 -15457 2576
rect -15523 2038 -15507 2564
rect -15473 2038 -15457 2564
rect -15523 2026 -15457 2038
rect -15427 2564 -15365 2576
rect -15427 2038 -15411 2564
rect -15377 2038 -15365 2564
rect -15427 2026 -15365 2038
rect -15335 2564 -15277 2576
rect -15335 2038 -15323 2564
rect -15289 2038 -15277 2564
rect -15335 2026 -15277 2038
rect -14931 2564 -14873 2576
rect -14931 2038 -14919 2564
rect -14885 2038 -14873 2564
rect -14931 2026 -14873 2038
rect -14843 2564 -14781 2576
rect -14843 2038 -14831 2564
rect -14797 2038 -14781 2564
rect -14843 2026 -14781 2038
rect -14751 2564 -14685 2576
rect -14751 2038 -14735 2564
rect -14701 2038 -14685 2564
rect -14751 2026 -14685 2038
rect -14655 2564 -14589 2576
rect -14655 2038 -14639 2564
rect -14605 2038 -14589 2564
rect -14655 2026 -14589 2038
rect -14559 2564 -14493 2576
rect -14559 2038 -14543 2564
rect -14509 2038 -14493 2564
rect -14559 2026 -14493 2038
rect -14463 2564 -14397 2576
rect -14463 2038 -14447 2564
rect -14413 2038 -14397 2564
rect -14463 2026 -14397 2038
rect -14367 2564 -14301 2576
rect -14367 2038 -14351 2564
rect -14317 2038 -14301 2564
rect -14367 2026 -14301 2038
rect -14271 2564 -14205 2576
rect -14271 2038 -14255 2564
rect -14221 2038 -14205 2564
rect -14271 2026 -14205 2038
rect -14175 2564 -14109 2576
rect -14175 2038 -14159 2564
rect -14125 2038 -14109 2564
rect -14175 2026 -14109 2038
rect -14079 2564 -14013 2576
rect -14079 2038 -14063 2564
rect -14029 2038 -14013 2564
rect -14079 2026 -14013 2038
rect -13983 2564 -13917 2576
rect -13983 2038 -13967 2564
rect -13933 2038 -13917 2564
rect -13983 2026 -13917 2038
rect -13887 2564 -13821 2576
rect -13887 2038 -13871 2564
rect -13837 2038 -13821 2564
rect -13887 2026 -13821 2038
rect -13791 2564 -13725 2576
rect -13791 2038 -13775 2564
rect -13741 2038 -13725 2564
rect -13791 2026 -13725 2038
rect -13695 2564 -13633 2576
rect -13695 2038 -13679 2564
rect -13645 2038 -13633 2564
rect -13695 2026 -13633 2038
rect -13603 2564 -13545 2576
rect -13603 2038 -13591 2564
rect -13557 2038 -13545 2564
rect -13603 2026 -13545 2038
rect -13372 2564 -13314 2576
rect -13372 2038 -13360 2564
rect -13326 2038 -13314 2564
rect -13372 2026 -13314 2038
rect -13284 2564 -13222 2576
rect -13284 2038 -13272 2564
rect -13238 2038 -13222 2564
rect -13284 2026 -13222 2038
rect -13192 2564 -13126 2576
rect -13192 2038 -13176 2564
rect -13142 2038 -13126 2564
rect -13192 2026 -13126 2038
rect -13096 2564 -13030 2576
rect -13096 2038 -13080 2564
rect -13046 2038 -13030 2564
rect -13096 2026 -13030 2038
rect -13000 2564 -12934 2576
rect -13000 2038 -12984 2564
rect -12950 2038 -12934 2564
rect -13000 2026 -12934 2038
rect -12904 2564 -12838 2576
rect -12904 2038 -12888 2564
rect -12854 2038 -12838 2564
rect -12904 2026 -12838 2038
rect -12808 2564 -12742 2576
rect -12808 2038 -12792 2564
rect -12758 2038 -12742 2564
rect -12808 2026 -12742 2038
rect -12712 2564 -12646 2576
rect -12712 2038 -12696 2564
rect -12662 2038 -12646 2564
rect -12712 2026 -12646 2038
rect -12616 2564 -12550 2576
rect -12616 2038 -12600 2564
rect -12566 2038 -12550 2564
rect -12616 2026 -12550 2038
rect -12520 2564 -12454 2576
rect -12520 2038 -12504 2564
rect -12470 2038 -12454 2564
rect -12520 2026 -12454 2038
rect -12424 2564 -12358 2576
rect -12424 2038 -12408 2564
rect -12374 2038 -12358 2564
rect -12424 2026 -12358 2038
rect -12328 2564 -12262 2576
rect -12328 2038 -12312 2564
rect -12278 2038 -12262 2564
rect -12328 2026 -12262 2038
rect -12232 2564 -12166 2576
rect -12232 2038 -12216 2564
rect -12182 2038 -12166 2564
rect -12232 2026 -12166 2038
rect -12136 2564 -12074 2576
rect -12136 2038 -12120 2564
rect -12086 2038 -12074 2564
rect -12136 2026 -12074 2038
rect -12044 2564 -11986 2576
rect -12044 2038 -12032 2564
rect -11998 2038 -11986 2564
rect -12044 2026 -11986 2038
rect -11640 2564 -11582 2576
rect -11640 2038 -11628 2564
rect -11594 2038 -11582 2564
rect -11640 2026 -11582 2038
rect -11552 2564 -11490 2576
rect -11552 2038 -11540 2564
rect -11506 2038 -11490 2564
rect -11552 2026 -11490 2038
rect -11460 2564 -11394 2576
rect -11460 2038 -11444 2564
rect -11410 2038 -11394 2564
rect -11460 2026 -11394 2038
rect -11364 2564 -11298 2576
rect -11364 2038 -11348 2564
rect -11314 2038 -11298 2564
rect -11364 2026 -11298 2038
rect -11268 2564 -11202 2576
rect -11268 2038 -11252 2564
rect -11218 2038 -11202 2564
rect -11268 2026 -11202 2038
rect -11172 2564 -11106 2576
rect -11172 2038 -11156 2564
rect -11122 2038 -11106 2564
rect -11172 2026 -11106 2038
rect -11076 2564 -11010 2576
rect -11076 2038 -11060 2564
rect -11026 2038 -11010 2564
rect -11076 2026 -11010 2038
rect -10980 2564 -10914 2576
rect -10980 2038 -10964 2564
rect -10930 2038 -10914 2564
rect -10980 2026 -10914 2038
rect -10884 2564 -10818 2576
rect -10884 2038 -10868 2564
rect -10834 2038 -10818 2564
rect -10884 2026 -10818 2038
rect -10788 2564 -10722 2576
rect -10788 2038 -10772 2564
rect -10738 2038 -10722 2564
rect -10788 2026 -10722 2038
rect -10692 2564 -10626 2576
rect -10692 2038 -10676 2564
rect -10642 2038 -10626 2564
rect -10692 2026 -10626 2038
rect -10596 2564 -10530 2576
rect -10596 2038 -10580 2564
rect -10546 2038 -10530 2564
rect -10596 2026 -10530 2038
rect -10500 2564 -10434 2576
rect -10500 2038 -10484 2564
rect -10450 2038 -10434 2564
rect -10500 2026 -10434 2038
rect -10404 2564 -10342 2576
rect -10404 2038 -10388 2564
rect -10354 2038 -10342 2564
rect -10404 2026 -10342 2038
rect -10312 2564 -10254 2576
rect -10312 2038 -10300 2564
rect -10266 2038 -10254 2564
rect -10312 2026 -10254 2038
rect -10081 2564 -10023 2576
rect -10081 2038 -10069 2564
rect -10035 2038 -10023 2564
rect -10081 2026 -10023 2038
rect -9993 2564 -9931 2576
rect -9993 2038 -9981 2564
rect -9947 2038 -9931 2564
rect -9993 2026 -9931 2038
rect -9901 2564 -9835 2576
rect -9901 2038 -9885 2564
rect -9851 2038 -9835 2564
rect -9901 2026 -9835 2038
rect -9805 2564 -9739 2576
rect -9805 2038 -9789 2564
rect -9755 2038 -9739 2564
rect -9805 2026 -9739 2038
rect -9709 2564 -9643 2576
rect -9709 2038 -9693 2564
rect -9659 2038 -9643 2564
rect -9709 2026 -9643 2038
rect -9613 2564 -9547 2576
rect -9613 2038 -9597 2564
rect -9563 2038 -9547 2564
rect -9613 2026 -9547 2038
rect -9517 2564 -9451 2576
rect -9517 2038 -9501 2564
rect -9467 2038 -9451 2564
rect -9517 2026 -9451 2038
rect -9421 2564 -9355 2576
rect -9421 2038 -9405 2564
rect -9371 2038 -9355 2564
rect -9421 2026 -9355 2038
rect -9325 2564 -9259 2576
rect -9325 2038 -9309 2564
rect -9275 2038 -9259 2564
rect -9325 2026 -9259 2038
rect -9229 2564 -9163 2576
rect -9229 2038 -9213 2564
rect -9179 2038 -9163 2564
rect -9229 2026 -9163 2038
rect -9133 2564 -9067 2576
rect -9133 2038 -9117 2564
rect -9083 2038 -9067 2564
rect -9133 2026 -9067 2038
rect -9037 2564 -8971 2576
rect -9037 2038 -9021 2564
rect -8987 2038 -8971 2564
rect -9037 2026 -8971 2038
rect -8941 2564 -8875 2576
rect -8941 2038 -8925 2564
rect -8891 2038 -8875 2564
rect -8941 2026 -8875 2038
rect -8845 2564 -8783 2576
rect -8845 2038 -8829 2564
rect -8795 2038 -8783 2564
rect -8845 2026 -8783 2038
rect -8753 2564 -8695 2576
rect -8753 2038 -8741 2564
rect -8707 2038 -8695 2564
rect -8753 2026 -8695 2038
rect -8350 2564 -8292 2576
rect -8350 2038 -8338 2564
rect -8304 2038 -8292 2564
rect -8350 2026 -8292 2038
rect -8262 2564 -8200 2576
rect -8262 2038 -8250 2564
rect -8216 2038 -8200 2564
rect -8262 2026 -8200 2038
rect -8170 2564 -8104 2576
rect -8170 2038 -8154 2564
rect -8120 2038 -8104 2564
rect -8170 2026 -8104 2038
rect -8074 2564 -8008 2576
rect -8074 2038 -8058 2564
rect -8024 2038 -8008 2564
rect -8074 2026 -8008 2038
rect -7978 2564 -7912 2576
rect -7978 2038 -7962 2564
rect -7928 2038 -7912 2564
rect -7978 2026 -7912 2038
rect -7882 2564 -7816 2576
rect -7882 2038 -7866 2564
rect -7832 2038 -7816 2564
rect -7882 2026 -7816 2038
rect -7786 2564 -7720 2576
rect -7786 2038 -7770 2564
rect -7736 2038 -7720 2564
rect -7786 2026 -7720 2038
rect -7690 2564 -7624 2576
rect -7690 2038 -7674 2564
rect -7640 2038 -7624 2564
rect -7690 2026 -7624 2038
rect -7594 2564 -7528 2576
rect -7594 2038 -7578 2564
rect -7544 2038 -7528 2564
rect -7594 2026 -7528 2038
rect -7498 2564 -7432 2576
rect -7498 2038 -7482 2564
rect -7448 2038 -7432 2564
rect -7498 2026 -7432 2038
rect -7402 2564 -7336 2576
rect -7402 2038 -7386 2564
rect -7352 2038 -7336 2564
rect -7402 2026 -7336 2038
rect -7306 2564 -7240 2576
rect -7306 2038 -7290 2564
rect -7256 2038 -7240 2564
rect -7306 2026 -7240 2038
rect -7210 2564 -7144 2576
rect -7210 2038 -7194 2564
rect -7160 2038 -7144 2564
rect -7210 2026 -7144 2038
rect -7114 2564 -7052 2576
rect -7114 2038 -7098 2564
rect -7064 2038 -7052 2564
rect -7114 2026 -7052 2038
rect -7022 2564 -6964 2576
rect -7022 2038 -7010 2564
rect -6976 2038 -6964 2564
rect -7022 2026 -6964 2038
rect -6791 2564 -6733 2576
rect -6791 2038 -6779 2564
rect -6745 2038 -6733 2564
rect -6791 2026 -6733 2038
rect -6703 2564 -6641 2576
rect -6703 2038 -6691 2564
rect -6657 2038 -6641 2564
rect -6703 2026 -6641 2038
rect -6611 2564 -6545 2576
rect -6611 2038 -6595 2564
rect -6561 2038 -6545 2564
rect -6611 2026 -6545 2038
rect -6515 2564 -6449 2576
rect -6515 2038 -6499 2564
rect -6465 2038 -6449 2564
rect -6515 2026 -6449 2038
rect -6419 2564 -6353 2576
rect -6419 2038 -6403 2564
rect -6369 2038 -6353 2564
rect -6419 2026 -6353 2038
rect -6323 2564 -6257 2576
rect -6323 2038 -6307 2564
rect -6273 2038 -6257 2564
rect -6323 2026 -6257 2038
rect -6227 2564 -6161 2576
rect -6227 2038 -6211 2564
rect -6177 2038 -6161 2564
rect -6227 2026 -6161 2038
rect -6131 2564 -6065 2576
rect -6131 2038 -6115 2564
rect -6081 2038 -6065 2564
rect -6131 2026 -6065 2038
rect -6035 2564 -5969 2576
rect -6035 2038 -6019 2564
rect -5985 2038 -5969 2564
rect -6035 2026 -5969 2038
rect -5939 2564 -5873 2576
rect -5939 2038 -5923 2564
rect -5889 2038 -5873 2564
rect -5939 2026 -5873 2038
rect -5843 2564 -5777 2576
rect -5843 2038 -5827 2564
rect -5793 2038 -5777 2564
rect -5843 2026 -5777 2038
rect -5747 2564 -5681 2576
rect -5747 2038 -5731 2564
rect -5697 2038 -5681 2564
rect -5747 2026 -5681 2038
rect -5651 2564 -5585 2576
rect -5651 2038 -5635 2564
rect -5601 2038 -5585 2564
rect -5651 2026 -5585 2038
rect -5555 2564 -5493 2576
rect -5555 2038 -5539 2564
rect -5505 2038 -5493 2564
rect -5555 2026 -5493 2038
rect -5463 2564 -5405 2576
rect -5463 2038 -5451 2564
rect -5417 2038 -5405 2564
rect -5463 2026 -5405 2038
rect -5059 2564 -5001 2576
rect -5059 2038 -5047 2564
rect -5013 2038 -5001 2564
rect -5059 2026 -5001 2038
rect -4971 2564 -4909 2576
rect -4971 2038 -4959 2564
rect -4925 2038 -4909 2564
rect -4971 2026 -4909 2038
rect -4879 2564 -4813 2576
rect -4879 2038 -4863 2564
rect -4829 2038 -4813 2564
rect -4879 2026 -4813 2038
rect -4783 2564 -4717 2576
rect -4783 2038 -4767 2564
rect -4733 2038 -4717 2564
rect -4783 2026 -4717 2038
rect -4687 2564 -4621 2576
rect -4687 2038 -4671 2564
rect -4637 2038 -4621 2564
rect -4687 2026 -4621 2038
rect -4591 2564 -4525 2576
rect -4591 2038 -4575 2564
rect -4541 2038 -4525 2564
rect -4591 2026 -4525 2038
rect -4495 2564 -4429 2576
rect -4495 2038 -4479 2564
rect -4445 2038 -4429 2564
rect -4495 2026 -4429 2038
rect -4399 2564 -4333 2576
rect -4399 2038 -4383 2564
rect -4349 2038 -4333 2564
rect -4399 2026 -4333 2038
rect -4303 2564 -4237 2576
rect -4303 2038 -4287 2564
rect -4253 2038 -4237 2564
rect -4303 2026 -4237 2038
rect -4207 2564 -4141 2576
rect -4207 2038 -4191 2564
rect -4157 2038 -4141 2564
rect -4207 2026 -4141 2038
rect -4111 2564 -4045 2576
rect -4111 2038 -4095 2564
rect -4061 2038 -4045 2564
rect -4111 2026 -4045 2038
rect -4015 2564 -3949 2576
rect -4015 2038 -3999 2564
rect -3965 2038 -3949 2564
rect -4015 2026 -3949 2038
rect -3919 2564 -3853 2576
rect -3919 2038 -3903 2564
rect -3869 2038 -3853 2564
rect -3919 2026 -3853 2038
rect -3823 2564 -3761 2576
rect -3823 2038 -3807 2564
rect -3773 2038 -3761 2564
rect -3823 2026 -3761 2038
rect -3731 2564 -3673 2576
rect -3731 2038 -3719 2564
rect -3685 2038 -3673 2564
rect -3731 2026 -3673 2038
rect -3500 2564 -3442 2576
rect -3500 2038 -3488 2564
rect -3454 2038 -3442 2564
rect -3500 2026 -3442 2038
rect -3412 2564 -3350 2576
rect -3412 2038 -3400 2564
rect -3366 2038 -3350 2564
rect -3412 2026 -3350 2038
rect -3320 2564 -3254 2576
rect -3320 2038 -3304 2564
rect -3270 2038 -3254 2564
rect -3320 2026 -3254 2038
rect -3224 2564 -3158 2576
rect -3224 2038 -3208 2564
rect -3174 2038 -3158 2564
rect -3224 2026 -3158 2038
rect -3128 2564 -3062 2576
rect -3128 2038 -3112 2564
rect -3078 2038 -3062 2564
rect -3128 2026 -3062 2038
rect -3032 2564 -2966 2576
rect -3032 2038 -3016 2564
rect -2982 2038 -2966 2564
rect -3032 2026 -2966 2038
rect -2936 2564 -2870 2576
rect -2936 2038 -2920 2564
rect -2886 2038 -2870 2564
rect -2936 2026 -2870 2038
rect -2840 2564 -2774 2576
rect -2840 2038 -2824 2564
rect -2790 2038 -2774 2564
rect -2840 2026 -2774 2038
rect -2744 2564 -2678 2576
rect -2744 2038 -2728 2564
rect -2694 2038 -2678 2564
rect -2744 2026 -2678 2038
rect -2648 2564 -2582 2576
rect -2648 2038 -2632 2564
rect -2598 2038 -2582 2564
rect -2648 2026 -2582 2038
rect -2552 2564 -2486 2576
rect -2552 2038 -2536 2564
rect -2502 2038 -2486 2564
rect -2552 2026 -2486 2038
rect -2456 2564 -2390 2576
rect -2456 2038 -2440 2564
rect -2406 2038 -2390 2564
rect -2456 2026 -2390 2038
rect -2360 2564 -2294 2576
rect -2360 2038 -2344 2564
rect -2310 2038 -2294 2564
rect -2360 2026 -2294 2038
rect -2264 2564 -2202 2576
rect -2264 2038 -2248 2564
rect -2214 2038 -2202 2564
rect -2264 2026 -2202 2038
rect -2172 2564 -2114 2576
rect -2172 2038 -2160 2564
rect -2126 2038 -2114 2564
rect -2172 2026 -2114 2038
rect -1768 2564 -1710 2576
rect -1768 2038 -1756 2564
rect -1722 2038 -1710 2564
rect -1768 2026 -1710 2038
rect -1680 2564 -1618 2576
rect -1680 2038 -1668 2564
rect -1634 2038 -1618 2564
rect -1680 2026 -1618 2038
rect -1588 2564 -1522 2576
rect -1588 2038 -1572 2564
rect -1538 2038 -1522 2564
rect -1588 2026 -1522 2038
rect -1492 2564 -1426 2576
rect -1492 2038 -1476 2564
rect -1442 2038 -1426 2564
rect -1492 2026 -1426 2038
rect -1396 2564 -1330 2576
rect -1396 2038 -1380 2564
rect -1346 2038 -1330 2564
rect -1396 2026 -1330 2038
rect -1300 2564 -1234 2576
rect -1300 2038 -1284 2564
rect -1250 2038 -1234 2564
rect -1300 2026 -1234 2038
rect -1204 2564 -1138 2576
rect -1204 2038 -1188 2564
rect -1154 2038 -1138 2564
rect -1204 2026 -1138 2038
rect -1108 2564 -1042 2576
rect -1108 2038 -1092 2564
rect -1058 2038 -1042 2564
rect -1108 2026 -1042 2038
rect -1012 2564 -946 2576
rect -1012 2038 -996 2564
rect -962 2038 -946 2564
rect -1012 2026 -946 2038
rect -916 2564 -850 2576
rect -916 2038 -900 2564
rect -866 2038 -850 2564
rect -916 2026 -850 2038
rect -820 2564 -754 2576
rect -820 2038 -804 2564
rect -770 2038 -754 2564
rect -820 2026 -754 2038
rect -724 2564 -658 2576
rect -724 2038 -708 2564
rect -674 2038 -658 2564
rect -724 2026 -658 2038
rect -628 2564 -562 2576
rect -628 2038 -612 2564
rect -578 2038 -562 2564
rect -628 2026 -562 2038
rect -532 2564 -470 2576
rect -532 2038 -516 2564
rect -482 2038 -470 2564
rect -532 2026 -470 2038
rect -440 2564 -382 2576
rect -440 2038 -428 2564
rect -394 2038 -382 2564
rect -440 2026 -382 2038
rect -209 2564 -151 2576
rect -209 2038 -197 2564
rect -163 2038 -151 2564
rect -209 2026 -151 2038
rect -121 2564 -59 2576
rect -121 2038 -109 2564
rect -75 2038 -59 2564
rect -121 2026 -59 2038
rect -29 2564 37 2576
rect -29 2038 -13 2564
rect 21 2038 37 2564
rect -29 2026 37 2038
rect 67 2564 133 2576
rect 67 2038 83 2564
rect 117 2038 133 2564
rect 67 2026 133 2038
rect 163 2564 229 2576
rect 163 2038 179 2564
rect 213 2038 229 2564
rect 163 2026 229 2038
rect 259 2564 325 2576
rect 259 2038 275 2564
rect 309 2038 325 2564
rect 259 2026 325 2038
rect 355 2564 421 2576
rect 355 2038 371 2564
rect 405 2038 421 2564
rect 355 2026 421 2038
rect 451 2564 517 2576
rect 451 2038 467 2564
rect 501 2038 517 2564
rect 451 2026 517 2038
rect 547 2564 613 2576
rect 547 2038 563 2564
rect 597 2038 613 2564
rect 547 2026 613 2038
rect 643 2564 709 2576
rect 643 2038 659 2564
rect 693 2038 709 2564
rect 643 2026 709 2038
rect 739 2564 805 2576
rect 739 2038 755 2564
rect 789 2038 805 2564
rect 739 2026 805 2038
rect 835 2564 901 2576
rect 835 2038 851 2564
rect 885 2038 901 2564
rect 835 2026 901 2038
rect 931 2564 997 2576
rect 931 2038 947 2564
rect 981 2038 997 2564
rect 931 2026 997 2038
rect 1027 2564 1089 2576
rect 1027 2038 1043 2564
rect 1077 2038 1089 2564
rect 1027 2026 1089 2038
rect 1119 2564 1177 2576
rect 1119 2038 1131 2564
rect 1165 2038 1177 2564
rect 1119 2026 1177 2038
rect 11773 1997 11835 2009
rect 11773 1765 11785 1997
rect 11819 1765 11835 1997
rect 11773 1753 11835 1765
rect 11865 1997 11931 2009
rect 11865 1765 11881 1997
rect 11915 1765 11931 1997
rect 11865 1753 11931 1765
rect 11961 1997 12027 2009
rect 11961 1765 11977 1997
rect 12011 1765 12027 1997
rect 11961 1753 12027 1765
rect 12057 1997 12123 2009
rect 12057 1765 12073 1997
rect 12107 1765 12123 1997
rect 12057 1753 12123 1765
rect 12153 1997 12219 2009
rect 12153 1765 12169 1997
rect 12203 1765 12219 1997
rect 12153 1753 12219 1765
rect 12249 1997 12315 2009
rect 12249 1765 12265 1997
rect 12299 1765 12315 1997
rect 12249 1753 12315 1765
rect 12345 1997 12411 2009
rect 12345 1765 12361 1997
rect 12395 1765 12411 1997
rect 12345 1753 12411 1765
rect 12441 1997 12507 2009
rect 12441 1765 12457 1997
rect 12491 1765 12507 1997
rect 12441 1753 12507 1765
rect 12537 1997 12603 2009
rect 12537 1765 12553 1997
rect 12587 1765 12603 1997
rect 12537 1753 12603 1765
rect 12633 1997 12699 2009
rect 12633 1765 12649 1997
rect 12683 1765 12699 1997
rect 12633 1753 12699 1765
rect 12729 1997 12791 2009
rect 12729 1765 12745 1997
rect 12779 1765 12791 1997
rect 12923 1893 13137 1905
rect 12729 1753 12791 1765
rect -24597 863 -24535 875
rect -24597 673 -24585 863
rect -24551 673 -24535 863
rect -24597 661 -24535 673
rect -24505 863 -24439 875
rect -24505 673 -24489 863
rect -24455 673 -24439 863
rect -24505 661 -24439 673
rect -24409 863 -24343 875
rect -24409 673 -24393 863
rect -24359 673 -24343 863
rect -24409 661 -24343 673
rect -24313 863 -24247 875
rect -24313 673 -24297 863
rect -24263 673 -24247 863
rect -24313 661 -24247 673
rect -24217 863 -24151 875
rect -24217 673 -24201 863
rect -24167 673 -24151 863
rect -24217 661 -24151 673
rect -24121 863 -24055 875
rect -24121 673 -24105 863
rect -24071 673 -24055 863
rect -24121 661 -24055 673
rect -24025 863 -23963 875
rect -24025 673 -24009 863
rect -23975 673 -23963 863
rect -24025 661 -23963 673
rect -23488 863 -23426 875
rect -23488 673 -23476 863
rect -23442 673 -23426 863
rect -23488 661 -23426 673
rect -23396 863 -23330 875
rect -23396 673 -23380 863
rect -23346 673 -23330 863
rect -23396 661 -23330 673
rect -23300 863 -23234 875
rect -23300 673 -23284 863
rect -23250 673 -23234 863
rect -23300 661 -23234 673
rect -23204 863 -23138 875
rect -23204 673 -23188 863
rect -23154 673 -23138 863
rect -23204 661 -23138 673
rect -23108 863 -23042 875
rect -23108 673 -23092 863
rect -23058 673 -23042 863
rect -23108 661 -23042 673
rect -23012 863 -22946 875
rect -23012 673 -22996 863
rect -22962 673 -22946 863
rect -23012 661 -22946 673
rect -22916 863 -22854 875
rect -22916 673 -22900 863
rect -22866 673 -22854 863
rect -22916 661 -22854 673
rect -22606 863 -22544 875
rect -22606 673 -22594 863
rect -22560 673 -22544 863
rect -22606 661 -22544 673
rect -22514 863 -22448 875
rect -22514 673 -22498 863
rect -22464 673 -22448 863
rect -22514 661 -22448 673
rect -22418 863 -22352 875
rect -22418 673 -22402 863
rect -22368 673 -22352 863
rect -22418 661 -22352 673
rect -22322 863 -22256 875
rect -22322 673 -22306 863
rect -22272 673 -22256 863
rect -22322 661 -22256 673
rect -22226 863 -22160 875
rect -22226 673 -22210 863
rect -22176 673 -22160 863
rect -22226 661 -22160 673
rect -22130 863 -22064 875
rect -22130 673 -22114 863
rect -22080 673 -22064 863
rect -22130 661 -22064 673
rect -22034 863 -21972 875
rect -22034 673 -22018 863
rect -21984 673 -21972 863
rect -22034 661 -21972 673
rect -21306 863 -21244 875
rect -21306 673 -21294 863
rect -21260 673 -21244 863
rect -21306 661 -21244 673
rect -21214 863 -21148 875
rect -21214 673 -21198 863
rect -21164 673 -21148 863
rect -21214 661 -21148 673
rect -21118 863 -21052 875
rect -21118 673 -21102 863
rect -21068 673 -21052 863
rect -21118 661 -21052 673
rect -21022 863 -20956 875
rect -21022 673 -21006 863
rect -20972 673 -20956 863
rect -21022 661 -20956 673
rect -20926 863 -20860 875
rect -20926 673 -20910 863
rect -20876 673 -20860 863
rect -20926 661 -20860 673
rect -20830 863 -20764 875
rect -20830 673 -20814 863
rect -20780 673 -20764 863
rect -20830 661 -20764 673
rect -20734 863 -20672 875
rect -20734 673 -20718 863
rect -20684 673 -20672 863
rect -20734 661 -20672 673
rect -20197 863 -20135 875
rect -20197 673 -20185 863
rect -20151 673 -20135 863
rect -20197 661 -20135 673
rect -20105 863 -20039 875
rect -20105 673 -20089 863
rect -20055 673 -20039 863
rect -20105 661 -20039 673
rect -20009 863 -19943 875
rect -20009 673 -19993 863
rect -19959 673 -19943 863
rect -20009 661 -19943 673
rect -19913 863 -19847 875
rect -19913 673 -19897 863
rect -19863 673 -19847 863
rect -19913 661 -19847 673
rect -19817 863 -19751 875
rect -19817 673 -19801 863
rect -19767 673 -19751 863
rect -19817 661 -19751 673
rect -19721 863 -19655 875
rect -19721 673 -19705 863
rect -19671 673 -19655 863
rect -19721 661 -19655 673
rect -19625 863 -19563 875
rect -19625 673 -19609 863
rect -19575 673 -19563 863
rect -19625 661 -19563 673
rect -19315 863 -19253 875
rect -19315 673 -19303 863
rect -19269 673 -19253 863
rect -19315 661 -19253 673
rect -19223 863 -19157 875
rect -19223 673 -19207 863
rect -19173 673 -19157 863
rect -19223 661 -19157 673
rect -19127 863 -19061 875
rect -19127 673 -19111 863
rect -19077 673 -19061 863
rect -19127 661 -19061 673
rect -19031 863 -18965 875
rect -19031 673 -19015 863
rect -18981 673 -18965 863
rect -19031 661 -18965 673
rect -18935 863 -18869 875
rect -18935 673 -18919 863
rect -18885 673 -18869 863
rect -18935 661 -18869 673
rect -18839 863 -18773 875
rect -18839 673 -18823 863
rect -18789 673 -18773 863
rect -18839 661 -18773 673
rect -18743 863 -18681 875
rect -18743 673 -18727 863
rect -18693 673 -18681 863
rect -18743 661 -18681 673
rect -18015 863 -17953 875
rect -18015 673 -18003 863
rect -17969 673 -17953 863
rect -18015 661 -17953 673
rect -17923 863 -17857 875
rect -17923 673 -17907 863
rect -17873 673 -17857 863
rect -17923 661 -17857 673
rect -17827 863 -17761 875
rect -17827 673 -17811 863
rect -17777 673 -17761 863
rect -17827 661 -17761 673
rect -17731 863 -17665 875
rect -17731 673 -17715 863
rect -17681 673 -17665 863
rect -17731 661 -17665 673
rect -17635 863 -17569 875
rect -17635 673 -17619 863
rect -17585 673 -17569 863
rect -17635 661 -17569 673
rect -17539 863 -17473 875
rect -17539 673 -17523 863
rect -17489 673 -17473 863
rect -17539 661 -17473 673
rect -17443 863 -17381 875
rect -17443 673 -17427 863
rect -17393 673 -17381 863
rect -17443 661 -17381 673
rect -16906 863 -16844 875
rect -16906 673 -16894 863
rect -16860 673 -16844 863
rect -16906 661 -16844 673
rect -16814 863 -16748 875
rect -16814 673 -16798 863
rect -16764 673 -16748 863
rect -16814 661 -16748 673
rect -16718 863 -16652 875
rect -16718 673 -16702 863
rect -16668 673 -16652 863
rect -16718 661 -16652 673
rect -16622 863 -16556 875
rect -16622 673 -16606 863
rect -16572 673 -16556 863
rect -16622 661 -16556 673
rect -16526 863 -16460 875
rect -16526 673 -16510 863
rect -16476 673 -16460 863
rect -16526 661 -16460 673
rect -16430 863 -16364 875
rect -16430 673 -16414 863
rect -16380 673 -16364 863
rect -16430 661 -16364 673
rect -16334 863 -16272 875
rect -16334 673 -16318 863
rect -16284 673 -16272 863
rect -16334 661 -16272 673
rect -16024 863 -15962 875
rect -16024 673 -16012 863
rect -15978 673 -15962 863
rect -16024 661 -15962 673
rect -15932 863 -15866 875
rect -15932 673 -15916 863
rect -15882 673 -15866 863
rect -15932 661 -15866 673
rect -15836 863 -15770 875
rect -15836 673 -15820 863
rect -15786 673 -15770 863
rect -15836 661 -15770 673
rect -15740 863 -15674 875
rect -15740 673 -15724 863
rect -15690 673 -15674 863
rect -15740 661 -15674 673
rect -15644 863 -15578 875
rect -15644 673 -15628 863
rect -15594 673 -15578 863
rect -15644 661 -15578 673
rect -15548 863 -15482 875
rect -15548 673 -15532 863
rect -15498 673 -15482 863
rect -15548 661 -15482 673
rect -15452 863 -15390 875
rect -15452 673 -15436 863
rect -15402 673 -15390 863
rect -15452 661 -15390 673
rect -14724 863 -14662 875
rect -14724 673 -14712 863
rect -14678 673 -14662 863
rect -14724 661 -14662 673
rect -14632 863 -14566 875
rect -14632 673 -14616 863
rect -14582 673 -14566 863
rect -14632 661 -14566 673
rect -14536 863 -14470 875
rect -14536 673 -14520 863
rect -14486 673 -14470 863
rect -14536 661 -14470 673
rect -14440 863 -14374 875
rect -14440 673 -14424 863
rect -14390 673 -14374 863
rect -14440 661 -14374 673
rect -14344 863 -14278 875
rect -14344 673 -14328 863
rect -14294 673 -14278 863
rect -14344 661 -14278 673
rect -14248 863 -14182 875
rect -14248 673 -14232 863
rect -14198 673 -14182 863
rect -14248 661 -14182 673
rect -14152 863 -14090 875
rect -14152 673 -14136 863
rect -14102 673 -14090 863
rect -14152 661 -14090 673
rect -13615 863 -13553 875
rect -13615 673 -13603 863
rect -13569 673 -13553 863
rect -13615 661 -13553 673
rect -13523 863 -13457 875
rect -13523 673 -13507 863
rect -13473 673 -13457 863
rect -13523 661 -13457 673
rect -13427 863 -13361 875
rect -13427 673 -13411 863
rect -13377 673 -13361 863
rect -13427 661 -13361 673
rect -13331 863 -13265 875
rect -13331 673 -13315 863
rect -13281 673 -13265 863
rect -13331 661 -13265 673
rect -13235 863 -13169 875
rect -13235 673 -13219 863
rect -13185 673 -13169 863
rect -13235 661 -13169 673
rect -13139 863 -13073 875
rect -13139 673 -13123 863
rect -13089 673 -13073 863
rect -13139 661 -13073 673
rect -13043 863 -12981 875
rect -13043 673 -13027 863
rect -12993 673 -12981 863
rect -13043 661 -12981 673
rect -12733 863 -12671 875
rect -12733 673 -12721 863
rect -12687 673 -12671 863
rect -12733 661 -12671 673
rect -12641 863 -12575 875
rect -12641 673 -12625 863
rect -12591 673 -12575 863
rect -12641 661 -12575 673
rect -12545 863 -12479 875
rect -12545 673 -12529 863
rect -12495 673 -12479 863
rect -12545 661 -12479 673
rect -12449 863 -12383 875
rect -12449 673 -12433 863
rect -12399 673 -12383 863
rect -12449 661 -12383 673
rect -12353 863 -12287 875
rect -12353 673 -12337 863
rect -12303 673 -12287 863
rect -12353 661 -12287 673
rect -12257 863 -12191 875
rect -12257 673 -12241 863
rect -12207 673 -12191 863
rect -12257 661 -12191 673
rect -12161 863 -12099 875
rect -12161 673 -12145 863
rect -12111 673 -12099 863
rect -12161 661 -12099 673
rect -11433 863 -11371 875
rect -11433 673 -11421 863
rect -11387 673 -11371 863
rect -11433 661 -11371 673
rect -11341 863 -11275 875
rect -11341 673 -11325 863
rect -11291 673 -11275 863
rect -11341 661 -11275 673
rect -11245 863 -11179 875
rect -11245 673 -11229 863
rect -11195 673 -11179 863
rect -11245 661 -11179 673
rect -11149 863 -11083 875
rect -11149 673 -11133 863
rect -11099 673 -11083 863
rect -11149 661 -11083 673
rect -11053 863 -10987 875
rect -11053 673 -11037 863
rect -11003 673 -10987 863
rect -11053 661 -10987 673
rect -10957 863 -10891 875
rect -10957 673 -10941 863
rect -10907 673 -10891 863
rect -10957 661 -10891 673
rect -10861 863 -10799 875
rect -10861 673 -10845 863
rect -10811 673 -10799 863
rect -10861 661 -10799 673
rect -10324 863 -10262 875
rect -10324 673 -10312 863
rect -10278 673 -10262 863
rect -10324 661 -10262 673
rect -10232 863 -10166 875
rect -10232 673 -10216 863
rect -10182 673 -10166 863
rect -10232 661 -10166 673
rect -10136 863 -10070 875
rect -10136 673 -10120 863
rect -10086 673 -10070 863
rect -10136 661 -10070 673
rect -10040 863 -9974 875
rect -10040 673 -10024 863
rect -9990 673 -9974 863
rect -10040 661 -9974 673
rect -9944 863 -9878 875
rect -9944 673 -9928 863
rect -9894 673 -9878 863
rect -9944 661 -9878 673
rect -9848 863 -9782 875
rect -9848 673 -9832 863
rect -9798 673 -9782 863
rect -9848 661 -9782 673
rect -9752 863 -9690 875
rect -9752 673 -9736 863
rect -9702 673 -9690 863
rect -9752 661 -9690 673
rect -9442 863 -9380 875
rect -9442 673 -9430 863
rect -9396 673 -9380 863
rect -9442 661 -9380 673
rect -9350 863 -9284 875
rect -9350 673 -9334 863
rect -9300 673 -9284 863
rect -9350 661 -9284 673
rect -9254 863 -9188 875
rect -9254 673 -9238 863
rect -9204 673 -9188 863
rect -9254 661 -9188 673
rect -9158 863 -9092 875
rect -9158 673 -9142 863
rect -9108 673 -9092 863
rect -9158 661 -9092 673
rect -9062 863 -8996 875
rect -9062 673 -9046 863
rect -9012 673 -8996 863
rect -9062 661 -8996 673
rect -8966 863 -8900 875
rect -8966 673 -8950 863
rect -8916 673 -8900 863
rect -8966 661 -8900 673
rect -8870 863 -8808 875
rect -8870 673 -8854 863
rect -8820 673 -8808 863
rect -8870 661 -8808 673
rect -8143 863 -8081 875
rect -8143 673 -8131 863
rect -8097 673 -8081 863
rect -8143 661 -8081 673
rect -8051 863 -7985 875
rect -8051 673 -8035 863
rect -8001 673 -7985 863
rect -8051 661 -7985 673
rect -7955 863 -7889 875
rect -7955 673 -7939 863
rect -7905 673 -7889 863
rect -7955 661 -7889 673
rect -7859 863 -7793 875
rect -7859 673 -7843 863
rect -7809 673 -7793 863
rect -7859 661 -7793 673
rect -7763 863 -7697 875
rect -7763 673 -7747 863
rect -7713 673 -7697 863
rect -7763 661 -7697 673
rect -7667 863 -7601 875
rect -7667 673 -7651 863
rect -7617 673 -7601 863
rect -7667 661 -7601 673
rect -7571 863 -7509 875
rect -7571 673 -7555 863
rect -7521 673 -7509 863
rect -7571 661 -7509 673
rect -7034 863 -6972 875
rect -7034 673 -7022 863
rect -6988 673 -6972 863
rect -7034 661 -6972 673
rect -6942 863 -6876 875
rect -6942 673 -6926 863
rect -6892 673 -6876 863
rect -6942 661 -6876 673
rect -6846 863 -6780 875
rect -6846 673 -6830 863
rect -6796 673 -6780 863
rect -6846 661 -6780 673
rect -6750 863 -6684 875
rect -6750 673 -6734 863
rect -6700 673 -6684 863
rect -6750 661 -6684 673
rect -6654 863 -6588 875
rect -6654 673 -6638 863
rect -6604 673 -6588 863
rect -6654 661 -6588 673
rect -6558 863 -6492 875
rect -6558 673 -6542 863
rect -6508 673 -6492 863
rect -6558 661 -6492 673
rect -6462 863 -6400 875
rect -6462 673 -6446 863
rect -6412 673 -6400 863
rect -6462 661 -6400 673
rect -6152 863 -6090 875
rect -6152 673 -6140 863
rect -6106 673 -6090 863
rect -6152 661 -6090 673
rect -6060 863 -5994 875
rect -6060 673 -6044 863
rect -6010 673 -5994 863
rect -6060 661 -5994 673
rect -5964 863 -5898 875
rect -5964 673 -5948 863
rect -5914 673 -5898 863
rect -5964 661 -5898 673
rect -5868 863 -5802 875
rect -5868 673 -5852 863
rect -5818 673 -5802 863
rect -5868 661 -5802 673
rect -5772 863 -5706 875
rect -5772 673 -5756 863
rect -5722 673 -5706 863
rect -5772 661 -5706 673
rect -5676 863 -5610 875
rect -5676 673 -5660 863
rect -5626 673 -5610 863
rect -5676 661 -5610 673
rect -5580 863 -5518 875
rect -5580 673 -5564 863
rect -5530 673 -5518 863
rect -5580 661 -5518 673
rect -4852 863 -4790 875
rect -4852 673 -4840 863
rect -4806 673 -4790 863
rect -4852 661 -4790 673
rect -4760 863 -4694 875
rect -4760 673 -4744 863
rect -4710 673 -4694 863
rect -4760 661 -4694 673
rect -4664 863 -4598 875
rect -4664 673 -4648 863
rect -4614 673 -4598 863
rect -4664 661 -4598 673
rect -4568 863 -4502 875
rect -4568 673 -4552 863
rect -4518 673 -4502 863
rect -4568 661 -4502 673
rect -4472 863 -4406 875
rect -4472 673 -4456 863
rect -4422 673 -4406 863
rect -4472 661 -4406 673
rect -4376 863 -4310 875
rect -4376 673 -4360 863
rect -4326 673 -4310 863
rect -4376 661 -4310 673
rect -4280 863 -4218 875
rect -4280 673 -4264 863
rect -4230 673 -4218 863
rect -4280 661 -4218 673
rect -3743 863 -3681 875
rect -3743 673 -3731 863
rect -3697 673 -3681 863
rect -3743 661 -3681 673
rect -3651 863 -3585 875
rect -3651 673 -3635 863
rect -3601 673 -3585 863
rect -3651 661 -3585 673
rect -3555 863 -3489 875
rect -3555 673 -3539 863
rect -3505 673 -3489 863
rect -3555 661 -3489 673
rect -3459 863 -3393 875
rect -3459 673 -3443 863
rect -3409 673 -3393 863
rect -3459 661 -3393 673
rect -3363 863 -3297 875
rect -3363 673 -3347 863
rect -3313 673 -3297 863
rect -3363 661 -3297 673
rect -3267 863 -3201 875
rect -3267 673 -3251 863
rect -3217 673 -3201 863
rect -3267 661 -3201 673
rect -3171 863 -3109 875
rect -3171 673 -3155 863
rect -3121 673 -3109 863
rect -3171 661 -3109 673
rect -2861 863 -2799 875
rect -2861 673 -2849 863
rect -2815 673 -2799 863
rect -2861 661 -2799 673
rect -2769 863 -2703 875
rect -2769 673 -2753 863
rect -2719 673 -2703 863
rect -2769 661 -2703 673
rect -2673 863 -2607 875
rect -2673 673 -2657 863
rect -2623 673 -2607 863
rect -2673 661 -2607 673
rect -2577 863 -2511 875
rect -2577 673 -2561 863
rect -2527 673 -2511 863
rect -2577 661 -2511 673
rect -2481 863 -2415 875
rect -2481 673 -2465 863
rect -2431 673 -2415 863
rect -2481 661 -2415 673
rect -2385 863 -2319 875
rect -2385 673 -2369 863
rect -2335 673 -2319 863
rect -2385 661 -2319 673
rect -2289 863 -2227 875
rect -2289 673 -2273 863
rect -2239 673 -2227 863
rect -2289 661 -2227 673
rect -1561 863 -1499 875
rect -1561 673 -1549 863
rect -1515 673 -1499 863
rect -1561 661 -1499 673
rect -1469 863 -1403 875
rect -1469 673 -1453 863
rect -1419 673 -1403 863
rect -1469 661 -1403 673
rect -1373 863 -1307 875
rect -1373 673 -1357 863
rect -1323 673 -1307 863
rect -1373 661 -1307 673
rect -1277 863 -1211 875
rect -1277 673 -1261 863
rect -1227 673 -1211 863
rect -1277 661 -1211 673
rect -1181 863 -1115 875
rect -1181 673 -1165 863
rect -1131 673 -1115 863
rect -1181 661 -1115 673
rect -1085 863 -1019 875
rect -1085 673 -1069 863
rect -1035 673 -1019 863
rect -1085 661 -1019 673
rect -989 863 -927 875
rect -989 673 -973 863
rect -939 673 -927 863
rect -989 661 -927 673
rect -452 863 -390 875
rect -452 673 -440 863
rect -406 673 -390 863
rect -452 661 -390 673
rect -360 863 -294 875
rect -360 673 -344 863
rect -310 673 -294 863
rect -360 661 -294 673
rect -264 863 -198 875
rect -264 673 -248 863
rect -214 673 -198 863
rect -264 661 -198 673
rect -168 863 -102 875
rect -168 673 -152 863
rect -118 673 -102 863
rect -168 661 -102 673
rect -72 863 -6 875
rect -72 673 -56 863
rect -22 673 -6 863
rect -72 661 -6 673
rect 24 863 90 875
rect 24 673 40 863
rect 74 673 90 863
rect 24 661 90 673
rect 120 863 182 875
rect 120 673 136 863
rect 170 673 182 863
rect 120 661 182 673
rect 430 863 492 875
rect 430 673 442 863
rect 476 673 492 863
rect 430 661 492 673
rect 522 863 588 875
rect 522 673 538 863
rect 572 673 588 863
rect 522 661 588 673
rect 618 863 684 875
rect 618 673 634 863
rect 668 673 684 863
rect 618 661 684 673
rect 714 863 780 875
rect 714 673 730 863
rect 764 673 780 863
rect 714 661 780 673
rect 810 863 876 875
rect 810 673 826 863
rect 860 673 876 863
rect 810 661 876 673
rect 906 863 972 875
rect 906 673 922 863
rect 956 673 972 863
rect 906 661 972 673
rect 1002 863 1064 875
rect 1002 673 1018 863
rect 1052 673 1064 863
rect 1002 661 1064 673
rect 12923 1859 12935 1893
rect 13125 1859 13137 1893
rect 12923 1843 13137 1859
rect 12923 1797 13137 1813
rect 12923 1763 12935 1797
rect 13129 1763 13137 1797
rect 12923 1747 13137 1763
rect 12923 1701 13137 1717
rect 12923 1667 12935 1701
rect 13125 1667 13137 1701
rect 12923 1651 13137 1667
rect 12923 1605 13137 1621
rect 12923 1571 12935 1605
rect 13129 1571 13137 1605
rect 12923 1559 13137 1571
rect 7138 343 7200 355
rect 7138 45 7150 343
rect 7184 45 7200 343
rect 7138 33 7200 45
rect 7230 343 7296 355
rect 7230 45 7246 343
rect 7280 45 7296 343
rect 7230 33 7296 45
rect 7326 343 7392 355
rect 7326 45 7342 343
rect 7376 45 7392 343
rect 7326 33 7392 45
rect 7422 343 7488 355
rect 7422 45 7438 343
rect 7472 45 7488 343
rect 7422 33 7488 45
rect 7518 343 7584 355
rect 7518 45 7534 343
rect 7568 45 7584 343
rect 7518 33 7584 45
rect 7614 343 7680 355
rect 7614 45 7630 343
rect 7664 45 7680 343
rect 7614 33 7680 45
rect 7710 343 7776 355
rect 7710 45 7726 343
rect 7760 45 7776 343
rect 7710 33 7776 45
rect 7806 343 7872 355
rect 7806 45 7822 343
rect 7856 45 7872 343
rect 7806 33 7872 45
rect 7902 343 7964 355
rect 7902 45 7918 343
rect 7952 45 7964 343
rect 7902 33 7964 45
rect 8086 343 8148 355
rect 8086 45 8098 343
rect 8132 45 8148 343
rect 8086 33 8148 45
rect 8178 343 8244 355
rect 8178 45 8194 343
rect 8228 45 8244 343
rect 8178 33 8244 45
rect 8274 343 8340 355
rect 8274 45 8290 343
rect 8324 45 8340 343
rect 8274 33 8340 45
rect 8370 343 8436 355
rect 8370 45 8386 343
rect 8420 45 8436 343
rect 8370 33 8436 45
rect 8466 343 8532 355
rect 8466 45 8482 343
rect 8516 45 8532 343
rect 8466 33 8532 45
rect 8562 343 8628 355
rect 8562 45 8578 343
rect 8612 45 8628 343
rect 8562 33 8628 45
rect 8658 343 8724 355
rect 8658 45 8674 343
rect 8708 45 8724 343
rect 8658 33 8724 45
rect 8754 343 8820 355
rect 8754 45 8770 343
rect 8804 45 8820 343
rect 8754 33 8820 45
rect 8850 343 8912 355
rect 8850 45 8866 343
rect 8900 45 8912 343
rect 8850 33 8912 45
rect 9022 343 9084 355
rect 9022 45 9034 343
rect 9068 45 9084 343
rect 9022 33 9084 45
rect 9114 343 9180 355
rect 9114 45 9130 343
rect 9164 45 9180 343
rect 9114 33 9180 45
rect 9210 343 9276 355
rect 9210 45 9226 343
rect 9260 45 9276 343
rect 9210 33 9276 45
rect 9306 343 9372 355
rect 9306 45 9322 343
rect 9356 45 9372 343
rect 9306 33 9372 45
rect 9402 343 9468 355
rect 9402 45 9418 343
rect 9452 45 9468 343
rect 9402 33 9468 45
rect 9498 343 9564 355
rect 9498 45 9514 343
rect 9548 45 9564 343
rect 9498 33 9564 45
rect 9594 343 9660 355
rect 9594 45 9610 343
rect 9644 45 9660 343
rect 9594 33 9660 45
rect 9690 343 9756 355
rect 9690 45 9706 343
rect 9740 45 9756 343
rect 9690 33 9756 45
rect 9786 343 9848 355
rect 9786 45 9802 343
rect 9836 45 9848 343
rect 9786 33 9848 45
rect 9953 344 10015 356
rect 9953 46 9965 344
rect 9999 46 10015 344
rect 9953 34 10015 46
rect 10045 344 10111 356
rect 10045 46 10061 344
rect 10095 46 10111 344
rect 10045 34 10111 46
rect 10141 344 10207 356
rect 10141 46 10157 344
rect 10191 46 10207 344
rect 10141 34 10207 46
rect 10237 344 10303 356
rect 10237 46 10253 344
rect 10287 46 10303 344
rect 10237 34 10303 46
rect 10333 344 10399 356
rect 10333 46 10349 344
rect 10383 46 10399 344
rect 10333 34 10399 46
rect 10429 344 10495 356
rect 10429 46 10445 344
rect 10479 46 10495 344
rect 10429 34 10495 46
rect 10525 344 10591 356
rect 10525 46 10541 344
rect 10575 46 10591 344
rect 10525 34 10591 46
rect 10621 344 10687 356
rect 10621 46 10637 344
rect 10671 46 10687 344
rect 10621 34 10687 46
rect 10717 344 10779 356
rect 10717 46 10733 344
rect 10767 46 10779 344
rect 10717 34 10779 46
rect 10880 343 10942 355
rect 10880 45 10892 343
rect 10926 45 10942 343
rect 10880 33 10942 45
rect 10972 343 11038 355
rect 10972 45 10988 343
rect 11022 45 11038 343
rect 10972 33 11038 45
rect 11068 343 11134 355
rect 11068 45 11084 343
rect 11118 45 11134 343
rect 11068 33 11134 45
rect 11164 343 11230 355
rect 11164 45 11180 343
rect 11214 45 11230 343
rect 11164 33 11230 45
rect 11260 343 11326 355
rect 11260 45 11276 343
rect 11310 45 11326 343
rect 11260 33 11326 45
rect 11356 343 11422 355
rect 11356 45 11372 343
rect 11406 45 11422 343
rect 11356 33 11422 45
rect 11452 343 11518 355
rect 11452 45 11468 343
rect 11502 45 11518 343
rect 11452 33 11518 45
rect 11548 343 11614 355
rect 11548 45 11564 343
rect 11598 45 11614 343
rect 11548 33 11614 45
rect 11644 343 11706 355
rect 11644 45 11660 343
rect 11694 45 11706 343
rect 11644 33 11706 45
rect 5658 -617 5872 -605
rect 5658 -651 5670 -617
rect 5860 -651 5872 -617
rect 6098 -617 6312 -605
rect 5658 -667 5872 -651
rect 5658 -713 5872 -697
rect 5658 -747 5670 -713
rect 5864 -747 5872 -713
rect 5658 -763 5872 -747
rect 5658 -809 5872 -793
rect 5658 -843 5670 -809
rect 5860 -843 5872 -809
rect 5658 -859 5872 -843
rect 5658 -905 5872 -889
rect 5658 -939 5670 -905
rect 5864 -939 5872 -905
rect 6098 -651 6110 -617
rect 6300 -651 6312 -617
rect 6538 -617 6752 -605
rect 6098 -667 6312 -651
rect 6098 -713 6312 -697
rect 6098 -747 6110 -713
rect 6304 -747 6312 -713
rect 6098 -763 6312 -747
rect 6098 -809 6312 -793
rect 6098 -843 6110 -809
rect 6300 -843 6312 -809
rect 6098 -859 6312 -843
rect 6098 -905 6312 -889
rect 5658 -951 5872 -939
rect 6098 -939 6110 -905
rect 6304 -939 6312 -905
rect 6538 -651 6550 -617
rect 6740 -651 6752 -617
rect 6538 -667 6752 -651
rect 6538 -713 6752 -697
rect 6538 -747 6550 -713
rect 6744 -747 6752 -713
rect 6538 -763 6752 -747
rect 6538 -809 6752 -793
rect 6538 -843 6550 -809
rect 6740 -843 6752 -809
rect 6538 -859 6752 -843
rect 6538 -905 6752 -889
rect 6098 -951 6312 -939
rect 6538 -939 6550 -905
rect 6744 -939 6752 -905
rect 6538 -951 6752 -939
rect 7138 -1321 7200 -1309
rect 7138 -1619 7150 -1321
rect 7184 -1619 7200 -1321
rect 7138 -1631 7200 -1619
rect 7230 -1321 7296 -1309
rect 7230 -1619 7246 -1321
rect 7280 -1619 7296 -1321
rect 7230 -1631 7296 -1619
rect 7326 -1321 7392 -1309
rect 7326 -1619 7342 -1321
rect 7376 -1619 7392 -1321
rect 7326 -1631 7392 -1619
rect 7422 -1321 7488 -1309
rect 7422 -1619 7438 -1321
rect 7472 -1619 7488 -1321
rect 7422 -1631 7488 -1619
rect 7518 -1321 7584 -1309
rect 7518 -1619 7534 -1321
rect 7568 -1619 7584 -1321
rect 7518 -1631 7584 -1619
rect 7614 -1321 7680 -1309
rect 7614 -1619 7630 -1321
rect 7664 -1619 7680 -1321
rect 7614 -1631 7680 -1619
rect 7710 -1321 7776 -1309
rect 7710 -1619 7726 -1321
rect 7760 -1619 7776 -1321
rect 7710 -1631 7776 -1619
rect 7806 -1321 7872 -1309
rect 7806 -1619 7822 -1321
rect 7856 -1619 7872 -1321
rect 7806 -1631 7872 -1619
rect 7902 -1321 7964 -1309
rect 7902 -1619 7918 -1321
rect 7952 -1619 7964 -1321
rect 7902 -1631 7964 -1619
rect 8086 -1321 8148 -1309
rect 8086 -1619 8098 -1321
rect 8132 -1619 8148 -1321
rect 8086 -1631 8148 -1619
rect 8178 -1321 8244 -1309
rect 8178 -1619 8194 -1321
rect 8228 -1619 8244 -1321
rect 8178 -1631 8244 -1619
rect 8274 -1321 8340 -1309
rect 8274 -1619 8290 -1321
rect 8324 -1619 8340 -1321
rect 8274 -1631 8340 -1619
rect 8370 -1321 8436 -1309
rect 8370 -1619 8386 -1321
rect 8420 -1619 8436 -1321
rect 8370 -1631 8436 -1619
rect 8466 -1321 8532 -1309
rect 8466 -1619 8482 -1321
rect 8516 -1619 8532 -1321
rect 8466 -1631 8532 -1619
rect 8562 -1321 8628 -1309
rect 8562 -1619 8578 -1321
rect 8612 -1619 8628 -1321
rect 8562 -1631 8628 -1619
rect 8658 -1321 8724 -1309
rect 8658 -1619 8674 -1321
rect 8708 -1619 8724 -1321
rect 8658 -1631 8724 -1619
rect 8754 -1321 8820 -1309
rect 8754 -1619 8770 -1321
rect 8804 -1619 8820 -1321
rect 8754 -1631 8820 -1619
rect 8850 -1321 8912 -1309
rect 8850 -1619 8866 -1321
rect 8900 -1619 8912 -1321
rect 8850 -1631 8912 -1619
rect 9022 -1321 9084 -1309
rect 9022 -1619 9034 -1321
rect 9068 -1619 9084 -1321
rect 9022 -1631 9084 -1619
rect 9114 -1321 9180 -1309
rect 9114 -1619 9130 -1321
rect 9164 -1619 9180 -1321
rect 9114 -1631 9180 -1619
rect 9210 -1321 9276 -1309
rect 9210 -1619 9226 -1321
rect 9260 -1619 9276 -1321
rect 9210 -1631 9276 -1619
rect 9306 -1321 9372 -1309
rect 9306 -1619 9322 -1321
rect 9356 -1619 9372 -1321
rect 9306 -1631 9372 -1619
rect 9402 -1321 9468 -1309
rect 9402 -1619 9418 -1321
rect 9452 -1619 9468 -1321
rect 9402 -1631 9468 -1619
rect 9498 -1321 9564 -1309
rect 9498 -1619 9514 -1321
rect 9548 -1619 9564 -1321
rect 9498 -1631 9564 -1619
rect 9594 -1321 9660 -1309
rect 9594 -1619 9610 -1321
rect 9644 -1619 9660 -1321
rect 9594 -1631 9660 -1619
rect 9690 -1321 9756 -1309
rect 9690 -1619 9706 -1321
rect 9740 -1619 9756 -1321
rect 9690 -1631 9756 -1619
rect 9786 -1321 9848 -1309
rect 9786 -1619 9802 -1321
rect 9836 -1619 9848 -1321
rect 9786 -1631 9848 -1619
rect 9953 -1321 10015 -1309
rect 9953 -1619 9965 -1321
rect 9999 -1619 10015 -1321
rect 9953 -1631 10015 -1619
rect 10045 -1321 10111 -1309
rect 10045 -1619 10061 -1321
rect 10095 -1619 10111 -1321
rect 10045 -1631 10111 -1619
rect 10141 -1321 10207 -1309
rect 10141 -1619 10157 -1321
rect 10191 -1619 10207 -1321
rect 10141 -1631 10207 -1619
rect 10237 -1321 10303 -1309
rect 10237 -1619 10253 -1321
rect 10287 -1619 10303 -1321
rect 10237 -1631 10303 -1619
rect 10333 -1321 10399 -1309
rect 10333 -1619 10349 -1321
rect 10383 -1619 10399 -1321
rect 10333 -1631 10399 -1619
rect 10429 -1321 10495 -1309
rect 10429 -1619 10445 -1321
rect 10479 -1619 10495 -1321
rect 10429 -1631 10495 -1619
rect 10525 -1321 10591 -1309
rect 10525 -1619 10541 -1321
rect 10575 -1619 10591 -1321
rect 10525 -1631 10591 -1619
rect 10621 -1321 10687 -1309
rect 10621 -1619 10637 -1321
rect 10671 -1619 10687 -1321
rect 10621 -1631 10687 -1619
rect 10717 -1321 10779 -1309
rect 10717 -1619 10733 -1321
rect 10767 -1619 10779 -1321
rect 10717 -1631 10779 -1619
rect 10880 -1321 10942 -1309
rect 10880 -1619 10892 -1321
rect 10926 -1619 10942 -1321
rect 10880 -1631 10942 -1619
rect 10972 -1321 11038 -1309
rect 10972 -1619 10988 -1321
rect 11022 -1619 11038 -1321
rect 10972 -1631 11038 -1619
rect 11068 -1321 11134 -1309
rect 11068 -1619 11084 -1321
rect 11118 -1619 11134 -1321
rect 11068 -1631 11134 -1619
rect 11164 -1321 11230 -1309
rect 11164 -1619 11180 -1321
rect 11214 -1619 11230 -1321
rect 11164 -1631 11230 -1619
rect 11260 -1321 11326 -1309
rect 11260 -1619 11276 -1321
rect 11310 -1619 11326 -1321
rect 11260 -1631 11326 -1619
rect 11356 -1321 11422 -1309
rect 11356 -1619 11372 -1321
rect 11406 -1619 11422 -1321
rect 11356 -1631 11422 -1619
rect 11452 -1321 11518 -1309
rect 11452 -1619 11468 -1321
rect 11502 -1619 11518 -1321
rect 11452 -1631 11518 -1619
rect 11548 -1321 11614 -1309
rect 11548 -1619 11564 -1321
rect 11598 -1619 11614 -1321
rect 11548 -1631 11614 -1619
rect 11644 -1321 11706 -1309
rect 11644 -1619 11660 -1321
rect 11694 -1619 11706 -1321
rect 11644 -1631 11706 -1619
rect -23628 -2319 -23414 -2307
rect -24447 -2425 -24385 -2413
rect -24447 -2615 -24435 -2425
rect -24401 -2615 -24385 -2425
rect -24447 -2627 -24385 -2615
rect -24355 -2425 -24289 -2413
rect -24355 -2615 -24339 -2425
rect -24305 -2615 -24289 -2425
rect -24355 -2627 -24289 -2615
rect -24259 -2425 -24193 -2413
rect -24259 -2615 -24243 -2425
rect -24209 -2615 -24193 -2425
rect -24259 -2627 -24193 -2615
rect -24163 -2425 -24097 -2413
rect -24163 -2615 -24147 -2425
rect -24113 -2615 -24097 -2425
rect -24163 -2627 -24097 -2615
rect -24067 -2425 -24001 -2413
rect -24067 -2615 -24051 -2425
rect -24017 -2615 -24001 -2425
rect -24067 -2627 -24001 -2615
rect -23971 -2425 -23905 -2413
rect -23971 -2615 -23955 -2425
rect -23921 -2615 -23905 -2425
rect -23971 -2627 -23905 -2615
rect -23875 -2425 -23813 -2413
rect -23875 -2615 -23859 -2425
rect -23825 -2615 -23813 -2425
rect -23628 -2353 -23616 -2319
rect -23426 -2353 -23414 -2319
rect -23628 -2369 -23414 -2353
rect -21608 -2319 -21394 -2307
rect -23628 -2415 -23414 -2399
rect -23628 -2449 -23616 -2415
rect -23422 -2449 -23414 -2415
rect -23628 -2465 -23414 -2449
rect -22410 -2425 -22348 -2413
rect -23628 -2511 -23414 -2495
rect -23628 -2545 -23616 -2511
rect -23426 -2545 -23414 -2511
rect -23628 -2561 -23414 -2545
rect -23628 -2607 -23414 -2591
rect -23875 -2627 -23813 -2615
rect -23628 -2641 -23616 -2607
rect -23422 -2641 -23414 -2607
rect -22410 -2615 -22398 -2425
rect -22364 -2615 -22348 -2425
rect -22410 -2627 -22348 -2615
rect -22318 -2425 -22252 -2413
rect -22318 -2615 -22302 -2425
rect -22268 -2615 -22252 -2425
rect -22318 -2627 -22252 -2615
rect -22222 -2425 -22156 -2413
rect -22222 -2615 -22206 -2425
rect -22172 -2615 -22156 -2425
rect -22222 -2627 -22156 -2615
rect -22126 -2425 -22060 -2413
rect -22126 -2615 -22110 -2425
rect -22076 -2615 -22060 -2425
rect -22126 -2627 -22060 -2615
rect -22030 -2425 -21964 -2413
rect -22030 -2615 -22014 -2425
rect -21980 -2615 -21964 -2425
rect -22030 -2627 -21964 -2615
rect -21934 -2425 -21868 -2413
rect -21934 -2615 -21918 -2425
rect -21884 -2615 -21868 -2425
rect -21934 -2627 -21868 -2615
rect -21838 -2425 -21776 -2413
rect -21838 -2615 -21822 -2425
rect -21788 -2615 -21776 -2425
rect -21608 -2353 -21596 -2319
rect -21406 -2353 -21394 -2319
rect -21608 -2369 -21394 -2353
rect -19867 -2319 -19653 -2307
rect -21608 -2415 -21394 -2399
rect -21608 -2449 -21596 -2415
rect -21402 -2449 -21394 -2415
rect -21608 -2465 -21394 -2449
rect -20680 -2425 -20618 -2413
rect -21608 -2511 -21394 -2495
rect -21608 -2545 -21596 -2511
rect -21406 -2545 -21394 -2511
rect -21608 -2561 -21394 -2545
rect -21608 -2607 -21394 -2591
rect -21838 -2627 -21776 -2615
rect -23628 -2653 -23414 -2641
rect -21608 -2641 -21596 -2607
rect -21402 -2641 -21394 -2607
rect -20680 -2615 -20668 -2425
rect -20634 -2615 -20618 -2425
rect -20680 -2627 -20618 -2615
rect -20588 -2425 -20522 -2413
rect -20588 -2615 -20572 -2425
rect -20538 -2615 -20522 -2425
rect -20588 -2627 -20522 -2615
rect -20492 -2425 -20426 -2413
rect -20492 -2615 -20476 -2425
rect -20442 -2615 -20426 -2425
rect -20492 -2627 -20426 -2615
rect -20396 -2425 -20330 -2413
rect -20396 -2615 -20380 -2425
rect -20346 -2615 -20330 -2425
rect -20396 -2627 -20330 -2615
rect -20300 -2425 -20234 -2413
rect -20300 -2615 -20284 -2425
rect -20250 -2615 -20234 -2425
rect -20300 -2627 -20234 -2615
rect -20204 -2425 -20138 -2413
rect -20204 -2615 -20188 -2425
rect -20154 -2615 -20138 -2425
rect -20204 -2627 -20138 -2615
rect -20108 -2425 -20046 -2413
rect -20108 -2615 -20092 -2425
rect -20058 -2615 -20046 -2425
rect -19867 -2353 -19855 -2319
rect -19665 -2353 -19653 -2319
rect -19867 -2369 -19653 -2353
rect -18088 -2319 -17874 -2307
rect -19867 -2415 -19653 -2399
rect -19867 -2449 -19855 -2415
rect -19661 -2449 -19653 -2415
rect -19867 -2465 -19653 -2449
rect -18920 -2425 -18858 -2413
rect -19867 -2511 -19653 -2495
rect -19867 -2545 -19855 -2511
rect -19665 -2545 -19653 -2511
rect -19867 -2561 -19653 -2545
rect -19867 -2607 -19653 -2591
rect -20108 -2627 -20046 -2615
rect -21608 -2653 -21394 -2641
rect -19867 -2641 -19855 -2607
rect -19661 -2641 -19653 -2607
rect -18920 -2615 -18908 -2425
rect -18874 -2615 -18858 -2425
rect -18920 -2627 -18858 -2615
rect -18828 -2425 -18762 -2413
rect -18828 -2615 -18812 -2425
rect -18778 -2615 -18762 -2425
rect -18828 -2627 -18762 -2615
rect -18732 -2425 -18666 -2413
rect -18732 -2615 -18716 -2425
rect -18682 -2615 -18666 -2425
rect -18732 -2627 -18666 -2615
rect -18636 -2425 -18570 -2413
rect -18636 -2615 -18620 -2425
rect -18586 -2615 -18570 -2425
rect -18636 -2627 -18570 -2615
rect -18540 -2425 -18474 -2413
rect -18540 -2615 -18524 -2425
rect -18490 -2615 -18474 -2425
rect -18540 -2627 -18474 -2615
rect -18444 -2425 -18378 -2413
rect -18444 -2615 -18428 -2425
rect -18394 -2615 -18378 -2425
rect -18444 -2627 -18378 -2615
rect -18348 -2425 -18286 -2413
rect -18348 -2615 -18332 -2425
rect -18298 -2615 -18286 -2425
rect -18088 -2353 -18076 -2319
rect -17886 -2353 -17874 -2319
rect -18088 -2369 -17874 -2353
rect -18088 -2415 -17874 -2399
rect -18088 -2449 -18076 -2415
rect -17882 -2449 -17874 -2415
rect -18088 -2465 -17874 -2449
rect -18088 -2511 -17874 -2495
rect -18088 -2545 -18076 -2511
rect -17886 -2545 -17874 -2511
rect -18088 -2561 -17874 -2545
rect -18088 -2607 -17874 -2591
rect -18348 -2627 -18286 -2615
rect -19867 -2653 -19653 -2641
rect -18088 -2641 -18076 -2607
rect -17882 -2641 -17874 -2607
rect -18088 -2653 -17874 -2641
rect 11773 -2531 11835 -2519
rect 11773 -2763 11785 -2531
rect 11819 -2763 11835 -2531
rect 11773 -2775 11835 -2763
rect 11865 -2531 11931 -2519
rect 11865 -2763 11881 -2531
rect 11915 -2763 11931 -2531
rect 11865 -2775 11931 -2763
rect 11961 -2531 12027 -2519
rect 11961 -2763 11977 -2531
rect 12011 -2763 12027 -2531
rect 11961 -2775 12027 -2763
rect 12057 -2531 12123 -2519
rect 12057 -2763 12073 -2531
rect 12107 -2763 12123 -2531
rect 12057 -2775 12123 -2763
rect 12153 -2531 12219 -2519
rect 12153 -2763 12169 -2531
rect 12203 -2763 12219 -2531
rect 12153 -2775 12219 -2763
rect 12249 -2531 12315 -2519
rect 12249 -2763 12265 -2531
rect 12299 -2763 12315 -2531
rect 12249 -2775 12315 -2763
rect 12345 -2531 12411 -2519
rect 12345 -2763 12361 -2531
rect 12395 -2763 12411 -2531
rect 12345 -2775 12411 -2763
rect 12441 -2531 12507 -2519
rect 12441 -2763 12457 -2531
rect 12491 -2763 12507 -2531
rect 12441 -2775 12507 -2763
rect 12537 -2531 12603 -2519
rect 12537 -2763 12553 -2531
rect 12587 -2763 12603 -2531
rect 12537 -2775 12603 -2763
rect 12633 -2531 12699 -2519
rect 12633 -2763 12649 -2531
rect 12683 -2763 12699 -2531
rect 12633 -2775 12699 -2763
rect 12729 -2531 12791 -2519
rect 12729 -2763 12745 -2531
rect 12779 -2763 12791 -2531
rect 12923 -2635 13137 -2623
rect 12729 -2775 12791 -2763
rect -20737 -3996 -20679 -3984
rect -23584 -4131 -23370 -4119
rect -24396 -4237 -24334 -4225
rect -24396 -4427 -24384 -4237
rect -24350 -4427 -24334 -4237
rect -24396 -4439 -24334 -4427
rect -24304 -4237 -24238 -4225
rect -24304 -4427 -24288 -4237
rect -24254 -4427 -24238 -4237
rect -24304 -4439 -24238 -4427
rect -24208 -4237 -24142 -4225
rect -24208 -4427 -24192 -4237
rect -24158 -4427 -24142 -4237
rect -24208 -4439 -24142 -4427
rect -24112 -4237 -24046 -4225
rect -24112 -4427 -24096 -4237
rect -24062 -4427 -24046 -4237
rect -24112 -4439 -24046 -4427
rect -24016 -4237 -23950 -4225
rect -24016 -4427 -24000 -4237
rect -23966 -4427 -23950 -4237
rect -24016 -4439 -23950 -4427
rect -23920 -4237 -23854 -4225
rect -23920 -4427 -23904 -4237
rect -23870 -4427 -23854 -4237
rect -23920 -4439 -23854 -4427
rect -23824 -4237 -23762 -4225
rect -23824 -4427 -23808 -4237
rect -23774 -4427 -23762 -4237
rect -23584 -4165 -23572 -4131
rect -23382 -4165 -23370 -4131
rect -23584 -4181 -23370 -4165
rect -21846 -4131 -21632 -4119
rect -23584 -4227 -23370 -4211
rect -23584 -4261 -23572 -4227
rect -23378 -4261 -23370 -4227
rect -23584 -4277 -23370 -4261
rect -22660 -4237 -22598 -4225
rect -23584 -4323 -23370 -4307
rect -23584 -4357 -23572 -4323
rect -23382 -4357 -23370 -4323
rect -23584 -4373 -23370 -4357
rect -23584 -4419 -23370 -4403
rect -23824 -4439 -23762 -4427
rect -23584 -4453 -23572 -4419
rect -23378 -4453 -23370 -4419
rect -22660 -4427 -22648 -4237
rect -22614 -4427 -22598 -4237
rect -22660 -4439 -22598 -4427
rect -22568 -4237 -22502 -4225
rect -22568 -4427 -22552 -4237
rect -22518 -4427 -22502 -4237
rect -22568 -4439 -22502 -4427
rect -22472 -4237 -22406 -4225
rect -22472 -4427 -22456 -4237
rect -22422 -4427 -22406 -4237
rect -22472 -4439 -22406 -4427
rect -22376 -4237 -22310 -4225
rect -22376 -4427 -22360 -4237
rect -22326 -4427 -22310 -4237
rect -22376 -4439 -22310 -4427
rect -22280 -4237 -22214 -4225
rect -22280 -4427 -22264 -4237
rect -22230 -4427 -22214 -4237
rect -22280 -4439 -22214 -4427
rect -22184 -4237 -22118 -4225
rect -22184 -4427 -22168 -4237
rect -22134 -4427 -22118 -4237
rect -22184 -4439 -22118 -4427
rect -22088 -4237 -22026 -4225
rect -22088 -4427 -22072 -4237
rect -22038 -4427 -22026 -4237
rect -21846 -4165 -21834 -4131
rect -21644 -4165 -21632 -4131
rect -21846 -4181 -21632 -4165
rect -21846 -4227 -21632 -4211
rect -21846 -4261 -21834 -4227
rect -21640 -4261 -21632 -4227
rect -21846 -4277 -21632 -4261
rect -21846 -4323 -21632 -4307
rect -21846 -4357 -21834 -4323
rect -21644 -4357 -21632 -4323
rect -21846 -4373 -21632 -4357
rect -21846 -4419 -21632 -4403
rect -22088 -4439 -22026 -4427
rect -23584 -4465 -23370 -4453
rect -21846 -4453 -21834 -4419
rect -21640 -4453 -21632 -4419
rect -21846 -4465 -21632 -4453
rect -20737 -4522 -20725 -3996
rect -20691 -4522 -20679 -3996
rect -20737 -4534 -20679 -4522
rect -20649 -3996 -20587 -3984
rect -20649 -4522 -20637 -3996
rect -20603 -4522 -20587 -3996
rect -20649 -4534 -20587 -4522
rect -20557 -3996 -20491 -3984
rect -20557 -4522 -20541 -3996
rect -20507 -4522 -20491 -3996
rect -20557 -4534 -20491 -4522
rect -20461 -3996 -20395 -3984
rect -20461 -4522 -20445 -3996
rect -20411 -4522 -20395 -3996
rect -20461 -4534 -20395 -4522
rect -20365 -3996 -20299 -3984
rect -20365 -4522 -20349 -3996
rect -20315 -4522 -20299 -3996
rect -20365 -4534 -20299 -4522
rect -20269 -3996 -20203 -3984
rect -20269 -4522 -20253 -3996
rect -20219 -4522 -20203 -3996
rect -20269 -4534 -20203 -4522
rect -20173 -3996 -20107 -3984
rect -20173 -4522 -20157 -3996
rect -20123 -4522 -20107 -3996
rect -20173 -4534 -20107 -4522
rect -20077 -3996 -20011 -3984
rect -20077 -4522 -20061 -3996
rect -20027 -4522 -20011 -3996
rect -20077 -4534 -20011 -4522
rect -19981 -3996 -19915 -3984
rect -19981 -4522 -19965 -3996
rect -19931 -4522 -19915 -3996
rect -19981 -4534 -19915 -4522
rect -19885 -3996 -19819 -3984
rect -19885 -4522 -19869 -3996
rect -19835 -4522 -19819 -3996
rect -19885 -4534 -19819 -4522
rect -19789 -3996 -19723 -3984
rect -19789 -4522 -19773 -3996
rect -19739 -4522 -19723 -3996
rect -19789 -4534 -19723 -4522
rect -19693 -3996 -19627 -3984
rect -19693 -4522 -19677 -3996
rect -19643 -4522 -19627 -3996
rect -19693 -4534 -19627 -4522
rect -19597 -3996 -19531 -3984
rect -19597 -4522 -19581 -3996
rect -19547 -4522 -19531 -3996
rect -19597 -4534 -19531 -4522
rect -19501 -3996 -19439 -3984
rect -19501 -4522 -19485 -3996
rect -19451 -4522 -19439 -3996
rect -19501 -4534 -19439 -4522
rect -19409 -3996 -19351 -3984
rect -19409 -4522 -19397 -3996
rect -19363 -4522 -19351 -3996
rect -19409 -4534 -19351 -4522
rect -19178 -3996 -19120 -3984
rect -19178 -4522 -19166 -3996
rect -19132 -4522 -19120 -3996
rect -19178 -4534 -19120 -4522
rect -19090 -3996 -19028 -3984
rect -19090 -4522 -19078 -3996
rect -19044 -4522 -19028 -3996
rect -19090 -4534 -19028 -4522
rect -18998 -3996 -18932 -3984
rect -18998 -4522 -18982 -3996
rect -18948 -4522 -18932 -3996
rect -18998 -4534 -18932 -4522
rect -18902 -3996 -18836 -3984
rect -18902 -4522 -18886 -3996
rect -18852 -4522 -18836 -3996
rect -18902 -4534 -18836 -4522
rect -18806 -3996 -18740 -3984
rect -18806 -4522 -18790 -3996
rect -18756 -4522 -18740 -3996
rect -18806 -4534 -18740 -4522
rect -18710 -3996 -18644 -3984
rect -18710 -4522 -18694 -3996
rect -18660 -4522 -18644 -3996
rect -18710 -4534 -18644 -4522
rect -18614 -3996 -18548 -3984
rect -18614 -4522 -18598 -3996
rect -18564 -4522 -18548 -3996
rect -18614 -4534 -18548 -4522
rect -18518 -3996 -18452 -3984
rect -18518 -4522 -18502 -3996
rect -18468 -4522 -18452 -3996
rect -18518 -4534 -18452 -4522
rect -18422 -3996 -18356 -3984
rect -18422 -4522 -18406 -3996
rect -18372 -4522 -18356 -3996
rect -18422 -4534 -18356 -4522
rect -18326 -3996 -18260 -3984
rect -18326 -4522 -18310 -3996
rect -18276 -4522 -18260 -3996
rect -18326 -4534 -18260 -4522
rect -18230 -3996 -18164 -3984
rect -18230 -4522 -18214 -3996
rect -18180 -4522 -18164 -3996
rect -18230 -4534 -18164 -4522
rect -18134 -3996 -18068 -3984
rect -18134 -4522 -18118 -3996
rect -18084 -4522 -18068 -3996
rect -18134 -4534 -18068 -4522
rect -18038 -3996 -17972 -3984
rect -18038 -4522 -18022 -3996
rect -17988 -4522 -17972 -3996
rect -18038 -4534 -17972 -4522
rect -17942 -3996 -17880 -3984
rect -17942 -4522 -17926 -3996
rect -17892 -4522 -17880 -3996
rect -17942 -4534 -17880 -4522
rect -17850 -3996 -17792 -3984
rect -17850 -4522 -17838 -3996
rect -17804 -4522 -17792 -3996
rect -17850 -4534 -17792 -4522
rect -17446 -3996 -17388 -3984
rect -17446 -4522 -17434 -3996
rect -17400 -4522 -17388 -3996
rect -17446 -4534 -17388 -4522
rect -17358 -3996 -17296 -3984
rect -17358 -4522 -17346 -3996
rect -17312 -4522 -17296 -3996
rect -17358 -4534 -17296 -4522
rect -17266 -3996 -17200 -3984
rect -17266 -4522 -17250 -3996
rect -17216 -4522 -17200 -3996
rect -17266 -4534 -17200 -4522
rect -17170 -3996 -17104 -3984
rect -17170 -4522 -17154 -3996
rect -17120 -4522 -17104 -3996
rect -17170 -4534 -17104 -4522
rect -17074 -3996 -17008 -3984
rect -17074 -4522 -17058 -3996
rect -17024 -4522 -17008 -3996
rect -17074 -4534 -17008 -4522
rect -16978 -3996 -16912 -3984
rect -16978 -4522 -16962 -3996
rect -16928 -4522 -16912 -3996
rect -16978 -4534 -16912 -4522
rect -16882 -3996 -16816 -3984
rect -16882 -4522 -16866 -3996
rect -16832 -4522 -16816 -3996
rect -16882 -4534 -16816 -4522
rect -16786 -3996 -16720 -3984
rect -16786 -4522 -16770 -3996
rect -16736 -4522 -16720 -3996
rect -16786 -4534 -16720 -4522
rect -16690 -3996 -16624 -3984
rect -16690 -4522 -16674 -3996
rect -16640 -4522 -16624 -3996
rect -16690 -4534 -16624 -4522
rect -16594 -3996 -16528 -3984
rect -16594 -4522 -16578 -3996
rect -16544 -4522 -16528 -3996
rect -16594 -4534 -16528 -4522
rect -16498 -3996 -16432 -3984
rect -16498 -4522 -16482 -3996
rect -16448 -4522 -16432 -3996
rect -16498 -4534 -16432 -4522
rect -16402 -3996 -16336 -3984
rect -16402 -4522 -16386 -3996
rect -16352 -4522 -16336 -3996
rect -16402 -4534 -16336 -4522
rect -16306 -3996 -16240 -3984
rect -16306 -4522 -16290 -3996
rect -16256 -4522 -16240 -3996
rect -16306 -4534 -16240 -4522
rect -16210 -3996 -16148 -3984
rect -16210 -4522 -16194 -3996
rect -16160 -4522 -16148 -3996
rect -16210 -4534 -16148 -4522
rect -16118 -3996 -16060 -3984
rect -16118 -4522 -16106 -3996
rect -16072 -4522 -16060 -3996
rect -16118 -4534 -16060 -4522
rect -15887 -3996 -15829 -3984
rect -15887 -4522 -15875 -3996
rect -15841 -4522 -15829 -3996
rect -15887 -4534 -15829 -4522
rect -15799 -3996 -15737 -3984
rect -15799 -4522 -15787 -3996
rect -15753 -4522 -15737 -3996
rect -15799 -4534 -15737 -4522
rect -15707 -3996 -15641 -3984
rect -15707 -4522 -15691 -3996
rect -15657 -4522 -15641 -3996
rect -15707 -4534 -15641 -4522
rect -15611 -3996 -15545 -3984
rect -15611 -4522 -15595 -3996
rect -15561 -4522 -15545 -3996
rect -15611 -4534 -15545 -4522
rect -15515 -3996 -15449 -3984
rect -15515 -4522 -15499 -3996
rect -15465 -4522 -15449 -3996
rect -15515 -4534 -15449 -4522
rect -15419 -3996 -15353 -3984
rect -15419 -4522 -15403 -3996
rect -15369 -4522 -15353 -3996
rect -15419 -4534 -15353 -4522
rect -15323 -3996 -15257 -3984
rect -15323 -4522 -15307 -3996
rect -15273 -4522 -15257 -3996
rect -15323 -4534 -15257 -4522
rect -15227 -3996 -15161 -3984
rect -15227 -4522 -15211 -3996
rect -15177 -4522 -15161 -3996
rect -15227 -4534 -15161 -4522
rect -15131 -3996 -15065 -3984
rect -15131 -4522 -15115 -3996
rect -15081 -4522 -15065 -3996
rect -15131 -4534 -15065 -4522
rect -15035 -3996 -14969 -3984
rect -15035 -4522 -15019 -3996
rect -14985 -4522 -14969 -3996
rect -15035 -4534 -14969 -4522
rect -14939 -3996 -14873 -3984
rect -14939 -4522 -14923 -3996
rect -14889 -4522 -14873 -3996
rect -14939 -4534 -14873 -4522
rect -14843 -3996 -14777 -3984
rect -14843 -4522 -14827 -3996
rect -14793 -4522 -14777 -3996
rect -14843 -4534 -14777 -4522
rect -14747 -3996 -14681 -3984
rect -14747 -4522 -14731 -3996
rect -14697 -4522 -14681 -3996
rect -14747 -4534 -14681 -4522
rect -14651 -3996 -14589 -3984
rect -14651 -4522 -14635 -3996
rect -14601 -4522 -14589 -3996
rect -14651 -4534 -14589 -4522
rect -14559 -3996 -14501 -3984
rect -14559 -4522 -14547 -3996
rect -14513 -4522 -14501 -3996
rect -14559 -4534 -14501 -4522
rect -14155 -3996 -14097 -3984
rect -14155 -4522 -14143 -3996
rect -14109 -4522 -14097 -3996
rect -14155 -4534 -14097 -4522
rect -14067 -3996 -14005 -3984
rect -14067 -4522 -14055 -3996
rect -14021 -4522 -14005 -3996
rect -14067 -4534 -14005 -4522
rect -13975 -3996 -13909 -3984
rect -13975 -4522 -13959 -3996
rect -13925 -4522 -13909 -3996
rect -13975 -4534 -13909 -4522
rect -13879 -3996 -13813 -3984
rect -13879 -4522 -13863 -3996
rect -13829 -4522 -13813 -3996
rect -13879 -4534 -13813 -4522
rect -13783 -3996 -13717 -3984
rect -13783 -4522 -13767 -3996
rect -13733 -4522 -13717 -3996
rect -13783 -4534 -13717 -4522
rect -13687 -3996 -13621 -3984
rect -13687 -4522 -13671 -3996
rect -13637 -4522 -13621 -3996
rect -13687 -4534 -13621 -4522
rect -13591 -3996 -13525 -3984
rect -13591 -4522 -13575 -3996
rect -13541 -4522 -13525 -3996
rect -13591 -4534 -13525 -4522
rect -13495 -3996 -13429 -3984
rect -13495 -4522 -13479 -3996
rect -13445 -4522 -13429 -3996
rect -13495 -4534 -13429 -4522
rect -13399 -3996 -13333 -3984
rect -13399 -4522 -13383 -3996
rect -13349 -4522 -13333 -3996
rect -13399 -4534 -13333 -4522
rect -13303 -3996 -13237 -3984
rect -13303 -4522 -13287 -3996
rect -13253 -4522 -13237 -3996
rect -13303 -4534 -13237 -4522
rect -13207 -3996 -13141 -3984
rect -13207 -4522 -13191 -3996
rect -13157 -4522 -13141 -3996
rect -13207 -4534 -13141 -4522
rect -13111 -3996 -13045 -3984
rect -13111 -4522 -13095 -3996
rect -13061 -4522 -13045 -3996
rect -13111 -4534 -13045 -4522
rect -13015 -3996 -12949 -3984
rect -13015 -4522 -12999 -3996
rect -12965 -4522 -12949 -3996
rect -13015 -4534 -12949 -4522
rect -12919 -3996 -12857 -3984
rect -12919 -4522 -12903 -3996
rect -12869 -4522 -12857 -3996
rect -12919 -4534 -12857 -4522
rect -12827 -3996 -12769 -3984
rect -12827 -4522 -12815 -3996
rect -12781 -4522 -12769 -3996
rect -12827 -4534 -12769 -4522
rect -12596 -3996 -12538 -3984
rect -12596 -4522 -12584 -3996
rect -12550 -4522 -12538 -3996
rect -12596 -4534 -12538 -4522
rect -12508 -3996 -12446 -3984
rect -12508 -4522 -12496 -3996
rect -12462 -4522 -12446 -3996
rect -12508 -4534 -12446 -4522
rect -12416 -3996 -12350 -3984
rect -12416 -4522 -12400 -3996
rect -12366 -4522 -12350 -3996
rect -12416 -4534 -12350 -4522
rect -12320 -3996 -12254 -3984
rect -12320 -4522 -12304 -3996
rect -12270 -4522 -12254 -3996
rect -12320 -4534 -12254 -4522
rect -12224 -3996 -12158 -3984
rect -12224 -4522 -12208 -3996
rect -12174 -4522 -12158 -3996
rect -12224 -4534 -12158 -4522
rect -12128 -3996 -12062 -3984
rect -12128 -4522 -12112 -3996
rect -12078 -4522 -12062 -3996
rect -12128 -4534 -12062 -4522
rect -12032 -3996 -11966 -3984
rect -12032 -4522 -12016 -3996
rect -11982 -4522 -11966 -3996
rect -12032 -4534 -11966 -4522
rect -11936 -3996 -11870 -3984
rect -11936 -4522 -11920 -3996
rect -11886 -4522 -11870 -3996
rect -11936 -4534 -11870 -4522
rect -11840 -3996 -11774 -3984
rect -11840 -4522 -11824 -3996
rect -11790 -4522 -11774 -3996
rect -11840 -4534 -11774 -4522
rect -11744 -3996 -11678 -3984
rect -11744 -4522 -11728 -3996
rect -11694 -4522 -11678 -3996
rect -11744 -4534 -11678 -4522
rect -11648 -3996 -11582 -3984
rect -11648 -4522 -11632 -3996
rect -11598 -4522 -11582 -3996
rect -11648 -4534 -11582 -4522
rect -11552 -3996 -11486 -3984
rect -11552 -4522 -11536 -3996
rect -11502 -4522 -11486 -3996
rect -11552 -4534 -11486 -4522
rect -11456 -3996 -11390 -3984
rect -11456 -4522 -11440 -3996
rect -11406 -4522 -11390 -3996
rect -11456 -4534 -11390 -4522
rect -11360 -3996 -11298 -3984
rect -11360 -4522 -11344 -3996
rect -11310 -4522 -11298 -3996
rect -11360 -4534 -11298 -4522
rect -11268 -3996 -11210 -3984
rect -11268 -4522 -11256 -3996
rect -11222 -4522 -11210 -3996
rect -11268 -4534 -11210 -4522
rect -10864 -3996 -10806 -3984
rect -10864 -4522 -10852 -3996
rect -10818 -4522 -10806 -3996
rect -10864 -4534 -10806 -4522
rect -10776 -3996 -10714 -3984
rect -10776 -4522 -10764 -3996
rect -10730 -4522 -10714 -3996
rect -10776 -4534 -10714 -4522
rect -10684 -3996 -10618 -3984
rect -10684 -4522 -10668 -3996
rect -10634 -4522 -10618 -3996
rect -10684 -4534 -10618 -4522
rect -10588 -3996 -10522 -3984
rect -10588 -4522 -10572 -3996
rect -10538 -4522 -10522 -3996
rect -10588 -4534 -10522 -4522
rect -10492 -3996 -10426 -3984
rect -10492 -4522 -10476 -3996
rect -10442 -4522 -10426 -3996
rect -10492 -4534 -10426 -4522
rect -10396 -3996 -10330 -3984
rect -10396 -4522 -10380 -3996
rect -10346 -4522 -10330 -3996
rect -10396 -4534 -10330 -4522
rect -10300 -3996 -10234 -3984
rect -10300 -4522 -10284 -3996
rect -10250 -4522 -10234 -3996
rect -10300 -4534 -10234 -4522
rect -10204 -3996 -10138 -3984
rect -10204 -4522 -10188 -3996
rect -10154 -4522 -10138 -3996
rect -10204 -4534 -10138 -4522
rect -10108 -3996 -10042 -3984
rect -10108 -4522 -10092 -3996
rect -10058 -4522 -10042 -3996
rect -10108 -4534 -10042 -4522
rect -10012 -3996 -9946 -3984
rect -10012 -4522 -9996 -3996
rect -9962 -4522 -9946 -3996
rect -10012 -4534 -9946 -4522
rect -9916 -3996 -9850 -3984
rect -9916 -4522 -9900 -3996
rect -9866 -4522 -9850 -3996
rect -9916 -4534 -9850 -4522
rect -9820 -3996 -9754 -3984
rect -9820 -4522 -9804 -3996
rect -9770 -4522 -9754 -3996
rect -9820 -4534 -9754 -4522
rect -9724 -3996 -9658 -3984
rect -9724 -4522 -9708 -3996
rect -9674 -4522 -9658 -3996
rect -9724 -4534 -9658 -4522
rect -9628 -3996 -9566 -3984
rect -9628 -4522 -9612 -3996
rect -9578 -4522 -9566 -3996
rect -9628 -4534 -9566 -4522
rect -9536 -3996 -9478 -3984
rect -9536 -4522 -9524 -3996
rect -9490 -4522 -9478 -3996
rect -9536 -4534 -9478 -4522
rect -9305 -3996 -9247 -3984
rect -9305 -4522 -9293 -3996
rect -9259 -4522 -9247 -3996
rect -9305 -4534 -9247 -4522
rect -9217 -3996 -9155 -3984
rect -9217 -4522 -9205 -3996
rect -9171 -4522 -9155 -3996
rect -9217 -4534 -9155 -4522
rect -9125 -3996 -9059 -3984
rect -9125 -4522 -9109 -3996
rect -9075 -4522 -9059 -3996
rect -9125 -4534 -9059 -4522
rect -9029 -3996 -8963 -3984
rect -9029 -4522 -9013 -3996
rect -8979 -4522 -8963 -3996
rect -9029 -4534 -8963 -4522
rect -8933 -3996 -8867 -3984
rect -8933 -4522 -8917 -3996
rect -8883 -4522 -8867 -3996
rect -8933 -4534 -8867 -4522
rect -8837 -3996 -8771 -3984
rect -8837 -4522 -8821 -3996
rect -8787 -4522 -8771 -3996
rect -8837 -4534 -8771 -4522
rect -8741 -3996 -8675 -3984
rect -8741 -4522 -8725 -3996
rect -8691 -4522 -8675 -3996
rect -8741 -4534 -8675 -4522
rect -8645 -3996 -8579 -3984
rect -8645 -4522 -8629 -3996
rect -8595 -4522 -8579 -3996
rect -8645 -4534 -8579 -4522
rect -8549 -3996 -8483 -3984
rect -8549 -4522 -8533 -3996
rect -8499 -4522 -8483 -3996
rect -8549 -4534 -8483 -4522
rect -8453 -3996 -8387 -3984
rect -8453 -4522 -8437 -3996
rect -8403 -4522 -8387 -3996
rect -8453 -4534 -8387 -4522
rect -8357 -3996 -8291 -3984
rect -8357 -4522 -8341 -3996
rect -8307 -4522 -8291 -3996
rect -8357 -4534 -8291 -4522
rect -8261 -3996 -8195 -3984
rect -8261 -4522 -8245 -3996
rect -8211 -4522 -8195 -3996
rect -8261 -4534 -8195 -4522
rect -8165 -3996 -8099 -3984
rect -8165 -4522 -8149 -3996
rect -8115 -4522 -8099 -3996
rect -8165 -4534 -8099 -4522
rect -8069 -3996 -8007 -3984
rect -8069 -4522 -8053 -3996
rect -8019 -4522 -8007 -3996
rect -8069 -4534 -8007 -4522
rect -7977 -3996 -7919 -3984
rect -7977 -4522 -7965 -3996
rect -7931 -4522 -7919 -3996
rect 12923 -2669 12935 -2635
rect 13125 -2669 13137 -2635
rect 12923 -2685 13137 -2669
rect 12923 -2731 13137 -2715
rect 12923 -2765 12935 -2731
rect 13129 -2765 13137 -2731
rect 12923 -2781 13137 -2765
rect 12923 -2827 13137 -2811
rect 12923 -2861 12935 -2827
rect 13125 -2861 13137 -2827
rect 12923 -2877 13137 -2861
rect 12923 -2923 13137 -2907
rect 12923 -2957 12935 -2923
rect 13129 -2957 13137 -2923
rect 12923 -2969 13137 -2957
rect 7138 -4185 7200 -4173
rect 7138 -4483 7150 -4185
rect 7184 -4483 7200 -4185
rect 7138 -4495 7200 -4483
rect 7230 -4185 7296 -4173
rect 7230 -4483 7246 -4185
rect 7280 -4483 7296 -4185
rect 7230 -4495 7296 -4483
rect 7326 -4185 7392 -4173
rect 7326 -4483 7342 -4185
rect 7376 -4483 7392 -4185
rect 7326 -4495 7392 -4483
rect 7422 -4185 7488 -4173
rect 7422 -4483 7438 -4185
rect 7472 -4483 7488 -4185
rect 7422 -4495 7488 -4483
rect 7518 -4185 7584 -4173
rect 7518 -4483 7534 -4185
rect 7568 -4483 7584 -4185
rect 7518 -4495 7584 -4483
rect 7614 -4185 7680 -4173
rect 7614 -4483 7630 -4185
rect 7664 -4483 7680 -4185
rect 7614 -4495 7680 -4483
rect 7710 -4185 7776 -4173
rect 7710 -4483 7726 -4185
rect 7760 -4483 7776 -4185
rect 7710 -4495 7776 -4483
rect 7806 -4185 7872 -4173
rect 7806 -4483 7822 -4185
rect 7856 -4483 7872 -4185
rect 7806 -4495 7872 -4483
rect 7902 -4185 7964 -4173
rect 7902 -4483 7918 -4185
rect 7952 -4483 7964 -4185
rect 7902 -4495 7964 -4483
rect 8086 -4185 8148 -4173
rect 8086 -4483 8098 -4185
rect 8132 -4483 8148 -4185
rect 8086 -4495 8148 -4483
rect 8178 -4185 8244 -4173
rect 8178 -4483 8194 -4185
rect 8228 -4483 8244 -4185
rect 8178 -4495 8244 -4483
rect 8274 -4185 8340 -4173
rect 8274 -4483 8290 -4185
rect 8324 -4483 8340 -4185
rect 8274 -4495 8340 -4483
rect 8370 -4185 8436 -4173
rect 8370 -4483 8386 -4185
rect 8420 -4483 8436 -4185
rect 8370 -4495 8436 -4483
rect 8466 -4185 8532 -4173
rect 8466 -4483 8482 -4185
rect 8516 -4483 8532 -4185
rect 8466 -4495 8532 -4483
rect 8562 -4185 8628 -4173
rect 8562 -4483 8578 -4185
rect 8612 -4483 8628 -4185
rect 8562 -4495 8628 -4483
rect 8658 -4185 8724 -4173
rect 8658 -4483 8674 -4185
rect 8708 -4483 8724 -4185
rect 8658 -4495 8724 -4483
rect 8754 -4185 8820 -4173
rect 8754 -4483 8770 -4185
rect 8804 -4483 8820 -4185
rect 8754 -4495 8820 -4483
rect 8850 -4185 8912 -4173
rect 8850 -4483 8866 -4185
rect 8900 -4483 8912 -4185
rect 8850 -4495 8912 -4483
rect 9022 -4185 9084 -4173
rect 9022 -4483 9034 -4185
rect 9068 -4483 9084 -4185
rect 9022 -4495 9084 -4483
rect 9114 -4185 9180 -4173
rect 9114 -4483 9130 -4185
rect 9164 -4483 9180 -4185
rect 9114 -4495 9180 -4483
rect 9210 -4185 9276 -4173
rect 9210 -4483 9226 -4185
rect 9260 -4483 9276 -4185
rect 9210 -4495 9276 -4483
rect 9306 -4185 9372 -4173
rect 9306 -4483 9322 -4185
rect 9356 -4483 9372 -4185
rect 9306 -4495 9372 -4483
rect 9402 -4185 9468 -4173
rect 9402 -4483 9418 -4185
rect 9452 -4483 9468 -4185
rect 9402 -4495 9468 -4483
rect 9498 -4185 9564 -4173
rect 9498 -4483 9514 -4185
rect 9548 -4483 9564 -4185
rect 9498 -4495 9564 -4483
rect 9594 -4185 9660 -4173
rect 9594 -4483 9610 -4185
rect 9644 -4483 9660 -4185
rect 9594 -4495 9660 -4483
rect 9690 -4185 9756 -4173
rect 9690 -4483 9706 -4185
rect 9740 -4483 9756 -4185
rect 9690 -4495 9756 -4483
rect 9786 -4185 9848 -4173
rect 9786 -4483 9802 -4185
rect 9836 -4483 9848 -4185
rect 9786 -4495 9848 -4483
rect 9953 -4184 10015 -4172
rect 9953 -4482 9965 -4184
rect 9999 -4482 10015 -4184
rect 9953 -4494 10015 -4482
rect 10045 -4184 10111 -4172
rect 10045 -4482 10061 -4184
rect 10095 -4482 10111 -4184
rect 10045 -4494 10111 -4482
rect 10141 -4184 10207 -4172
rect 10141 -4482 10157 -4184
rect 10191 -4482 10207 -4184
rect 10141 -4494 10207 -4482
rect 10237 -4184 10303 -4172
rect 10237 -4482 10253 -4184
rect 10287 -4482 10303 -4184
rect 10237 -4494 10303 -4482
rect 10333 -4184 10399 -4172
rect 10333 -4482 10349 -4184
rect 10383 -4482 10399 -4184
rect 10333 -4494 10399 -4482
rect 10429 -4184 10495 -4172
rect 10429 -4482 10445 -4184
rect 10479 -4482 10495 -4184
rect 10429 -4494 10495 -4482
rect 10525 -4184 10591 -4172
rect 10525 -4482 10541 -4184
rect 10575 -4482 10591 -4184
rect 10525 -4494 10591 -4482
rect 10621 -4184 10687 -4172
rect 10621 -4482 10637 -4184
rect 10671 -4482 10687 -4184
rect 10621 -4494 10687 -4482
rect 10717 -4184 10779 -4172
rect 10717 -4482 10733 -4184
rect 10767 -4482 10779 -4184
rect 10717 -4494 10779 -4482
rect 10880 -4185 10942 -4173
rect 10880 -4483 10892 -4185
rect 10926 -4483 10942 -4185
rect 10880 -4495 10942 -4483
rect 10972 -4185 11038 -4173
rect 10972 -4483 10988 -4185
rect 11022 -4483 11038 -4185
rect 10972 -4495 11038 -4483
rect 11068 -4185 11134 -4173
rect 11068 -4483 11084 -4185
rect 11118 -4483 11134 -4185
rect 11068 -4495 11134 -4483
rect 11164 -4185 11230 -4173
rect 11164 -4483 11180 -4185
rect 11214 -4483 11230 -4185
rect 11164 -4495 11230 -4483
rect 11260 -4185 11326 -4173
rect 11260 -4483 11276 -4185
rect 11310 -4483 11326 -4185
rect 11260 -4495 11326 -4483
rect 11356 -4185 11422 -4173
rect 11356 -4483 11372 -4185
rect 11406 -4483 11422 -4185
rect 11356 -4495 11422 -4483
rect 11452 -4185 11518 -4173
rect 11452 -4483 11468 -4185
rect 11502 -4483 11518 -4185
rect 11452 -4495 11518 -4483
rect 11548 -4185 11614 -4173
rect 11548 -4483 11564 -4185
rect 11598 -4483 11614 -4185
rect 11548 -4495 11614 -4483
rect 11644 -4185 11706 -4173
rect 11644 -4483 11660 -4185
rect 11694 -4483 11706 -4185
rect 11644 -4495 11706 -4483
rect -7977 -4534 -7919 -4522
rect 5658 -5045 5872 -5033
rect 5658 -5079 5670 -5045
rect 5860 -5079 5872 -5045
rect 6098 -5045 6312 -5033
rect 5658 -5095 5872 -5079
rect 5658 -5141 5872 -5125
rect 5658 -5175 5670 -5141
rect 5864 -5175 5872 -5141
rect 5658 -5191 5872 -5175
rect 5658 -5237 5872 -5221
rect 5658 -5271 5670 -5237
rect 5860 -5271 5872 -5237
rect 5658 -5287 5872 -5271
rect 5658 -5333 5872 -5317
rect 5658 -5367 5670 -5333
rect 5864 -5367 5872 -5333
rect 6098 -5079 6110 -5045
rect 6300 -5079 6312 -5045
rect 6538 -5045 6752 -5033
rect 6098 -5095 6312 -5079
rect 6098 -5141 6312 -5125
rect 6098 -5175 6110 -5141
rect 6304 -5175 6312 -5141
rect 6098 -5191 6312 -5175
rect 6098 -5237 6312 -5221
rect 6098 -5271 6110 -5237
rect 6300 -5271 6312 -5237
rect 6098 -5287 6312 -5271
rect 6098 -5333 6312 -5317
rect 5658 -5379 5872 -5367
rect 6098 -5367 6110 -5333
rect 6304 -5367 6312 -5333
rect 6538 -5079 6550 -5045
rect 6740 -5079 6752 -5045
rect 6538 -5095 6752 -5079
rect 6538 -5141 6752 -5125
rect 6538 -5175 6550 -5141
rect 6744 -5175 6752 -5141
rect 6538 -5191 6752 -5175
rect 6538 -5237 6752 -5221
rect 6538 -5271 6550 -5237
rect 6740 -5271 6752 -5237
rect 6538 -5287 6752 -5271
rect 6538 -5333 6752 -5317
rect 6098 -5379 6312 -5367
rect 6538 -5367 6550 -5333
rect 6744 -5367 6752 -5333
rect 6538 -5379 6752 -5367
rect -23586 -5423 -23372 -5411
rect -24396 -5529 -24334 -5517
rect -24396 -5719 -24384 -5529
rect -24350 -5719 -24334 -5529
rect -24396 -5731 -24334 -5719
rect -24304 -5529 -24238 -5517
rect -24304 -5719 -24288 -5529
rect -24254 -5719 -24238 -5529
rect -24304 -5731 -24238 -5719
rect -24208 -5529 -24142 -5517
rect -24208 -5719 -24192 -5529
rect -24158 -5719 -24142 -5529
rect -24208 -5731 -24142 -5719
rect -24112 -5529 -24046 -5517
rect -24112 -5719 -24096 -5529
rect -24062 -5719 -24046 -5529
rect -24112 -5731 -24046 -5719
rect -24016 -5529 -23950 -5517
rect -24016 -5719 -24000 -5529
rect -23966 -5719 -23950 -5529
rect -24016 -5731 -23950 -5719
rect -23920 -5529 -23854 -5517
rect -23920 -5719 -23904 -5529
rect -23870 -5719 -23854 -5529
rect -23920 -5731 -23854 -5719
rect -23824 -5529 -23762 -5517
rect -23824 -5719 -23808 -5529
rect -23774 -5719 -23762 -5529
rect -23586 -5457 -23574 -5423
rect -23384 -5457 -23372 -5423
rect -23586 -5473 -23372 -5457
rect -21852 -5423 -21638 -5411
rect -23586 -5519 -23372 -5503
rect -23586 -5553 -23574 -5519
rect -23380 -5553 -23372 -5519
rect -23586 -5569 -23372 -5553
rect -22660 -5529 -22598 -5517
rect -23586 -5615 -23372 -5599
rect -23586 -5649 -23574 -5615
rect -23384 -5649 -23372 -5615
rect -23586 -5665 -23372 -5649
rect -23586 -5711 -23372 -5695
rect -23824 -5731 -23762 -5719
rect -23586 -5745 -23574 -5711
rect -23380 -5745 -23372 -5711
rect -22660 -5719 -22648 -5529
rect -22614 -5719 -22598 -5529
rect -22660 -5731 -22598 -5719
rect -22568 -5529 -22502 -5517
rect -22568 -5719 -22552 -5529
rect -22518 -5719 -22502 -5529
rect -22568 -5731 -22502 -5719
rect -22472 -5529 -22406 -5517
rect -22472 -5719 -22456 -5529
rect -22422 -5719 -22406 -5529
rect -22472 -5731 -22406 -5719
rect -22376 -5529 -22310 -5517
rect -22376 -5719 -22360 -5529
rect -22326 -5719 -22310 -5529
rect -22376 -5731 -22310 -5719
rect -22280 -5529 -22214 -5517
rect -22280 -5719 -22264 -5529
rect -22230 -5719 -22214 -5529
rect -22280 -5731 -22214 -5719
rect -22184 -5529 -22118 -5517
rect -22184 -5719 -22168 -5529
rect -22134 -5719 -22118 -5529
rect -22184 -5731 -22118 -5719
rect -22088 -5529 -22026 -5517
rect -22088 -5719 -22072 -5529
rect -22038 -5719 -22026 -5529
rect -21852 -5457 -21840 -5423
rect -21650 -5457 -21638 -5423
rect -21852 -5473 -21638 -5457
rect -21852 -5519 -21638 -5503
rect -21852 -5553 -21840 -5519
rect -21646 -5553 -21638 -5519
rect -21852 -5569 -21638 -5553
rect -21852 -5615 -21638 -5599
rect -21852 -5649 -21840 -5615
rect -21650 -5649 -21638 -5615
rect -21852 -5665 -21638 -5649
rect -21852 -5711 -21638 -5695
rect -22088 -5731 -22026 -5719
rect -23586 -5757 -23372 -5745
rect -21852 -5745 -21840 -5711
rect -21646 -5745 -21638 -5711
rect -21852 -5757 -21638 -5745
rect -20530 -5697 -20468 -5685
rect -20530 -5887 -20518 -5697
rect -20484 -5887 -20468 -5697
rect -20530 -5899 -20468 -5887
rect -20438 -5697 -20372 -5685
rect -20438 -5887 -20422 -5697
rect -20388 -5887 -20372 -5697
rect -20438 -5899 -20372 -5887
rect -20342 -5697 -20276 -5685
rect -20342 -5887 -20326 -5697
rect -20292 -5887 -20276 -5697
rect -20342 -5899 -20276 -5887
rect -20246 -5697 -20180 -5685
rect -20246 -5887 -20230 -5697
rect -20196 -5887 -20180 -5697
rect -20246 -5899 -20180 -5887
rect -20150 -5697 -20084 -5685
rect -20150 -5887 -20134 -5697
rect -20100 -5887 -20084 -5697
rect -20150 -5899 -20084 -5887
rect -20054 -5697 -19988 -5685
rect -20054 -5887 -20038 -5697
rect -20004 -5887 -19988 -5697
rect -20054 -5899 -19988 -5887
rect -19958 -5697 -19896 -5685
rect -19958 -5887 -19942 -5697
rect -19908 -5887 -19896 -5697
rect -19958 -5899 -19896 -5887
rect -19421 -5697 -19359 -5685
rect -19421 -5887 -19409 -5697
rect -19375 -5887 -19359 -5697
rect -19421 -5899 -19359 -5887
rect -19329 -5697 -19263 -5685
rect -19329 -5887 -19313 -5697
rect -19279 -5887 -19263 -5697
rect -19329 -5899 -19263 -5887
rect -19233 -5697 -19167 -5685
rect -19233 -5887 -19217 -5697
rect -19183 -5887 -19167 -5697
rect -19233 -5899 -19167 -5887
rect -19137 -5697 -19071 -5685
rect -19137 -5887 -19121 -5697
rect -19087 -5887 -19071 -5697
rect -19137 -5899 -19071 -5887
rect -19041 -5697 -18975 -5685
rect -19041 -5887 -19025 -5697
rect -18991 -5887 -18975 -5697
rect -19041 -5899 -18975 -5887
rect -18945 -5697 -18879 -5685
rect -18945 -5887 -18929 -5697
rect -18895 -5887 -18879 -5697
rect -18945 -5899 -18879 -5887
rect -18849 -5697 -18787 -5685
rect -18849 -5887 -18833 -5697
rect -18799 -5887 -18787 -5697
rect -18849 -5899 -18787 -5887
rect -18539 -5697 -18477 -5685
rect -18539 -5887 -18527 -5697
rect -18493 -5887 -18477 -5697
rect -18539 -5899 -18477 -5887
rect -18447 -5697 -18381 -5685
rect -18447 -5887 -18431 -5697
rect -18397 -5887 -18381 -5697
rect -18447 -5899 -18381 -5887
rect -18351 -5697 -18285 -5685
rect -18351 -5887 -18335 -5697
rect -18301 -5887 -18285 -5697
rect -18351 -5899 -18285 -5887
rect -18255 -5697 -18189 -5685
rect -18255 -5887 -18239 -5697
rect -18205 -5887 -18189 -5697
rect -18255 -5899 -18189 -5887
rect -18159 -5697 -18093 -5685
rect -18159 -5887 -18143 -5697
rect -18109 -5887 -18093 -5697
rect -18159 -5899 -18093 -5887
rect -18063 -5697 -17997 -5685
rect -18063 -5887 -18047 -5697
rect -18013 -5887 -17997 -5697
rect -18063 -5899 -17997 -5887
rect -17967 -5697 -17905 -5685
rect -17967 -5887 -17951 -5697
rect -17917 -5887 -17905 -5697
rect -17967 -5899 -17905 -5887
rect -17239 -5697 -17177 -5685
rect -17239 -5887 -17227 -5697
rect -17193 -5887 -17177 -5697
rect -17239 -5899 -17177 -5887
rect -17147 -5697 -17081 -5685
rect -17147 -5887 -17131 -5697
rect -17097 -5887 -17081 -5697
rect -17147 -5899 -17081 -5887
rect -17051 -5697 -16985 -5685
rect -17051 -5887 -17035 -5697
rect -17001 -5887 -16985 -5697
rect -17051 -5899 -16985 -5887
rect -16955 -5697 -16889 -5685
rect -16955 -5887 -16939 -5697
rect -16905 -5887 -16889 -5697
rect -16955 -5899 -16889 -5887
rect -16859 -5697 -16793 -5685
rect -16859 -5887 -16843 -5697
rect -16809 -5887 -16793 -5697
rect -16859 -5899 -16793 -5887
rect -16763 -5697 -16697 -5685
rect -16763 -5887 -16747 -5697
rect -16713 -5887 -16697 -5697
rect -16763 -5899 -16697 -5887
rect -16667 -5697 -16605 -5685
rect -16667 -5887 -16651 -5697
rect -16617 -5887 -16605 -5697
rect -16667 -5899 -16605 -5887
rect -16130 -5697 -16068 -5685
rect -16130 -5887 -16118 -5697
rect -16084 -5887 -16068 -5697
rect -16130 -5899 -16068 -5887
rect -16038 -5697 -15972 -5685
rect -16038 -5887 -16022 -5697
rect -15988 -5887 -15972 -5697
rect -16038 -5899 -15972 -5887
rect -15942 -5697 -15876 -5685
rect -15942 -5887 -15926 -5697
rect -15892 -5887 -15876 -5697
rect -15942 -5899 -15876 -5887
rect -15846 -5697 -15780 -5685
rect -15846 -5887 -15830 -5697
rect -15796 -5887 -15780 -5697
rect -15846 -5899 -15780 -5887
rect -15750 -5697 -15684 -5685
rect -15750 -5887 -15734 -5697
rect -15700 -5887 -15684 -5697
rect -15750 -5899 -15684 -5887
rect -15654 -5697 -15588 -5685
rect -15654 -5887 -15638 -5697
rect -15604 -5887 -15588 -5697
rect -15654 -5899 -15588 -5887
rect -15558 -5697 -15496 -5685
rect -15558 -5887 -15542 -5697
rect -15508 -5887 -15496 -5697
rect -15558 -5899 -15496 -5887
rect -15248 -5697 -15186 -5685
rect -15248 -5887 -15236 -5697
rect -15202 -5887 -15186 -5697
rect -15248 -5899 -15186 -5887
rect -15156 -5697 -15090 -5685
rect -15156 -5887 -15140 -5697
rect -15106 -5887 -15090 -5697
rect -15156 -5899 -15090 -5887
rect -15060 -5697 -14994 -5685
rect -15060 -5887 -15044 -5697
rect -15010 -5887 -14994 -5697
rect -15060 -5899 -14994 -5887
rect -14964 -5697 -14898 -5685
rect -14964 -5887 -14948 -5697
rect -14914 -5887 -14898 -5697
rect -14964 -5899 -14898 -5887
rect -14868 -5697 -14802 -5685
rect -14868 -5887 -14852 -5697
rect -14818 -5887 -14802 -5697
rect -14868 -5899 -14802 -5887
rect -14772 -5697 -14706 -5685
rect -14772 -5887 -14756 -5697
rect -14722 -5887 -14706 -5697
rect -14772 -5899 -14706 -5887
rect -14676 -5697 -14614 -5685
rect -14676 -5887 -14660 -5697
rect -14626 -5887 -14614 -5697
rect -14676 -5899 -14614 -5887
rect -13948 -5697 -13886 -5685
rect -13948 -5887 -13936 -5697
rect -13902 -5887 -13886 -5697
rect -13948 -5899 -13886 -5887
rect -13856 -5697 -13790 -5685
rect -13856 -5887 -13840 -5697
rect -13806 -5887 -13790 -5697
rect -13856 -5899 -13790 -5887
rect -13760 -5697 -13694 -5685
rect -13760 -5887 -13744 -5697
rect -13710 -5887 -13694 -5697
rect -13760 -5899 -13694 -5887
rect -13664 -5697 -13598 -5685
rect -13664 -5887 -13648 -5697
rect -13614 -5887 -13598 -5697
rect -13664 -5899 -13598 -5887
rect -13568 -5697 -13502 -5685
rect -13568 -5887 -13552 -5697
rect -13518 -5887 -13502 -5697
rect -13568 -5899 -13502 -5887
rect -13472 -5697 -13406 -5685
rect -13472 -5887 -13456 -5697
rect -13422 -5887 -13406 -5697
rect -13472 -5899 -13406 -5887
rect -13376 -5697 -13314 -5685
rect -13376 -5887 -13360 -5697
rect -13326 -5887 -13314 -5697
rect -13376 -5899 -13314 -5887
rect -12839 -5697 -12777 -5685
rect -12839 -5887 -12827 -5697
rect -12793 -5887 -12777 -5697
rect -12839 -5899 -12777 -5887
rect -12747 -5697 -12681 -5685
rect -12747 -5887 -12731 -5697
rect -12697 -5887 -12681 -5697
rect -12747 -5899 -12681 -5887
rect -12651 -5697 -12585 -5685
rect -12651 -5887 -12635 -5697
rect -12601 -5887 -12585 -5697
rect -12651 -5899 -12585 -5887
rect -12555 -5697 -12489 -5685
rect -12555 -5887 -12539 -5697
rect -12505 -5887 -12489 -5697
rect -12555 -5899 -12489 -5887
rect -12459 -5697 -12393 -5685
rect -12459 -5887 -12443 -5697
rect -12409 -5887 -12393 -5697
rect -12459 -5899 -12393 -5887
rect -12363 -5697 -12297 -5685
rect -12363 -5887 -12347 -5697
rect -12313 -5887 -12297 -5697
rect -12363 -5899 -12297 -5887
rect -12267 -5697 -12205 -5685
rect -12267 -5887 -12251 -5697
rect -12217 -5887 -12205 -5697
rect -12267 -5899 -12205 -5887
rect -11957 -5697 -11895 -5685
rect -11957 -5887 -11945 -5697
rect -11911 -5887 -11895 -5697
rect -11957 -5899 -11895 -5887
rect -11865 -5697 -11799 -5685
rect -11865 -5887 -11849 -5697
rect -11815 -5887 -11799 -5697
rect -11865 -5899 -11799 -5887
rect -11769 -5697 -11703 -5685
rect -11769 -5887 -11753 -5697
rect -11719 -5887 -11703 -5697
rect -11769 -5899 -11703 -5887
rect -11673 -5697 -11607 -5685
rect -11673 -5887 -11657 -5697
rect -11623 -5887 -11607 -5697
rect -11673 -5899 -11607 -5887
rect -11577 -5697 -11511 -5685
rect -11577 -5887 -11561 -5697
rect -11527 -5887 -11511 -5697
rect -11577 -5899 -11511 -5887
rect -11481 -5697 -11415 -5685
rect -11481 -5887 -11465 -5697
rect -11431 -5887 -11415 -5697
rect -11481 -5899 -11415 -5887
rect -11385 -5697 -11323 -5685
rect -11385 -5887 -11369 -5697
rect -11335 -5887 -11323 -5697
rect -11385 -5899 -11323 -5887
rect -10657 -5697 -10595 -5685
rect -10657 -5887 -10645 -5697
rect -10611 -5887 -10595 -5697
rect -10657 -5899 -10595 -5887
rect -10565 -5697 -10499 -5685
rect -10565 -5887 -10549 -5697
rect -10515 -5887 -10499 -5697
rect -10565 -5899 -10499 -5887
rect -10469 -5697 -10403 -5685
rect -10469 -5887 -10453 -5697
rect -10419 -5887 -10403 -5697
rect -10469 -5899 -10403 -5887
rect -10373 -5697 -10307 -5685
rect -10373 -5887 -10357 -5697
rect -10323 -5887 -10307 -5697
rect -10373 -5899 -10307 -5887
rect -10277 -5697 -10211 -5685
rect -10277 -5887 -10261 -5697
rect -10227 -5887 -10211 -5697
rect -10277 -5899 -10211 -5887
rect -10181 -5697 -10115 -5685
rect -10181 -5887 -10165 -5697
rect -10131 -5887 -10115 -5697
rect -10181 -5899 -10115 -5887
rect -10085 -5697 -10023 -5685
rect -10085 -5887 -10069 -5697
rect -10035 -5887 -10023 -5697
rect -10085 -5899 -10023 -5887
rect -9548 -5697 -9486 -5685
rect -9548 -5887 -9536 -5697
rect -9502 -5887 -9486 -5697
rect -9548 -5899 -9486 -5887
rect -9456 -5697 -9390 -5685
rect -9456 -5887 -9440 -5697
rect -9406 -5887 -9390 -5697
rect -9456 -5899 -9390 -5887
rect -9360 -5697 -9294 -5685
rect -9360 -5887 -9344 -5697
rect -9310 -5887 -9294 -5697
rect -9360 -5899 -9294 -5887
rect -9264 -5697 -9198 -5685
rect -9264 -5887 -9248 -5697
rect -9214 -5887 -9198 -5697
rect -9264 -5899 -9198 -5887
rect -9168 -5697 -9102 -5685
rect -9168 -5887 -9152 -5697
rect -9118 -5887 -9102 -5697
rect -9168 -5899 -9102 -5887
rect -9072 -5697 -9006 -5685
rect -9072 -5887 -9056 -5697
rect -9022 -5887 -9006 -5697
rect -9072 -5899 -9006 -5887
rect -8976 -5697 -8914 -5685
rect -8976 -5887 -8960 -5697
rect -8926 -5887 -8914 -5697
rect -8976 -5899 -8914 -5887
rect -8666 -5697 -8604 -5685
rect -8666 -5887 -8654 -5697
rect -8620 -5887 -8604 -5697
rect -8666 -5899 -8604 -5887
rect -8574 -5697 -8508 -5685
rect -8574 -5887 -8558 -5697
rect -8524 -5887 -8508 -5697
rect -8574 -5899 -8508 -5887
rect -8478 -5697 -8412 -5685
rect -8478 -5887 -8462 -5697
rect -8428 -5887 -8412 -5697
rect -8478 -5899 -8412 -5887
rect -8382 -5697 -8316 -5685
rect -8382 -5887 -8366 -5697
rect -8332 -5887 -8316 -5697
rect -8382 -5899 -8316 -5887
rect -8286 -5697 -8220 -5685
rect -8286 -5887 -8270 -5697
rect -8236 -5887 -8220 -5697
rect -8286 -5899 -8220 -5887
rect -8190 -5697 -8124 -5685
rect -8190 -5887 -8174 -5697
rect -8140 -5887 -8124 -5697
rect -8190 -5899 -8124 -5887
rect -8094 -5697 -8032 -5685
rect -8094 -5887 -8078 -5697
rect -8044 -5887 -8032 -5697
rect -8094 -5899 -8032 -5887
rect 7138 -5749 7200 -5737
rect 7138 -6047 7150 -5749
rect 7184 -6047 7200 -5749
rect 7138 -6059 7200 -6047
rect 7230 -5749 7296 -5737
rect 7230 -6047 7246 -5749
rect 7280 -6047 7296 -5749
rect 7230 -6059 7296 -6047
rect 7326 -5749 7392 -5737
rect 7326 -6047 7342 -5749
rect 7376 -6047 7392 -5749
rect 7326 -6059 7392 -6047
rect 7422 -5749 7488 -5737
rect 7422 -6047 7438 -5749
rect 7472 -6047 7488 -5749
rect 7422 -6059 7488 -6047
rect 7518 -5749 7584 -5737
rect 7518 -6047 7534 -5749
rect 7568 -6047 7584 -5749
rect 7518 -6059 7584 -6047
rect 7614 -5749 7680 -5737
rect 7614 -6047 7630 -5749
rect 7664 -6047 7680 -5749
rect 7614 -6059 7680 -6047
rect 7710 -5749 7776 -5737
rect 7710 -6047 7726 -5749
rect 7760 -6047 7776 -5749
rect 7710 -6059 7776 -6047
rect 7806 -5749 7872 -5737
rect 7806 -6047 7822 -5749
rect 7856 -6047 7872 -5749
rect 7806 -6059 7872 -6047
rect 7902 -5749 7964 -5737
rect 7902 -6047 7918 -5749
rect 7952 -6047 7964 -5749
rect 7902 -6059 7964 -6047
rect 8086 -5749 8148 -5737
rect 8086 -6047 8098 -5749
rect 8132 -6047 8148 -5749
rect 8086 -6059 8148 -6047
rect 8178 -5749 8244 -5737
rect 8178 -6047 8194 -5749
rect 8228 -6047 8244 -5749
rect 8178 -6059 8244 -6047
rect 8274 -5749 8340 -5737
rect 8274 -6047 8290 -5749
rect 8324 -6047 8340 -5749
rect 8274 -6059 8340 -6047
rect 8370 -5749 8436 -5737
rect 8370 -6047 8386 -5749
rect 8420 -6047 8436 -5749
rect 8370 -6059 8436 -6047
rect 8466 -5749 8532 -5737
rect 8466 -6047 8482 -5749
rect 8516 -6047 8532 -5749
rect 8466 -6059 8532 -6047
rect 8562 -5749 8628 -5737
rect 8562 -6047 8578 -5749
rect 8612 -6047 8628 -5749
rect 8562 -6059 8628 -6047
rect 8658 -5749 8724 -5737
rect 8658 -6047 8674 -5749
rect 8708 -6047 8724 -5749
rect 8658 -6059 8724 -6047
rect 8754 -5749 8820 -5737
rect 8754 -6047 8770 -5749
rect 8804 -6047 8820 -5749
rect 8754 -6059 8820 -6047
rect 8850 -5749 8912 -5737
rect 8850 -6047 8866 -5749
rect 8900 -6047 8912 -5749
rect 8850 -6059 8912 -6047
rect 9022 -5749 9084 -5737
rect 9022 -6047 9034 -5749
rect 9068 -6047 9084 -5749
rect 9022 -6059 9084 -6047
rect 9114 -5749 9180 -5737
rect 9114 -6047 9130 -5749
rect 9164 -6047 9180 -5749
rect 9114 -6059 9180 -6047
rect 9210 -5749 9276 -5737
rect 9210 -6047 9226 -5749
rect 9260 -6047 9276 -5749
rect 9210 -6059 9276 -6047
rect 9306 -5749 9372 -5737
rect 9306 -6047 9322 -5749
rect 9356 -6047 9372 -5749
rect 9306 -6059 9372 -6047
rect 9402 -5749 9468 -5737
rect 9402 -6047 9418 -5749
rect 9452 -6047 9468 -5749
rect 9402 -6059 9468 -6047
rect 9498 -5749 9564 -5737
rect 9498 -6047 9514 -5749
rect 9548 -6047 9564 -5749
rect 9498 -6059 9564 -6047
rect 9594 -5749 9660 -5737
rect 9594 -6047 9610 -5749
rect 9644 -6047 9660 -5749
rect 9594 -6059 9660 -6047
rect 9690 -5749 9756 -5737
rect 9690 -6047 9706 -5749
rect 9740 -6047 9756 -5749
rect 9690 -6059 9756 -6047
rect 9786 -5749 9848 -5737
rect 9786 -6047 9802 -5749
rect 9836 -6047 9848 -5749
rect 9786 -6059 9848 -6047
rect 9953 -5749 10015 -5737
rect 9953 -6047 9965 -5749
rect 9999 -6047 10015 -5749
rect 9953 -6059 10015 -6047
rect 10045 -5749 10111 -5737
rect 10045 -6047 10061 -5749
rect 10095 -6047 10111 -5749
rect 10045 -6059 10111 -6047
rect 10141 -5749 10207 -5737
rect 10141 -6047 10157 -5749
rect 10191 -6047 10207 -5749
rect 10141 -6059 10207 -6047
rect 10237 -5749 10303 -5737
rect 10237 -6047 10253 -5749
rect 10287 -6047 10303 -5749
rect 10237 -6059 10303 -6047
rect 10333 -5749 10399 -5737
rect 10333 -6047 10349 -5749
rect 10383 -6047 10399 -5749
rect 10333 -6059 10399 -6047
rect 10429 -5749 10495 -5737
rect 10429 -6047 10445 -5749
rect 10479 -6047 10495 -5749
rect 10429 -6059 10495 -6047
rect 10525 -5749 10591 -5737
rect 10525 -6047 10541 -5749
rect 10575 -6047 10591 -5749
rect 10525 -6059 10591 -6047
rect 10621 -5749 10687 -5737
rect 10621 -6047 10637 -5749
rect 10671 -6047 10687 -5749
rect 10621 -6059 10687 -6047
rect 10717 -5749 10779 -5737
rect 10717 -6047 10733 -5749
rect 10767 -6047 10779 -5749
rect 10717 -6059 10779 -6047
rect 10880 -5749 10942 -5737
rect 10880 -6047 10892 -5749
rect 10926 -6047 10942 -5749
rect 10880 -6059 10942 -6047
rect 10972 -5749 11038 -5737
rect 10972 -6047 10988 -5749
rect 11022 -6047 11038 -5749
rect 10972 -6059 11038 -6047
rect 11068 -5749 11134 -5737
rect 11068 -6047 11084 -5749
rect 11118 -6047 11134 -5749
rect 11068 -6059 11134 -6047
rect 11164 -5749 11230 -5737
rect 11164 -6047 11180 -5749
rect 11214 -6047 11230 -5749
rect 11164 -6059 11230 -6047
rect 11260 -5749 11326 -5737
rect 11260 -6047 11276 -5749
rect 11310 -6047 11326 -5749
rect 11260 -6059 11326 -6047
rect 11356 -5749 11422 -5737
rect 11356 -6047 11372 -5749
rect 11406 -6047 11422 -5749
rect 11356 -6059 11422 -6047
rect 11452 -5749 11518 -5737
rect 11452 -6047 11468 -5749
rect 11502 -6047 11518 -5749
rect 11452 -6059 11518 -6047
rect 11548 -5749 11614 -5737
rect 11548 -6047 11564 -5749
rect 11598 -6047 11614 -5749
rect 11548 -6059 11614 -6047
rect 11644 -5749 11706 -5737
rect 11644 -6047 11660 -5749
rect 11694 -6047 11706 -5749
rect 11644 -6059 11706 -6047
rect -20737 -7261 -20679 -7249
rect -23584 -7396 -23370 -7384
rect -24396 -7502 -24334 -7490
rect -24396 -7692 -24384 -7502
rect -24350 -7692 -24334 -7502
rect -24396 -7704 -24334 -7692
rect -24304 -7502 -24238 -7490
rect -24304 -7692 -24288 -7502
rect -24254 -7692 -24238 -7502
rect -24304 -7704 -24238 -7692
rect -24208 -7502 -24142 -7490
rect -24208 -7692 -24192 -7502
rect -24158 -7692 -24142 -7502
rect -24208 -7704 -24142 -7692
rect -24112 -7502 -24046 -7490
rect -24112 -7692 -24096 -7502
rect -24062 -7692 -24046 -7502
rect -24112 -7704 -24046 -7692
rect -24016 -7502 -23950 -7490
rect -24016 -7692 -24000 -7502
rect -23966 -7692 -23950 -7502
rect -24016 -7704 -23950 -7692
rect -23920 -7502 -23854 -7490
rect -23920 -7692 -23904 -7502
rect -23870 -7692 -23854 -7502
rect -23920 -7704 -23854 -7692
rect -23824 -7502 -23762 -7490
rect -23824 -7692 -23808 -7502
rect -23774 -7692 -23762 -7502
rect -23584 -7430 -23572 -7396
rect -23382 -7430 -23370 -7396
rect -23584 -7446 -23370 -7430
rect -21850 -7396 -21636 -7384
rect -23584 -7492 -23370 -7476
rect -23584 -7526 -23572 -7492
rect -23378 -7526 -23370 -7492
rect -23584 -7542 -23370 -7526
rect -22659 -7502 -22597 -7490
rect -23584 -7588 -23370 -7572
rect -23584 -7622 -23572 -7588
rect -23382 -7622 -23370 -7588
rect -23584 -7638 -23370 -7622
rect -23584 -7684 -23370 -7668
rect -23824 -7704 -23762 -7692
rect -23584 -7718 -23572 -7684
rect -23378 -7718 -23370 -7684
rect -22659 -7692 -22647 -7502
rect -22613 -7692 -22597 -7502
rect -22659 -7704 -22597 -7692
rect -22567 -7502 -22501 -7490
rect -22567 -7692 -22551 -7502
rect -22517 -7692 -22501 -7502
rect -22567 -7704 -22501 -7692
rect -22471 -7502 -22405 -7490
rect -22471 -7692 -22455 -7502
rect -22421 -7692 -22405 -7502
rect -22471 -7704 -22405 -7692
rect -22375 -7502 -22309 -7490
rect -22375 -7692 -22359 -7502
rect -22325 -7692 -22309 -7502
rect -22375 -7704 -22309 -7692
rect -22279 -7502 -22213 -7490
rect -22279 -7692 -22263 -7502
rect -22229 -7692 -22213 -7502
rect -22279 -7704 -22213 -7692
rect -22183 -7502 -22117 -7490
rect -22183 -7692 -22167 -7502
rect -22133 -7692 -22117 -7502
rect -22183 -7704 -22117 -7692
rect -22087 -7502 -22025 -7490
rect -22087 -7692 -22071 -7502
rect -22037 -7692 -22025 -7502
rect -21850 -7430 -21838 -7396
rect -21648 -7430 -21636 -7396
rect -21850 -7446 -21636 -7430
rect -21850 -7492 -21636 -7476
rect -21850 -7526 -21838 -7492
rect -21644 -7526 -21636 -7492
rect -21850 -7542 -21636 -7526
rect -21850 -7588 -21636 -7572
rect -21850 -7622 -21838 -7588
rect -21648 -7622 -21636 -7588
rect -21850 -7638 -21636 -7622
rect -21850 -7684 -21636 -7668
rect -22087 -7704 -22025 -7692
rect -23584 -7730 -23370 -7718
rect -21850 -7718 -21838 -7684
rect -21644 -7718 -21636 -7684
rect -21850 -7730 -21636 -7718
rect -20737 -7787 -20725 -7261
rect -20691 -7787 -20679 -7261
rect -20737 -7799 -20679 -7787
rect -20649 -7261 -20587 -7249
rect -20649 -7787 -20637 -7261
rect -20603 -7787 -20587 -7261
rect -20649 -7799 -20587 -7787
rect -20557 -7261 -20491 -7249
rect -20557 -7787 -20541 -7261
rect -20507 -7787 -20491 -7261
rect -20557 -7799 -20491 -7787
rect -20461 -7261 -20395 -7249
rect -20461 -7787 -20445 -7261
rect -20411 -7787 -20395 -7261
rect -20461 -7799 -20395 -7787
rect -20365 -7261 -20299 -7249
rect -20365 -7787 -20349 -7261
rect -20315 -7787 -20299 -7261
rect -20365 -7799 -20299 -7787
rect -20269 -7261 -20203 -7249
rect -20269 -7787 -20253 -7261
rect -20219 -7787 -20203 -7261
rect -20269 -7799 -20203 -7787
rect -20173 -7261 -20107 -7249
rect -20173 -7787 -20157 -7261
rect -20123 -7787 -20107 -7261
rect -20173 -7799 -20107 -7787
rect -20077 -7261 -20011 -7249
rect -20077 -7787 -20061 -7261
rect -20027 -7787 -20011 -7261
rect -20077 -7799 -20011 -7787
rect -19981 -7261 -19915 -7249
rect -19981 -7787 -19965 -7261
rect -19931 -7787 -19915 -7261
rect -19981 -7799 -19915 -7787
rect -19885 -7261 -19819 -7249
rect -19885 -7787 -19869 -7261
rect -19835 -7787 -19819 -7261
rect -19885 -7799 -19819 -7787
rect -19789 -7261 -19723 -7249
rect -19789 -7787 -19773 -7261
rect -19739 -7787 -19723 -7261
rect -19789 -7799 -19723 -7787
rect -19693 -7261 -19627 -7249
rect -19693 -7787 -19677 -7261
rect -19643 -7787 -19627 -7261
rect -19693 -7799 -19627 -7787
rect -19597 -7261 -19531 -7249
rect -19597 -7787 -19581 -7261
rect -19547 -7787 -19531 -7261
rect -19597 -7799 -19531 -7787
rect -19501 -7261 -19439 -7249
rect -19501 -7787 -19485 -7261
rect -19451 -7787 -19439 -7261
rect -19501 -7799 -19439 -7787
rect -19409 -7261 -19351 -7249
rect -19409 -7787 -19397 -7261
rect -19363 -7787 -19351 -7261
rect -19409 -7799 -19351 -7787
rect -19178 -7261 -19120 -7249
rect -19178 -7787 -19166 -7261
rect -19132 -7787 -19120 -7261
rect -19178 -7799 -19120 -7787
rect -19090 -7261 -19028 -7249
rect -19090 -7787 -19078 -7261
rect -19044 -7787 -19028 -7261
rect -19090 -7799 -19028 -7787
rect -18998 -7261 -18932 -7249
rect -18998 -7787 -18982 -7261
rect -18948 -7787 -18932 -7261
rect -18998 -7799 -18932 -7787
rect -18902 -7261 -18836 -7249
rect -18902 -7787 -18886 -7261
rect -18852 -7787 -18836 -7261
rect -18902 -7799 -18836 -7787
rect -18806 -7261 -18740 -7249
rect -18806 -7787 -18790 -7261
rect -18756 -7787 -18740 -7261
rect -18806 -7799 -18740 -7787
rect -18710 -7261 -18644 -7249
rect -18710 -7787 -18694 -7261
rect -18660 -7787 -18644 -7261
rect -18710 -7799 -18644 -7787
rect -18614 -7261 -18548 -7249
rect -18614 -7787 -18598 -7261
rect -18564 -7787 -18548 -7261
rect -18614 -7799 -18548 -7787
rect -18518 -7261 -18452 -7249
rect -18518 -7787 -18502 -7261
rect -18468 -7787 -18452 -7261
rect -18518 -7799 -18452 -7787
rect -18422 -7261 -18356 -7249
rect -18422 -7787 -18406 -7261
rect -18372 -7787 -18356 -7261
rect -18422 -7799 -18356 -7787
rect -18326 -7261 -18260 -7249
rect -18326 -7787 -18310 -7261
rect -18276 -7787 -18260 -7261
rect -18326 -7799 -18260 -7787
rect -18230 -7261 -18164 -7249
rect -18230 -7787 -18214 -7261
rect -18180 -7787 -18164 -7261
rect -18230 -7799 -18164 -7787
rect -18134 -7261 -18068 -7249
rect -18134 -7787 -18118 -7261
rect -18084 -7787 -18068 -7261
rect -18134 -7799 -18068 -7787
rect -18038 -7261 -17972 -7249
rect -18038 -7787 -18022 -7261
rect -17988 -7787 -17972 -7261
rect -18038 -7799 -17972 -7787
rect -17942 -7261 -17880 -7249
rect -17942 -7787 -17926 -7261
rect -17892 -7787 -17880 -7261
rect -17942 -7799 -17880 -7787
rect -17850 -7261 -17792 -7249
rect -17850 -7787 -17838 -7261
rect -17804 -7787 -17792 -7261
rect -17850 -7799 -17792 -7787
rect -17446 -7261 -17388 -7249
rect -17446 -7787 -17434 -7261
rect -17400 -7787 -17388 -7261
rect -17446 -7799 -17388 -7787
rect -17358 -7261 -17296 -7249
rect -17358 -7787 -17346 -7261
rect -17312 -7787 -17296 -7261
rect -17358 -7799 -17296 -7787
rect -17266 -7261 -17200 -7249
rect -17266 -7787 -17250 -7261
rect -17216 -7787 -17200 -7261
rect -17266 -7799 -17200 -7787
rect -17170 -7261 -17104 -7249
rect -17170 -7787 -17154 -7261
rect -17120 -7787 -17104 -7261
rect -17170 -7799 -17104 -7787
rect -17074 -7261 -17008 -7249
rect -17074 -7787 -17058 -7261
rect -17024 -7787 -17008 -7261
rect -17074 -7799 -17008 -7787
rect -16978 -7261 -16912 -7249
rect -16978 -7787 -16962 -7261
rect -16928 -7787 -16912 -7261
rect -16978 -7799 -16912 -7787
rect -16882 -7261 -16816 -7249
rect -16882 -7787 -16866 -7261
rect -16832 -7787 -16816 -7261
rect -16882 -7799 -16816 -7787
rect -16786 -7261 -16720 -7249
rect -16786 -7787 -16770 -7261
rect -16736 -7787 -16720 -7261
rect -16786 -7799 -16720 -7787
rect -16690 -7261 -16624 -7249
rect -16690 -7787 -16674 -7261
rect -16640 -7787 -16624 -7261
rect -16690 -7799 -16624 -7787
rect -16594 -7261 -16528 -7249
rect -16594 -7787 -16578 -7261
rect -16544 -7787 -16528 -7261
rect -16594 -7799 -16528 -7787
rect -16498 -7261 -16432 -7249
rect -16498 -7787 -16482 -7261
rect -16448 -7787 -16432 -7261
rect -16498 -7799 -16432 -7787
rect -16402 -7261 -16336 -7249
rect -16402 -7787 -16386 -7261
rect -16352 -7787 -16336 -7261
rect -16402 -7799 -16336 -7787
rect -16306 -7261 -16240 -7249
rect -16306 -7787 -16290 -7261
rect -16256 -7787 -16240 -7261
rect -16306 -7799 -16240 -7787
rect -16210 -7261 -16148 -7249
rect -16210 -7787 -16194 -7261
rect -16160 -7787 -16148 -7261
rect -16210 -7799 -16148 -7787
rect -16118 -7261 -16060 -7249
rect -16118 -7787 -16106 -7261
rect -16072 -7787 -16060 -7261
rect -16118 -7799 -16060 -7787
rect -15887 -7261 -15829 -7249
rect -15887 -7787 -15875 -7261
rect -15841 -7787 -15829 -7261
rect -15887 -7799 -15829 -7787
rect -15799 -7261 -15737 -7249
rect -15799 -7787 -15787 -7261
rect -15753 -7787 -15737 -7261
rect -15799 -7799 -15737 -7787
rect -15707 -7261 -15641 -7249
rect -15707 -7787 -15691 -7261
rect -15657 -7787 -15641 -7261
rect -15707 -7799 -15641 -7787
rect -15611 -7261 -15545 -7249
rect -15611 -7787 -15595 -7261
rect -15561 -7787 -15545 -7261
rect -15611 -7799 -15545 -7787
rect -15515 -7261 -15449 -7249
rect -15515 -7787 -15499 -7261
rect -15465 -7787 -15449 -7261
rect -15515 -7799 -15449 -7787
rect -15419 -7261 -15353 -7249
rect -15419 -7787 -15403 -7261
rect -15369 -7787 -15353 -7261
rect -15419 -7799 -15353 -7787
rect -15323 -7261 -15257 -7249
rect -15323 -7787 -15307 -7261
rect -15273 -7787 -15257 -7261
rect -15323 -7799 -15257 -7787
rect -15227 -7261 -15161 -7249
rect -15227 -7787 -15211 -7261
rect -15177 -7787 -15161 -7261
rect -15227 -7799 -15161 -7787
rect -15131 -7261 -15065 -7249
rect -15131 -7787 -15115 -7261
rect -15081 -7787 -15065 -7261
rect -15131 -7799 -15065 -7787
rect -15035 -7261 -14969 -7249
rect -15035 -7787 -15019 -7261
rect -14985 -7787 -14969 -7261
rect -15035 -7799 -14969 -7787
rect -14939 -7261 -14873 -7249
rect -14939 -7787 -14923 -7261
rect -14889 -7787 -14873 -7261
rect -14939 -7799 -14873 -7787
rect -14843 -7261 -14777 -7249
rect -14843 -7787 -14827 -7261
rect -14793 -7787 -14777 -7261
rect -14843 -7799 -14777 -7787
rect -14747 -7261 -14681 -7249
rect -14747 -7787 -14731 -7261
rect -14697 -7787 -14681 -7261
rect -14747 -7799 -14681 -7787
rect -14651 -7261 -14589 -7249
rect -14651 -7787 -14635 -7261
rect -14601 -7787 -14589 -7261
rect -14651 -7799 -14589 -7787
rect -14559 -7261 -14501 -7249
rect -14559 -7787 -14547 -7261
rect -14513 -7787 -14501 -7261
rect -14559 -7799 -14501 -7787
rect -14155 -7261 -14097 -7249
rect -14155 -7787 -14143 -7261
rect -14109 -7787 -14097 -7261
rect -14155 -7799 -14097 -7787
rect -14067 -7261 -14005 -7249
rect -14067 -7787 -14055 -7261
rect -14021 -7787 -14005 -7261
rect -14067 -7799 -14005 -7787
rect -13975 -7261 -13909 -7249
rect -13975 -7787 -13959 -7261
rect -13925 -7787 -13909 -7261
rect -13975 -7799 -13909 -7787
rect -13879 -7261 -13813 -7249
rect -13879 -7787 -13863 -7261
rect -13829 -7787 -13813 -7261
rect -13879 -7799 -13813 -7787
rect -13783 -7261 -13717 -7249
rect -13783 -7787 -13767 -7261
rect -13733 -7787 -13717 -7261
rect -13783 -7799 -13717 -7787
rect -13687 -7261 -13621 -7249
rect -13687 -7787 -13671 -7261
rect -13637 -7787 -13621 -7261
rect -13687 -7799 -13621 -7787
rect -13591 -7261 -13525 -7249
rect -13591 -7787 -13575 -7261
rect -13541 -7787 -13525 -7261
rect -13591 -7799 -13525 -7787
rect -13495 -7261 -13429 -7249
rect -13495 -7787 -13479 -7261
rect -13445 -7787 -13429 -7261
rect -13495 -7799 -13429 -7787
rect -13399 -7261 -13333 -7249
rect -13399 -7787 -13383 -7261
rect -13349 -7787 -13333 -7261
rect -13399 -7799 -13333 -7787
rect -13303 -7261 -13237 -7249
rect -13303 -7787 -13287 -7261
rect -13253 -7787 -13237 -7261
rect -13303 -7799 -13237 -7787
rect -13207 -7261 -13141 -7249
rect -13207 -7787 -13191 -7261
rect -13157 -7787 -13141 -7261
rect -13207 -7799 -13141 -7787
rect -13111 -7261 -13045 -7249
rect -13111 -7787 -13095 -7261
rect -13061 -7787 -13045 -7261
rect -13111 -7799 -13045 -7787
rect -13015 -7261 -12949 -7249
rect -13015 -7787 -12999 -7261
rect -12965 -7787 -12949 -7261
rect -13015 -7799 -12949 -7787
rect -12919 -7261 -12857 -7249
rect -12919 -7787 -12903 -7261
rect -12869 -7787 -12857 -7261
rect -12919 -7799 -12857 -7787
rect -12827 -7261 -12769 -7249
rect -12827 -7787 -12815 -7261
rect -12781 -7787 -12769 -7261
rect -12827 -7799 -12769 -7787
rect -12596 -7261 -12538 -7249
rect -12596 -7787 -12584 -7261
rect -12550 -7787 -12538 -7261
rect -12596 -7799 -12538 -7787
rect -12508 -7261 -12446 -7249
rect -12508 -7787 -12496 -7261
rect -12462 -7787 -12446 -7261
rect -12508 -7799 -12446 -7787
rect -12416 -7261 -12350 -7249
rect -12416 -7787 -12400 -7261
rect -12366 -7787 -12350 -7261
rect -12416 -7799 -12350 -7787
rect -12320 -7261 -12254 -7249
rect -12320 -7787 -12304 -7261
rect -12270 -7787 -12254 -7261
rect -12320 -7799 -12254 -7787
rect -12224 -7261 -12158 -7249
rect -12224 -7787 -12208 -7261
rect -12174 -7787 -12158 -7261
rect -12224 -7799 -12158 -7787
rect -12128 -7261 -12062 -7249
rect -12128 -7787 -12112 -7261
rect -12078 -7787 -12062 -7261
rect -12128 -7799 -12062 -7787
rect -12032 -7261 -11966 -7249
rect -12032 -7787 -12016 -7261
rect -11982 -7787 -11966 -7261
rect -12032 -7799 -11966 -7787
rect -11936 -7261 -11870 -7249
rect -11936 -7787 -11920 -7261
rect -11886 -7787 -11870 -7261
rect -11936 -7799 -11870 -7787
rect -11840 -7261 -11774 -7249
rect -11840 -7787 -11824 -7261
rect -11790 -7787 -11774 -7261
rect -11840 -7799 -11774 -7787
rect -11744 -7261 -11678 -7249
rect -11744 -7787 -11728 -7261
rect -11694 -7787 -11678 -7261
rect -11744 -7799 -11678 -7787
rect -11648 -7261 -11582 -7249
rect -11648 -7787 -11632 -7261
rect -11598 -7787 -11582 -7261
rect -11648 -7799 -11582 -7787
rect -11552 -7261 -11486 -7249
rect -11552 -7787 -11536 -7261
rect -11502 -7787 -11486 -7261
rect -11552 -7799 -11486 -7787
rect -11456 -7261 -11390 -7249
rect -11456 -7787 -11440 -7261
rect -11406 -7787 -11390 -7261
rect -11456 -7799 -11390 -7787
rect -11360 -7261 -11298 -7249
rect -11360 -7787 -11344 -7261
rect -11310 -7787 -11298 -7261
rect -11360 -7799 -11298 -7787
rect -11268 -7261 -11210 -7249
rect -11268 -7787 -11256 -7261
rect -11222 -7787 -11210 -7261
rect -11268 -7799 -11210 -7787
rect -10864 -7261 -10806 -7249
rect -10864 -7787 -10852 -7261
rect -10818 -7787 -10806 -7261
rect -10864 -7799 -10806 -7787
rect -10776 -7261 -10714 -7249
rect -10776 -7787 -10764 -7261
rect -10730 -7787 -10714 -7261
rect -10776 -7799 -10714 -7787
rect -10684 -7261 -10618 -7249
rect -10684 -7787 -10668 -7261
rect -10634 -7787 -10618 -7261
rect -10684 -7799 -10618 -7787
rect -10588 -7261 -10522 -7249
rect -10588 -7787 -10572 -7261
rect -10538 -7787 -10522 -7261
rect -10588 -7799 -10522 -7787
rect -10492 -7261 -10426 -7249
rect -10492 -7787 -10476 -7261
rect -10442 -7787 -10426 -7261
rect -10492 -7799 -10426 -7787
rect -10396 -7261 -10330 -7249
rect -10396 -7787 -10380 -7261
rect -10346 -7787 -10330 -7261
rect -10396 -7799 -10330 -7787
rect -10300 -7261 -10234 -7249
rect -10300 -7787 -10284 -7261
rect -10250 -7787 -10234 -7261
rect -10300 -7799 -10234 -7787
rect -10204 -7261 -10138 -7249
rect -10204 -7787 -10188 -7261
rect -10154 -7787 -10138 -7261
rect -10204 -7799 -10138 -7787
rect -10108 -7261 -10042 -7249
rect -10108 -7787 -10092 -7261
rect -10058 -7787 -10042 -7261
rect -10108 -7799 -10042 -7787
rect -10012 -7261 -9946 -7249
rect -10012 -7787 -9996 -7261
rect -9962 -7787 -9946 -7261
rect -10012 -7799 -9946 -7787
rect -9916 -7261 -9850 -7249
rect -9916 -7787 -9900 -7261
rect -9866 -7787 -9850 -7261
rect -9916 -7799 -9850 -7787
rect -9820 -7261 -9754 -7249
rect -9820 -7787 -9804 -7261
rect -9770 -7787 -9754 -7261
rect -9820 -7799 -9754 -7787
rect -9724 -7261 -9658 -7249
rect -9724 -7787 -9708 -7261
rect -9674 -7787 -9658 -7261
rect -9724 -7799 -9658 -7787
rect -9628 -7261 -9566 -7249
rect -9628 -7787 -9612 -7261
rect -9578 -7787 -9566 -7261
rect -9628 -7799 -9566 -7787
rect -9536 -7261 -9478 -7249
rect -9536 -7787 -9524 -7261
rect -9490 -7787 -9478 -7261
rect -9536 -7799 -9478 -7787
rect -9305 -7261 -9247 -7249
rect -9305 -7787 -9293 -7261
rect -9259 -7787 -9247 -7261
rect -9305 -7799 -9247 -7787
rect -9217 -7261 -9155 -7249
rect -9217 -7787 -9205 -7261
rect -9171 -7787 -9155 -7261
rect -9217 -7799 -9155 -7787
rect -9125 -7261 -9059 -7249
rect -9125 -7787 -9109 -7261
rect -9075 -7787 -9059 -7261
rect -9125 -7799 -9059 -7787
rect -9029 -7261 -8963 -7249
rect -9029 -7787 -9013 -7261
rect -8979 -7787 -8963 -7261
rect -9029 -7799 -8963 -7787
rect -8933 -7261 -8867 -7249
rect -8933 -7787 -8917 -7261
rect -8883 -7787 -8867 -7261
rect -8933 -7799 -8867 -7787
rect -8837 -7261 -8771 -7249
rect -8837 -7787 -8821 -7261
rect -8787 -7787 -8771 -7261
rect -8837 -7799 -8771 -7787
rect -8741 -7261 -8675 -7249
rect -8741 -7787 -8725 -7261
rect -8691 -7787 -8675 -7261
rect -8741 -7799 -8675 -7787
rect -8645 -7261 -8579 -7249
rect -8645 -7787 -8629 -7261
rect -8595 -7787 -8579 -7261
rect -8645 -7799 -8579 -7787
rect -8549 -7261 -8483 -7249
rect -8549 -7787 -8533 -7261
rect -8499 -7787 -8483 -7261
rect -8549 -7799 -8483 -7787
rect -8453 -7261 -8387 -7249
rect -8453 -7787 -8437 -7261
rect -8403 -7787 -8387 -7261
rect -8453 -7799 -8387 -7787
rect -8357 -7261 -8291 -7249
rect -8357 -7787 -8341 -7261
rect -8307 -7787 -8291 -7261
rect -8357 -7799 -8291 -7787
rect -8261 -7261 -8195 -7249
rect -8261 -7787 -8245 -7261
rect -8211 -7787 -8195 -7261
rect -8261 -7799 -8195 -7787
rect -8165 -7261 -8099 -7249
rect -8165 -7787 -8149 -7261
rect -8115 -7787 -8099 -7261
rect -8165 -7799 -8099 -7787
rect -8069 -7261 -8007 -7249
rect -8069 -7787 -8053 -7261
rect -8019 -7787 -8007 -7261
rect -8069 -7799 -8007 -7787
rect -7977 -7261 -7919 -7249
rect -7977 -7787 -7965 -7261
rect -7931 -7787 -7919 -7261
rect 11773 -6959 11835 -6947
rect 11773 -7191 11785 -6959
rect 11819 -7191 11835 -6959
rect 11773 -7203 11835 -7191
rect 11865 -6959 11931 -6947
rect 11865 -7191 11881 -6959
rect 11915 -7191 11931 -6959
rect 11865 -7203 11931 -7191
rect 11961 -6959 12027 -6947
rect 11961 -7191 11977 -6959
rect 12011 -7191 12027 -6959
rect 11961 -7203 12027 -7191
rect 12057 -6959 12123 -6947
rect 12057 -7191 12073 -6959
rect 12107 -7191 12123 -6959
rect 12057 -7203 12123 -7191
rect 12153 -6959 12219 -6947
rect 12153 -7191 12169 -6959
rect 12203 -7191 12219 -6959
rect 12153 -7203 12219 -7191
rect 12249 -6959 12315 -6947
rect 12249 -7191 12265 -6959
rect 12299 -7191 12315 -6959
rect 12249 -7203 12315 -7191
rect 12345 -6959 12411 -6947
rect 12345 -7191 12361 -6959
rect 12395 -7191 12411 -6959
rect 12345 -7203 12411 -7191
rect 12441 -6959 12507 -6947
rect 12441 -7191 12457 -6959
rect 12491 -7191 12507 -6959
rect 12441 -7203 12507 -7191
rect 12537 -6959 12603 -6947
rect 12537 -7191 12553 -6959
rect 12587 -7191 12603 -6959
rect 12537 -7203 12603 -7191
rect 12633 -6959 12699 -6947
rect 12633 -7191 12649 -6959
rect 12683 -7191 12699 -6959
rect 12633 -7203 12699 -7191
rect 12729 -6959 12791 -6947
rect 12729 -7191 12745 -6959
rect 12779 -7191 12791 -6959
rect 12923 -7063 13137 -7051
rect 12729 -7203 12791 -7191
rect -7977 -7799 -7919 -7787
rect 12923 -7097 12935 -7063
rect 13125 -7097 13137 -7063
rect 12923 -7113 13137 -7097
rect 12923 -7159 13137 -7143
rect 12923 -7193 12935 -7159
rect 13129 -7193 13137 -7159
rect 12923 -7209 13137 -7193
rect 12923 -7255 13137 -7239
rect 12923 -7289 12935 -7255
rect 13125 -7289 13137 -7255
rect 12923 -7305 13137 -7289
rect 12923 -7351 13137 -7335
rect 12923 -7385 12935 -7351
rect 13129 -7385 13137 -7351
rect 12923 -7397 13137 -7385
rect -23583 -8688 -23369 -8676
rect -24396 -8794 -24334 -8782
rect -24396 -8984 -24384 -8794
rect -24350 -8984 -24334 -8794
rect -24396 -8996 -24334 -8984
rect -24304 -8794 -24238 -8782
rect -24304 -8984 -24288 -8794
rect -24254 -8984 -24238 -8794
rect -24304 -8996 -24238 -8984
rect -24208 -8794 -24142 -8782
rect -24208 -8984 -24192 -8794
rect -24158 -8984 -24142 -8794
rect -24208 -8996 -24142 -8984
rect -24112 -8794 -24046 -8782
rect -24112 -8984 -24096 -8794
rect -24062 -8984 -24046 -8794
rect -24112 -8996 -24046 -8984
rect -24016 -8794 -23950 -8782
rect -24016 -8984 -24000 -8794
rect -23966 -8984 -23950 -8794
rect -24016 -8996 -23950 -8984
rect -23920 -8794 -23854 -8782
rect -23920 -8984 -23904 -8794
rect -23870 -8984 -23854 -8794
rect -23920 -8996 -23854 -8984
rect -23824 -8794 -23762 -8782
rect -23824 -8984 -23808 -8794
rect -23774 -8984 -23762 -8794
rect -23583 -8722 -23571 -8688
rect -23381 -8722 -23369 -8688
rect -23583 -8738 -23369 -8722
rect -21846 -8688 -21632 -8676
rect -23583 -8784 -23369 -8768
rect -23583 -8818 -23571 -8784
rect -23377 -8818 -23369 -8784
rect -23583 -8834 -23369 -8818
rect -22660 -8794 -22598 -8782
rect -23583 -8880 -23369 -8864
rect -23583 -8914 -23571 -8880
rect -23381 -8914 -23369 -8880
rect -23583 -8930 -23369 -8914
rect -23583 -8976 -23369 -8960
rect -23824 -8996 -23762 -8984
rect -23583 -9010 -23571 -8976
rect -23377 -9010 -23369 -8976
rect -22660 -8984 -22648 -8794
rect -22614 -8984 -22598 -8794
rect -22660 -8996 -22598 -8984
rect -22568 -8794 -22502 -8782
rect -22568 -8984 -22552 -8794
rect -22518 -8984 -22502 -8794
rect -22568 -8996 -22502 -8984
rect -22472 -8794 -22406 -8782
rect -22472 -8984 -22456 -8794
rect -22422 -8984 -22406 -8794
rect -22472 -8996 -22406 -8984
rect -22376 -8794 -22310 -8782
rect -22376 -8984 -22360 -8794
rect -22326 -8984 -22310 -8794
rect -22376 -8996 -22310 -8984
rect -22280 -8794 -22214 -8782
rect -22280 -8984 -22264 -8794
rect -22230 -8984 -22214 -8794
rect -22280 -8996 -22214 -8984
rect -22184 -8794 -22118 -8782
rect -22184 -8984 -22168 -8794
rect -22134 -8984 -22118 -8794
rect -22184 -8996 -22118 -8984
rect -22088 -8794 -22026 -8782
rect -22088 -8984 -22072 -8794
rect -22038 -8984 -22026 -8794
rect -21846 -8722 -21834 -8688
rect -21644 -8722 -21632 -8688
rect -21846 -8738 -21632 -8722
rect 7138 -8613 7200 -8601
rect -21846 -8784 -21632 -8768
rect -21846 -8818 -21834 -8784
rect -21640 -8818 -21632 -8784
rect -21846 -8834 -21632 -8818
rect -21846 -8880 -21632 -8864
rect -21846 -8914 -21834 -8880
rect -21644 -8914 -21632 -8880
rect -21846 -8930 -21632 -8914
rect 7138 -8911 7150 -8613
rect 7184 -8911 7200 -8613
rect 7138 -8923 7200 -8911
rect 7230 -8613 7296 -8601
rect 7230 -8911 7246 -8613
rect 7280 -8911 7296 -8613
rect 7230 -8923 7296 -8911
rect 7326 -8613 7392 -8601
rect 7326 -8911 7342 -8613
rect 7376 -8911 7392 -8613
rect 7326 -8923 7392 -8911
rect 7422 -8613 7488 -8601
rect 7422 -8911 7438 -8613
rect 7472 -8911 7488 -8613
rect 7422 -8923 7488 -8911
rect 7518 -8613 7584 -8601
rect 7518 -8911 7534 -8613
rect 7568 -8911 7584 -8613
rect 7518 -8923 7584 -8911
rect 7614 -8613 7680 -8601
rect 7614 -8911 7630 -8613
rect 7664 -8911 7680 -8613
rect 7614 -8923 7680 -8911
rect 7710 -8613 7776 -8601
rect 7710 -8911 7726 -8613
rect 7760 -8911 7776 -8613
rect 7710 -8923 7776 -8911
rect 7806 -8613 7872 -8601
rect 7806 -8911 7822 -8613
rect 7856 -8911 7872 -8613
rect 7806 -8923 7872 -8911
rect 7902 -8613 7964 -8601
rect 7902 -8911 7918 -8613
rect 7952 -8911 7964 -8613
rect 7902 -8923 7964 -8911
rect 8086 -8613 8148 -8601
rect 8086 -8911 8098 -8613
rect 8132 -8911 8148 -8613
rect 8086 -8923 8148 -8911
rect 8178 -8613 8244 -8601
rect 8178 -8911 8194 -8613
rect 8228 -8911 8244 -8613
rect 8178 -8923 8244 -8911
rect 8274 -8613 8340 -8601
rect 8274 -8911 8290 -8613
rect 8324 -8911 8340 -8613
rect 8274 -8923 8340 -8911
rect 8370 -8613 8436 -8601
rect 8370 -8911 8386 -8613
rect 8420 -8911 8436 -8613
rect 8370 -8923 8436 -8911
rect 8466 -8613 8532 -8601
rect 8466 -8911 8482 -8613
rect 8516 -8911 8532 -8613
rect 8466 -8923 8532 -8911
rect 8562 -8613 8628 -8601
rect 8562 -8911 8578 -8613
rect 8612 -8911 8628 -8613
rect 8562 -8923 8628 -8911
rect 8658 -8613 8724 -8601
rect 8658 -8911 8674 -8613
rect 8708 -8911 8724 -8613
rect 8658 -8923 8724 -8911
rect 8754 -8613 8820 -8601
rect 8754 -8911 8770 -8613
rect 8804 -8911 8820 -8613
rect 8754 -8923 8820 -8911
rect 8850 -8613 8912 -8601
rect 8850 -8911 8866 -8613
rect 8900 -8911 8912 -8613
rect 8850 -8923 8912 -8911
rect 9022 -8613 9084 -8601
rect 9022 -8911 9034 -8613
rect 9068 -8911 9084 -8613
rect 9022 -8923 9084 -8911
rect 9114 -8613 9180 -8601
rect 9114 -8911 9130 -8613
rect 9164 -8911 9180 -8613
rect 9114 -8923 9180 -8911
rect 9210 -8613 9276 -8601
rect 9210 -8911 9226 -8613
rect 9260 -8911 9276 -8613
rect 9210 -8923 9276 -8911
rect 9306 -8613 9372 -8601
rect 9306 -8911 9322 -8613
rect 9356 -8911 9372 -8613
rect 9306 -8923 9372 -8911
rect 9402 -8613 9468 -8601
rect 9402 -8911 9418 -8613
rect 9452 -8911 9468 -8613
rect 9402 -8923 9468 -8911
rect 9498 -8613 9564 -8601
rect 9498 -8911 9514 -8613
rect 9548 -8911 9564 -8613
rect 9498 -8923 9564 -8911
rect 9594 -8613 9660 -8601
rect 9594 -8911 9610 -8613
rect 9644 -8911 9660 -8613
rect 9594 -8923 9660 -8911
rect 9690 -8613 9756 -8601
rect 9690 -8911 9706 -8613
rect 9740 -8911 9756 -8613
rect 9690 -8923 9756 -8911
rect 9786 -8613 9848 -8601
rect 9786 -8911 9802 -8613
rect 9836 -8911 9848 -8613
rect 9786 -8923 9848 -8911
rect 9953 -8612 10015 -8600
rect 9953 -8910 9965 -8612
rect 9999 -8910 10015 -8612
rect 9953 -8922 10015 -8910
rect 10045 -8612 10111 -8600
rect 10045 -8910 10061 -8612
rect 10095 -8910 10111 -8612
rect 10045 -8922 10111 -8910
rect 10141 -8612 10207 -8600
rect 10141 -8910 10157 -8612
rect 10191 -8910 10207 -8612
rect 10141 -8922 10207 -8910
rect 10237 -8612 10303 -8600
rect 10237 -8910 10253 -8612
rect 10287 -8910 10303 -8612
rect 10237 -8922 10303 -8910
rect 10333 -8612 10399 -8600
rect 10333 -8910 10349 -8612
rect 10383 -8910 10399 -8612
rect 10333 -8922 10399 -8910
rect 10429 -8612 10495 -8600
rect 10429 -8910 10445 -8612
rect 10479 -8910 10495 -8612
rect 10429 -8922 10495 -8910
rect 10525 -8612 10591 -8600
rect 10525 -8910 10541 -8612
rect 10575 -8910 10591 -8612
rect 10525 -8922 10591 -8910
rect 10621 -8612 10687 -8600
rect 10621 -8910 10637 -8612
rect 10671 -8910 10687 -8612
rect 10621 -8922 10687 -8910
rect 10717 -8612 10779 -8600
rect 10717 -8910 10733 -8612
rect 10767 -8910 10779 -8612
rect 10717 -8922 10779 -8910
rect 10880 -8613 10942 -8601
rect 10880 -8911 10892 -8613
rect 10926 -8911 10942 -8613
rect 10880 -8923 10942 -8911
rect 10972 -8613 11038 -8601
rect 10972 -8911 10988 -8613
rect 11022 -8911 11038 -8613
rect 10972 -8923 11038 -8911
rect 11068 -8613 11134 -8601
rect 11068 -8911 11084 -8613
rect 11118 -8911 11134 -8613
rect 11068 -8923 11134 -8911
rect 11164 -8613 11230 -8601
rect 11164 -8911 11180 -8613
rect 11214 -8911 11230 -8613
rect 11164 -8923 11230 -8911
rect 11260 -8613 11326 -8601
rect 11260 -8911 11276 -8613
rect 11310 -8911 11326 -8613
rect 11260 -8923 11326 -8911
rect 11356 -8613 11422 -8601
rect 11356 -8911 11372 -8613
rect 11406 -8911 11422 -8613
rect 11356 -8923 11422 -8911
rect 11452 -8613 11518 -8601
rect 11452 -8911 11468 -8613
rect 11502 -8911 11518 -8613
rect 11452 -8923 11518 -8911
rect 11548 -8613 11614 -8601
rect 11548 -8911 11564 -8613
rect 11598 -8911 11614 -8613
rect 11548 -8923 11614 -8911
rect 11644 -8613 11706 -8601
rect 11644 -8911 11660 -8613
rect 11694 -8911 11706 -8613
rect 11644 -8923 11706 -8911
rect -21846 -8976 -21632 -8960
rect -22088 -8996 -22026 -8984
rect -23583 -9022 -23369 -9010
rect -21846 -9010 -21834 -8976
rect -21640 -9010 -21632 -8976
rect -21846 -9022 -21632 -9010
rect -20530 -8962 -20468 -8950
rect -20530 -9152 -20518 -8962
rect -20484 -9152 -20468 -8962
rect -20530 -9164 -20468 -9152
rect -20438 -8962 -20372 -8950
rect -20438 -9152 -20422 -8962
rect -20388 -9152 -20372 -8962
rect -20438 -9164 -20372 -9152
rect -20342 -8962 -20276 -8950
rect -20342 -9152 -20326 -8962
rect -20292 -9152 -20276 -8962
rect -20342 -9164 -20276 -9152
rect -20246 -8962 -20180 -8950
rect -20246 -9152 -20230 -8962
rect -20196 -9152 -20180 -8962
rect -20246 -9164 -20180 -9152
rect -20150 -8962 -20084 -8950
rect -20150 -9152 -20134 -8962
rect -20100 -9152 -20084 -8962
rect -20150 -9164 -20084 -9152
rect -20054 -8962 -19988 -8950
rect -20054 -9152 -20038 -8962
rect -20004 -9152 -19988 -8962
rect -20054 -9164 -19988 -9152
rect -19958 -8962 -19896 -8950
rect -19958 -9152 -19942 -8962
rect -19908 -9152 -19896 -8962
rect -19958 -9164 -19896 -9152
rect -19421 -8962 -19359 -8950
rect -19421 -9152 -19409 -8962
rect -19375 -9152 -19359 -8962
rect -19421 -9164 -19359 -9152
rect -19329 -8962 -19263 -8950
rect -19329 -9152 -19313 -8962
rect -19279 -9152 -19263 -8962
rect -19329 -9164 -19263 -9152
rect -19233 -8962 -19167 -8950
rect -19233 -9152 -19217 -8962
rect -19183 -9152 -19167 -8962
rect -19233 -9164 -19167 -9152
rect -19137 -8962 -19071 -8950
rect -19137 -9152 -19121 -8962
rect -19087 -9152 -19071 -8962
rect -19137 -9164 -19071 -9152
rect -19041 -8962 -18975 -8950
rect -19041 -9152 -19025 -8962
rect -18991 -9152 -18975 -8962
rect -19041 -9164 -18975 -9152
rect -18945 -8962 -18879 -8950
rect -18945 -9152 -18929 -8962
rect -18895 -9152 -18879 -8962
rect -18945 -9164 -18879 -9152
rect -18849 -8962 -18787 -8950
rect -18849 -9152 -18833 -8962
rect -18799 -9152 -18787 -8962
rect -18849 -9164 -18787 -9152
rect -18539 -8962 -18477 -8950
rect -18539 -9152 -18527 -8962
rect -18493 -9152 -18477 -8962
rect -18539 -9164 -18477 -9152
rect -18447 -8962 -18381 -8950
rect -18447 -9152 -18431 -8962
rect -18397 -9152 -18381 -8962
rect -18447 -9164 -18381 -9152
rect -18351 -8962 -18285 -8950
rect -18351 -9152 -18335 -8962
rect -18301 -9152 -18285 -8962
rect -18351 -9164 -18285 -9152
rect -18255 -8962 -18189 -8950
rect -18255 -9152 -18239 -8962
rect -18205 -9152 -18189 -8962
rect -18255 -9164 -18189 -9152
rect -18159 -8962 -18093 -8950
rect -18159 -9152 -18143 -8962
rect -18109 -9152 -18093 -8962
rect -18159 -9164 -18093 -9152
rect -18063 -8962 -17997 -8950
rect -18063 -9152 -18047 -8962
rect -18013 -9152 -17997 -8962
rect -18063 -9164 -17997 -9152
rect -17967 -8962 -17905 -8950
rect -17967 -9152 -17951 -8962
rect -17917 -9152 -17905 -8962
rect -17967 -9164 -17905 -9152
rect -17239 -8962 -17177 -8950
rect -17239 -9152 -17227 -8962
rect -17193 -9152 -17177 -8962
rect -17239 -9164 -17177 -9152
rect -17147 -8962 -17081 -8950
rect -17147 -9152 -17131 -8962
rect -17097 -9152 -17081 -8962
rect -17147 -9164 -17081 -9152
rect -17051 -8962 -16985 -8950
rect -17051 -9152 -17035 -8962
rect -17001 -9152 -16985 -8962
rect -17051 -9164 -16985 -9152
rect -16955 -8962 -16889 -8950
rect -16955 -9152 -16939 -8962
rect -16905 -9152 -16889 -8962
rect -16955 -9164 -16889 -9152
rect -16859 -8962 -16793 -8950
rect -16859 -9152 -16843 -8962
rect -16809 -9152 -16793 -8962
rect -16859 -9164 -16793 -9152
rect -16763 -8962 -16697 -8950
rect -16763 -9152 -16747 -8962
rect -16713 -9152 -16697 -8962
rect -16763 -9164 -16697 -9152
rect -16667 -8962 -16605 -8950
rect -16667 -9152 -16651 -8962
rect -16617 -9152 -16605 -8962
rect -16667 -9164 -16605 -9152
rect -16130 -8962 -16068 -8950
rect -16130 -9152 -16118 -8962
rect -16084 -9152 -16068 -8962
rect -16130 -9164 -16068 -9152
rect -16038 -8962 -15972 -8950
rect -16038 -9152 -16022 -8962
rect -15988 -9152 -15972 -8962
rect -16038 -9164 -15972 -9152
rect -15942 -8962 -15876 -8950
rect -15942 -9152 -15926 -8962
rect -15892 -9152 -15876 -8962
rect -15942 -9164 -15876 -9152
rect -15846 -8962 -15780 -8950
rect -15846 -9152 -15830 -8962
rect -15796 -9152 -15780 -8962
rect -15846 -9164 -15780 -9152
rect -15750 -8962 -15684 -8950
rect -15750 -9152 -15734 -8962
rect -15700 -9152 -15684 -8962
rect -15750 -9164 -15684 -9152
rect -15654 -8962 -15588 -8950
rect -15654 -9152 -15638 -8962
rect -15604 -9152 -15588 -8962
rect -15654 -9164 -15588 -9152
rect -15558 -8962 -15496 -8950
rect -15558 -9152 -15542 -8962
rect -15508 -9152 -15496 -8962
rect -15558 -9164 -15496 -9152
rect -15248 -8962 -15186 -8950
rect -15248 -9152 -15236 -8962
rect -15202 -9152 -15186 -8962
rect -15248 -9164 -15186 -9152
rect -15156 -8962 -15090 -8950
rect -15156 -9152 -15140 -8962
rect -15106 -9152 -15090 -8962
rect -15156 -9164 -15090 -9152
rect -15060 -8962 -14994 -8950
rect -15060 -9152 -15044 -8962
rect -15010 -9152 -14994 -8962
rect -15060 -9164 -14994 -9152
rect -14964 -8962 -14898 -8950
rect -14964 -9152 -14948 -8962
rect -14914 -9152 -14898 -8962
rect -14964 -9164 -14898 -9152
rect -14868 -8962 -14802 -8950
rect -14868 -9152 -14852 -8962
rect -14818 -9152 -14802 -8962
rect -14868 -9164 -14802 -9152
rect -14772 -8962 -14706 -8950
rect -14772 -9152 -14756 -8962
rect -14722 -9152 -14706 -8962
rect -14772 -9164 -14706 -9152
rect -14676 -8962 -14614 -8950
rect -14676 -9152 -14660 -8962
rect -14626 -9152 -14614 -8962
rect -14676 -9164 -14614 -9152
rect -13948 -8962 -13886 -8950
rect -13948 -9152 -13936 -8962
rect -13902 -9152 -13886 -8962
rect -13948 -9164 -13886 -9152
rect -13856 -8962 -13790 -8950
rect -13856 -9152 -13840 -8962
rect -13806 -9152 -13790 -8962
rect -13856 -9164 -13790 -9152
rect -13760 -8962 -13694 -8950
rect -13760 -9152 -13744 -8962
rect -13710 -9152 -13694 -8962
rect -13760 -9164 -13694 -9152
rect -13664 -8962 -13598 -8950
rect -13664 -9152 -13648 -8962
rect -13614 -9152 -13598 -8962
rect -13664 -9164 -13598 -9152
rect -13568 -8962 -13502 -8950
rect -13568 -9152 -13552 -8962
rect -13518 -9152 -13502 -8962
rect -13568 -9164 -13502 -9152
rect -13472 -8962 -13406 -8950
rect -13472 -9152 -13456 -8962
rect -13422 -9152 -13406 -8962
rect -13472 -9164 -13406 -9152
rect -13376 -8962 -13314 -8950
rect -13376 -9152 -13360 -8962
rect -13326 -9152 -13314 -8962
rect -13376 -9164 -13314 -9152
rect -12839 -8962 -12777 -8950
rect -12839 -9152 -12827 -8962
rect -12793 -9152 -12777 -8962
rect -12839 -9164 -12777 -9152
rect -12747 -8962 -12681 -8950
rect -12747 -9152 -12731 -8962
rect -12697 -9152 -12681 -8962
rect -12747 -9164 -12681 -9152
rect -12651 -8962 -12585 -8950
rect -12651 -9152 -12635 -8962
rect -12601 -9152 -12585 -8962
rect -12651 -9164 -12585 -9152
rect -12555 -8962 -12489 -8950
rect -12555 -9152 -12539 -8962
rect -12505 -9152 -12489 -8962
rect -12555 -9164 -12489 -9152
rect -12459 -8962 -12393 -8950
rect -12459 -9152 -12443 -8962
rect -12409 -9152 -12393 -8962
rect -12459 -9164 -12393 -9152
rect -12363 -8962 -12297 -8950
rect -12363 -9152 -12347 -8962
rect -12313 -9152 -12297 -8962
rect -12363 -9164 -12297 -9152
rect -12267 -8962 -12205 -8950
rect -12267 -9152 -12251 -8962
rect -12217 -9152 -12205 -8962
rect -12267 -9164 -12205 -9152
rect -11957 -8962 -11895 -8950
rect -11957 -9152 -11945 -8962
rect -11911 -9152 -11895 -8962
rect -11957 -9164 -11895 -9152
rect -11865 -8962 -11799 -8950
rect -11865 -9152 -11849 -8962
rect -11815 -9152 -11799 -8962
rect -11865 -9164 -11799 -9152
rect -11769 -8962 -11703 -8950
rect -11769 -9152 -11753 -8962
rect -11719 -9152 -11703 -8962
rect -11769 -9164 -11703 -9152
rect -11673 -8962 -11607 -8950
rect -11673 -9152 -11657 -8962
rect -11623 -9152 -11607 -8962
rect -11673 -9164 -11607 -9152
rect -11577 -8962 -11511 -8950
rect -11577 -9152 -11561 -8962
rect -11527 -9152 -11511 -8962
rect -11577 -9164 -11511 -9152
rect -11481 -8962 -11415 -8950
rect -11481 -9152 -11465 -8962
rect -11431 -9152 -11415 -8962
rect -11481 -9164 -11415 -9152
rect -11385 -8962 -11323 -8950
rect -11385 -9152 -11369 -8962
rect -11335 -9152 -11323 -8962
rect -11385 -9164 -11323 -9152
rect -10657 -8962 -10595 -8950
rect -10657 -9152 -10645 -8962
rect -10611 -9152 -10595 -8962
rect -10657 -9164 -10595 -9152
rect -10565 -8962 -10499 -8950
rect -10565 -9152 -10549 -8962
rect -10515 -9152 -10499 -8962
rect -10565 -9164 -10499 -9152
rect -10469 -8962 -10403 -8950
rect -10469 -9152 -10453 -8962
rect -10419 -9152 -10403 -8962
rect -10469 -9164 -10403 -9152
rect -10373 -8962 -10307 -8950
rect -10373 -9152 -10357 -8962
rect -10323 -9152 -10307 -8962
rect -10373 -9164 -10307 -9152
rect -10277 -8962 -10211 -8950
rect -10277 -9152 -10261 -8962
rect -10227 -9152 -10211 -8962
rect -10277 -9164 -10211 -9152
rect -10181 -8962 -10115 -8950
rect -10181 -9152 -10165 -8962
rect -10131 -9152 -10115 -8962
rect -10181 -9164 -10115 -9152
rect -10085 -8962 -10023 -8950
rect -10085 -9152 -10069 -8962
rect -10035 -9152 -10023 -8962
rect -10085 -9164 -10023 -9152
rect -9548 -8962 -9486 -8950
rect -9548 -9152 -9536 -8962
rect -9502 -9152 -9486 -8962
rect -9548 -9164 -9486 -9152
rect -9456 -8962 -9390 -8950
rect -9456 -9152 -9440 -8962
rect -9406 -9152 -9390 -8962
rect -9456 -9164 -9390 -9152
rect -9360 -8962 -9294 -8950
rect -9360 -9152 -9344 -8962
rect -9310 -9152 -9294 -8962
rect -9360 -9164 -9294 -9152
rect -9264 -8962 -9198 -8950
rect -9264 -9152 -9248 -8962
rect -9214 -9152 -9198 -8962
rect -9264 -9164 -9198 -9152
rect -9168 -8962 -9102 -8950
rect -9168 -9152 -9152 -8962
rect -9118 -9152 -9102 -8962
rect -9168 -9164 -9102 -9152
rect -9072 -8962 -9006 -8950
rect -9072 -9152 -9056 -8962
rect -9022 -9152 -9006 -8962
rect -9072 -9164 -9006 -9152
rect -8976 -8962 -8914 -8950
rect -8976 -9152 -8960 -8962
rect -8926 -9152 -8914 -8962
rect -8976 -9164 -8914 -9152
rect -8666 -8962 -8604 -8950
rect -8666 -9152 -8654 -8962
rect -8620 -9152 -8604 -8962
rect -8666 -9164 -8604 -9152
rect -8574 -8962 -8508 -8950
rect -8574 -9152 -8558 -8962
rect -8524 -9152 -8508 -8962
rect -8574 -9164 -8508 -9152
rect -8478 -8962 -8412 -8950
rect -8478 -9152 -8462 -8962
rect -8428 -9152 -8412 -8962
rect -8478 -9164 -8412 -9152
rect -8382 -8962 -8316 -8950
rect -8382 -9152 -8366 -8962
rect -8332 -9152 -8316 -8962
rect -8382 -9164 -8316 -9152
rect -8286 -8962 -8220 -8950
rect -8286 -9152 -8270 -8962
rect -8236 -9152 -8220 -8962
rect -8286 -9164 -8220 -9152
rect -8190 -8962 -8124 -8950
rect -8190 -9152 -8174 -8962
rect -8140 -9152 -8124 -8962
rect -8190 -9164 -8124 -9152
rect -8094 -8962 -8032 -8950
rect -8094 -9152 -8078 -8962
rect -8044 -9152 -8032 -8962
rect -8094 -9164 -8032 -9152
rect 5658 -9673 5872 -9661
rect 5658 -9707 5670 -9673
rect 5860 -9707 5872 -9673
rect 6098 -9673 6312 -9661
rect 5658 -9723 5872 -9707
rect 5658 -9769 5872 -9753
rect 5658 -9803 5670 -9769
rect 5864 -9803 5872 -9769
rect 5658 -9819 5872 -9803
rect 5658 -9865 5872 -9849
rect 5658 -9899 5670 -9865
rect 5860 -9899 5872 -9865
rect 5658 -9915 5872 -9899
rect 5658 -9961 5872 -9945
rect 5658 -9995 5670 -9961
rect 5864 -9995 5872 -9961
rect 6098 -9707 6110 -9673
rect 6300 -9707 6312 -9673
rect 6538 -9673 6752 -9661
rect 6098 -9723 6312 -9707
rect 6098 -9769 6312 -9753
rect 6098 -9803 6110 -9769
rect 6304 -9803 6312 -9769
rect 6098 -9819 6312 -9803
rect 6098 -9865 6312 -9849
rect 6098 -9899 6110 -9865
rect 6300 -9899 6312 -9865
rect 6098 -9915 6312 -9899
rect 6098 -9961 6312 -9945
rect 5658 -10007 5872 -9995
rect 6098 -9995 6110 -9961
rect 6304 -9995 6312 -9961
rect 6538 -9707 6550 -9673
rect 6740 -9707 6752 -9673
rect 6538 -9723 6752 -9707
rect 6538 -9769 6752 -9753
rect 6538 -9803 6550 -9769
rect 6744 -9803 6752 -9769
rect 6538 -9819 6752 -9803
rect 6538 -9865 6752 -9849
rect 6538 -9899 6550 -9865
rect 6740 -9899 6752 -9865
rect 6538 -9915 6752 -9899
rect 6538 -9961 6752 -9945
rect 6098 -10007 6312 -9995
rect 6538 -9995 6550 -9961
rect 6744 -9995 6752 -9961
rect 6538 -10007 6752 -9995
rect 7138 -10377 7200 -10365
rect -20737 -10525 -20679 -10513
rect -23583 -10660 -23369 -10648
rect -24396 -10766 -24334 -10754
rect -24396 -10956 -24384 -10766
rect -24350 -10956 -24334 -10766
rect -24396 -10968 -24334 -10956
rect -24304 -10766 -24238 -10754
rect -24304 -10956 -24288 -10766
rect -24254 -10956 -24238 -10766
rect -24304 -10968 -24238 -10956
rect -24208 -10766 -24142 -10754
rect -24208 -10956 -24192 -10766
rect -24158 -10956 -24142 -10766
rect -24208 -10968 -24142 -10956
rect -24112 -10766 -24046 -10754
rect -24112 -10956 -24096 -10766
rect -24062 -10956 -24046 -10766
rect -24112 -10968 -24046 -10956
rect -24016 -10766 -23950 -10754
rect -24016 -10956 -24000 -10766
rect -23966 -10956 -23950 -10766
rect -24016 -10968 -23950 -10956
rect -23920 -10766 -23854 -10754
rect -23920 -10956 -23904 -10766
rect -23870 -10956 -23854 -10766
rect -23920 -10968 -23854 -10956
rect -23824 -10766 -23762 -10754
rect -23824 -10956 -23808 -10766
rect -23774 -10956 -23762 -10766
rect -23583 -10694 -23571 -10660
rect -23381 -10694 -23369 -10660
rect -23583 -10710 -23369 -10694
rect -21850 -10660 -21636 -10648
rect -23583 -10756 -23369 -10740
rect -23583 -10790 -23571 -10756
rect -23377 -10790 -23369 -10756
rect -23583 -10806 -23369 -10790
rect -22659 -10766 -22597 -10754
rect -23583 -10852 -23369 -10836
rect -23583 -10886 -23571 -10852
rect -23381 -10886 -23369 -10852
rect -23583 -10902 -23369 -10886
rect -23583 -10948 -23369 -10932
rect -23824 -10968 -23762 -10956
rect -23583 -10982 -23571 -10948
rect -23377 -10982 -23369 -10948
rect -22659 -10956 -22647 -10766
rect -22613 -10956 -22597 -10766
rect -22659 -10968 -22597 -10956
rect -22567 -10766 -22501 -10754
rect -22567 -10956 -22551 -10766
rect -22517 -10956 -22501 -10766
rect -22567 -10968 -22501 -10956
rect -22471 -10766 -22405 -10754
rect -22471 -10956 -22455 -10766
rect -22421 -10956 -22405 -10766
rect -22471 -10968 -22405 -10956
rect -22375 -10766 -22309 -10754
rect -22375 -10956 -22359 -10766
rect -22325 -10956 -22309 -10766
rect -22375 -10968 -22309 -10956
rect -22279 -10766 -22213 -10754
rect -22279 -10956 -22263 -10766
rect -22229 -10956 -22213 -10766
rect -22279 -10968 -22213 -10956
rect -22183 -10766 -22117 -10754
rect -22183 -10956 -22167 -10766
rect -22133 -10956 -22117 -10766
rect -22183 -10968 -22117 -10956
rect -22087 -10766 -22025 -10754
rect -22087 -10956 -22071 -10766
rect -22037 -10956 -22025 -10766
rect -21850 -10694 -21838 -10660
rect -21648 -10694 -21636 -10660
rect -21850 -10710 -21636 -10694
rect -21850 -10756 -21636 -10740
rect -21850 -10790 -21838 -10756
rect -21644 -10790 -21636 -10756
rect -21850 -10806 -21636 -10790
rect -21850 -10852 -21636 -10836
rect -21850 -10886 -21838 -10852
rect -21648 -10886 -21636 -10852
rect -21850 -10902 -21636 -10886
rect -21850 -10948 -21636 -10932
rect -22087 -10968 -22025 -10956
rect -23583 -10994 -23369 -10982
rect -21850 -10982 -21838 -10948
rect -21644 -10982 -21636 -10948
rect -21850 -10994 -21636 -10982
rect -20737 -11051 -20725 -10525
rect -20691 -11051 -20679 -10525
rect -20737 -11063 -20679 -11051
rect -20649 -10525 -20587 -10513
rect -20649 -11051 -20637 -10525
rect -20603 -11051 -20587 -10525
rect -20649 -11063 -20587 -11051
rect -20557 -10525 -20491 -10513
rect -20557 -11051 -20541 -10525
rect -20507 -11051 -20491 -10525
rect -20557 -11063 -20491 -11051
rect -20461 -10525 -20395 -10513
rect -20461 -11051 -20445 -10525
rect -20411 -11051 -20395 -10525
rect -20461 -11063 -20395 -11051
rect -20365 -10525 -20299 -10513
rect -20365 -11051 -20349 -10525
rect -20315 -11051 -20299 -10525
rect -20365 -11063 -20299 -11051
rect -20269 -10525 -20203 -10513
rect -20269 -11051 -20253 -10525
rect -20219 -11051 -20203 -10525
rect -20269 -11063 -20203 -11051
rect -20173 -10525 -20107 -10513
rect -20173 -11051 -20157 -10525
rect -20123 -11051 -20107 -10525
rect -20173 -11063 -20107 -11051
rect -20077 -10525 -20011 -10513
rect -20077 -11051 -20061 -10525
rect -20027 -11051 -20011 -10525
rect -20077 -11063 -20011 -11051
rect -19981 -10525 -19915 -10513
rect -19981 -11051 -19965 -10525
rect -19931 -11051 -19915 -10525
rect -19981 -11063 -19915 -11051
rect -19885 -10525 -19819 -10513
rect -19885 -11051 -19869 -10525
rect -19835 -11051 -19819 -10525
rect -19885 -11063 -19819 -11051
rect -19789 -10525 -19723 -10513
rect -19789 -11051 -19773 -10525
rect -19739 -11051 -19723 -10525
rect -19789 -11063 -19723 -11051
rect -19693 -10525 -19627 -10513
rect -19693 -11051 -19677 -10525
rect -19643 -11051 -19627 -10525
rect -19693 -11063 -19627 -11051
rect -19597 -10525 -19531 -10513
rect -19597 -11051 -19581 -10525
rect -19547 -11051 -19531 -10525
rect -19597 -11063 -19531 -11051
rect -19501 -10525 -19439 -10513
rect -19501 -11051 -19485 -10525
rect -19451 -11051 -19439 -10525
rect -19501 -11063 -19439 -11051
rect -19409 -10525 -19351 -10513
rect -19409 -11051 -19397 -10525
rect -19363 -11051 -19351 -10525
rect -19409 -11063 -19351 -11051
rect -19178 -10525 -19120 -10513
rect -19178 -11051 -19166 -10525
rect -19132 -11051 -19120 -10525
rect -19178 -11063 -19120 -11051
rect -19090 -10525 -19028 -10513
rect -19090 -11051 -19078 -10525
rect -19044 -11051 -19028 -10525
rect -19090 -11063 -19028 -11051
rect -18998 -10525 -18932 -10513
rect -18998 -11051 -18982 -10525
rect -18948 -11051 -18932 -10525
rect -18998 -11063 -18932 -11051
rect -18902 -10525 -18836 -10513
rect -18902 -11051 -18886 -10525
rect -18852 -11051 -18836 -10525
rect -18902 -11063 -18836 -11051
rect -18806 -10525 -18740 -10513
rect -18806 -11051 -18790 -10525
rect -18756 -11051 -18740 -10525
rect -18806 -11063 -18740 -11051
rect -18710 -10525 -18644 -10513
rect -18710 -11051 -18694 -10525
rect -18660 -11051 -18644 -10525
rect -18710 -11063 -18644 -11051
rect -18614 -10525 -18548 -10513
rect -18614 -11051 -18598 -10525
rect -18564 -11051 -18548 -10525
rect -18614 -11063 -18548 -11051
rect -18518 -10525 -18452 -10513
rect -18518 -11051 -18502 -10525
rect -18468 -11051 -18452 -10525
rect -18518 -11063 -18452 -11051
rect -18422 -10525 -18356 -10513
rect -18422 -11051 -18406 -10525
rect -18372 -11051 -18356 -10525
rect -18422 -11063 -18356 -11051
rect -18326 -10525 -18260 -10513
rect -18326 -11051 -18310 -10525
rect -18276 -11051 -18260 -10525
rect -18326 -11063 -18260 -11051
rect -18230 -10525 -18164 -10513
rect -18230 -11051 -18214 -10525
rect -18180 -11051 -18164 -10525
rect -18230 -11063 -18164 -11051
rect -18134 -10525 -18068 -10513
rect -18134 -11051 -18118 -10525
rect -18084 -11051 -18068 -10525
rect -18134 -11063 -18068 -11051
rect -18038 -10525 -17972 -10513
rect -18038 -11051 -18022 -10525
rect -17988 -11051 -17972 -10525
rect -18038 -11063 -17972 -11051
rect -17942 -10525 -17880 -10513
rect -17942 -11051 -17926 -10525
rect -17892 -11051 -17880 -10525
rect -17942 -11063 -17880 -11051
rect -17850 -10525 -17792 -10513
rect -17850 -11051 -17838 -10525
rect -17804 -11051 -17792 -10525
rect -17850 -11063 -17792 -11051
rect -17446 -10525 -17388 -10513
rect -17446 -11051 -17434 -10525
rect -17400 -11051 -17388 -10525
rect -17446 -11063 -17388 -11051
rect -17358 -10525 -17296 -10513
rect -17358 -11051 -17346 -10525
rect -17312 -11051 -17296 -10525
rect -17358 -11063 -17296 -11051
rect -17266 -10525 -17200 -10513
rect -17266 -11051 -17250 -10525
rect -17216 -11051 -17200 -10525
rect -17266 -11063 -17200 -11051
rect -17170 -10525 -17104 -10513
rect -17170 -11051 -17154 -10525
rect -17120 -11051 -17104 -10525
rect -17170 -11063 -17104 -11051
rect -17074 -10525 -17008 -10513
rect -17074 -11051 -17058 -10525
rect -17024 -11051 -17008 -10525
rect -17074 -11063 -17008 -11051
rect -16978 -10525 -16912 -10513
rect -16978 -11051 -16962 -10525
rect -16928 -11051 -16912 -10525
rect -16978 -11063 -16912 -11051
rect -16882 -10525 -16816 -10513
rect -16882 -11051 -16866 -10525
rect -16832 -11051 -16816 -10525
rect -16882 -11063 -16816 -11051
rect -16786 -10525 -16720 -10513
rect -16786 -11051 -16770 -10525
rect -16736 -11051 -16720 -10525
rect -16786 -11063 -16720 -11051
rect -16690 -10525 -16624 -10513
rect -16690 -11051 -16674 -10525
rect -16640 -11051 -16624 -10525
rect -16690 -11063 -16624 -11051
rect -16594 -10525 -16528 -10513
rect -16594 -11051 -16578 -10525
rect -16544 -11051 -16528 -10525
rect -16594 -11063 -16528 -11051
rect -16498 -10525 -16432 -10513
rect -16498 -11051 -16482 -10525
rect -16448 -11051 -16432 -10525
rect -16498 -11063 -16432 -11051
rect -16402 -10525 -16336 -10513
rect -16402 -11051 -16386 -10525
rect -16352 -11051 -16336 -10525
rect -16402 -11063 -16336 -11051
rect -16306 -10525 -16240 -10513
rect -16306 -11051 -16290 -10525
rect -16256 -11051 -16240 -10525
rect -16306 -11063 -16240 -11051
rect -16210 -10525 -16148 -10513
rect -16210 -11051 -16194 -10525
rect -16160 -11051 -16148 -10525
rect -16210 -11063 -16148 -11051
rect -16118 -10525 -16060 -10513
rect -16118 -11051 -16106 -10525
rect -16072 -11051 -16060 -10525
rect -16118 -11063 -16060 -11051
rect -15887 -10525 -15829 -10513
rect -15887 -11051 -15875 -10525
rect -15841 -11051 -15829 -10525
rect -15887 -11063 -15829 -11051
rect -15799 -10525 -15737 -10513
rect -15799 -11051 -15787 -10525
rect -15753 -11051 -15737 -10525
rect -15799 -11063 -15737 -11051
rect -15707 -10525 -15641 -10513
rect -15707 -11051 -15691 -10525
rect -15657 -11051 -15641 -10525
rect -15707 -11063 -15641 -11051
rect -15611 -10525 -15545 -10513
rect -15611 -11051 -15595 -10525
rect -15561 -11051 -15545 -10525
rect -15611 -11063 -15545 -11051
rect -15515 -10525 -15449 -10513
rect -15515 -11051 -15499 -10525
rect -15465 -11051 -15449 -10525
rect -15515 -11063 -15449 -11051
rect -15419 -10525 -15353 -10513
rect -15419 -11051 -15403 -10525
rect -15369 -11051 -15353 -10525
rect -15419 -11063 -15353 -11051
rect -15323 -10525 -15257 -10513
rect -15323 -11051 -15307 -10525
rect -15273 -11051 -15257 -10525
rect -15323 -11063 -15257 -11051
rect -15227 -10525 -15161 -10513
rect -15227 -11051 -15211 -10525
rect -15177 -11051 -15161 -10525
rect -15227 -11063 -15161 -11051
rect -15131 -10525 -15065 -10513
rect -15131 -11051 -15115 -10525
rect -15081 -11051 -15065 -10525
rect -15131 -11063 -15065 -11051
rect -15035 -10525 -14969 -10513
rect -15035 -11051 -15019 -10525
rect -14985 -11051 -14969 -10525
rect -15035 -11063 -14969 -11051
rect -14939 -10525 -14873 -10513
rect -14939 -11051 -14923 -10525
rect -14889 -11051 -14873 -10525
rect -14939 -11063 -14873 -11051
rect -14843 -10525 -14777 -10513
rect -14843 -11051 -14827 -10525
rect -14793 -11051 -14777 -10525
rect -14843 -11063 -14777 -11051
rect -14747 -10525 -14681 -10513
rect -14747 -11051 -14731 -10525
rect -14697 -11051 -14681 -10525
rect -14747 -11063 -14681 -11051
rect -14651 -10525 -14589 -10513
rect -14651 -11051 -14635 -10525
rect -14601 -11051 -14589 -10525
rect -14651 -11063 -14589 -11051
rect -14559 -10525 -14501 -10513
rect -14559 -11051 -14547 -10525
rect -14513 -11051 -14501 -10525
rect -14559 -11063 -14501 -11051
rect -14155 -10525 -14097 -10513
rect -14155 -11051 -14143 -10525
rect -14109 -11051 -14097 -10525
rect -14155 -11063 -14097 -11051
rect -14067 -10525 -14005 -10513
rect -14067 -11051 -14055 -10525
rect -14021 -11051 -14005 -10525
rect -14067 -11063 -14005 -11051
rect -13975 -10525 -13909 -10513
rect -13975 -11051 -13959 -10525
rect -13925 -11051 -13909 -10525
rect -13975 -11063 -13909 -11051
rect -13879 -10525 -13813 -10513
rect -13879 -11051 -13863 -10525
rect -13829 -11051 -13813 -10525
rect -13879 -11063 -13813 -11051
rect -13783 -10525 -13717 -10513
rect -13783 -11051 -13767 -10525
rect -13733 -11051 -13717 -10525
rect -13783 -11063 -13717 -11051
rect -13687 -10525 -13621 -10513
rect -13687 -11051 -13671 -10525
rect -13637 -11051 -13621 -10525
rect -13687 -11063 -13621 -11051
rect -13591 -10525 -13525 -10513
rect -13591 -11051 -13575 -10525
rect -13541 -11051 -13525 -10525
rect -13591 -11063 -13525 -11051
rect -13495 -10525 -13429 -10513
rect -13495 -11051 -13479 -10525
rect -13445 -11051 -13429 -10525
rect -13495 -11063 -13429 -11051
rect -13399 -10525 -13333 -10513
rect -13399 -11051 -13383 -10525
rect -13349 -11051 -13333 -10525
rect -13399 -11063 -13333 -11051
rect -13303 -10525 -13237 -10513
rect -13303 -11051 -13287 -10525
rect -13253 -11051 -13237 -10525
rect -13303 -11063 -13237 -11051
rect -13207 -10525 -13141 -10513
rect -13207 -11051 -13191 -10525
rect -13157 -11051 -13141 -10525
rect -13207 -11063 -13141 -11051
rect -13111 -10525 -13045 -10513
rect -13111 -11051 -13095 -10525
rect -13061 -11051 -13045 -10525
rect -13111 -11063 -13045 -11051
rect -13015 -10525 -12949 -10513
rect -13015 -11051 -12999 -10525
rect -12965 -11051 -12949 -10525
rect -13015 -11063 -12949 -11051
rect -12919 -10525 -12857 -10513
rect -12919 -11051 -12903 -10525
rect -12869 -11051 -12857 -10525
rect -12919 -11063 -12857 -11051
rect -12827 -10525 -12769 -10513
rect -12827 -11051 -12815 -10525
rect -12781 -11051 -12769 -10525
rect -12827 -11063 -12769 -11051
rect -12596 -10525 -12538 -10513
rect -12596 -11051 -12584 -10525
rect -12550 -11051 -12538 -10525
rect -12596 -11063 -12538 -11051
rect -12508 -10525 -12446 -10513
rect -12508 -11051 -12496 -10525
rect -12462 -11051 -12446 -10525
rect -12508 -11063 -12446 -11051
rect -12416 -10525 -12350 -10513
rect -12416 -11051 -12400 -10525
rect -12366 -11051 -12350 -10525
rect -12416 -11063 -12350 -11051
rect -12320 -10525 -12254 -10513
rect -12320 -11051 -12304 -10525
rect -12270 -11051 -12254 -10525
rect -12320 -11063 -12254 -11051
rect -12224 -10525 -12158 -10513
rect -12224 -11051 -12208 -10525
rect -12174 -11051 -12158 -10525
rect -12224 -11063 -12158 -11051
rect -12128 -10525 -12062 -10513
rect -12128 -11051 -12112 -10525
rect -12078 -11051 -12062 -10525
rect -12128 -11063 -12062 -11051
rect -12032 -10525 -11966 -10513
rect -12032 -11051 -12016 -10525
rect -11982 -11051 -11966 -10525
rect -12032 -11063 -11966 -11051
rect -11936 -10525 -11870 -10513
rect -11936 -11051 -11920 -10525
rect -11886 -11051 -11870 -10525
rect -11936 -11063 -11870 -11051
rect -11840 -10525 -11774 -10513
rect -11840 -11051 -11824 -10525
rect -11790 -11051 -11774 -10525
rect -11840 -11063 -11774 -11051
rect -11744 -10525 -11678 -10513
rect -11744 -11051 -11728 -10525
rect -11694 -11051 -11678 -10525
rect -11744 -11063 -11678 -11051
rect -11648 -10525 -11582 -10513
rect -11648 -11051 -11632 -10525
rect -11598 -11051 -11582 -10525
rect -11648 -11063 -11582 -11051
rect -11552 -10525 -11486 -10513
rect -11552 -11051 -11536 -10525
rect -11502 -11051 -11486 -10525
rect -11552 -11063 -11486 -11051
rect -11456 -10525 -11390 -10513
rect -11456 -11051 -11440 -10525
rect -11406 -11051 -11390 -10525
rect -11456 -11063 -11390 -11051
rect -11360 -10525 -11298 -10513
rect -11360 -11051 -11344 -10525
rect -11310 -11051 -11298 -10525
rect -11360 -11063 -11298 -11051
rect -11268 -10525 -11210 -10513
rect -11268 -11051 -11256 -10525
rect -11222 -11051 -11210 -10525
rect -11268 -11063 -11210 -11051
rect -10864 -10525 -10806 -10513
rect -10864 -11051 -10852 -10525
rect -10818 -11051 -10806 -10525
rect -10864 -11063 -10806 -11051
rect -10776 -10525 -10714 -10513
rect -10776 -11051 -10764 -10525
rect -10730 -11051 -10714 -10525
rect -10776 -11063 -10714 -11051
rect -10684 -10525 -10618 -10513
rect -10684 -11051 -10668 -10525
rect -10634 -11051 -10618 -10525
rect -10684 -11063 -10618 -11051
rect -10588 -10525 -10522 -10513
rect -10588 -11051 -10572 -10525
rect -10538 -11051 -10522 -10525
rect -10588 -11063 -10522 -11051
rect -10492 -10525 -10426 -10513
rect -10492 -11051 -10476 -10525
rect -10442 -11051 -10426 -10525
rect -10492 -11063 -10426 -11051
rect -10396 -10525 -10330 -10513
rect -10396 -11051 -10380 -10525
rect -10346 -11051 -10330 -10525
rect -10396 -11063 -10330 -11051
rect -10300 -10525 -10234 -10513
rect -10300 -11051 -10284 -10525
rect -10250 -11051 -10234 -10525
rect -10300 -11063 -10234 -11051
rect -10204 -10525 -10138 -10513
rect -10204 -11051 -10188 -10525
rect -10154 -11051 -10138 -10525
rect -10204 -11063 -10138 -11051
rect -10108 -10525 -10042 -10513
rect -10108 -11051 -10092 -10525
rect -10058 -11051 -10042 -10525
rect -10108 -11063 -10042 -11051
rect -10012 -10525 -9946 -10513
rect -10012 -11051 -9996 -10525
rect -9962 -11051 -9946 -10525
rect -10012 -11063 -9946 -11051
rect -9916 -10525 -9850 -10513
rect -9916 -11051 -9900 -10525
rect -9866 -11051 -9850 -10525
rect -9916 -11063 -9850 -11051
rect -9820 -10525 -9754 -10513
rect -9820 -11051 -9804 -10525
rect -9770 -11051 -9754 -10525
rect -9820 -11063 -9754 -11051
rect -9724 -10525 -9658 -10513
rect -9724 -11051 -9708 -10525
rect -9674 -11051 -9658 -10525
rect -9724 -11063 -9658 -11051
rect -9628 -10525 -9566 -10513
rect -9628 -11051 -9612 -10525
rect -9578 -11051 -9566 -10525
rect -9628 -11063 -9566 -11051
rect -9536 -10525 -9478 -10513
rect -9536 -11051 -9524 -10525
rect -9490 -11051 -9478 -10525
rect -9536 -11063 -9478 -11051
rect -9305 -10525 -9247 -10513
rect -9305 -11051 -9293 -10525
rect -9259 -11051 -9247 -10525
rect -9305 -11063 -9247 -11051
rect -9217 -10525 -9155 -10513
rect -9217 -11051 -9205 -10525
rect -9171 -11051 -9155 -10525
rect -9217 -11063 -9155 -11051
rect -9125 -10525 -9059 -10513
rect -9125 -11051 -9109 -10525
rect -9075 -11051 -9059 -10525
rect -9125 -11063 -9059 -11051
rect -9029 -10525 -8963 -10513
rect -9029 -11051 -9013 -10525
rect -8979 -11051 -8963 -10525
rect -9029 -11063 -8963 -11051
rect -8933 -10525 -8867 -10513
rect -8933 -11051 -8917 -10525
rect -8883 -11051 -8867 -10525
rect -8933 -11063 -8867 -11051
rect -8837 -10525 -8771 -10513
rect -8837 -11051 -8821 -10525
rect -8787 -11051 -8771 -10525
rect -8837 -11063 -8771 -11051
rect -8741 -10525 -8675 -10513
rect -8741 -11051 -8725 -10525
rect -8691 -11051 -8675 -10525
rect -8741 -11063 -8675 -11051
rect -8645 -10525 -8579 -10513
rect -8645 -11051 -8629 -10525
rect -8595 -11051 -8579 -10525
rect -8645 -11063 -8579 -11051
rect -8549 -10525 -8483 -10513
rect -8549 -11051 -8533 -10525
rect -8499 -11051 -8483 -10525
rect -8549 -11063 -8483 -11051
rect -8453 -10525 -8387 -10513
rect -8453 -11051 -8437 -10525
rect -8403 -11051 -8387 -10525
rect -8453 -11063 -8387 -11051
rect -8357 -10525 -8291 -10513
rect -8357 -11051 -8341 -10525
rect -8307 -11051 -8291 -10525
rect -8357 -11063 -8291 -11051
rect -8261 -10525 -8195 -10513
rect -8261 -11051 -8245 -10525
rect -8211 -11051 -8195 -10525
rect -8261 -11063 -8195 -11051
rect -8165 -10525 -8099 -10513
rect -8165 -11051 -8149 -10525
rect -8115 -11051 -8099 -10525
rect -8165 -11063 -8099 -11051
rect -8069 -10525 -8007 -10513
rect -8069 -11051 -8053 -10525
rect -8019 -11051 -8007 -10525
rect -8069 -11063 -8007 -11051
rect -7977 -10525 -7919 -10513
rect -7977 -11051 -7965 -10525
rect -7931 -11051 -7919 -10525
rect 7138 -10675 7150 -10377
rect 7184 -10675 7200 -10377
rect 7138 -10687 7200 -10675
rect 7230 -10377 7296 -10365
rect 7230 -10675 7246 -10377
rect 7280 -10675 7296 -10377
rect 7230 -10687 7296 -10675
rect 7326 -10377 7392 -10365
rect 7326 -10675 7342 -10377
rect 7376 -10675 7392 -10377
rect 7326 -10687 7392 -10675
rect 7422 -10377 7488 -10365
rect 7422 -10675 7438 -10377
rect 7472 -10675 7488 -10377
rect 7422 -10687 7488 -10675
rect 7518 -10377 7584 -10365
rect 7518 -10675 7534 -10377
rect 7568 -10675 7584 -10377
rect 7518 -10687 7584 -10675
rect 7614 -10377 7680 -10365
rect 7614 -10675 7630 -10377
rect 7664 -10675 7680 -10377
rect 7614 -10687 7680 -10675
rect 7710 -10377 7776 -10365
rect 7710 -10675 7726 -10377
rect 7760 -10675 7776 -10377
rect 7710 -10687 7776 -10675
rect 7806 -10377 7872 -10365
rect 7806 -10675 7822 -10377
rect 7856 -10675 7872 -10377
rect 7806 -10687 7872 -10675
rect 7902 -10377 7964 -10365
rect 7902 -10675 7918 -10377
rect 7952 -10675 7964 -10377
rect 7902 -10687 7964 -10675
rect 8086 -10377 8148 -10365
rect 8086 -10675 8098 -10377
rect 8132 -10675 8148 -10377
rect 8086 -10687 8148 -10675
rect 8178 -10377 8244 -10365
rect 8178 -10675 8194 -10377
rect 8228 -10675 8244 -10377
rect 8178 -10687 8244 -10675
rect 8274 -10377 8340 -10365
rect 8274 -10675 8290 -10377
rect 8324 -10675 8340 -10377
rect 8274 -10687 8340 -10675
rect 8370 -10377 8436 -10365
rect 8370 -10675 8386 -10377
rect 8420 -10675 8436 -10377
rect 8370 -10687 8436 -10675
rect 8466 -10377 8532 -10365
rect 8466 -10675 8482 -10377
rect 8516 -10675 8532 -10377
rect 8466 -10687 8532 -10675
rect 8562 -10377 8628 -10365
rect 8562 -10675 8578 -10377
rect 8612 -10675 8628 -10377
rect 8562 -10687 8628 -10675
rect 8658 -10377 8724 -10365
rect 8658 -10675 8674 -10377
rect 8708 -10675 8724 -10377
rect 8658 -10687 8724 -10675
rect 8754 -10377 8820 -10365
rect 8754 -10675 8770 -10377
rect 8804 -10675 8820 -10377
rect 8754 -10687 8820 -10675
rect 8850 -10377 8912 -10365
rect 8850 -10675 8866 -10377
rect 8900 -10675 8912 -10377
rect 8850 -10687 8912 -10675
rect 9022 -10377 9084 -10365
rect 9022 -10675 9034 -10377
rect 9068 -10675 9084 -10377
rect 9022 -10687 9084 -10675
rect 9114 -10377 9180 -10365
rect 9114 -10675 9130 -10377
rect 9164 -10675 9180 -10377
rect 9114 -10687 9180 -10675
rect 9210 -10377 9276 -10365
rect 9210 -10675 9226 -10377
rect 9260 -10675 9276 -10377
rect 9210 -10687 9276 -10675
rect 9306 -10377 9372 -10365
rect 9306 -10675 9322 -10377
rect 9356 -10675 9372 -10377
rect 9306 -10687 9372 -10675
rect 9402 -10377 9468 -10365
rect 9402 -10675 9418 -10377
rect 9452 -10675 9468 -10377
rect 9402 -10687 9468 -10675
rect 9498 -10377 9564 -10365
rect 9498 -10675 9514 -10377
rect 9548 -10675 9564 -10377
rect 9498 -10687 9564 -10675
rect 9594 -10377 9660 -10365
rect 9594 -10675 9610 -10377
rect 9644 -10675 9660 -10377
rect 9594 -10687 9660 -10675
rect 9690 -10377 9756 -10365
rect 9690 -10675 9706 -10377
rect 9740 -10675 9756 -10377
rect 9690 -10687 9756 -10675
rect 9786 -10377 9848 -10365
rect 9786 -10675 9802 -10377
rect 9836 -10675 9848 -10377
rect 9786 -10687 9848 -10675
rect 9953 -10377 10015 -10365
rect 9953 -10675 9965 -10377
rect 9999 -10675 10015 -10377
rect 9953 -10687 10015 -10675
rect 10045 -10377 10111 -10365
rect 10045 -10675 10061 -10377
rect 10095 -10675 10111 -10377
rect 10045 -10687 10111 -10675
rect 10141 -10377 10207 -10365
rect 10141 -10675 10157 -10377
rect 10191 -10675 10207 -10377
rect 10141 -10687 10207 -10675
rect 10237 -10377 10303 -10365
rect 10237 -10675 10253 -10377
rect 10287 -10675 10303 -10377
rect 10237 -10687 10303 -10675
rect 10333 -10377 10399 -10365
rect 10333 -10675 10349 -10377
rect 10383 -10675 10399 -10377
rect 10333 -10687 10399 -10675
rect 10429 -10377 10495 -10365
rect 10429 -10675 10445 -10377
rect 10479 -10675 10495 -10377
rect 10429 -10687 10495 -10675
rect 10525 -10377 10591 -10365
rect 10525 -10675 10541 -10377
rect 10575 -10675 10591 -10377
rect 10525 -10687 10591 -10675
rect 10621 -10377 10687 -10365
rect 10621 -10675 10637 -10377
rect 10671 -10675 10687 -10377
rect 10621 -10687 10687 -10675
rect 10717 -10377 10779 -10365
rect 10717 -10675 10733 -10377
rect 10767 -10675 10779 -10377
rect 10717 -10687 10779 -10675
rect 10880 -10377 10942 -10365
rect 10880 -10675 10892 -10377
rect 10926 -10675 10942 -10377
rect 10880 -10687 10942 -10675
rect 10972 -10377 11038 -10365
rect 10972 -10675 10988 -10377
rect 11022 -10675 11038 -10377
rect 10972 -10687 11038 -10675
rect 11068 -10377 11134 -10365
rect 11068 -10675 11084 -10377
rect 11118 -10675 11134 -10377
rect 11068 -10687 11134 -10675
rect 11164 -10377 11230 -10365
rect 11164 -10675 11180 -10377
rect 11214 -10675 11230 -10377
rect 11164 -10687 11230 -10675
rect 11260 -10377 11326 -10365
rect 11260 -10675 11276 -10377
rect 11310 -10675 11326 -10377
rect 11260 -10687 11326 -10675
rect 11356 -10377 11422 -10365
rect 11356 -10675 11372 -10377
rect 11406 -10675 11422 -10377
rect 11356 -10687 11422 -10675
rect 11452 -10377 11518 -10365
rect 11452 -10675 11468 -10377
rect 11502 -10675 11518 -10377
rect 11452 -10687 11518 -10675
rect 11548 -10377 11614 -10365
rect 11548 -10675 11564 -10377
rect 11598 -10675 11614 -10377
rect 11548 -10687 11614 -10675
rect 11644 -10377 11706 -10365
rect 11644 -10675 11660 -10377
rect 11694 -10675 11706 -10377
rect 11644 -10687 11706 -10675
rect -7977 -11063 -7919 -11051
rect 11773 -11587 11835 -11575
rect 11773 -11819 11785 -11587
rect 11819 -11819 11835 -11587
rect 11773 -11831 11835 -11819
rect 11865 -11587 11931 -11575
rect 11865 -11819 11881 -11587
rect 11915 -11819 11931 -11587
rect 11865 -11831 11931 -11819
rect 11961 -11587 12027 -11575
rect 11961 -11819 11977 -11587
rect 12011 -11819 12027 -11587
rect 11961 -11831 12027 -11819
rect 12057 -11587 12123 -11575
rect 12057 -11819 12073 -11587
rect 12107 -11819 12123 -11587
rect 12057 -11831 12123 -11819
rect 12153 -11587 12219 -11575
rect 12153 -11819 12169 -11587
rect 12203 -11819 12219 -11587
rect 12153 -11831 12219 -11819
rect 12249 -11587 12315 -11575
rect 12249 -11819 12265 -11587
rect 12299 -11819 12315 -11587
rect 12249 -11831 12315 -11819
rect 12345 -11587 12411 -11575
rect 12345 -11819 12361 -11587
rect 12395 -11819 12411 -11587
rect 12345 -11831 12411 -11819
rect 12441 -11587 12507 -11575
rect 12441 -11819 12457 -11587
rect 12491 -11819 12507 -11587
rect 12441 -11831 12507 -11819
rect 12537 -11587 12603 -11575
rect 12537 -11819 12553 -11587
rect 12587 -11819 12603 -11587
rect 12537 -11831 12603 -11819
rect 12633 -11587 12699 -11575
rect 12633 -11819 12649 -11587
rect 12683 -11819 12699 -11587
rect 12633 -11831 12699 -11819
rect 12729 -11587 12791 -11575
rect 12729 -11819 12745 -11587
rect 12779 -11819 12791 -11587
rect 12923 -11691 13137 -11679
rect 12729 -11831 12791 -11819
rect -23583 -11952 -23369 -11940
rect -24396 -12058 -24334 -12046
rect -24396 -12248 -24384 -12058
rect -24350 -12248 -24334 -12058
rect -24396 -12260 -24334 -12248
rect -24304 -12058 -24238 -12046
rect -24304 -12248 -24288 -12058
rect -24254 -12248 -24238 -12058
rect -24304 -12260 -24238 -12248
rect -24208 -12058 -24142 -12046
rect -24208 -12248 -24192 -12058
rect -24158 -12248 -24142 -12058
rect -24208 -12260 -24142 -12248
rect -24112 -12058 -24046 -12046
rect -24112 -12248 -24096 -12058
rect -24062 -12248 -24046 -12058
rect -24112 -12260 -24046 -12248
rect -24016 -12058 -23950 -12046
rect -24016 -12248 -24000 -12058
rect -23966 -12248 -23950 -12058
rect -24016 -12260 -23950 -12248
rect -23920 -12058 -23854 -12046
rect -23920 -12248 -23904 -12058
rect -23870 -12248 -23854 -12058
rect -23920 -12260 -23854 -12248
rect -23824 -12058 -23762 -12046
rect -23824 -12248 -23808 -12058
rect -23774 -12248 -23762 -12058
rect -23583 -11986 -23571 -11952
rect -23381 -11986 -23369 -11952
rect -23583 -12002 -23369 -11986
rect -21854 -11952 -21640 -11940
rect -23583 -12048 -23369 -12032
rect -23583 -12082 -23571 -12048
rect -23377 -12082 -23369 -12048
rect -23583 -12098 -23369 -12082
rect -22659 -12058 -22597 -12046
rect -23583 -12144 -23369 -12128
rect -23583 -12178 -23571 -12144
rect -23381 -12178 -23369 -12144
rect -23583 -12194 -23369 -12178
rect -23583 -12240 -23369 -12224
rect -23824 -12260 -23762 -12248
rect -23583 -12274 -23571 -12240
rect -23377 -12274 -23369 -12240
rect -22659 -12248 -22647 -12058
rect -22613 -12248 -22597 -12058
rect -22659 -12260 -22597 -12248
rect -22567 -12058 -22501 -12046
rect -22567 -12248 -22551 -12058
rect -22517 -12248 -22501 -12058
rect -22567 -12260 -22501 -12248
rect -22471 -12058 -22405 -12046
rect -22471 -12248 -22455 -12058
rect -22421 -12248 -22405 -12058
rect -22471 -12260 -22405 -12248
rect -22375 -12058 -22309 -12046
rect -22375 -12248 -22359 -12058
rect -22325 -12248 -22309 -12058
rect -22375 -12260 -22309 -12248
rect -22279 -12058 -22213 -12046
rect -22279 -12248 -22263 -12058
rect -22229 -12248 -22213 -12058
rect -22279 -12260 -22213 -12248
rect -22183 -12058 -22117 -12046
rect -22183 -12248 -22167 -12058
rect -22133 -12248 -22117 -12058
rect -22183 -12260 -22117 -12248
rect -22087 -12058 -22025 -12046
rect -22087 -12248 -22071 -12058
rect -22037 -12248 -22025 -12058
rect -21854 -11986 -21842 -11952
rect -21652 -11986 -21640 -11952
rect -21854 -12002 -21640 -11986
rect -21854 -12048 -21640 -12032
rect -21854 -12082 -21842 -12048
rect -21648 -12082 -21640 -12048
rect -21854 -12098 -21640 -12082
rect -21854 -12144 -21640 -12128
rect -21854 -12178 -21842 -12144
rect -21652 -12178 -21640 -12144
rect -21854 -12194 -21640 -12178
rect -21854 -12240 -21640 -12224
rect -22087 -12260 -22025 -12248
rect -23583 -12286 -23369 -12274
rect -21854 -12274 -21842 -12240
rect -21648 -12274 -21640 -12240
rect -21854 -12286 -21640 -12274
rect -20530 -12226 -20468 -12214
rect -20530 -12416 -20518 -12226
rect -20484 -12416 -20468 -12226
rect -20530 -12428 -20468 -12416
rect -20438 -12226 -20372 -12214
rect -20438 -12416 -20422 -12226
rect -20388 -12416 -20372 -12226
rect -20438 -12428 -20372 -12416
rect -20342 -12226 -20276 -12214
rect -20342 -12416 -20326 -12226
rect -20292 -12416 -20276 -12226
rect -20342 -12428 -20276 -12416
rect -20246 -12226 -20180 -12214
rect -20246 -12416 -20230 -12226
rect -20196 -12416 -20180 -12226
rect -20246 -12428 -20180 -12416
rect -20150 -12226 -20084 -12214
rect -20150 -12416 -20134 -12226
rect -20100 -12416 -20084 -12226
rect -20150 -12428 -20084 -12416
rect -20054 -12226 -19988 -12214
rect -20054 -12416 -20038 -12226
rect -20004 -12416 -19988 -12226
rect -20054 -12428 -19988 -12416
rect -19958 -12226 -19896 -12214
rect -19958 -12416 -19942 -12226
rect -19908 -12416 -19896 -12226
rect -19958 -12428 -19896 -12416
rect -19421 -12226 -19359 -12214
rect -19421 -12416 -19409 -12226
rect -19375 -12416 -19359 -12226
rect -19421 -12428 -19359 -12416
rect -19329 -12226 -19263 -12214
rect -19329 -12416 -19313 -12226
rect -19279 -12416 -19263 -12226
rect -19329 -12428 -19263 -12416
rect -19233 -12226 -19167 -12214
rect -19233 -12416 -19217 -12226
rect -19183 -12416 -19167 -12226
rect -19233 -12428 -19167 -12416
rect -19137 -12226 -19071 -12214
rect -19137 -12416 -19121 -12226
rect -19087 -12416 -19071 -12226
rect -19137 -12428 -19071 -12416
rect -19041 -12226 -18975 -12214
rect -19041 -12416 -19025 -12226
rect -18991 -12416 -18975 -12226
rect -19041 -12428 -18975 -12416
rect -18945 -12226 -18879 -12214
rect -18945 -12416 -18929 -12226
rect -18895 -12416 -18879 -12226
rect -18945 -12428 -18879 -12416
rect -18849 -12226 -18787 -12214
rect -18849 -12416 -18833 -12226
rect -18799 -12416 -18787 -12226
rect -18849 -12428 -18787 -12416
rect -18539 -12226 -18477 -12214
rect -18539 -12416 -18527 -12226
rect -18493 -12416 -18477 -12226
rect -18539 -12428 -18477 -12416
rect -18447 -12226 -18381 -12214
rect -18447 -12416 -18431 -12226
rect -18397 -12416 -18381 -12226
rect -18447 -12428 -18381 -12416
rect -18351 -12226 -18285 -12214
rect -18351 -12416 -18335 -12226
rect -18301 -12416 -18285 -12226
rect -18351 -12428 -18285 -12416
rect -18255 -12226 -18189 -12214
rect -18255 -12416 -18239 -12226
rect -18205 -12416 -18189 -12226
rect -18255 -12428 -18189 -12416
rect -18159 -12226 -18093 -12214
rect -18159 -12416 -18143 -12226
rect -18109 -12416 -18093 -12226
rect -18159 -12428 -18093 -12416
rect -18063 -12226 -17997 -12214
rect -18063 -12416 -18047 -12226
rect -18013 -12416 -17997 -12226
rect -18063 -12428 -17997 -12416
rect -17967 -12226 -17905 -12214
rect -17967 -12416 -17951 -12226
rect -17917 -12416 -17905 -12226
rect -17967 -12428 -17905 -12416
rect -17239 -12226 -17177 -12214
rect -17239 -12416 -17227 -12226
rect -17193 -12416 -17177 -12226
rect -17239 -12428 -17177 -12416
rect -17147 -12226 -17081 -12214
rect -17147 -12416 -17131 -12226
rect -17097 -12416 -17081 -12226
rect -17147 -12428 -17081 -12416
rect -17051 -12226 -16985 -12214
rect -17051 -12416 -17035 -12226
rect -17001 -12416 -16985 -12226
rect -17051 -12428 -16985 -12416
rect -16955 -12226 -16889 -12214
rect -16955 -12416 -16939 -12226
rect -16905 -12416 -16889 -12226
rect -16955 -12428 -16889 -12416
rect -16859 -12226 -16793 -12214
rect -16859 -12416 -16843 -12226
rect -16809 -12416 -16793 -12226
rect -16859 -12428 -16793 -12416
rect -16763 -12226 -16697 -12214
rect -16763 -12416 -16747 -12226
rect -16713 -12416 -16697 -12226
rect -16763 -12428 -16697 -12416
rect -16667 -12226 -16605 -12214
rect -16667 -12416 -16651 -12226
rect -16617 -12416 -16605 -12226
rect -16667 -12428 -16605 -12416
rect -16130 -12226 -16068 -12214
rect -16130 -12416 -16118 -12226
rect -16084 -12416 -16068 -12226
rect -16130 -12428 -16068 -12416
rect -16038 -12226 -15972 -12214
rect -16038 -12416 -16022 -12226
rect -15988 -12416 -15972 -12226
rect -16038 -12428 -15972 -12416
rect -15942 -12226 -15876 -12214
rect -15942 -12416 -15926 -12226
rect -15892 -12416 -15876 -12226
rect -15942 -12428 -15876 -12416
rect -15846 -12226 -15780 -12214
rect -15846 -12416 -15830 -12226
rect -15796 -12416 -15780 -12226
rect -15846 -12428 -15780 -12416
rect -15750 -12226 -15684 -12214
rect -15750 -12416 -15734 -12226
rect -15700 -12416 -15684 -12226
rect -15750 -12428 -15684 -12416
rect -15654 -12226 -15588 -12214
rect -15654 -12416 -15638 -12226
rect -15604 -12416 -15588 -12226
rect -15654 -12428 -15588 -12416
rect -15558 -12226 -15496 -12214
rect -15558 -12416 -15542 -12226
rect -15508 -12416 -15496 -12226
rect -15558 -12428 -15496 -12416
rect -15248 -12226 -15186 -12214
rect -15248 -12416 -15236 -12226
rect -15202 -12416 -15186 -12226
rect -15248 -12428 -15186 -12416
rect -15156 -12226 -15090 -12214
rect -15156 -12416 -15140 -12226
rect -15106 -12416 -15090 -12226
rect -15156 -12428 -15090 -12416
rect -15060 -12226 -14994 -12214
rect -15060 -12416 -15044 -12226
rect -15010 -12416 -14994 -12226
rect -15060 -12428 -14994 -12416
rect -14964 -12226 -14898 -12214
rect -14964 -12416 -14948 -12226
rect -14914 -12416 -14898 -12226
rect -14964 -12428 -14898 -12416
rect -14868 -12226 -14802 -12214
rect -14868 -12416 -14852 -12226
rect -14818 -12416 -14802 -12226
rect -14868 -12428 -14802 -12416
rect -14772 -12226 -14706 -12214
rect -14772 -12416 -14756 -12226
rect -14722 -12416 -14706 -12226
rect -14772 -12428 -14706 -12416
rect -14676 -12226 -14614 -12214
rect -14676 -12416 -14660 -12226
rect -14626 -12416 -14614 -12226
rect -14676 -12428 -14614 -12416
rect -13948 -12226 -13886 -12214
rect -13948 -12416 -13936 -12226
rect -13902 -12416 -13886 -12226
rect -13948 -12428 -13886 -12416
rect -13856 -12226 -13790 -12214
rect -13856 -12416 -13840 -12226
rect -13806 -12416 -13790 -12226
rect -13856 -12428 -13790 -12416
rect -13760 -12226 -13694 -12214
rect -13760 -12416 -13744 -12226
rect -13710 -12416 -13694 -12226
rect -13760 -12428 -13694 -12416
rect -13664 -12226 -13598 -12214
rect -13664 -12416 -13648 -12226
rect -13614 -12416 -13598 -12226
rect -13664 -12428 -13598 -12416
rect -13568 -12226 -13502 -12214
rect -13568 -12416 -13552 -12226
rect -13518 -12416 -13502 -12226
rect -13568 -12428 -13502 -12416
rect -13472 -12226 -13406 -12214
rect -13472 -12416 -13456 -12226
rect -13422 -12416 -13406 -12226
rect -13472 -12428 -13406 -12416
rect -13376 -12226 -13314 -12214
rect -13376 -12416 -13360 -12226
rect -13326 -12416 -13314 -12226
rect -13376 -12428 -13314 -12416
rect -12839 -12226 -12777 -12214
rect -12839 -12416 -12827 -12226
rect -12793 -12416 -12777 -12226
rect -12839 -12428 -12777 -12416
rect -12747 -12226 -12681 -12214
rect -12747 -12416 -12731 -12226
rect -12697 -12416 -12681 -12226
rect -12747 -12428 -12681 -12416
rect -12651 -12226 -12585 -12214
rect -12651 -12416 -12635 -12226
rect -12601 -12416 -12585 -12226
rect -12651 -12428 -12585 -12416
rect -12555 -12226 -12489 -12214
rect -12555 -12416 -12539 -12226
rect -12505 -12416 -12489 -12226
rect -12555 -12428 -12489 -12416
rect -12459 -12226 -12393 -12214
rect -12459 -12416 -12443 -12226
rect -12409 -12416 -12393 -12226
rect -12459 -12428 -12393 -12416
rect -12363 -12226 -12297 -12214
rect -12363 -12416 -12347 -12226
rect -12313 -12416 -12297 -12226
rect -12363 -12428 -12297 -12416
rect -12267 -12226 -12205 -12214
rect -12267 -12416 -12251 -12226
rect -12217 -12416 -12205 -12226
rect -12267 -12428 -12205 -12416
rect -11957 -12226 -11895 -12214
rect -11957 -12416 -11945 -12226
rect -11911 -12416 -11895 -12226
rect -11957 -12428 -11895 -12416
rect -11865 -12226 -11799 -12214
rect -11865 -12416 -11849 -12226
rect -11815 -12416 -11799 -12226
rect -11865 -12428 -11799 -12416
rect -11769 -12226 -11703 -12214
rect -11769 -12416 -11753 -12226
rect -11719 -12416 -11703 -12226
rect -11769 -12428 -11703 -12416
rect -11673 -12226 -11607 -12214
rect -11673 -12416 -11657 -12226
rect -11623 -12416 -11607 -12226
rect -11673 -12428 -11607 -12416
rect -11577 -12226 -11511 -12214
rect -11577 -12416 -11561 -12226
rect -11527 -12416 -11511 -12226
rect -11577 -12428 -11511 -12416
rect -11481 -12226 -11415 -12214
rect -11481 -12416 -11465 -12226
rect -11431 -12416 -11415 -12226
rect -11481 -12428 -11415 -12416
rect -11385 -12226 -11323 -12214
rect -11385 -12416 -11369 -12226
rect -11335 -12416 -11323 -12226
rect -11385 -12428 -11323 -12416
rect -10657 -12226 -10595 -12214
rect -10657 -12416 -10645 -12226
rect -10611 -12416 -10595 -12226
rect -10657 -12428 -10595 -12416
rect -10565 -12226 -10499 -12214
rect -10565 -12416 -10549 -12226
rect -10515 -12416 -10499 -12226
rect -10565 -12428 -10499 -12416
rect -10469 -12226 -10403 -12214
rect -10469 -12416 -10453 -12226
rect -10419 -12416 -10403 -12226
rect -10469 -12428 -10403 -12416
rect -10373 -12226 -10307 -12214
rect -10373 -12416 -10357 -12226
rect -10323 -12416 -10307 -12226
rect -10373 -12428 -10307 -12416
rect -10277 -12226 -10211 -12214
rect -10277 -12416 -10261 -12226
rect -10227 -12416 -10211 -12226
rect -10277 -12428 -10211 -12416
rect -10181 -12226 -10115 -12214
rect -10181 -12416 -10165 -12226
rect -10131 -12416 -10115 -12226
rect -10181 -12428 -10115 -12416
rect -10085 -12226 -10023 -12214
rect -10085 -12416 -10069 -12226
rect -10035 -12416 -10023 -12226
rect -10085 -12428 -10023 -12416
rect -9548 -12226 -9486 -12214
rect -9548 -12416 -9536 -12226
rect -9502 -12416 -9486 -12226
rect -9548 -12428 -9486 -12416
rect -9456 -12226 -9390 -12214
rect -9456 -12416 -9440 -12226
rect -9406 -12416 -9390 -12226
rect -9456 -12428 -9390 -12416
rect -9360 -12226 -9294 -12214
rect -9360 -12416 -9344 -12226
rect -9310 -12416 -9294 -12226
rect -9360 -12428 -9294 -12416
rect -9264 -12226 -9198 -12214
rect -9264 -12416 -9248 -12226
rect -9214 -12416 -9198 -12226
rect -9264 -12428 -9198 -12416
rect -9168 -12226 -9102 -12214
rect -9168 -12416 -9152 -12226
rect -9118 -12416 -9102 -12226
rect -9168 -12428 -9102 -12416
rect -9072 -12226 -9006 -12214
rect -9072 -12416 -9056 -12226
rect -9022 -12416 -9006 -12226
rect -9072 -12428 -9006 -12416
rect -8976 -12226 -8914 -12214
rect -8976 -12416 -8960 -12226
rect -8926 -12416 -8914 -12226
rect -8976 -12428 -8914 -12416
rect -8666 -12226 -8604 -12214
rect -8666 -12416 -8654 -12226
rect -8620 -12416 -8604 -12226
rect -8666 -12428 -8604 -12416
rect -8574 -12226 -8508 -12214
rect -8574 -12416 -8558 -12226
rect -8524 -12416 -8508 -12226
rect -8574 -12428 -8508 -12416
rect -8478 -12226 -8412 -12214
rect -8478 -12416 -8462 -12226
rect -8428 -12416 -8412 -12226
rect -8478 -12428 -8412 -12416
rect -8382 -12226 -8316 -12214
rect -8382 -12416 -8366 -12226
rect -8332 -12416 -8316 -12226
rect -8382 -12428 -8316 -12416
rect -8286 -12226 -8220 -12214
rect -8286 -12416 -8270 -12226
rect -8236 -12416 -8220 -12226
rect -8286 -12428 -8220 -12416
rect -8190 -12226 -8124 -12214
rect -8190 -12416 -8174 -12226
rect -8140 -12416 -8124 -12226
rect -8190 -12428 -8124 -12416
rect -8094 -12226 -8032 -12214
rect -8094 -12416 -8078 -12226
rect -8044 -12416 -8032 -12226
rect -8094 -12428 -8032 -12416
rect 12923 -11725 12935 -11691
rect 13125 -11725 13137 -11691
rect 12923 -11741 13137 -11725
rect 12923 -11787 13137 -11771
rect 12923 -11821 12935 -11787
rect 13129 -11821 13137 -11787
rect 12923 -11837 13137 -11821
rect 12923 -11883 13137 -11867
rect 12923 -11917 12935 -11883
rect 13125 -11917 13137 -11883
rect 12923 -11933 13137 -11917
rect 12923 -11979 13137 -11963
rect 12923 -12013 12935 -11979
rect 13129 -12013 13137 -11979
rect 12923 -12025 13137 -12013
rect 7138 -13241 7200 -13229
rect 7138 -13539 7150 -13241
rect 7184 -13539 7200 -13241
rect 7138 -13551 7200 -13539
rect 7230 -13241 7296 -13229
rect 7230 -13539 7246 -13241
rect 7280 -13539 7296 -13241
rect 7230 -13551 7296 -13539
rect 7326 -13241 7392 -13229
rect 7326 -13539 7342 -13241
rect 7376 -13539 7392 -13241
rect 7326 -13551 7392 -13539
rect 7422 -13241 7488 -13229
rect 7422 -13539 7438 -13241
rect 7472 -13539 7488 -13241
rect 7422 -13551 7488 -13539
rect 7518 -13241 7584 -13229
rect 7518 -13539 7534 -13241
rect 7568 -13539 7584 -13241
rect 7518 -13551 7584 -13539
rect 7614 -13241 7680 -13229
rect 7614 -13539 7630 -13241
rect 7664 -13539 7680 -13241
rect 7614 -13551 7680 -13539
rect 7710 -13241 7776 -13229
rect 7710 -13539 7726 -13241
rect 7760 -13539 7776 -13241
rect 7710 -13551 7776 -13539
rect 7806 -13241 7872 -13229
rect 7806 -13539 7822 -13241
rect 7856 -13539 7872 -13241
rect 7806 -13551 7872 -13539
rect 7902 -13241 7964 -13229
rect 7902 -13539 7918 -13241
rect 7952 -13539 7964 -13241
rect 7902 -13551 7964 -13539
rect 8086 -13241 8148 -13229
rect 8086 -13539 8098 -13241
rect 8132 -13539 8148 -13241
rect 8086 -13551 8148 -13539
rect 8178 -13241 8244 -13229
rect 8178 -13539 8194 -13241
rect 8228 -13539 8244 -13241
rect 8178 -13551 8244 -13539
rect 8274 -13241 8340 -13229
rect 8274 -13539 8290 -13241
rect 8324 -13539 8340 -13241
rect 8274 -13551 8340 -13539
rect 8370 -13241 8436 -13229
rect 8370 -13539 8386 -13241
rect 8420 -13539 8436 -13241
rect 8370 -13551 8436 -13539
rect 8466 -13241 8532 -13229
rect 8466 -13539 8482 -13241
rect 8516 -13539 8532 -13241
rect 8466 -13551 8532 -13539
rect 8562 -13241 8628 -13229
rect 8562 -13539 8578 -13241
rect 8612 -13539 8628 -13241
rect 8562 -13551 8628 -13539
rect 8658 -13241 8724 -13229
rect 8658 -13539 8674 -13241
rect 8708 -13539 8724 -13241
rect 8658 -13551 8724 -13539
rect 8754 -13241 8820 -13229
rect 8754 -13539 8770 -13241
rect 8804 -13539 8820 -13241
rect 8754 -13551 8820 -13539
rect 8850 -13241 8912 -13229
rect 8850 -13539 8866 -13241
rect 8900 -13539 8912 -13241
rect 8850 -13551 8912 -13539
rect 9022 -13241 9084 -13229
rect 9022 -13539 9034 -13241
rect 9068 -13539 9084 -13241
rect 9022 -13551 9084 -13539
rect 9114 -13241 9180 -13229
rect 9114 -13539 9130 -13241
rect 9164 -13539 9180 -13241
rect 9114 -13551 9180 -13539
rect 9210 -13241 9276 -13229
rect 9210 -13539 9226 -13241
rect 9260 -13539 9276 -13241
rect 9210 -13551 9276 -13539
rect 9306 -13241 9372 -13229
rect 9306 -13539 9322 -13241
rect 9356 -13539 9372 -13241
rect 9306 -13551 9372 -13539
rect 9402 -13241 9468 -13229
rect 9402 -13539 9418 -13241
rect 9452 -13539 9468 -13241
rect 9402 -13551 9468 -13539
rect 9498 -13241 9564 -13229
rect 9498 -13539 9514 -13241
rect 9548 -13539 9564 -13241
rect 9498 -13551 9564 -13539
rect 9594 -13241 9660 -13229
rect 9594 -13539 9610 -13241
rect 9644 -13539 9660 -13241
rect 9594 -13551 9660 -13539
rect 9690 -13241 9756 -13229
rect 9690 -13539 9706 -13241
rect 9740 -13539 9756 -13241
rect 9690 -13551 9756 -13539
rect 9786 -13241 9848 -13229
rect 9786 -13539 9802 -13241
rect 9836 -13539 9848 -13241
rect 9786 -13551 9848 -13539
rect 9953 -13240 10015 -13228
rect 9953 -13538 9965 -13240
rect 9999 -13538 10015 -13240
rect 9953 -13550 10015 -13538
rect 10045 -13240 10111 -13228
rect 10045 -13538 10061 -13240
rect 10095 -13538 10111 -13240
rect 10045 -13550 10111 -13538
rect 10141 -13240 10207 -13228
rect 10141 -13538 10157 -13240
rect 10191 -13538 10207 -13240
rect 10141 -13550 10207 -13538
rect 10237 -13240 10303 -13228
rect 10237 -13538 10253 -13240
rect 10287 -13538 10303 -13240
rect 10237 -13550 10303 -13538
rect 10333 -13240 10399 -13228
rect 10333 -13538 10349 -13240
rect 10383 -13538 10399 -13240
rect 10333 -13550 10399 -13538
rect 10429 -13240 10495 -13228
rect 10429 -13538 10445 -13240
rect 10479 -13538 10495 -13240
rect 10429 -13550 10495 -13538
rect 10525 -13240 10591 -13228
rect 10525 -13538 10541 -13240
rect 10575 -13538 10591 -13240
rect 10525 -13550 10591 -13538
rect 10621 -13240 10687 -13228
rect 10621 -13538 10637 -13240
rect 10671 -13538 10687 -13240
rect 10621 -13550 10687 -13538
rect 10717 -13240 10779 -13228
rect 10717 -13538 10733 -13240
rect 10767 -13538 10779 -13240
rect 10717 -13550 10779 -13538
rect 10880 -13241 10942 -13229
rect 10880 -13539 10892 -13241
rect 10926 -13539 10942 -13241
rect 10880 -13551 10942 -13539
rect 10972 -13241 11038 -13229
rect 10972 -13539 10988 -13241
rect 11022 -13539 11038 -13241
rect 10972 -13551 11038 -13539
rect 11068 -13241 11134 -13229
rect 11068 -13539 11084 -13241
rect 11118 -13539 11134 -13241
rect 11068 -13551 11134 -13539
rect 11164 -13241 11230 -13229
rect 11164 -13539 11180 -13241
rect 11214 -13539 11230 -13241
rect 11164 -13551 11230 -13539
rect 11260 -13241 11326 -13229
rect 11260 -13539 11276 -13241
rect 11310 -13539 11326 -13241
rect 11260 -13551 11326 -13539
rect 11356 -13241 11422 -13229
rect 11356 -13539 11372 -13241
rect 11406 -13539 11422 -13241
rect 11356 -13551 11422 -13539
rect 11452 -13241 11518 -13229
rect 11452 -13539 11468 -13241
rect 11502 -13539 11518 -13241
rect 11452 -13551 11518 -13539
rect 11548 -13241 11614 -13229
rect 11548 -13539 11564 -13241
rect 11598 -13539 11614 -13241
rect 11548 -13551 11614 -13539
rect 11644 -13241 11706 -13229
rect 11644 -13539 11660 -13241
rect 11694 -13539 11706 -13241
rect 11644 -13551 11706 -13539
rect -2112 -13830 -2050 -13818
rect -2112 -14020 -2100 -13830
rect -2066 -14020 -2050 -13830
rect -2112 -14032 -2050 -14020
rect -2020 -13826 -1954 -13818
rect -2020 -14020 -2004 -13826
rect -1970 -14020 -1954 -13826
rect -2020 -14032 -1954 -14020
rect -1924 -13830 -1858 -13818
rect -1924 -14020 -1908 -13830
rect -1874 -14020 -1858 -13830
rect -1924 -14032 -1858 -14020
rect -1828 -13826 -1766 -13818
rect -1828 -14020 -1812 -13826
rect -1778 -14020 -1766 -13826
rect -1828 -14032 -1766 -14020
rect -12316 -14105 -11766 -14093
rect -12316 -14139 -12304 -14105
rect -11778 -14139 -11766 -14105
rect -12316 -14151 -11766 -14139
rect -17677 -14511 -17421 -14499
rect -17677 -14545 -17665 -14511
rect -17433 -14545 -17421 -14511
rect -17677 -14561 -17421 -14545
rect -17677 -14607 -17421 -14591
rect -17677 -14641 -17665 -14607
rect -17433 -14641 -17421 -14607
rect -17677 -14657 -17421 -14641
rect -17677 -14703 -17421 -14687
rect -17677 -14737 -17665 -14703
rect -17433 -14737 -17421 -14703
rect -17677 -14753 -17421 -14737
rect -17677 -14799 -17421 -14783
rect -17677 -14833 -17665 -14799
rect -17433 -14833 -17421 -14799
rect -17677 -14849 -17421 -14833
rect -17677 -14895 -17421 -14879
rect -24449 -14928 -24235 -14916
rect -24449 -14962 -24437 -14928
rect -24247 -14962 -24235 -14928
rect -24449 -14978 -24235 -14962
rect -24449 -15024 -24235 -15008
rect -24449 -15058 -24437 -15024
rect -24247 -15058 -24235 -15024
rect -24449 -15074 -24235 -15058
rect -24449 -15120 -24235 -15104
rect -24449 -15154 -24437 -15120
rect -24247 -15154 -24235 -15120
rect -24449 -15170 -24235 -15154
rect -24449 -15216 -24235 -15200
rect -24449 -15250 -24437 -15216
rect -24247 -15250 -24235 -15216
rect -24449 -15266 -24235 -15250
rect -24449 -15312 -24235 -15296
rect -24449 -15346 -24437 -15312
rect -24247 -15346 -24235 -15312
rect -24449 -15362 -24235 -15346
rect -17677 -14929 -17665 -14895
rect -17433 -14929 -17421 -14895
rect -17677 -14945 -17421 -14929
rect -17677 -14991 -17421 -14975
rect -17677 -15025 -17665 -14991
rect -17433 -15025 -17421 -14991
rect -17677 -15041 -17421 -15025
rect -17677 -15087 -17421 -15071
rect -24449 -15408 -24235 -15392
rect -24449 -15442 -24437 -15408
rect -24247 -15442 -24235 -15408
rect -24449 -15458 -24235 -15442
rect -24449 -15504 -24235 -15488
rect -17677 -15121 -17665 -15087
rect -17433 -15121 -17421 -15087
rect -17677 -15137 -17421 -15121
rect -17677 -15183 -17421 -15167
rect -17677 -15217 -17665 -15183
rect -17433 -15217 -17421 -15183
rect -17677 -15233 -17421 -15217
rect -17677 -15279 -17421 -15263
rect -17677 -15313 -17665 -15279
rect -17433 -15313 -17421 -15279
rect -17677 -15329 -17421 -15313
rect -17677 -15375 -17421 -15359
rect -17677 -15409 -17665 -15375
rect -17433 -15409 -17421 -15375
rect -17677 -15425 -17421 -15409
rect -12316 -14193 -11766 -14181
rect -12316 -14227 -12304 -14193
rect -11778 -14227 -11766 -14193
rect -12316 -14243 -11766 -14227
rect -12316 -14289 -11766 -14273
rect -12316 -14323 -12304 -14289
rect -11778 -14323 -11766 -14289
rect -12316 -14339 -11766 -14323
rect -12316 -14385 -11766 -14369
rect -12316 -14419 -12304 -14385
rect -11778 -14419 -11766 -14385
rect -12316 -14435 -11766 -14419
rect -12316 -14481 -11766 -14465
rect -12316 -14515 -12304 -14481
rect -11778 -14515 -11766 -14481
rect -12316 -14531 -11766 -14515
rect -12316 -14577 -11766 -14561
rect -12316 -14611 -12304 -14577
rect -11778 -14611 -11766 -14577
rect -12316 -14627 -11766 -14611
rect -12316 -14673 -11766 -14657
rect -12316 -14707 -12304 -14673
rect -11778 -14707 -11766 -14673
rect -12316 -14723 -11766 -14707
rect -12316 -14769 -11766 -14753
rect -12316 -14803 -12304 -14769
rect -11778 -14803 -11766 -14769
rect -12316 -14819 -11766 -14803
rect -12316 -14865 -11766 -14849
rect -12316 -14899 -12304 -14865
rect -11778 -14899 -11766 -14865
rect -12316 -14915 -11766 -14899
rect -12316 -14961 -11766 -14945
rect -12316 -14995 -12304 -14961
rect -11778 -14995 -11766 -14961
rect -12316 -15011 -11766 -14995
rect -12316 -15057 -11766 -15041
rect -12316 -15091 -12304 -15057
rect -11778 -15091 -11766 -15057
rect -12316 -15107 -11766 -15091
rect -12316 -15153 -11766 -15137
rect -12316 -15187 -12304 -15153
rect -11778 -15187 -11766 -15153
rect -12316 -15203 -11766 -15187
rect -12316 -15249 -11766 -15233
rect -12316 -15283 -12304 -15249
rect -11778 -15283 -11766 -15249
rect -12316 -15299 -11766 -15283
rect -12316 -15345 -11766 -15329
rect -12316 -15379 -12304 -15345
rect -11778 -15379 -11766 -15345
rect -12316 -15391 -11766 -15379
rect -4828 -14215 -4766 -14203
rect -4828 -14405 -4816 -14215
rect -4782 -14405 -4766 -14215
rect -4828 -14417 -4766 -14405
rect -4736 -14215 -4670 -14203
rect -4736 -14409 -4720 -14215
rect -4686 -14409 -4670 -14215
rect -4736 -14417 -4670 -14409
rect -4640 -14215 -4574 -14203
rect -4640 -14405 -4624 -14215
rect -4590 -14405 -4574 -14215
rect -4640 -14417 -4574 -14405
rect -4544 -14215 -4482 -14203
rect -4544 -14409 -4528 -14215
rect -4494 -14409 -4482 -14215
rect -2112 -14209 -2050 -14197
rect -4544 -14417 -4482 -14409
rect -2112 -14399 -2100 -14209
rect -2066 -14399 -2050 -14209
rect -2112 -14411 -2050 -14399
rect -2020 -14205 -1954 -14197
rect -2020 -14399 -2004 -14205
rect -1970 -14399 -1954 -14205
rect -2020 -14411 -1954 -14399
rect -1924 -14209 -1858 -14197
rect -1924 -14399 -1908 -14209
rect -1874 -14399 -1858 -14209
rect -1924 -14411 -1858 -14399
rect -1828 -14205 -1766 -14197
rect -1828 -14399 -1812 -14205
rect -1778 -14399 -1766 -14205
rect 5658 -14201 5872 -14189
rect -1828 -14411 -1766 -14399
rect 5658 -14235 5670 -14201
rect 5860 -14235 5872 -14201
rect 6098 -14201 6312 -14189
rect 5658 -14251 5872 -14235
rect 5658 -14297 5872 -14281
rect 5658 -14331 5670 -14297
rect 5864 -14331 5872 -14297
rect 5658 -14347 5872 -14331
rect 5658 -14393 5872 -14377
rect 5658 -14427 5670 -14393
rect 5860 -14427 5872 -14393
rect 5658 -14443 5872 -14427
rect 5658 -14489 5872 -14473
rect 5658 -14523 5670 -14489
rect 5864 -14523 5872 -14489
rect 6098 -14235 6110 -14201
rect 6300 -14235 6312 -14201
rect 6538 -14201 6752 -14189
rect 6098 -14251 6312 -14235
rect 6098 -14297 6312 -14281
rect 6098 -14331 6110 -14297
rect 6304 -14331 6312 -14297
rect 6098 -14347 6312 -14331
rect 6098 -14393 6312 -14377
rect 6098 -14427 6110 -14393
rect 6300 -14427 6312 -14393
rect 6098 -14443 6312 -14427
rect 6098 -14489 6312 -14473
rect 5658 -14535 5872 -14523
rect 6098 -14523 6110 -14489
rect 6304 -14523 6312 -14489
rect 6538 -14235 6550 -14201
rect 6740 -14235 6752 -14201
rect 6538 -14251 6752 -14235
rect 6538 -14297 6752 -14281
rect 6538 -14331 6550 -14297
rect 6744 -14331 6752 -14297
rect 6538 -14347 6752 -14331
rect 6538 -14393 6752 -14377
rect 6538 -14427 6550 -14393
rect 6740 -14427 6752 -14393
rect 6538 -14443 6752 -14427
rect 6538 -14489 6752 -14473
rect 6098 -14535 6312 -14523
rect 6538 -14523 6550 -14489
rect 6744 -14523 6752 -14489
rect 6538 -14535 6752 -14523
rect -4828 -14655 -4766 -14643
rect -4828 -14845 -4816 -14655
rect -4782 -14845 -4766 -14655
rect -4828 -14857 -4766 -14845
rect -4736 -14655 -4670 -14643
rect -4736 -14849 -4720 -14655
rect -4686 -14849 -4670 -14655
rect -4736 -14857 -4670 -14849
rect -4640 -14655 -4574 -14643
rect -4640 -14845 -4624 -14655
rect -4590 -14845 -4574 -14655
rect -4640 -14857 -4574 -14845
rect -4544 -14655 -4482 -14643
rect -4544 -14849 -4528 -14655
rect -4494 -14849 -4482 -14655
rect -2112 -14649 -2050 -14637
rect -4544 -14857 -4482 -14849
rect -2112 -14839 -2100 -14649
rect -2066 -14839 -2050 -14649
rect -2112 -14851 -2050 -14839
rect -2020 -14645 -1954 -14637
rect -2020 -14839 -2004 -14645
rect -1970 -14839 -1954 -14645
rect -2020 -14851 -1954 -14839
rect -1924 -14649 -1858 -14637
rect -1924 -14839 -1908 -14649
rect -1874 -14839 -1858 -14649
rect -1924 -14851 -1858 -14839
rect -1828 -14645 -1766 -14637
rect -1828 -14839 -1812 -14645
rect -1778 -14839 -1766 -14645
rect -1828 -14851 -1766 -14839
rect 7138 -14905 7200 -14893
rect -4828 -15034 -4766 -15022
rect -4828 -15224 -4816 -15034
rect -4782 -15224 -4766 -15034
rect -4828 -15236 -4766 -15224
rect -4736 -15034 -4670 -15022
rect -4736 -15228 -4720 -15034
rect -4686 -15228 -4670 -15034
rect -4736 -15236 -4670 -15228
rect -4640 -15034 -4574 -15022
rect -4640 -15224 -4624 -15034
rect -4590 -15224 -4574 -15034
rect -4640 -15236 -4574 -15224
rect -4544 -15034 -4482 -15022
rect -4544 -15228 -4528 -15034
rect -4494 -15228 -4482 -15034
rect -2112 -15028 -2050 -15016
rect -4544 -15236 -4482 -15228
rect -2112 -15218 -2100 -15028
rect -2066 -15218 -2050 -15028
rect -2112 -15230 -2050 -15218
rect -2020 -15024 -1954 -15016
rect -2020 -15218 -2004 -15024
rect -1970 -15218 -1954 -15024
rect -2020 -15230 -1954 -15218
rect -1924 -15028 -1858 -15016
rect -1924 -15218 -1908 -15028
rect -1874 -15218 -1858 -15028
rect -1924 -15230 -1858 -15218
rect -1828 -15024 -1766 -15016
rect -1828 -15218 -1812 -15024
rect -1778 -15218 -1766 -15024
rect -1828 -15230 -1766 -15218
rect 7138 -15203 7150 -14905
rect 7184 -15203 7200 -14905
rect 7138 -15215 7200 -15203
rect 7230 -14905 7296 -14893
rect 7230 -15203 7246 -14905
rect 7280 -15203 7296 -14905
rect 7230 -15215 7296 -15203
rect 7326 -14905 7392 -14893
rect 7326 -15203 7342 -14905
rect 7376 -15203 7392 -14905
rect 7326 -15215 7392 -15203
rect 7422 -14905 7488 -14893
rect 7422 -15203 7438 -14905
rect 7472 -15203 7488 -14905
rect 7422 -15215 7488 -15203
rect 7518 -14905 7584 -14893
rect 7518 -15203 7534 -14905
rect 7568 -15203 7584 -14905
rect 7518 -15215 7584 -15203
rect 7614 -14905 7680 -14893
rect 7614 -15203 7630 -14905
rect 7664 -15203 7680 -14905
rect 7614 -15215 7680 -15203
rect 7710 -14905 7776 -14893
rect 7710 -15203 7726 -14905
rect 7760 -15203 7776 -14905
rect 7710 -15215 7776 -15203
rect 7806 -14905 7872 -14893
rect 7806 -15203 7822 -14905
rect 7856 -15203 7872 -14905
rect 7806 -15215 7872 -15203
rect 7902 -14905 7964 -14893
rect 7902 -15203 7918 -14905
rect 7952 -15203 7964 -14905
rect 7902 -15215 7964 -15203
rect 8086 -14905 8148 -14893
rect 8086 -15203 8098 -14905
rect 8132 -15203 8148 -14905
rect 8086 -15215 8148 -15203
rect 8178 -14905 8244 -14893
rect 8178 -15203 8194 -14905
rect 8228 -15203 8244 -14905
rect 8178 -15215 8244 -15203
rect 8274 -14905 8340 -14893
rect 8274 -15203 8290 -14905
rect 8324 -15203 8340 -14905
rect 8274 -15215 8340 -15203
rect 8370 -14905 8436 -14893
rect 8370 -15203 8386 -14905
rect 8420 -15203 8436 -14905
rect 8370 -15215 8436 -15203
rect 8466 -14905 8532 -14893
rect 8466 -15203 8482 -14905
rect 8516 -15203 8532 -14905
rect 8466 -15215 8532 -15203
rect 8562 -14905 8628 -14893
rect 8562 -15203 8578 -14905
rect 8612 -15203 8628 -14905
rect 8562 -15215 8628 -15203
rect 8658 -14905 8724 -14893
rect 8658 -15203 8674 -14905
rect 8708 -15203 8724 -14905
rect 8658 -15215 8724 -15203
rect 8754 -14905 8820 -14893
rect 8754 -15203 8770 -14905
rect 8804 -15203 8820 -14905
rect 8754 -15215 8820 -15203
rect 8850 -14905 8912 -14893
rect 8850 -15203 8866 -14905
rect 8900 -15203 8912 -14905
rect 8850 -15215 8912 -15203
rect 9022 -14905 9084 -14893
rect 9022 -15203 9034 -14905
rect 9068 -15203 9084 -14905
rect 9022 -15215 9084 -15203
rect 9114 -14905 9180 -14893
rect 9114 -15203 9130 -14905
rect 9164 -15203 9180 -14905
rect 9114 -15215 9180 -15203
rect 9210 -14905 9276 -14893
rect 9210 -15203 9226 -14905
rect 9260 -15203 9276 -14905
rect 9210 -15215 9276 -15203
rect 9306 -14905 9372 -14893
rect 9306 -15203 9322 -14905
rect 9356 -15203 9372 -14905
rect 9306 -15215 9372 -15203
rect 9402 -14905 9468 -14893
rect 9402 -15203 9418 -14905
rect 9452 -15203 9468 -14905
rect 9402 -15215 9468 -15203
rect 9498 -14905 9564 -14893
rect 9498 -15203 9514 -14905
rect 9548 -15203 9564 -14905
rect 9498 -15215 9564 -15203
rect 9594 -14905 9660 -14893
rect 9594 -15203 9610 -14905
rect 9644 -15203 9660 -14905
rect 9594 -15215 9660 -15203
rect 9690 -14905 9756 -14893
rect 9690 -15203 9706 -14905
rect 9740 -15203 9756 -14905
rect 9690 -15215 9756 -15203
rect 9786 -14905 9848 -14893
rect 9786 -15203 9802 -14905
rect 9836 -15203 9848 -14905
rect 9786 -15215 9848 -15203
rect 9953 -14905 10015 -14893
rect 9953 -15203 9965 -14905
rect 9999 -15203 10015 -14905
rect 9953 -15215 10015 -15203
rect 10045 -14905 10111 -14893
rect 10045 -15203 10061 -14905
rect 10095 -15203 10111 -14905
rect 10045 -15215 10111 -15203
rect 10141 -14905 10207 -14893
rect 10141 -15203 10157 -14905
rect 10191 -15203 10207 -14905
rect 10141 -15215 10207 -15203
rect 10237 -14905 10303 -14893
rect 10237 -15203 10253 -14905
rect 10287 -15203 10303 -14905
rect 10237 -15215 10303 -15203
rect 10333 -14905 10399 -14893
rect 10333 -15203 10349 -14905
rect 10383 -15203 10399 -14905
rect 10333 -15215 10399 -15203
rect 10429 -14905 10495 -14893
rect 10429 -15203 10445 -14905
rect 10479 -15203 10495 -14905
rect 10429 -15215 10495 -15203
rect 10525 -14905 10591 -14893
rect 10525 -15203 10541 -14905
rect 10575 -15203 10591 -14905
rect 10525 -15215 10591 -15203
rect 10621 -14905 10687 -14893
rect 10621 -15203 10637 -14905
rect 10671 -15203 10687 -14905
rect 10621 -15215 10687 -15203
rect 10717 -14905 10779 -14893
rect 10717 -15203 10733 -14905
rect 10767 -15203 10779 -14905
rect 10717 -15215 10779 -15203
rect 10880 -14905 10942 -14893
rect 10880 -15203 10892 -14905
rect 10926 -15203 10942 -14905
rect 10880 -15215 10942 -15203
rect 10972 -14905 11038 -14893
rect 10972 -15203 10988 -14905
rect 11022 -15203 11038 -14905
rect 10972 -15215 11038 -15203
rect 11068 -14905 11134 -14893
rect 11068 -15203 11084 -14905
rect 11118 -15203 11134 -14905
rect 11068 -15215 11134 -15203
rect 11164 -14905 11230 -14893
rect 11164 -15203 11180 -14905
rect 11214 -15203 11230 -14905
rect 11164 -15215 11230 -15203
rect 11260 -14905 11326 -14893
rect 11260 -15203 11276 -14905
rect 11310 -15203 11326 -14905
rect 11260 -15215 11326 -15203
rect 11356 -14905 11422 -14893
rect 11356 -15203 11372 -14905
rect 11406 -15203 11422 -14905
rect 11356 -15215 11422 -15203
rect 11452 -14905 11518 -14893
rect 11452 -15203 11468 -14905
rect 11502 -15203 11518 -14905
rect 11452 -15215 11518 -15203
rect 11548 -14905 11614 -14893
rect 11548 -15203 11564 -14905
rect 11598 -15203 11614 -14905
rect 11548 -15215 11614 -15203
rect 11644 -14905 11706 -14893
rect 11644 -15203 11660 -14905
rect 11694 -15203 11706 -14905
rect 11644 -15215 11706 -15203
rect -8179 -15358 -8117 -15346
rect -12316 -15433 -11766 -15421
rect -24449 -15538 -24437 -15504
rect -24247 -15538 -24235 -15504
rect -17677 -15471 -17421 -15455
rect -17677 -15505 -17665 -15471
rect -17433 -15505 -17421 -15471
rect -12316 -15467 -12304 -15433
rect -11778 -15467 -11766 -15433
rect -12316 -15479 -11766 -15467
rect -17677 -15517 -17421 -15505
rect -24449 -15550 -24235 -15538
rect -8179 -15548 -8167 -15358
rect -8133 -15548 -8117 -15358
rect -8179 -15560 -8117 -15548
rect -8087 -15354 -8021 -15346
rect -8087 -15548 -8071 -15354
rect -8037 -15548 -8021 -15354
rect -8087 -15560 -8021 -15548
rect -7991 -15358 -7925 -15346
rect -7991 -15548 -7975 -15358
rect -7941 -15548 -7925 -15358
rect -7991 -15560 -7925 -15548
rect -7895 -15354 -7833 -15346
rect -7895 -15548 -7879 -15354
rect -7845 -15548 -7833 -15354
rect -7895 -15560 -7833 -15548
rect -4828 -15474 -4766 -15462
rect -4828 -15664 -4816 -15474
rect -4782 -15664 -4766 -15474
rect -4828 -15676 -4766 -15664
rect -4736 -15474 -4670 -15462
rect -4736 -15668 -4720 -15474
rect -4686 -15668 -4670 -15474
rect -4736 -15676 -4670 -15668
rect -4640 -15474 -4574 -15462
rect -4640 -15664 -4624 -15474
rect -4590 -15664 -4574 -15474
rect -4640 -15676 -4574 -15664
rect -4544 -15474 -4482 -15462
rect -4544 -15668 -4528 -15474
rect -4494 -15668 -4482 -15474
rect -2112 -15468 -2050 -15456
rect -4544 -15676 -4482 -15668
rect -2112 -15658 -2100 -15468
rect -2066 -15658 -2050 -15468
rect -2112 -15670 -2050 -15658
rect -2020 -15464 -1954 -15456
rect -2020 -15658 -2004 -15464
rect -1970 -15658 -1954 -15464
rect -2020 -15670 -1954 -15658
rect -1924 -15468 -1858 -15456
rect -1924 -15658 -1908 -15468
rect -1874 -15658 -1858 -15468
rect -1924 -15670 -1858 -15658
rect -1828 -15464 -1766 -15456
rect -1828 -15658 -1812 -15464
rect -1778 -15658 -1766 -15464
rect -1828 -15670 -1766 -15658
rect -17677 -15911 -17421 -15899
rect -17677 -15945 -17665 -15911
rect -17433 -15945 -17421 -15911
rect -17677 -15961 -17421 -15945
rect -8178 -15858 -8116 -15846
rect -17677 -16007 -17421 -15991
rect -17677 -16041 -17665 -16007
rect -17433 -16041 -17421 -16007
rect -17677 -16057 -17421 -16041
rect -8178 -16048 -8166 -15858
rect -8132 -16048 -8116 -15858
rect -8178 -16060 -8116 -16048
rect -8086 -15854 -8020 -15846
rect -8086 -16048 -8070 -15854
rect -8036 -16048 -8020 -15854
rect -8086 -16060 -8020 -16048
rect -7990 -15858 -7924 -15846
rect -7990 -16048 -7974 -15858
rect -7940 -16048 -7924 -15858
rect -7990 -16060 -7924 -16048
rect -7894 -15854 -7832 -15846
rect -7894 -16048 -7878 -15854
rect -7844 -16048 -7832 -15854
rect -7894 -16060 -7832 -16048
rect -4828 -15853 -4766 -15841
rect -4828 -16043 -4816 -15853
rect -4782 -16043 -4766 -15853
rect -4828 -16055 -4766 -16043
rect -4736 -15853 -4670 -15841
rect -4736 -16047 -4720 -15853
rect -4686 -16047 -4670 -15853
rect -4736 -16055 -4670 -16047
rect -4640 -15853 -4574 -15841
rect -4640 -16043 -4624 -15853
rect -4590 -16043 -4574 -15853
rect -4640 -16055 -4574 -16043
rect -4544 -15853 -4482 -15841
rect -4544 -16047 -4528 -15853
rect -4494 -16047 -4482 -15853
rect -2112 -15847 -2050 -15835
rect -4544 -16055 -4482 -16047
rect -24448 -16113 -24234 -16101
rect -24448 -16147 -24436 -16113
rect -24246 -16147 -24234 -16113
rect -24448 -16163 -24234 -16147
rect -24448 -16209 -24234 -16193
rect -24448 -16243 -24436 -16209
rect -24246 -16243 -24234 -16209
rect -24448 -16259 -24234 -16243
rect -24448 -16305 -24234 -16289
rect -24448 -16339 -24436 -16305
rect -24246 -16339 -24234 -16305
rect -24448 -16355 -24234 -16339
rect -24448 -16401 -24234 -16385
rect -24448 -16435 -24436 -16401
rect -24246 -16435 -24234 -16401
rect -24448 -16451 -24234 -16435
rect -24448 -16497 -24234 -16481
rect -24448 -16531 -24436 -16497
rect -24246 -16531 -24234 -16497
rect -24448 -16547 -24234 -16531
rect -17677 -16103 -17421 -16087
rect -17677 -16137 -17665 -16103
rect -17433 -16137 -17421 -16103
rect -17677 -16153 -17421 -16137
rect -2112 -16037 -2100 -15847
rect -2066 -16037 -2050 -15847
rect -2112 -16049 -2050 -16037
rect -2020 -15843 -1954 -15835
rect -2020 -16037 -2004 -15843
rect -1970 -16037 -1954 -15843
rect -2020 -16049 -1954 -16037
rect -1924 -15847 -1858 -15835
rect -1924 -16037 -1908 -15847
rect -1874 -16037 -1858 -15847
rect -1924 -16049 -1858 -16037
rect -1828 -15843 -1766 -15835
rect -1828 -16037 -1812 -15843
rect -1778 -16037 -1766 -15843
rect -1828 -16049 -1766 -16037
rect -17677 -16199 -17421 -16183
rect -17677 -16233 -17665 -16199
rect -17433 -16233 -17421 -16199
rect -17677 -16249 -17421 -16233
rect -17677 -16295 -17421 -16279
rect -17677 -16329 -17665 -16295
rect -17433 -16329 -17421 -16295
rect -17677 -16345 -17421 -16329
rect -17677 -16391 -17421 -16375
rect -17677 -16425 -17665 -16391
rect -17433 -16425 -17421 -16391
rect -17677 -16441 -17421 -16425
rect -17677 -16487 -17421 -16471
rect -24448 -16593 -24234 -16577
rect -24448 -16627 -24436 -16593
rect -24246 -16627 -24234 -16593
rect -24448 -16643 -24234 -16627
rect -24448 -16689 -24234 -16673
rect -24448 -16723 -24436 -16689
rect -24246 -16723 -24234 -16689
rect -24448 -16735 -24234 -16723
rect -17677 -16521 -17665 -16487
rect -17433 -16521 -17421 -16487
rect -17677 -16537 -17421 -16521
rect -8179 -16338 -8117 -16326
rect -8179 -16528 -8167 -16338
rect -8133 -16528 -8117 -16338
rect -8179 -16540 -8117 -16528
rect -8087 -16334 -8021 -16326
rect -8087 -16528 -8071 -16334
rect -8037 -16528 -8021 -16334
rect -8087 -16540 -8021 -16528
rect -7991 -16338 -7925 -16326
rect -7991 -16528 -7975 -16338
rect -7941 -16528 -7925 -16338
rect -7991 -16540 -7925 -16528
rect -7895 -16334 -7833 -16326
rect -7895 -16528 -7879 -16334
rect -7845 -16528 -7833 -16334
rect -7895 -16540 -7833 -16528
rect -4828 -16293 -4766 -16281
rect -4828 -16483 -4816 -16293
rect -4782 -16483 -4766 -16293
rect -4828 -16495 -4766 -16483
rect -4736 -16293 -4670 -16281
rect -4736 -16487 -4720 -16293
rect -4686 -16487 -4670 -16293
rect -4736 -16495 -4670 -16487
rect -4640 -16293 -4574 -16281
rect -4640 -16483 -4624 -16293
rect -4590 -16483 -4574 -16293
rect -4640 -16495 -4574 -16483
rect -4544 -16293 -4482 -16281
rect -4544 -16487 -4528 -16293
rect -4494 -16487 -4482 -16293
rect -2112 -16287 -2050 -16275
rect -4544 -16495 -4482 -16487
rect -2112 -16477 -2100 -16287
rect -2066 -16477 -2050 -16287
rect -2112 -16489 -2050 -16477
rect -2020 -16283 -1954 -16275
rect -2020 -16477 -2004 -16283
rect -1970 -16477 -1954 -16283
rect -2020 -16489 -1954 -16477
rect -1924 -16287 -1858 -16275
rect -1924 -16477 -1908 -16287
rect -1874 -16477 -1858 -16287
rect -1924 -16489 -1858 -16477
rect -1828 -16283 -1766 -16275
rect -1828 -16477 -1812 -16283
rect -1778 -16477 -1766 -16283
rect -1828 -16489 -1766 -16477
rect 11773 -16115 11835 -16103
rect 11773 -16347 11785 -16115
rect 11819 -16347 11835 -16115
rect 11773 -16359 11835 -16347
rect 11865 -16115 11931 -16103
rect 11865 -16347 11881 -16115
rect 11915 -16347 11931 -16115
rect 11865 -16359 11931 -16347
rect 11961 -16115 12027 -16103
rect 11961 -16347 11977 -16115
rect 12011 -16347 12027 -16115
rect 11961 -16359 12027 -16347
rect 12057 -16115 12123 -16103
rect 12057 -16347 12073 -16115
rect 12107 -16347 12123 -16115
rect 12057 -16359 12123 -16347
rect 12153 -16115 12219 -16103
rect 12153 -16347 12169 -16115
rect 12203 -16347 12219 -16115
rect 12153 -16359 12219 -16347
rect 12249 -16115 12315 -16103
rect 12249 -16347 12265 -16115
rect 12299 -16347 12315 -16115
rect 12249 -16359 12315 -16347
rect 12345 -16115 12411 -16103
rect 12345 -16347 12361 -16115
rect 12395 -16347 12411 -16115
rect 12345 -16359 12411 -16347
rect 12441 -16115 12507 -16103
rect 12441 -16347 12457 -16115
rect 12491 -16347 12507 -16115
rect 12441 -16359 12507 -16347
rect 12537 -16115 12603 -16103
rect 12537 -16347 12553 -16115
rect 12587 -16347 12603 -16115
rect 12537 -16359 12603 -16347
rect 12633 -16115 12699 -16103
rect 12633 -16347 12649 -16115
rect 12683 -16347 12699 -16115
rect 12633 -16359 12699 -16347
rect 12729 -16115 12791 -16103
rect 12729 -16347 12745 -16115
rect 12779 -16347 12791 -16115
rect 12923 -16219 13137 -16207
rect 12729 -16359 12791 -16347
rect -17677 -16583 -17421 -16567
rect -17677 -16617 -17665 -16583
rect -17433 -16617 -17421 -16583
rect -17677 -16633 -17421 -16617
rect -17677 -16679 -17421 -16663
rect -17677 -16713 -17665 -16679
rect -17433 -16713 -17421 -16679
rect -17677 -16729 -17421 -16713
rect -17677 -16775 -17421 -16759
rect -17677 -16809 -17665 -16775
rect -17433 -16809 -17421 -16775
rect -17677 -16825 -17421 -16809
rect -4828 -16672 -4766 -16660
rect -17677 -16871 -17421 -16855
rect -17677 -16905 -17665 -16871
rect -17433 -16905 -17421 -16871
rect -17677 -16917 -17421 -16905
rect -8179 -16838 -8117 -16826
rect -12314 -16921 -11764 -16909
rect -12314 -16955 -12302 -16921
rect -11776 -16955 -11764 -16921
rect -12314 -16967 -11764 -16955
rect -17677 -17311 -17421 -17299
rect -24443 -17326 -24229 -17314
rect -24443 -17360 -24431 -17326
rect -24241 -17360 -24229 -17326
rect -24443 -17376 -24229 -17360
rect -24443 -17422 -24229 -17406
rect -24443 -17456 -24431 -17422
rect -24241 -17456 -24229 -17422
rect -24443 -17472 -24229 -17456
rect -24443 -17518 -24229 -17502
rect -24443 -17552 -24431 -17518
rect -24241 -17552 -24229 -17518
rect -24443 -17568 -24229 -17552
rect -24443 -17614 -24229 -17598
rect -24443 -17648 -24431 -17614
rect -24241 -17648 -24229 -17614
rect -24443 -17664 -24229 -17648
rect -24443 -17710 -24229 -17694
rect -24443 -17744 -24431 -17710
rect -24241 -17744 -24229 -17710
rect -24443 -17760 -24229 -17744
rect -17677 -17345 -17665 -17311
rect -17433 -17345 -17421 -17311
rect -17677 -17361 -17421 -17345
rect -17677 -17407 -17421 -17391
rect -17677 -17441 -17665 -17407
rect -17433 -17441 -17421 -17407
rect -17677 -17457 -17421 -17441
rect -17677 -17503 -17421 -17487
rect -17677 -17537 -17665 -17503
rect -17433 -17537 -17421 -17503
rect -17677 -17553 -17421 -17537
rect -17677 -17599 -17421 -17583
rect -17677 -17633 -17665 -17599
rect -17433 -17633 -17421 -17599
rect -17677 -17649 -17421 -17633
rect -17677 -17695 -17421 -17679
rect -24443 -17806 -24229 -17790
rect -24443 -17840 -24431 -17806
rect -24241 -17840 -24229 -17806
rect -24443 -17856 -24229 -17840
rect -17677 -17729 -17665 -17695
rect -17433 -17729 -17421 -17695
rect -17677 -17745 -17421 -17729
rect -17677 -17791 -17421 -17775
rect -17677 -17825 -17665 -17791
rect -17433 -17825 -17421 -17791
rect -17677 -17841 -17421 -17825
rect -24443 -17902 -24229 -17886
rect -17677 -17887 -17421 -17871
rect -24443 -17936 -24431 -17902
rect -24241 -17936 -24229 -17902
rect -24443 -17948 -24229 -17936
rect -21618 -18046 -21556 -18034
rect -21618 -18236 -21606 -18046
rect -21572 -18236 -21556 -18046
rect -21618 -18248 -21556 -18236
rect -21526 -18042 -21460 -18034
rect -21526 -18236 -21510 -18042
rect -21476 -18236 -21460 -18042
rect -21526 -18248 -21460 -18236
rect -21430 -18046 -21364 -18034
rect -21430 -18236 -21414 -18046
rect -21380 -18236 -21364 -18046
rect -21430 -18248 -21364 -18236
rect -21334 -18042 -21272 -18034
rect -21334 -18236 -21318 -18042
rect -21284 -18236 -21272 -18042
rect -21334 -18248 -21272 -18236
rect -17677 -17921 -17665 -17887
rect -17433 -17921 -17421 -17887
rect -17677 -17937 -17421 -17921
rect -17677 -17983 -17421 -17967
rect -17677 -18017 -17665 -17983
rect -17433 -18017 -17421 -17983
rect -17677 -18033 -17421 -18017
rect -17677 -18079 -17421 -18063
rect -17677 -18113 -17665 -18079
rect -17433 -18113 -17421 -18079
rect -17677 -18129 -17421 -18113
rect -16027 -17917 -15965 -17905
rect -16027 -18107 -16015 -17917
rect -15981 -18107 -15965 -17917
rect -16027 -18119 -15965 -18107
rect -15935 -17913 -15869 -17905
rect -15935 -18107 -15919 -17913
rect -15885 -18107 -15869 -17913
rect -15935 -18119 -15869 -18107
rect -15839 -17917 -15773 -17905
rect -15839 -18107 -15823 -17917
rect -15789 -18107 -15773 -17917
rect -15839 -18119 -15773 -18107
rect -15743 -17913 -15681 -17905
rect -15743 -18107 -15727 -17913
rect -15693 -18107 -15681 -17913
rect -15743 -18119 -15681 -18107
rect -17677 -18175 -17421 -18159
rect -17677 -18209 -17665 -18175
rect -17433 -18209 -17421 -18175
rect -17677 -18225 -17421 -18209
rect -12314 -17009 -11764 -16997
rect -12314 -17043 -12302 -17009
rect -11776 -17043 -11764 -17009
rect -12314 -17059 -11764 -17043
rect -12314 -17105 -11764 -17089
rect -12314 -17139 -12302 -17105
rect -11776 -17139 -11764 -17105
rect -12314 -17155 -11764 -17139
rect -12314 -17201 -11764 -17185
rect -12314 -17235 -12302 -17201
rect -11776 -17235 -11764 -17201
rect -12314 -17251 -11764 -17235
rect -12314 -17297 -11764 -17281
rect -12314 -17331 -12302 -17297
rect -11776 -17331 -11764 -17297
rect -12314 -17347 -11764 -17331
rect -12314 -17393 -11764 -17377
rect -12314 -17427 -12302 -17393
rect -11776 -17427 -11764 -17393
rect -12314 -17443 -11764 -17427
rect -12314 -17489 -11764 -17473
rect -12314 -17523 -12302 -17489
rect -11776 -17523 -11764 -17489
rect -12314 -17539 -11764 -17523
rect -12314 -17585 -11764 -17569
rect -12314 -17619 -12302 -17585
rect -11776 -17619 -11764 -17585
rect -12314 -17635 -11764 -17619
rect -12314 -17681 -11764 -17665
rect -12314 -17715 -12302 -17681
rect -11776 -17715 -11764 -17681
rect -12314 -17731 -11764 -17715
rect -12314 -17777 -11764 -17761
rect -12314 -17811 -12302 -17777
rect -11776 -17811 -11764 -17777
rect -12314 -17827 -11764 -17811
rect -12314 -17873 -11764 -17857
rect -12314 -17907 -12302 -17873
rect -11776 -17907 -11764 -17873
rect -12314 -17923 -11764 -17907
rect -12314 -17969 -11764 -17953
rect -12314 -18003 -12302 -17969
rect -11776 -18003 -11764 -17969
rect -12314 -18019 -11764 -18003
rect -12314 -18065 -11764 -18049
rect -12314 -18099 -12302 -18065
rect -11776 -18099 -11764 -18065
rect -12314 -18115 -11764 -18099
rect -12314 -18161 -11764 -18145
rect -12314 -18195 -12302 -18161
rect -11776 -18195 -11764 -18161
rect -12314 -18207 -11764 -18195
rect -8179 -17028 -8167 -16838
rect -8133 -17028 -8117 -16838
rect -8179 -17040 -8117 -17028
rect -8087 -16834 -8021 -16826
rect -8087 -17028 -8071 -16834
rect -8037 -17028 -8021 -16834
rect -8087 -17040 -8021 -17028
rect -7991 -16838 -7925 -16826
rect -7991 -17028 -7975 -16838
rect -7941 -17028 -7925 -16838
rect -7991 -17040 -7925 -17028
rect -7895 -16834 -7833 -16826
rect -7895 -17028 -7879 -16834
rect -7845 -17028 -7833 -16834
rect -7895 -17040 -7833 -17028
rect -4828 -16862 -4816 -16672
rect -4782 -16862 -4766 -16672
rect -4828 -16874 -4766 -16862
rect -4736 -16672 -4670 -16660
rect -4736 -16866 -4720 -16672
rect -4686 -16866 -4670 -16672
rect -4736 -16874 -4670 -16866
rect -4640 -16672 -4574 -16660
rect -4640 -16862 -4624 -16672
rect -4590 -16862 -4574 -16672
rect -4640 -16874 -4574 -16862
rect -4544 -16672 -4482 -16660
rect -4544 -16866 -4528 -16672
rect -4494 -16866 -4482 -16672
rect -2112 -16666 -2050 -16654
rect -4544 -16874 -4482 -16866
rect -2112 -16856 -2100 -16666
rect -2066 -16856 -2050 -16666
rect -2112 -16868 -2050 -16856
rect -2020 -16662 -1954 -16654
rect -2020 -16856 -2004 -16662
rect -1970 -16856 -1954 -16662
rect -2020 -16868 -1954 -16856
rect -1924 -16666 -1858 -16654
rect -1924 -16856 -1908 -16666
rect -1874 -16856 -1858 -16666
rect -1924 -16868 -1858 -16856
rect -1828 -16662 -1766 -16654
rect -1828 -16856 -1812 -16662
rect -1778 -16856 -1766 -16662
rect -1828 -16868 -1766 -16856
rect -4828 -17112 -4766 -17100
rect -8179 -17318 -8117 -17306
rect -8179 -17508 -8167 -17318
rect -8133 -17508 -8117 -17318
rect -8179 -17520 -8117 -17508
rect -8087 -17314 -8021 -17306
rect -8087 -17508 -8071 -17314
rect -8037 -17508 -8021 -17314
rect -8087 -17520 -8021 -17508
rect -7991 -17318 -7925 -17306
rect -7991 -17508 -7975 -17318
rect -7941 -17508 -7925 -17318
rect -7991 -17520 -7925 -17508
rect -7895 -17314 -7833 -17306
rect -7895 -17508 -7879 -17314
rect -7845 -17508 -7833 -17314
rect -4828 -17302 -4816 -17112
rect -4782 -17302 -4766 -17112
rect -4828 -17314 -4766 -17302
rect -4736 -17112 -4670 -17100
rect -4736 -17306 -4720 -17112
rect -4686 -17306 -4670 -17112
rect -4736 -17314 -4670 -17306
rect -4640 -17112 -4574 -17100
rect -4640 -17302 -4624 -17112
rect -4590 -17302 -4574 -17112
rect -4640 -17314 -4574 -17302
rect -4544 -17112 -4482 -17100
rect -4544 -17306 -4528 -17112
rect -4494 -17306 -4482 -17112
rect -2112 -17106 -2050 -17094
rect -4544 -17314 -4482 -17306
rect -7895 -17520 -7833 -17508
rect -2112 -17296 -2100 -17106
rect -2066 -17296 -2050 -17106
rect -2112 -17308 -2050 -17296
rect -2020 -17102 -1954 -17094
rect -2020 -17296 -2004 -17102
rect -1970 -17296 -1954 -17102
rect -2020 -17308 -1954 -17296
rect -1924 -17106 -1858 -17094
rect -1924 -17296 -1908 -17106
rect -1874 -17296 -1858 -17106
rect -1924 -17308 -1858 -17296
rect -1828 -17102 -1766 -17094
rect -1828 -17296 -1812 -17102
rect -1778 -17296 -1766 -17102
rect -1828 -17308 -1766 -17296
rect -4828 -17491 -4766 -17479
rect -4828 -17681 -4816 -17491
rect -4782 -17681 -4766 -17491
rect -4828 -17693 -4766 -17681
rect -4736 -17491 -4670 -17479
rect -4736 -17685 -4720 -17491
rect -4686 -17685 -4670 -17491
rect -4736 -17693 -4670 -17685
rect -4640 -17491 -4574 -17479
rect -4640 -17681 -4624 -17491
rect -4590 -17681 -4574 -17491
rect -4640 -17693 -4574 -17681
rect -4544 -17491 -4482 -17479
rect -4544 -17685 -4528 -17491
rect -4494 -17685 -4482 -17491
rect -2112 -17485 -2050 -17473
rect -4544 -17693 -4482 -17685
rect -2112 -17675 -2100 -17485
rect -2066 -17675 -2050 -17485
rect -2112 -17687 -2050 -17675
rect -2020 -17481 -1954 -17473
rect -2020 -17675 -2004 -17481
rect -1970 -17675 -1954 -17481
rect -2020 -17687 -1954 -17675
rect -1924 -17485 -1858 -17473
rect -1924 -17675 -1908 -17485
rect -1874 -17675 -1858 -17485
rect -1924 -17687 -1858 -17675
rect -1828 -17481 -1766 -17473
rect -1828 -17675 -1812 -17481
rect -1778 -17675 -1766 -17481
rect -1828 -17687 -1766 -17675
rect -8179 -17778 -8117 -17766
rect -8179 -17968 -8167 -17778
rect -8133 -17968 -8117 -17778
rect -8179 -17980 -8117 -17968
rect -8087 -17774 -8021 -17766
rect -8087 -17968 -8071 -17774
rect -8037 -17968 -8021 -17774
rect -8087 -17980 -8021 -17968
rect -7991 -17778 -7925 -17766
rect -7991 -17968 -7975 -17778
rect -7941 -17968 -7925 -17778
rect -7991 -17980 -7925 -17968
rect -7895 -17774 -7833 -17766
rect -7895 -17968 -7879 -17774
rect -7845 -17968 -7833 -17774
rect -7895 -17980 -7833 -17968
rect 12923 -16253 12935 -16219
rect 13125 -16253 13137 -16219
rect 12923 -16269 13137 -16253
rect 12923 -16315 13137 -16299
rect 12923 -16349 12935 -16315
rect 13129 -16349 13137 -16315
rect 12923 -16365 13137 -16349
rect 12923 -16411 13137 -16395
rect 12923 -16445 12935 -16411
rect 13125 -16445 13137 -16411
rect 12923 -16461 13137 -16445
rect 12923 -16507 13137 -16491
rect 12923 -16541 12935 -16507
rect 13129 -16541 13137 -16507
rect 12923 -16553 13137 -16541
rect 7138 -17769 7200 -17757
rect -4828 -17931 -4766 -17919
rect -4828 -18121 -4816 -17931
rect -4782 -18121 -4766 -17931
rect -4828 -18133 -4766 -18121
rect -4736 -17931 -4670 -17919
rect -4736 -18125 -4720 -17931
rect -4686 -18125 -4670 -17931
rect -4736 -18133 -4670 -18125
rect -4640 -17931 -4574 -17919
rect -4640 -18121 -4624 -17931
rect -4590 -18121 -4574 -17931
rect -4640 -18133 -4574 -18121
rect -4544 -17931 -4482 -17919
rect -4544 -18125 -4528 -17931
rect -4494 -18125 -4482 -17931
rect -2112 -17925 -2050 -17913
rect -4544 -18133 -4482 -18125
rect -2112 -18115 -2100 -17925
rect -2066 -18115 -2050 -17925
rect -2112 -18127 -2050 -18115
rect -2020 -17921 -1954 -17913
rect -2020 -18115 -2004 -17921
rect -1970 -18115 -1954 -17921
rect -2020 -18127 -1954 -18115
rect -1924 -17925 -1858 -17913
rect -1924 -18115 -1908 -17925
rect -1874 -18115 -1858 -17925
rect -1924 -18127 -1858 -18115
rect -1828 -17921 -1766 -17913
rect -1828 -18115 -1812 -17921
rect -1778 -18115 -1766 -17921
rect -1828 -18127 -1766 -18115
rect 7138 -18067 7150 -17769
rect 7184 -18067 7200 -17769
rect 7138 -18079 7200 -18067
rect 7230 -17769 7296 -17757
rect 7230 -18067 7246 -17769
rect 7280 -18067 7296 -17769
rect 7230 -18079 7296 -18067
rect 7326 -17769 7392 -17757
rect 7326 -18067 7342 -17769
rect 7376 -18067 7392 -17769
rect 7326 -18079 7392 -18067
rect 7422 -17769 7488 -17757
rect 7422 -18067 7438 -17769
rect 7472 -18067 7488 -17769
rect 7422 -18079 7488 -18067
rect 7518 -17769 7584 -17757
rect 7518 -18067 7534 -17769
rect 7568 -18067 7584 -17769
rect 7518 -18079 7584 -18067
rect 7614 -17769 7680 -17757
rect 7614 -18067 7630 -17769
rect 7664 -18067 7680 -17769
rect 7614 -18079 7680 -18067
rect 7710 -17769 7776 -17757
rect 7710 -18067 7726 -17769
rect 7760 -18067 7776 -17769
rect 7710 -18079 7776 -18067
rect 7806 -17769 7872 -17757
rect 7806 -18067 7822 -17769
rect 7856 -18067 7872 -17769
rect 7806 -18079 7872 -18067
rect 7902 -17769 7964 -17757
rect 7902 -18067 7918 -17769
rect 7952 -18067 7964 -17769
rect 7902 -18079 7964 -18067
rect 8086 -17769 8148 -17757
rect 8086 -18067 8098 -17769
rect 8132 -18067 8148 -17769
rect 8086 -18079 8148 -18067
rect 8178 -17769 8244 -17757
rect 8178 -18067 8194 -17769
rect 8228 -18067 8244 -17769
rect 8178 -18079 8244 -18067
rect 8274 -17769 8340 -17757
rect 8274 -18067 8290 -17769
rect 8324 -18067 8340 -17769
rect 8274 -18079 8340 -18067
rect 8370 -17769 8436 -17757
rect 8370 -18067 8386 -17769
rect 8420 -18067 8436 -17769
rect 8370 -18079 8436 -18067
rect 8466 -17769 8532 -17757
rect 8466 -18067 8482 -17769
rect 8516 -18067 8532 -17769
rect 8466 -18079 8532 -18067
rect 8562 -17769 8628 -17757
rect 8562 -18067 8578 -17769
rect 8612 -18067 8628 -17769
rect 8562 -18079 8628 -18067
rect 8658 -17769 8724 -17757
rect 8658 -18067 8674 -17769
rect 8708 -18067 8724 -17769
rect 8658 -18079 8724 -18067
rect 8754 -17769 8820 -17757
rect 8754 -18067 8770 -17769
rect 8804 -18067 8820 -17769
rect 8754 -18079 8820 -18067
rect 8850 -17769 8912 -17757
rect 8850 -18067 8866 -17769
rect 8900 -18067 8912 -17769
rect 8850 -18079 8912 -18067
rect 9022 -17769 9084 -17757
rect 9022 -18067 9034 -17769
rect 9068 -18067 9084 -17769
rect 9022 -18079 9084 -18067
rect 9114 -17769 9180 -17757
rect 9114 -18067 9130 -17769
rect 9164 -18067 9180 -17769
rect 9114 -18079 9180 -18067
rect 9210 -17769 9276 -17757
rect 9210 -18067 9226 -17769
rect 9260 -18067 9276 -17769
rect 9210 -18079 9276 -18067
rect 9306 -17769 9372 -17757
rect 9306 -18067 9322 -17769
rect 9356 -18067 9372 -17769
rect 9306 -18079 9372 -18067
rect 9402 -17769 9468 -17757
rect 9402 -18067 9418 -17769
rect 9452 -18067 9468 -17769
rect 9402 -18079 9468 -18067
rect 9498 -17769 9564 -17757
rect 9498 -18067 9514 -17769
rect 9548 -18067 9564 -17769
rect 9498 -18079 9564 -18067
rect 9594 -17769 9660 -17757
rect 9594 -18067 9610 -17769
rect 9644 -18067 9660 -17769
rect 9594 -18079 9660 -18067
rect 9690 -17769 9756 -17757
rect 9690 -18067 9706 -17769
rect 9740 -18067 9756 -17769
rect 9690 -18079 9756 -18067
rect 9786 -17769 9848 -17757
rect 9786 -18067 9802 -17769
rect 9836 -18067 9848 -17769
rect 9786 -18079 9848 -18067
rect 9953 -17768 10015 -17756
rect 9953 -18066 9965 -17768
rect 9999 -18066 10015 -17768
rect 9953 -18078 10015 -18066
rect 10045 -17768 10111 -17756
rect 10045 -18066 10061 -17768
rect 10095 -18066 10111 -17768
rect 10045 -18078 10111 -18066
rect 10141 -17768 10207 -17756
rect 10141 -18066 10157 -17768
rect 10191 -18066 10207 -17768
rect 10141 -18078 10207 -18066
rect 10237 -17768 10303 -17756
rect 10237 -18066 10253 -17768
rect 10287 -18066 10303 -17768
rect 10237 -18078 10303 -18066
rect 10333 -17768 10399 -17756
rect 10333 -18066 10349 -17768
rect 10383 -18066 10399 -17768
rect 10333 -18078 10399 -18066
rect 10429 -17768 10495 -17756
rect 10429 -18066 10445 -17768
rect 10479 -18066 10495 -17768
rect 10429 -18078 10495 -18066
rect 10525 -17768 10591 -17756
rect 10525 -18066 10541 -17768
rect 10575 -18066 10591 -17768
rect 10525 -18078 10591 -18066
rect 10621 -17768 10687 -17756
rect 10621 -18066 10637 -17768
rect 10671 -18066 10687 -17768
rect 10621 -18078 10687 -18066
rect 10717 -17768 10779 -17756
rect 15763 -17679 15825 -17667
rect 10717 -18066 10733 -17768
rect 10767 -18066 10779 -17768
rect 10717 -18078 10779 -18066
rect 10880 -17769 10942 -17757
rect 10880 -18067 10892 -17769
rect 10926 -18067 10942 -17769
rect 10880 -18079 10942 -18067
rect 10972 -17769 11038 -17757
rect 10972 -18067 10988 -17769
rect 11022 -18067 11038 -17769
rect 10972 -18079 11038 -18067
rect 11068 -17769 11134 -17757
rect 11068 -18067 11084 -17769
rect 11118 -18067 11134 -17769
rect 11068 -18079 11134 -18067
rect 11164 -17769 11230 -17757
rect 11164 -18067 11180 -17769
rect 11214 -18067 11230 -17769
rect 11164 -18079 11230 -18067
rect 11260 -17769 11326 -17757
rect 11260 -18067 11276 -17769
rect 11310 -18067 11326 -17769
rect 11260 -18079 11326 -18067
rect 11356 -17769 11422 -17757
rect 11356 -18067 11372 -17769
rect 11406 -18067 11422 -17769
rect 11356 -18079 11422 -18067
rect 11452 -17769 11518 -17757
rect 11452 -18067 11468 -17769
rect 11502 -18067 11518 -17769
rect 11452 -18079 11518 -18067
rect 11548 -17769 11614 -17757
rect 11548 -18067 11564 -17769
rect 11598 -18067 11614 -17769
rect 11548 -18079 11614 -18067
rect 11644 -17769 11706 -17757
rect 11644 -18067 11660 -17769
rect 11694 -18067 11706 -17769
rect 11644 -18079 11706 -18067
rect -12314 -18249 -11764 -18237
rect -17677 -18271 -17421 -18255
rect -17677 -18305 -17665 -18271
rect -17433 -18305 -17421 -18271
rect -12314 -18283 -12302 -18249
rect -11776 -18283 -11764 -18249
rect -12314 -18295 -11764 -18283
rect -17677 -18317 -17421 -18305
rect -8193 -18238 -8131 -18226
rect -24428 -18445 -24214 -18433
rect -24428 -18479 -24416 -18445
rect -24226 -18479 -24214 -18445
rect -24428 -18495 -24214 -18479
rect -24428 -18541 -24214 -18525
rect -24428 -18575 -24416 -18541
rect -24226 -18575 -24214 -18541
rect -24428 -18591 -24214 -18575
rect -24428 -18637 -24214 -18621
rect -24428 -18671 -24416 -18637
rect -24226 -18671 -24214 -18637
rect -24428 -18687 -24214 -18671
rect -24428 -18733 -24214 -18717
rect -24428 -18767 -24416 -18733
rect -24226 -18767 -24214 -18733
rect -24428 -18783 -24214 -18767
rect -24428 -18829 -24214 -18813
rect -24428 -18863 -24416 -18829
rect -24226 -18863 -24214 -18829
rect -24428 -18879 -24214 -18863
rect -16026 -18417 -15964 -18405
rect -21617 -18546 -21555 -18534
rect -21617 -18736 -21605 -18546
rect -21571 -18736 -21555 -18546
rect -21617 -18748 -21555 -18736
rect -21525 -18542 -21459 -18534
rect -21525 -18736 -21509 -18542
rect -21475 -18736 -21459 -18542
rect -21525 -18748 -21459 -18736
rect -21429 -18546 -21363 -18534
rect -21429 -18736 -21413 -18546
rect -21379 -18736 -21363 -18546
rect -21429 -18748 -21363 -18736
rect -21333 -18542 -21271 -18534
rect -21333 -18736 -21317 -18542
rect -21283 -18736 -21271 -18542
rect -21333 -18748 -21271 -18736
rect -16026 -18607 -16014 -18417
rect -15980 -18607 -15964 -18417
rect -16026 -18619 -15964 -18607
rect -15934 -18413 -15868 -18405
rect -15934 -18607 -15918 -18413
rect -15884 -18607 -15868 -18413
rect -15934 -18619 -15868 -18607
rect -15838 -18417 -15772 -18405
rect -15838 -18607 -15822 -18417
rect -15788 -18607 -15772 -18417
rect -15838 -18619 -15772 -18607
rect -15742 -18413 -15680 -18405
rect -15742 -18607 -15726 -18413
rect -15692 -18607 -15680 -18413
rect -15742 -18619 -15680 -18607
rect -8193 -18428 -8181 -18238
rect -8147 -18428 -8131 -18238
rect -8193 -18440 -8131 -18428
rect -8101 -18234 -8035 -18226
rect -8101 -18428 -8085 -18234
rect -8051 -18428 -8035 -18234
rect -8101 -18440 -8035 -18428
rect -8005 -18238 -7939 -18226
rect -8005 -18428 -7989 -18238
rect -7955 -18428 -7939 -18238
rect -8005 -18440 -7939 -18428
rect -7909 -18234 -7847 -18226
rect -7909 -18428 -7893 -18234
rect -7859 -18428 -7847 -18234
rect -7909 -18440 -7847 -18428
rect -4828 -18310 -4766 -18298
rect -4828 -18500 -4816 -18310
rect -4782 -18500 -4766 -18310
rect -4828 -18512 -4766 -18500
rect -4736 -18310 -4670 -18298
rect -4736 -18504 -4720 -18310
rect -4686 -18504 -4670 -18310
rect -4736 -18512 -4670 -18504
rect -4640 -18310 -4574 -18298
rect -4640 -18500 -4624 -18310
rect -4590 -18500 -4574 -18310
rect -4640 -18512 -4574 -18500
rect -4544 -18310 -4482 -18298
rect -4544 -18504 -4528 -18310
rect -4494 -18504 -4482 -18310
rect -2112 -18304 -2050 -18292
rect -4544 -18512 -4482 -18504
rect -2112 -18494 -2100 -18304
rect -2066 -18494 -2050 -18304
rect -2112 -18506 -2050 -18494
rect -2020 -18300 -1954 -18292
rect -2020 -18494 -2004 -18300
rect -1970 -18494 -1954 -18300
rect -2020 -18506 -1954 -18494
rect -1924 -18304 -1858 -18292
rect -1924 -18494 -1908 -18304
rect -1874 -18494 -1858 -18304
rect -1924 -18506 -1858 -18494
rect -1828 -18300 -1766 -18292
rect -1828 -18494 -1812 -18300
rect -1778 -18494 -1766 -18300
rect -1828 -18506 -1766 -18494
rect 15763 -18511 15775 -17679
rect 15809 -18511 15825 -17679
rect 15763 -18523 15825 -18511
rect 15855 -17679 15921 -17667
rect 15855 -18511 15871 -17679
rect 15905 -18511 15921 -17679
rect 15855 -18523 15921 -18511
rect 15951 -17679 16017 -17667
rect 15951 -18511 15967 -17679
rect 16001 -18511 16017 -17679
rect 15951 -18523 16017 -18511
rect 16047 -17679 16113 -17667
rect 16047 -18511 16063 -17679
rect 16097 -18511 16113 -17679
rect 16047 -18523 16113 -18511
rect 16143 -17679 16209 -17667
rect 16143 -18511 16159 -17679
rect 16193 -18511 16209 -17679
rect 16143 -18523 16209 -18511
rect 16239 -17679 16305 -17667
rect 16239 -18511 16255 -17679
rect 16289 -18511 16305 -17679
rect 16239 -18523 16305 -18511
rect 16335 -17679 16401 -17667
rect 16335 -18511 16351 -17679
rect 16385 -18511 16401 -17679
rect 16335 -18523 16401 -18511
rect 16431 -17679 16497 -17667
rect 16431 -18511 16447 -17679
rect 16481 -18511 16497 -17679
rect 16431 -18523 16497 -18511
rect 16527 -17679 16593 -17667
rect 16527 -18511 16543 -17679
rect 16577 -18511 16593 -17679
rect 16527 -18523 16593 -18511
rect 16623 -17679 16689 -17667
rect 16623 -18511 16639 -17679
rect 16673 -18511 16689 -17679
rect 16623 -18523 16689 -18511
rect 16719 -17679 16785 -17667
rect 16719 -18511 16735 -17679
rect 16769 -18511 16785 -17679
rect 16719 -18523 16785 -18511
rect 16815 -17679 16881 -17667
rect 16815 -18511 16831 -17679
rect 16865 -18511 16881 -17679
rect 16815 -18523 16881 -18511
rect 16911 -17679 16973 -17667
rect 16911 -18511 16927 -17679
rect 16961 -18511 16973 -17679
rect 18096 -18259 18310 -18247
rect 17294 -18287 17356 -18275
rect 17294 -18477 17306 -18287
rect 17340 -18477 17356 -18287
rect 17294 -18489 17356 -18477
rect 17386 -18287 17452 -18275
rect 17386 -18477 17402 -18287
rect 17436 -18477 17452 -18287
rect 17386 -18489 17452 -18477
rect 17482 -18287 17548 -18275
rect 17482 -18477 17498 -18287
rect 17532 -18477 17548 -18287
rect 17482 -18489 17548 -18477
rect 17578 -18287 17644 -18275
rect 17578 -18477 17594 -18287
rect 17628 -18477 17644 -18287
rect 17578 -18489 17644 -18477
rect 17674 -18287 17740 -18275
rect 17674 -18477 17690 -18287
rect 17724 -18477 17740 -18287
rect 17674 -18489 17740 -18477
rect 17770 -18287 17836 -18275
rect 17770 -18477 17786 -18287
rect 17820 -18477 17836 -18287
rect 17770 -18489 17836 -18477
rect 17866 -18287 17928 -18275
rect 17866 -18477 17882 -18287
rect 17916 -18477 17928 -18287
rect 17866 -18489 17928 -18477
rect 16911 -18523 16973 -18511
rect -17677 -18711 -17421 -18699
rect -17677 -18745 -17665 -18711
rect -17433 -18745 -17421 -18711
rect -17677 -18761 -17421 -18745
rect -24428 -18925 -24214 -18909
rect -24428 -18959 -24416 -18925
rect -24226 -18959 -24214 -18925
rect -24428 -18975 -24214 -18959
rect -17677 -18807 -17421 -18791
rect -17677 -18841 -17665 -18807
rect -17433 -18841 -17421 -18807
rect -17677 -18857 -17421 -18841
rect -8191 -18718 -8129 -18706
rect -17677 -18903 -17421 -18887
rect -17677 -18937 -17665 -18903
rect -17433 -18937 -17421 -18903
rect -17677 -18953 -17421 -18937
rect -24428 -19021 -24214 -19005
rect -17677 -18999 -17421 -18983
rect -24428 -19055 -24416 -19021
rect -24226 -19055 -24214 -19021
rect -24428 -19067 -24214 -19055
rect -21618 -19026 -21556 -19014
rect -21618 -19216 -21606 -19026
rect -21572 -19216 -21556 -19026
rect -21618 -19228 -21556 -19216
rect -21526 -19022 -21460 -19014
rect -21526 -19216 -21510 -19022
rect -21476 -19216 -21460 -19022
rect -21526 -19228 -21460 -19216
rect -21430 -19026 -21364 -19014
rect -21430 -19216 -21414 -19026
rect -21380 -19216 -21364 -19026
rect -21430 -19228 -21364 -19216
rect -21334 -19022 -21272 -19014
rect -21334 -19216 -21318 -19022
rect -21284 -19216 -21272 -19022
rect -21334 -19228 -21272 -19216
rect -17677 -19033 -17665 -18999
rect -17433 -19033 -17421 -18999
rect -17677 -19049 -17421 -19033
rect -17677 -19095 -17421 -19079
rect -17677 -19129 -17665 -19095
rect -17433 -19129 -17421 -19095
rect -17677 -19145 -17421 -19129
rect -16027 -18897 -15965 -18885
rect -17677 -19191 -17421 -19175
rect -17677 -19225 -17665 -19191
rect -17433 -19225 -17421 -19191
rect -16027 -19087 -16015 -18897
rect -15981 -19087 -15965 -18897
rect -16027 -19099 -15965 -19087
rect -15935 -18893 -15869 -18885
rect -15935 -19087 -15919 -18893
rect -15885 -19087 -15869 -18893
rect -15935 -19099 -15869 -19087
rect -15839 -18897 -15773 -18885
rect -15839 -19087 -15823 -18897
rect -15789 -19087 -15773 -18897
rect -15839 -19099 -15773 -19087
rect -15743 -18893 -15681 -18885
rect -15743 -19087 -15727 -18893
rect -15693 -19087 -15681 -18893
rect -15743 -19099 -15681 -19087
rect -8191 -18908 -8179 -18718
rect -8145 -18908 -8129 -18718
rect -8191 -18920 -8129 -18908
rect -8099 -18714 -8033 -18706
rect -8099 -18908 -8083 -18714
rect -8049 -18908 -8033 -18714
rect -8099 -18920 -8033 -18908
rect -8003 -18718 -7937 -18706
rect -8003 -18908 -7987 -18718
rect -7953 -18908 -7937 -18718
rect -8003 -18920 -7937 -18908
rect -7907 -18714 -7845 -18706
rect -7907 -18908 -7891 -18714
rect -7857 -18908 -7845 -18714
rect 18096 -18293 18108 -18259
rect 18298 -18293 18310 -18259
rect 18096 -18309 18310 -18293
rect 18096 -18355 18310 -18339
rect 18096 -18389 18108 -18355
rect 18302 -18389 18310 -18355
rect 18096 -18405 18310 -18389
rect 18096 -18451 18310 -18435
rect 18096 -18485 18108 -18451
rect 18298 -18485 18310 -18451
rect 18096 -18501 18310 -18485
rect 18096 -18547 18310 -18531
rect 18096 -18581 18108 -18547
rect 18302 -18581 18310 -18547
rect -7907 -18920 -7845 -18908
rect -4828 -18750 -4766 -18738
rect -4828 -18940 -4816 -18750
rect -4782 -18940 -4766 -18750
rect -4828 -18952 -4766 -18940
rect -4736 -18750 -4670 -18738
rect -4736 -18944 -4720 -18750
rect -4686 -18944 -4670 -18750
rect -4736 -18952 -4670 -18944
rect -4640 -18750 -4574 -18738
rect -4640 -18940 -4624 -18750
rect -4590 -18940 -4574 -18750
rect -4640 -18952 -4574 -18940
rect -4544 -18750 -4482 -18738
rect -4544 -18944 -4528 -18750
rect -4494 -18944 -4482 -18750
rect -2112 -18744 -2050 -18732
rect -4544 -18952 -4482 -18944
rect -2112 -18934 -2100 -18744
rect -2066 -18934 -2050 -18744
rect -2112 -18946 -2050 -18934
rect -2020 -18740 -1954 -18732
rect -2020 -18934 -2004 -18740
rect -1970 -18934 -1954 -18740
rect -2020 -18946 -1954 -18934
rect -1924 -18744 -1858 -18732
rect -1924 -18934 -1908 -18744
rect -1874 -18934 -1858 -18744
rect -1924 -18946 -1858 -18934
rect -1828 -18740 -1766 -18732
rect -1828 -18934 -1812 -18740
rect -1778 -18934 -1766 -18740
rect 5658 -18729 5872 -18717
rect -1828 -18946 -1766 -18934
rect 5658 -18763 5670 -18729
rect 5860 -18763 5872 -18729
rect 6098 -18729 6312 -18717
rect 5658 -18779 5872 -18763
rect 5658 -18825 5872 -18809
rect 5658 -18859 5670 -18825
rect 5864 -18859 5872 -18825
rect 5658 -18875 5872 -18859
rect 5658 -18921 5872 -18905
rect 5658 -18955 5670 -18921
rect 5860 -18955 5872 -18921
rect 5658 -18971 5872 -18955
rect 5658 -19017 5872 -19001
rect 5658 -19051 5670 -19017
rect 5864 -19051 5872 -19017
rect 6098 -18763 6110 -18729
rect 6300 -18763 6312 -18729
rect 6538 -18729 6752 -18717
rect 6098 -18779 6312 -18763
rect 6098 -18825 6312 -18809
rect 6098 -18859 6110 -18825
rect 6304 -18859 6312 -18825
rect 6098 -18875 6312 -18859
rect 6098 -18921 6312 -18905
rect 6098 -18955 6110 -18921
rect 6300 -18955 6312 -18921
rect 6098 -18971 6312 -18955
rect 6098 -19017 6312 -19001
rect 5658 -19063 5872 -19051
rect 6098 -19051 6110 -19017
rect 6304 -19051 6312 -19017
rect 6538 -18763 6550 -18729
rect 6740 -18763 6752 -18729
rect 6538 -18779 6752 -18763
rect 6538 -18825 6752 -18809
rect 6538 -18859 6550 -18825
rect 6744 -18859 6752 -18825
rect 6538 -18875 6752 -18859
rect 6538 -18921 6752 -18905
rect 6538 -18955 6550 -18921
rect 6740 -18955 6752 -18921
rect 6538 -18971 6752 -18955
rect 6538 -19017 6752 -19001
rect 6098 -19063 6312 -19051
rect 6538 -19051 6550 -19017
rect 6744 -19051 6752 -19017
rect 6538 -19063 6752 -19051
rect -17677 -19241 -17421 -19225
rect -17677 -19287 -17421 -19271
rect -21618 -19526 -21556 -19514
rect -24426 -19639 -24212 -19627
rect -24426 -19673 -24414 -19639
rect -24224 -19673 -24212 -19639
rect -24426 -19689 -24212 -19673
rect -24426 -19735 -24212 -19719
rect -24426 -19769 -24414 -19735
rect -24224 -19769 -24212 -19735
rect -24426 -19785 -24212 -19769
rect -24426 -19831 -24212 -19815
rect -24426 -19865 -24414 -19831
rect -24224 -19865 -24212 -19831
rect -24426 -19881 -24212 -19865
rect -24426 -19927 -24212 -19911
rect -24426 -19961 -24414 -19927
rect -24224 -19961 -24212 -19927
rect -24426 -19977 -24212 -19961
rect -24426 -20023 -24212 -20007
rect -24426 -20057 -24414 -20023
rect -24224 -20057 -24212 -20023
rect -24426 -20073 -24212 -20057
rect -21618 -19716 -21606 -19526
rect -21572 -19716 -21556 -19526
rect -21618 -19728 -21556 -19716
rect -21526 -19522 -21460 -19514
rect -21526 -19716 -21510 -19522
rect -21476 -19716 -21460 -19522
rect -21526 -19728 -21460 -19716
rect -21430 -19526 -21364 -19514
rect -21430 -19716 -21414 -19526
rect -21380 -19716 -21364 -19526
rect -21430 -19728 -21364 -19716
rect -21334 -19522 -21272 -19514
rect -21334 -19716 -21318 -19522
rect -21284 -19716 -21272 -19522
rect -21334 -19728 -21272 -19716
rect -17677 -19321 -17665 -19287
rect -17433 -19321 -17421 -19287
rect -17677 -19337 -17421 -19321
rect -4828 -19129 -4766 -19117
rect -4828 -19319 -4816 -19129
rect -4782 -19319 -4766 -19129
rect -4828 -19331 -4766 -19319
rect -4736 -19129 -4670 -19117
rect -4736 -19323 -4720 -19129
rect -4686 -19323 -4670 -19129
rect -4736 -19331 -4670 -19323
rect -4640 -19129 -4574 -19117
rect -4640 -19319 -4624 -19129
rect -4590 -19319 -4574 -19129
rect -4640 -19331 -4574 -19319
rect -4544 -19129 -4482 -19117
rect -4544 -19323 -4528 -19129
rect -4494 -19323 -4482 -19129
rect -2112 -19123 -2050 -19111
rect -4544 -19331 -4482 -19323
rect -2112 -19313 -2100 -19123
rect -2066 -19313 -2050 -19123
rect -2112 -19325 -2050 -19313
rect -2020 -19119 -1954 -19111
rect -2020 -19313 -2004 -19119
rect -1970 -19313 -1954 -19119
rect -2020 -19325 -1954 -19313
rect -1924 -19123 -1858 -19111
rect -1924 -19313 -1908 -19123
rect -1874 -19313 -1858 -19123
rect -1924 -19325 -1858 -19313
rect -1828 -19119 -1766 -19111
rect -1828 -19313 -1812 -19119
rect -1778 -19313 -1766 -19119
rect -1828 -19325 -1766 -19313
rect 15763 -18661 15825 -18649
rect -17677 -19383 -17421 -19367
rect -17677 -19417 -17665 -19383
rect -17433 -19417 -17421 -19383
rect -17677 -19433 -17421 -19417
rect -17677 -19479 -17421 -19463
rect -17677 -19513 -17665 -19479
rect -17433 -19513 -17421 -19479
rect -17677 -19529 -17421 -19513
rect -17677 -19575 -17421 -19559
rect -17677 -19609 -17665 -19575
rect -17433 -19609 -17421 -19575
rect -17677 -19625 -17421 -19609
rect -16027 -19397 -15965 -19385
rect -16027 -19587 -16015 -19397
rect -15981 -19587 -15965 -19397
rect -16027 -19599 -15965 -19587
rect -15935 -19393 -15869 -19385
rect -15935 -19587 -15919 -19393
rect -15885 -19587 -15869 -19393
rect -15935 -19599 -15869 -19587
rect -15839 -19397 -15773 -19385
rect -15839 -19587 -15823 -19397
rect -15789 -19587 -15773 -19397
rect -15839 -19599 -15773 -19587
rect -15743 -19393 -15681 -19385
rect -15743 -19587 -15727 -19393
rect -15693 -19587 -15681 -19393
rect -15743 -19599 -15681 -19587
rect 7138 -19433 7200 -19421
rect -4828 -19569 -4766 -19557
rect -17677 -19671 -17421 -19655
rect -17677 -19705 -17665 -19671
rect -17433 -19705 -17421 -19671
rect -17677 -19717 -17421 -19705
rect -4828 -19759 -4816 -19569
rect -4782 -19759 -4766 -19569
rect -4828 -19771 -4766 -19759
rect -4736 -19569 -4670 -19557
rect -4736 -19763 -4720 -19569
rect -4686 -19763 -4670 -19569
rect -4736 -19771 -4670 -19763
rect -4640 -19569 -4574 -19557
rect -4640 -19759 -4624 -19569
rect -4590 -19759 -4574 -19569
rect -4640 -19771 -4574 -19759
rect -4544 -19569 -4482 -19557
rect -4544 -19763 -4528 -19569
rect -4494 -19763 -4482 -19569
rect -2112 -19563 -2050 -19551
rect -4544 -19771 -4482 -19763
rect -2112 -19753 -2100 -19563
rect -2066 -19753 -2050 -19563
rect -2112 -19765 -2050 -19753
rect -2020 -19559 -1954 -19551
rect -2020 -19753 -2004 -19559
rect -1970 -19753 -1954 -19559
rect -2020 -19765 -1954 -19753
rect -1924 -19563 -1858 -19551
rect -1924 -19753 -1908 -19563
rect -1874 -19753 -1858 -19563
rect -1924 -19765 -1858 -19753
rect -1828 -19559 -1766 -19551
rect -1828 -19753 -1812 -19559
rect -1778 -19753 -1766 -19559
rect -1828 -19765 -1766 -19753
rect 7138 -19731 7150 -19433
rect 7184 -19731 7200 -19433
rect 7138 -19743 7200 -19731
rect 7230 -19433 7296 -19421
rect 7230 -19731 7246 -19433
rect 7280 -19731 7296 -19433
rect 7230 -19743 7296 -19731
rect 7326 -19433 7392 -19421
rect 7326 -19731 7342 -19433
rect 7376 -19731 7392 -19433
rect 7326 -19743 7392 -19731
rect 7422 -19433 7488 -19421
rect 7422 -19731 7438 -19433
rect 7472 -19731 7488 -19433
rect 7422 -19743 7488 -19731
rect 7518 -19433 7584 -19421
rect 7518 -19731 7534 -19433
rect 7568 -19731 7584 -19433
rect 7518 -19743 7584 -19731
rect 7614 -19433 7680 -19421
rect 7614 -19731 7630 -19433
rect 7664 -19731 7680 -19433
rect 7614 -19743 7680 -19731
rect 7710 -19433 7776 -19421
rect 7710 -19731 7726 -19433
rect 7760 -19731 7776 -19433
rect 7710 -19743 7776 -19731
rect 7806 -19433 7872 -19421
rect 7806 -19731 7822 -19433
rect 7856 -19731 7872 -19433
rect 7806 -19743 7872 -19731
rect 7902 -19433 7964 -19421
rect 7902 -19731 7918 -19433
rect 7952 -19731 7964 -19433
rect 7902 -19743 7964 -19731
rect 8086 -19433 8148 -19421
rect 8086 -19731 8098 -19433
rect 8132 -19731 8148 -19433
rect 8086 -19743 8148 -19731
rect 8178 -19433 8244 -19421
rect 8178 -19731 8194 -19433
rect 8228 -19731 8244 -19433
rect 8178 -19743 8244 -19731
rect 8274 -19433 8340 -19421
rect 8274 -19731 8290 -19433
rect 8324 -19731 8340 -19433
rect 8274 -19743 8340 -19731
rect 8370 -19433 8436 -19421
rect 8370 -19731 8386 -19433
rect 8420 -19731 8436 -19433
rect 8370 -19743 8436 -19731
rect 8466 -19433 8532 -19421
rect 8466 -19731 8482 -19433
rect 8516 -19731 8532 -19433
rect 8466 -19743 8532 -19731
rect 8562 -19433 8628 -19421
rect 8562 -19731 8578 -19433
rect 8612 -19731 8628 -19433
rect 8562 -19743 8628 -19731
rect 8658 -19433 8724 -19421
rect 8658 -19731 8674 -19433
rect 8708 -19731 8724 -19433
rect 8658 -19743 8724 -19731
rect 8754 -19433 8820 -19421
rect 8754 -19731 8770 -19433
rect 8804 -19731 8820 -19433
rect 8754 -19743 8820 -19731
rect 8850 -19433 8912 -19421
rect 8850 -19731 8866 -19433
rect 8900 -19731 8912 -19433
rect 8850 -19743 8912 -19731
rect 9022 -19433 9084 -19421
rect 9022 -19731 9034 -19433
rect 9068 -19731 9084 -19433
rect 9022 -19743 9084 -19731
rect 9114 -19433 9180 -19421
rect 9114 -19731 9130 -19433
rect 9164 -19731 9180 -19433
rect 9114 -19743 9180 -19731
rect 9210 -19433 9276 -19421
rect 9210 -19731 9226 -19433
rect 9260 -19731 9276 -19433
rect 9210 -19743 9276 -19731
rect 9306 -19433 9372 -19421
rect 9306 -19731 9322 -19433
rect 9356 -19731 9372 -19433
rect 9306 -19743 9372 -19731
rect 9402 -19433 9468 -19421
rect 9402 -19731 9418 -19433
rect 9452 -19731 9468 -19433
rect 9402 -19743 9468 -19731
rect 9498 -19433 9564 -19421
rect 9498 -19731 9514 -19433
rect 9548 -19731 9564 -19433
rect 9498 -19743 9564 -19731
rect 9594 -19433 9660 -19421
rect 9594 -19731 9610 -19433
rect 9644 -19731 9660 -19433
rect 9594 -19743 9660 -19731
rect 9690 -19433 9756 -19421
rect 9690 -19731 9706 -19433
rect 9740 -19731 9756 -19433
rect 9690 -19743 9756 -19731
rect 9786 -19433 9848 -19421
rect 9786 -19731 9802 -19433
rect 9836 -19731 9848 -19433
rect 9786 -19743 9848 -19731
rect 9953 -19433 10015 -19421
rect 9953 -19731 9965 -19433
rect 9999 -19731 10015 -19433
rect 9953 -19743 10015 -19731
rect 10045 -19433 10111 -19421
rect 10045 -19731 10061 -19433
rect 10095 -19731 10111 -19433
rect 10045 -19743 10111 -19731
rect 10141 -19433 10207 -19421
rect 10141 -19731 10157 -19433
rect 10191 -19731 10207 -19433
rect 10141 -19743 10207 -19731
rect 10237 -19433 10303 -19421
rect 10237 -19731 10253 -19433
rect 10287 -19731 10303 -19433
rect 10237 -19743 10303 -19731
rect 10333 -19433 10399 -19421
rect 10333 -19731 10349 -19433
rect 10383 -19731 10399 -19433
rect 10333 -19743 10399 -19731
rect 10429 -19433 10495 -19421
rect 10429 -19731 10445 -19433
rect 10479 -19731 10495 -19433
rect 10429 -19743 10495 -19731
rect 10525 -19433 10591 -19421
rect 10525 -19731 10541 -19433
rect 10575 -19731 10591 -19433
rect 10525 -19743 10591 -19731
rect 10621 -19433 10687 -19421
rect 10621 -19731 10637 -19433
rect 10671 -19731 10687 -19433
rect 10621 -19743 10687 -19731
rect 10717 -19433 10779 -19421
rect 10717 -19731 10733 -19433
rect 10767 -19731 10779 -19433
rect 10717 -19743 10779 -19731
rect 10880 -19433 10942 -19421
rect 10880 -19731 10892 -19433
rect 10926 -19731 10942 -19433
rect 10880 -19743 10942 -19731
rect 10972 -19433 11038 -19421
rect 10972 -19731 10988 -19433
rect 11022 -19731 11038 -19433
rect 10972 -19743 11038 -19731
rect 11068 -19433 11134 -19421
rect 11068 -19731 11084 -19433
rect 11118 -19731 11134 -19433
rect 11068 -19743 11134 -19731
rect 11164 -19433 11230 -19421
rect 11164 -19731 11180 -19433
rect 11214 -19731 11230 -19433
rect 11164 -19743 11230 -19731
rect 11260 -19433 11326 -19421
rect 11260 -19731 11276 -19433
rect 11310 -19731 11326 -19433
rect 11260 -19743 11326 -19731
rect 11356 -19433 11422 -19421
rect 11356 -19731 11372 -19433
rect 11406 -19731 11422 -19433
rect 11356 -19743 11422 -19731
rect 11452 -19433 11518 -19421
rect 11452 -19731 11468 -19433
rect 11502 -19731 11518 -19433
rect 11452 -19743 11518 -19731
rect 11548 -19433 11614 -19421
rect 11548 -19731 11564 -19433
rect 11598 -19731 11614 -19433
rect 11548 -19743 11614 -19731
rect 11644 -19433 11706 -19421
rect 11644 -19731 11660 -19433
rect 11694 -19731 11706 -19433
rect 15763 -19493 15775 -18661
rect 15809 -19493 15825 -18661
rect 15763 -19505 15825 -19493
rect 15855 -18661 15921 -18649
rect 15855 -19493 15871 -18661
rect 15905 -19493 15921 -18661
rect 15855 -19505 15921 -19493
rect 15951 -18661 16017 -18649
rect 15951 -19493 15967 -18661
rect 16001 -19493 16017 -18661
rect 15951 -19505 16017 -19493
rect 16047 -18661 16113 -18649
rect 16047 -19493 16063 -18661
rect 16097 -19493 16113 -18661
rect 16047 -19505 16113 -19493
rect 16143 -18661 16209 -18649
rect 16143 -19493 16159 -18661
rect 16193 -19493 16209 -18661
rect 16143 -19505 16209 -19493
rect 16239 -18661 16305 -18649
rect 16239 -19493 16255 -18661
rect 16289 -19493 16305 -18661
rect 16239 -19505 16305 -19493
rect 16335 -18661 16401 -18649
rect 16335 -19493 16351 -18661
rect 16385 -19493 16401 -18661
rect 16335 -19505 16401 -19493
rect 16431 -18661 16497 -18649
rect 16431 -19493 16447 -18661
rect 16481 -19493 16497 -18661
rect 16431 -19505 16497 -19493
rect 16527 -18661 16593 -18649
rect 16527 -19493 16543 -18661
rect 16577 -19493 16593 -18661
rect 16527 -19505 16593 -19493
rect 16623 -18661 16689 -18649
rect 16623 -19493 16639 -18661
rect 16673 -19493 16689 -18661
rect 16623 -19505 16689 -19493
rect 16719 -18661 16785 -18649
rect 16719 -19493 16735 -18661
rect 16769 -19493 16785 -18661
rect 16719 -19505 16785 -19493
rect 16815 -18661 16881 -18649
rect 16815 -19493 16831 -18661
rect 16865 -19493 16881 -18661
rect 16815 -19505 16881 -19493
rect 16911 -18661 16973 -18649
rect 16911 -19493 16927 -18661
rect 16961 -19493 16973 -18661
rect 18096 -18593 18310 -18581
rect 16911 -19505 16973 -19493
rect 11644 -19743 11706 -19731
rect -16027 -19877 -15965 -19865
rect -24426 -20119 -24212 -20103
rect -24426 -20153 -24414 -20119
rect -24224 -20153 -24212 -20119
rect -24426 -20169 -24212 -20153
rect -24426 -20215 -24212 -20199
rect -21618 -20006 -21556 -19994
rect -21618 -20196 -21606 -20006
rect -21572 -20196 -21556 -20006
rect -21618 -20208 -21556 -20196
rect -21526 -20002 -21460 -19994
rect -21526 -20196 -21510 -20002
rect -21476 -20196 -21460 -20002
rect -21526 -20208 -21460 -20196
rect -21430 -20006 -21364 -19994
rect -21430 -20196 -21414 -20006
rect -21380 -20196 -21364 -20006
rect -21430 -20208 -21364 -20196
rect -21334 -20002 -21272 -19994
rect -21334 -20196 -21318 -20002
rect -21284 -20196 -21272 -20002
rect -21334 -20208 -21272 -20196
rect -16027 -20067 -16015 -19877
rect -15981 -20067 -15965 -19877
rect -16027 -20079 -15965 -20067
rect -15935 -19873 -15869 -19865
rect -15935 -20067 -15919 -19873
rect -15885 -20067 -15869 -19873
rect -15935 -20079 -15869 -20067
rect -15839 -19877 -15773 -19865
rect -15839 -20067 -15823 -19877
rect -15789 -20067 -15773 -19877
rect -15839 -20079 -15773 -20067
rect -15743 -19873 -15681 -19865
rect -15743 -20067 -15727 -19873
rect -15693 -20067 -15681 -19873
rect -12314 -19878 -11764 -19866
rect -15743 -20079 -15681 -20067
rect -12314 -19912 -12302 -19878
rect -11776 -19912 -11764 -19878
rect -12314 -19924 -11764 -19912
rect -17677 -20111 -17421 -20099
rect -17677 -20145 -17665 -20111
rect -17433 -20145 -17421 -20111
rect -17677 -20161 -17421 -20145
rect -17677 -20207 -17421 -20191
rect -24426 -20249 -24414 -20215
rect -24224 -20249 -24212 -20215
rect -24426 -20261 -24212 -20249
rect -17677 -20241 -17665 -20207
rect -17433 -20241 -17421 -20207
rect -17677 -20257 -17421 -20241
rect -17677 -20303 -17421 -20287
rect -17677 -20337 -17665 -20303
rect -17433 -20337 -17421 -20303
rect -17677 -20353 -17421 -20337
rect -17677 -20399 -17421 -20383
rect -17677 -20433 -17665 -20399
rect -17433 -20433 -17421 -20399
rect -21618 -20466 -21556 -20454
rect -21618 -20656 -21606 -20466
rect -21572 -20656 -21556 -20466
rect -21618 -20668 -21556 -20656
rect -21526 -20462 -21460 -20454
rect -21526 -20656 -21510 -20462
rect -21476 -20656 -21460 -20462
rect -21526 -20668 -21460 -20656
rect -21430 -20466 -21364 -20454
rect -21430 -20656 -21414 -20466
rect -21380 -20656 -21364 -20466
rect -21430 -20668 -21364 -20656
rect -21334 -20462 -21272 -20454
rect -21334 -20656 -21318 -20462
rect -21284 -20656 -21272 -20462
rect -17677 -20449 -17421 -20433
rect -21334 -20668 -21272 -20656
rect -17677 -20495 -17421 -20479
rect -17677 -20529 -17665 -20495
rect -17433 -20529 -17421 -20495
rect -17677 -20545 -17421 -20529
rect -16027 -20337 -15965 -20325
rect -17677 -20591 -17421 -20575
rect -17677 -20625 -17665 -20591
rect -17433 -20625 -17421 -20591
rect -17677 -20641 -17421 -20625
rect -17677 -20687 -17421 -20671
rect -24395 -20839 -24181 -20827
rect -24395 -20873 -24383 -20839
rect -24193 -20873 -24181 -20839
rect -24395 -20889 -24181 -20873
rect -24395 -20935 -24181 -20919
rect -24395 -20969 -24383 -20935
rect -24193 -20969 -24181 -20935
rect -24395 -20985 -24181 -20969
rect -24395 -21031 -24181 -21015
rect -24395 -21065 -24383 -21031
rect -24193 -21065 -24181 -21031
rect -24395 -21081 -24181 -21065
rect -24395 -21127 -24181 -21111
rect -24395 -21161 -24383 -21127
rect -24193 -21161 -24181 -21127
rect -24395 -21177 -24181 -21161
rect -24395 -21223 -24181 -21207
rect -24395 -21257 -24383 -21223
rect -24193 -21257 -24181 -21223
rect -24395 -21273 -24181 -21257
rect -21632 -20926 -21570 -20914
rect -21632 -21116 -21620 -20926
rect -21586 -21116 -21570 -20926
rect -21632 -21128 -21570 -21116
rect -21540 -20922 -21474 -20914
rect -21540 -21116 -21524 -20922
rect -21490 -21116 -21474 -20922
rect -21540 -21128 -21474 -21116
rect -21444 -20926 -21378 -20914
rect -21444 -21116 -21428 -20926
rect -21394 -21116 -21378 -20926
rect -21444 -21128 -21378 -21116
rect -21348 -20922 -21286 -20914
rect -21348 -21116 -21332 -20922
rect -21298 -21116 -21286 -20922
rect -21348 -21128 -21286 -21116
rect -17677 -20721 -17665 -20687
rect -17433 -20721 -17421 -20687
rect -17677 -20737 -17421 -20721
rect -16027 -20527 -16015 -20337
rect -15981 -20527 -15965 -20337
rect -16027 -20539 -15965 -20527
rect -15935 -20333 -15869 -20325
rect -15935 -20527 -15919 -20333
rect -15885 -20527 -15869 -20333
rect -15935 -20539 -15869 -20527
rect -15839 -20337 -15773 -20325
rect -15839 -20527 -15823 -20337
rect -15789 -20527 -15773 -20337
rect -15839 -20539 -15773 -20527
rect -15743 -20333 -15681 -20325
rect -15743 -20527 -15727 -20333
rect -15693 -20527 -15681 -20333
rect -15743 -20539 -15681 -20527
rect -17677 -20783 -17421 -20767
rect -17677 -20817 -17665 -20783
rect -17433 -20817 -17421 -20783
rect -17677 -20833 -17421 -20817
rect -17677 -20879 -17421 -20863
rect -17677 -20913 -17665 -20879
rect -17433 -20913 -17421 -20879
rect -17677 -20929 -17421 -20913
rect -17677 -20975 -17421 -20959
rect -17677 -21009 -17665 -20975
rect -17433 -21009 -17421 -20975
rect -17677 -21025 -17421 -21009
rect -16041 -20797 -15979 -20785
rect -16041 -20987 -16029 -20797
rect -15995 -20987 -15979 -20797
rect -16041 -20999 -15979 -20987
rect -15949 -20793 -15883 -20785
rect -15949 -20987 -15933 -20793
rect -15899 -20987 -15883 -20793
rect -15949 -20999 -15883 -20987
rect -15853 -20797 -15787 -20785
rect -15853 -20987 -15837 -20797
rect -15803 -20987 -15787 -20797
rect -15853 -20999 -15787 -20987
rect -15757 -20793 -15695 -20785
rect -15757 -20987 -15741 -20793
rect -15707 -20987 -15695 -20793
rect -15757 -20999 -15695 -20987
rect -17677 -21071 -17421 -21055
rect -17677 -21105 -17665 -21071
rect -17433 -21105 -17421 -21071
rect -17677 -21117 -17421 -21105
rect -12314 -19966 -11764 -19954
rect -12314 -20000 -12302 -19966
rect -11776 -20000 -11764 -19966
rect -12314 -20016 -11764 -20000
rect -12314 -20062 -11764 -20046
rect -12314 -20096 -12302 -20062
rect -11776 -20096 -11764 -20062
rect -12314 -20112 -11764 -20096
rect -12314 -20158 -11764 -20142
rect -12314 -20192 -12302 -20158
rect -11776 -20192 -11764 -20158
rect -12314 -20208 -11764 -20192
rect -12314 -20254 -11764 -20238
rect -12314 -20288 -12302 -20254
rect -11776 -20288 -11764 -20254
rect -12314 -20304 -11764 -20288
rect -12314 -20350 -11764 -20334
rect -12314 -20384 -12302 -20350
rect -11776 -20384 -11764 -20350
rect -12314 -20400 -11764 -20384
rect -12314 -20446 -11764 -20430
rect -12314 -20480 -12302 -20446
rect -11776 -20480 -11764 -20446
rect -12314 -20496 -11764 -20480
rect -12314 -20542 -11764 -20526
rect -12314 -20576 -12302 -20542
rect -11776 -20576 -11764 -20542
rect -12314 -20592 -11764 -20576
rect -12314 -20638 -11764 -20622
rect -12314 -20672 -12302 -20638
rect -11776 -20672 -11764 -20638
rect -12314 -20688 -11764 -20672
rect -12314 -20734 -11764 -20718
rect -12314 -20768 -12302 -20734
rect -11776 -20768 -11764 -20734
rect -12314 -20784 -11764 -20768
rect -12314 -20830 -11764 -20814
rect -12314 -20864 -12302 -20830
rect -11776 -20864 -11764 -20830
rect -12314 -20880 -11764 -20864
rect -12314 -20926 -11764 -20910
rect -12314 -20960 -12302 -20926
rect -11776 -20960 -11764 -20926
rect -12314 -20976 -11764 -20960
rect -12314 -21022 -11764 -21006
rect -12314 -21056 -12302 -21022
rect -11776 -21056 -11764 -21022
rect -12314 -21072 -11764 -21056
rect -12314 -21118 -11764 -21102
rect -12314 -21152 -12302 -21118
rect -11776 -21152 -11764 -21118
rect -12314 -21164 -11764 -21152
rect -4828 -19948 -4766 -19936
rect -4828 -20138 -4816 -19948
rect -4782 -20138 -4766 -19948
rect -4828 -20150 -4766 -20138
rect -4736 -19948 -4670 -19936
rect -4736 -20142 -4720 -19948
rect -4686 -20142 -4670 -19948
rect -4736 -20150 -4670 -20142
rect -4640 -19948 -4574 -19936
rect -4640 -20138 -4624 -19948
rect -4590 -20138 -4574 -19948
rect -4640 -20150 -4574 -20138
rect -4544 -19948 -4482 -19936
rect -4544 -20142 -4528 -19948
rect -4494 -20142 -4482 -19948
rect -2112 -19942 -2050 -19930
rect -4544 -20150 -4482 -20142
rect -2112 -20132 -2100 -19942
rect -2066 -20132 -2050 -19942
rect -2112 -20144 -2050 -20132
rect -2020 -19938 -1954 -19930
rect -2020 -20132 -2004 -19938
rect -1970 -20132 -1954 -19938
rect -2020 -20144 -1954 -20132
rect -1924 -19942 -1858 -19930
rect -1924 -20132 -1908 -19942
rect -1874 -20132 -1858 -19942
rect -1924 -20144 -1858 -20132
rect -1828 -19938 -1766 -19930
rect -1828 -20132 -1812 -19938
rect -1778 -20132 -1766 -19938
rect -1828 -20144 -1766 -20132
rect -4828 -20388 -4766 -20376
rect -4828 -20578 -4816 -20388
rect -4782 -20578 -4766 -20388
rect -4828 -20590 -4766 -20578
rect -4736 -20388 -4670 -20376
rect -4736 -20582 -4720 -20388
rect -4686 -20582 -4670 -20388
rect -4736 -20590 -4670 -20582
rect -4640 -20388 -4574 -20376
rect -4640 -20578 -4624 -20388
rect -4590 -20578 -4574 -20388
rect -4640 -20590 -4574 -20578
rect -4544 -20388 -4482 -20376
rect -4544 -20582 -4528 -20388
rect -4494 -20582 -4482 -20388
rect -2112 -20382 -2050 -20370
rect -4544 -20590 -4482 -20582
rect -2112 -20572 -2100 -20382
rect -2066 -20572 -2050 -20382
rect -2112 -20584 -2050 -20572
rect -2020 -20378 -1954 -20370
rect -2020 -20572 -2004 -20378
rect -1970 -20572 -1954 -20378
rect -2020 -20584 -1954 -20572
rect -1924 -20382 -1858 -20370
rect -1924 -20572 -1908 -20382
rect -1874 -20572 -1858 -20382
rect -1924 -20584 -1858 -20572
rect -1828 -20378 -1766 -20370
rect -1828 -20572 -1812 -20378
rect -1778 -20572 -1766 -20378
rect -1828 -20584 -1766 -20572
rect -4828 -20767 -4766 -20755
rect -4828 -20957 -4816 -20767
rect -4782 -20957 -4766 -20767
rect -4828 -20969 -4766 -20957
rect -4736 -20767 -4670 -20755
rect -4736 -20961 -4720 -20767
rect -4686 -20961 -4670 -20767
rect -4736 -20969 -4670 -20961
rect -4640 -20767 -4574 -20755
rect -4640 -20957 -4624 -20767
rect -4590 -20957 -4574 -20767
rect -4640 -20969 -4574 -20957
rect -4544 -20767 -4482 -20755
rect -4544 -20961 -4528 -20767
rect -4494 -20961 -4482 -20767
rect 11773 -20643 11835 -20631
rect 11773 -20875 11785 -20643
rect 11819 -20875 11835 -20643
rect 11773 -20887 11835 -20875
rect 11865 -20643 11931 -20631
rect 11865 -20875 11881 -20643
rect 11915 -20875 11931 -20643
rect 11865 -20887 11931 -20875
rect 11961 -20643 12027 -20631
rect 11961 -20875 11977 -20643
rect 12011 -20875 12027 -20643
rect 11961 -20887 12027 -20875
rect 12057 -20643 12123 -20631
rect 12057 -20875 12073 -20643
rect 12107 -20875 12123 -20643
rect 12057 -20887 12123 -20875
rect 12153 -20643 12219 -20631
rect 12153 -20875 12169 -20643
rect 12203 -20875 12219 -20643
rect 12153 -20887 12219 -20875
rect 12249 -20643 12315 -20631
rect 12249 -20875 12265 -20643
rect 12299 -20875 12315 -20643
rect 12249 -20887 12315 -20875
rect 12345 -20643 12411 -20631
rect 12345 -20875 12361 -20643
rect 12395 -20875 12411 -20643
rect 12345 -20887 12411 -20875
rect 12441 -20643 12507 -20631
rect 12441 -20875 12457 -20643
rect 12491 -20875 12507 -20643
rect 12441 -20887 12507 -20875
rect 12537 -20643 12603 -20631
rect 12537 -20875 12553 -20643
rect 12587 -20875 12603 -20643
rect 12537 -20887 12603 -20875
rect 12633 -20643 12699 -20631
rect 12633 -20875 12649 -20643
rect 12683 -20875 12699 -20643
rect 12633 -20887 12699 -20875
rect 12729 -20643 12791 -20631
rect 12729 -20875 12745 -20643
rect 12779 -20875 12791 -20643
rect 12923 -20747 13137 -20735
rect 12729 -20887 12791 -20875
rect -4544 -20969 -4482 -20961
rect -12314 -21206 -11764 -21194
rect -24395 -21319 -24181 -21303
rect -24395 -21353 -24383 -21319
rect -24193 -21353 -24181 -21319
rect -24395 -21369 -24181 -21353
rect -12314 -21240 -12302 -21206
rect -11776 -21240 -11764 -21206
rect -12314 -21252 -11764 -21240
rect -16039 -21277 -15977 -21265
rect -24395 -21415 -24181 -21399
rect -24395 -21449 -24383 -21415
rect -24193 -21449 -24181 -21415
rect -24395 -21461 -24181 -21449
rect -21630 -21406 -21568 -21394
rect -21630 -21596 -21618 -21406
rect -21584 -21596 -21568 -21406
rect -21630 -21608 -21568 -21596
rect -21538 -21402 -21472 -21394
rect -21538 -21596 -21522 -21402
rect -21488 -21596 -21472 -21402
rect -21538 -21608 -21472 -21596
rect -21442 -21406 -21376 -21394
rect -21442 -21596 -21426 -21406
rect -21392 -21596 -21376 -21406
rect -21442 -21608 -21376 -21596
rect -21346 -21402 -21284 -21394
rect -21346 -21596 -21330 -21402
rect -21296 -21596 -21284 -21402
rect -21346 -21608 -21284 -21596
rect -16039 -21467 -16027 -21277
rect -15993 -21467 -15977 -21277
rect -16039 -21479 -15977 -21467
rect -15947 -21273 -15881 -21265
rect -15947 -21467 -15931 -21273
rect -15897 -21467 -15881 -21273
rect -15947 -21479 -15881 -21467
rect -15851 -21277 -15785 -21265
rect -15851 -21467 -15835 -21277
rect -15801 -21467 -15785 -21277
rect -15851 -21479 -15785 -21467
rect -15755 -21273 -15693 -21265
rect -15755 -21467 -15739 -21273
rect -15705 -21467 -15693 -21273
rect -15755 -21479 -15693 -21467
rect -17677 -21511 -17421 -21499
rect -17677 -21545 -17665 -21511
rect -17433 -21545 -17421 -21511
rect -17677 -21561 -17421 -21545
rect -17677 -21607 -17421 -21591
rect -17677 -21641 -17665 -21607
rect -17433 -21641 -17421 -21607
rect -17677 -21657 -17421 -21641
rect -17677 -21703 -17421 -21687
rect -17677 -21737 -17665 -21703
rect -17433 -21737 -17421 -21703
rect -17677 -21753 -17421 -21737
rect -17677 -21799 -17421 -21783
rect -17677 -21833 -17665 -21799
rect -17433 -21833 -17421 -21799
rect -17677 -21849 -17421 -21833
rect -17677 -21895 -17421 -21879
rect -17677 -21929 -17665 -21895
rect -17433 -21929 -17421 -21895
rect -17677 -21945 -17421 -21929
rect -17677 -21991 -17421 -21975
rect -17677 -22025 -17665 -21991
rect -17433 -22025 -17421 -21991
rect -17677 -22041 -17421 -22025
rect -17677 -22087 -17421 -22071
rect -24396 -22142 -24182 -22130
rect -24396 -22176 -24384 -22142
rect -24194 -22176 -24182 -22142
rect -24396 -22192 -24182 -22176
rect -24396 -22238 -24182 -22222
rect -24396 -22272 -24384 -22238
rect -24194 -22272 -24182 -22238
rect -24396 -22288 -24182 -22272
rect -24396 -22334 -24182 -22318
rect -24396 -22368 -24384 -22334
rect -24194 -22368 -24182 -22334
rect -24396 -22384 -24182 -22368
rect -24396 -22430 -24182 -22414
rect -24396 -22464 -24384 -22430
rect -24194 -22464 -24182 -22430
rect -24396 -22480 -24182 -22464
rect -24396 -22526 -24182 -22510
rect -24396 -22560 -24384 -22526
rect -24194 -22560 -24182 -22526
rect -24396 -22576 -24182 -22560
rect -17677 -22121 -17665 -22087
rect -17433 -22121 -17421 -22087
rect -17677 -22137 -17421 -22121
rect -17677 -22183 -17421 -22167
rect -17677 -22217 -17665 -22183
rect -17433 -22217 -17421 -22183
rect -17677 -22233 -17421 -22217
rect 12923 -20781 12935 -20747
rect 13125 -20781 13137 -20747
rect 12923 -20797 13137 -20781
rect 12923 -20843 13137 -20827
rect 12923 -20877 12935 -20843
rect 13129 -20877 13137 -20843
rect 12923 -20893 13137 -20877
rect 12923 -20939 13137 -20923
rect 12923 -20973 12935 -20939
rect 13125 -20973 13137 -20939
rect 12923 -20989 13137 -20973
rect 12923 -21035 13137 -21019
rect 12923 -21069 12935 -21035
rect 13129 -21069 13137 -21035
rect 12923 -21081 13137 -21069
rect -17677 -22279 -17421 -22263
rect -17677 -22313 -17665 -22279
rect -17433 -22313 -17421 -22279
rect -17677 -22329 -17421 -22313
rect -17677 -22375 -17421 -22359
rect -17677 -22409 -17665 -22375
rect -17433 -22409 -17421 -22375
rect -17677 -22425 -17421 -22409
rect 7138 -22297 7200 -22285
rect -17677 -22471 -17421 -22455
rect -17677 -22505 -17665 -22471
rect -17433 -22505 -17421 -22471
rect -12314 -22457 -11764 -22445
rect -12314 -22491 -12302 -22457
rect -11776 -22491 -11764 -22457
rect -12314 -22503 -11764 -22491
rect -17677 -22517 -17421 -22505
rect -24396 -22622 -24182 -22606
rect -24396 -22656 -24384 -22622
rect -24194 -22656 -24182 -22622
rect -24396 -22672 -24182 -22656
rect -24396 -22718 -24182 -22702
rect -24396 -22752 -24384 -22718
rect -24194 -22752 -24182 -22718
rect -24396 -22764 -24182 -22752
rect -17677 -22911 -17421 -22899
rect -17677 -22945 -17665 -22911
rect -17433 -22945 -17421 -22911
rect -17677 -22961 -17421 -22945
rect -17677 -23007 -17421 -22991
rect -17677 -23041 -17665 -23007
rect -17433 -23041 -17421 -23007
rect -17677 -23057 -17421 -23041
rect -17677 -23103 -17421 -23087
rect -17677 -23137 -17665 -23103
rect -17433 -23137 -17421 -23103
rect -17677 -23153 -17421 -23137
rect -17677 -23199 -17421 -23183
rect -17677 -23233 -17665 -23199
rect -17433 -23233 -17421 -23199
rect -17677 -23249 -17421 -23233
rect -17677 -23295 -17421 -23279
rect -17677 -23329 -17665 -23295
rect -17433 -23329 -17421 -23295
rect -17677 -23345 -17421 -23329
rect -17677 -23391 -17421 -23375
rect -17677 -23425 -17665 -23391
rect -17433 -23425 -17421 -23391
rect -24396 -23451 -24182 -23439
rect -24396 -23485 -24384 -23451
rect -24194 -23485 -24182 -23451
rect -24396 -23501 -24182 -23485
rect -24396 -23547 -24182 -23531
rect -24396 -23581 -24384 -23547
rect -24194 -23581 -24182 -23547
rect -24396 -23597 -24182 -23581
rect -24396 -23643 -24182 -23627
rect -24396 -23677 -24384 -23643
rect -24194 -23677 -24182 -23643
rect -24396 -23693 -24182 -23677
rect -24396 -23739 -24182 -23723
rect -24396 -23773 -24384 -23739
rect -24194 -23773 -24182 -23739
rect -24396 -23789 -24182 -23773
rect -24396 -23835 -24182 -23819
rect -24396 -23869 -24384 -23835
rect -24194 -23869 -24182 -23835
rect -24396 -23885 -24182 -23869
rect -17677 -23441 -17421 -23425
rect -17677 -23487 -17421 -23471
rect -24396 -23931 -24182 -23915
rect -24396 -23965 -24384 -23931
rect -24194 -23965 -24182 -23931
rect -24396 -23981 -24182 -23965
rect -17677 -23521 -17665 -23487
rect -17433 -23521 -17421 -23487
rect -17677 -23537 -17421 -23521
rect -17677 -23583 -17421 -23567
rect -17677 -23617 -17665 -23583
rect -17433 -23617 -17421 -23583
rect -17677 -23633 -17421 -23617
rect -17677 -23679 -17421 -23663
rect -17677 -23713 -17665 -23679
rect -17433 -23713 -17421 -23679
rect -17677 -23729 -17421 -23713
rect -12314 -22545 -11764 -22533
rect -12314 -22579 -12302 -22545
rect -11776 -22579 -11764 -22545
rect -12314 -22595 -11764 -22579
rect -12314 -22641 -11764 -22625
rect -12314 -22675 -12302 -22641
rect -11776 -22675 -11764 -22641
rect -12314 -22691 -11764 -22675
rect -12314 -22737 -11764 -22721
rect -12314 -22771 -12302 -22737
rect -11776 -22771 -11764 -22737
rect -12314 -22787 -11764 -22771
rect -12314 -22833 -11764 -22817
rect -12314 -22867 -12302 -22833
rect -11776 -22867 -11764 -22833
rect -12314 -22883 -11764 -22867
rect -12314 -22929 -11764 -22913
rect -12314 -22963 -12302 -22929
rect -11776 -22963 -11764 -22929
rect -12314 -22979 -11764 -22963
rect -12314 -23025 -11764 -23009
rect -12314 -23059 -12302 -23025
rect -11776 -23059 -11764 -23025
rect -12314 -23075 -11764 -23059
rect -12314 -23121 -11764 -23105
rect -12314 -23155 -12302 -23121
rect -11776 -23155 -11764 -23121
rect -12314 -23171 -11764 -23155
rect -12314 -23217 -11764 -23201
rect -12314 -23251 -12302 -23217
rect -11776 -23251 -11764 -23217
rect -12314 -23267 -11764 -23251
rect -12314 -23313 -11764 -23297
rect -12314 -23347 -12302 -23313
rect -11776 -23347 -11764 -23313
rect -12314 -23363 -11764 -23347
rect -12314 -23409 -11764 -23393
rect -12314 -23443 -12302 -23409
rect -11776 -23443 -11764 -23409
rect -12314 -23459 -11764 -23443
rect -12314 -23505 -11764 -23489
rect -12314 -23539 -12302 -23505
rect -11776 -23539 -11764 -23505
rect -12314 -23555 -11764 -23539
rect -12314 -23601 -11764 -23585
rect -12314 -23635 -12302 -23601
rect -11776 -23635 -11764 -23601
rect -12314 -23651 -11764 -23635
rect -12314 -23697 -11764 -23681
rect -12314 -23731 -12302 -23697
rect -11776 -23731 -11764 -23697
rect -12314 -23743 -11764 -23731
rect 7138 -22595 7150 -22297
rect 7184 -22595 7200 -22297
rect 7138 -22607 7200 -22595
rect 7230 -22297 7296 -22285
rect 7230 -22595 7246 -22297
rect 7280 -22595 7296 -22297
rect 7230 -22607 7296 -22595
rect 7326 -22297 7392 -22285
rect 7326 -22595 7342 -22297
rect 7376 -22595 7392 -22297
rect 7326 -22607 7392 -22595
rect 7422 -22297 7488 -22285
rect 7422 -22595 7438 -22297
rect 7472 -22595 7488 -22297
rect 7422 -22607 7488 -22595
rect 7518 -22297 7584 -22285
rect 7518 -22595 7534 -22297
rect 7568 -22595 7584 -22297
rect 7518 -22607 7584 -22595
rect 7614 -22297 7680 -22285
rect 7614 -22595 7630 -22297
rect 7664 -22595 7680 -22297
rect 7614 -22607 7680 -22595
rect 7710 -22297 7776 -22285
rect 7710 -22595 7726 -22297
rect 7760 -22595 7776 -22297
rect 7710 -22607 7776 -22595
rect 7806 -22297 7872 -22285
rect 7806 -22595 7822 -22297
rect 7856 -22595 7872 -22297
rect 7806 -22607 7872 -22595
rect 7902 -22297 7964 -22285
rect 7902 -22595 7918 -22297
rect 7952 -22595 7964 -22297
rect 7902 -22607 7964 -22595
rect 8086 -22297 8148 -22285
rect 8086 -22595 8098 -22297
rect 8132 -22595 8148 -22297
rect 8086 -22607 8148 -22595
rect 8178 -22297 8244 -22285
rect 8178 -22595 8194 -22297
rect 8228 -22595 8244 -22297
rect 8178 -22607 8244 -22595
rect 8274 -22297 8340 -22285
rect 8274 -22595 8290 -22297
rect 8324 -22595 8340 -22297
rect 8274 -22607 8340 -22595
rect 8370 -22297 8436 -22285
rect 8370 -22595 8386 -22297
rect 8420 -22595 8436 -22297
rect 8370 -22607 8436 -22595
rect 8466 -22297 8532 -22285
rect 8466 -22595 8482 -22297
rect 8516 -22595 8532 -22297
rect 8466 -22607 8532 -22595
rect 8562 -22297 8628 -22285
rect 8562 -22595 8578 -22297
rect 8612 -22595 8628 -22297
rect 8562 -22607 8628 -22595
rect 8658 -22297 8724 -22285
rect 8658 -22595 8674 -22297
rect 8708 -22595 8724 -22297
rect 8658 -22607 8724 -22595
rect 8754 -22297 8820 -22285
rect 8754 -22595 8770 -22297
rect 8804 -22595 8820 -22297
rect 8754 -22607 8820 -22595
rect 8850 -22297 8912 -22285
rect 8850 -22595 8866 -22297
rect 8900 -22595 8912 -22297
rect 8850 -22607 8912 -22595
rect 9022 -22297 9084 -22285
rect 9022 -22595 9034 -22297
rect 9068 -22595 9084 -22297
rect 9022 -22607 9084 -22595
rect 9114 -22297 9180 -22285
rect 9114 -22595 9130 -22297
rect 9164 -22595 9180 -22297
rect 9114 -22607 9180 -22595
rect 9210 -22297 9276 -22285
rect 9210 -22595 9226 -22297
rect 9260 -22595 9276 -22297
rect 9210 -22607 9276 -22595
rect 9306 -22297 9372 -22285
rect 9306 -22595 9322 -22297
rect 9356 -22595 9372 -22297
rect 9306 -22607 9372 -22595
rect 9402 -22297 9468 -22285
rect 9402 -22595 9418 -22297
rect 9452 -22595 9468 -22297
rect 9402 -22607 9468 -22595
rect 9498 -22297 9564 -22285
rect 9498 -22595 9514 -22297
rect 9548 -22595 9564 -22297
rect 9498 -22607 9564 -22595
rect 9594 -22297 9660 -22285
rect 9594 -22595 9610 -22297
rect 9644 -22595 9660 -22297
rect 9594 -22607 9660 -22595
rect 9690 -22297 9756 -22285
rect 9690 -22595 9706 -22297
rect 9740 -22595 9756 -22297
rect 9690 -22607 9756 -22595
rect 9786 -22297 9848 -22285
rect 9786 -22595 9802 -22297
rect 9836 -22595 9848 -22297
rect 9786 -22607 9848 -22595
rect 9953 -22296 10015 -22284
rect 9953 -22594 9965 -22296
rect 9999 -22594 10015 -22296
rect 9953 -22606 10015 -22594
rect 10045 -22296 10111 -22284
rect 10045 -22594 10061 -22296
rect 10095 -22594 10111 -22296
rect 10045 -22606 10111 -22594
rect 10141 -22296 10207 -22284
rect 10141 -22594 10157 -22296
rect 10191 -22594 10207 -22296
rect 10141 -22606 10207 -22594
rect 10237 -22296 10303 -22284
rect 10237 -22594 10253 -22296
rect 10287 -22594 10303 -22296
rect 10237 -22606 10303 -22594
rect 10333 -22296 10399 -22284
rect 10333 -22594 10349 -22296
rect 10383 -22594 10399 -22296
rect 10333 -22606 10399 -22594
rect 10429 -22296 10495 -22284
rect 10429 -22594 10445 -22296
rect 10479 -22594 10495 -22296
rect 10429 -22606 10495 -22594
rect 10525 -22296 10591 -22284
rect 10525 -22594 10541 -22296
rect 10575 -22594 10591 -22296
rect 10525 -22606 10591 -22594
rect 10621 -22296 10687 -22284
rect 10621 -22594 10637 -22296
rect 10671 -22594 10687 -22296
rect 10621 -22606 10687 -22594
rect 10717 -22296 10779 -22284
rect 10717 -22594 10733 -22296
rect 10767 -22594 10779 -22296
rect 10717 -22606 10779 -22594
rect 10880 -22297 10942 -22285
rect 10880 -22595 10892 -22297
rect 10926 -22595 10942 -22297
rect 10880 -22607 10942 -22595
rect 10972 -22297 11038 -22285
rect 10972 -22595 10988 -22297
rect 11022 -22595 11038 -22297
rect 10972 -22607 11038 -22595
rect 11068 -22297 11134 -22285
rect 11068 -22595 11084 -22297
rect 11118 -22595 11134 -22297
rect 11068 -22607 11134 -22595
rect 11164 -22297 11230 -22285
rect 11164 -22595 11180 -22297
rect 11214 -22595 11230 -22297
rect 11164 -22607 11230 -22595
rect 11260 -22297 11326 -22285
rect 11260 -22595 11276 -22297
rect 11310 -22595 11326 -22297
rect 11260 -22607 11326 -22595
rect 11356 -22297 11422 -22285
rect 11356 -22595 11372 -22297
rect 11406 -22595 11422 -22297
rect 11356 -22607 11422 -22595
rect 11452 -22297 11518 -22285
rect 11452 -22595 11468 -22297
rect 11502 -22595 11518 -22297
rect 11452 -22607 11518 -22595
rect 11548 -22297 11614 -22285
rect 11548 -22595 11564 -22297
rect 11598 -22595 11614 -22297
rect 11548 -22607 11614 -22595
rect 11644 -22297 11706 -22285
rect 11644 -22595 11660 -22297
rect 11694 -22595 11706 -22297
rect 11644 -22607 11706 -22595
rect 5658 -23257 5872 -23245
rect 5658 -23291 5670 -23257
rect 5860 -23291 5872 -23257
rect 6098 -23257 6312 -23245
rect 5658 -23307 5872 -23291
rect 5658 -23353 5872 -23337
rect 5658 -23387 5670 -23353
rect 5864 -23387 5872 -23353
rect 5658 -23403 5872 -23387
rect 5658 -23449 5872 -23433
rect 5658 -23483 5670 -23449
rect 5860 -23483 5872 -23449
rect 5658 -23499 5872 -23483
rect 5658 -23545 5872 -23529
rect 5658 -23579 5670 -23545
rect 5864 -23579 5872 -23545
rect 6098 -23291 6110 -23257
rect 6300 -23291 6312 -23257
rect 6538 -23257 6752 -23245
rect 6098 -23307 6312 -23291
rect 6098 -23353 6312 -23337
rect 6098 -23387 6110 -23353
rect 6304 -23387 6312 -23353
rect 6098 -23403 6312 -23387
rect 6098 -23449 6312 -23433
rect 6098 -23483 6110 -23449
rect 6300 -23483 6312 -23449
rect 6098 -23499 6312 -23483
rect 6098 -23545 6312 -23529
rect 5658 -23591 5872 -23579
rect 6098 -23579 6110 -23545
rect 6304 -23579 6312 -23545
rect 6538 -23291 6550 -23257
rect 6740 -23291 6752 -23257
rect 6538 -23307 6752 -23291
rect 6538 -23353 6752 -23337
rect 6538 -23387 6550 -23353
rect 6744 -23387 6752 -23353
rect 6538 -23403 6752 -23387
rect 6538 -23449 6752 -23433
rect 6538 -23483 6550 -23449
rect 6740 -23483 6752 -23449
rect 6538 -23499 6752 -23483
rect 6538 -23545 6752 -23529
rect 6098 -23591 6312 -23579
rect 6538 -23579 6550 -23545
rect 6744 -23579 6752 -23545
rect 6538 -23591 6752 -23579
rect -17677 -23775 -17421 -23759
rect -17677 -23809 -17665 -23775
rect -17433 -23809 -17421 -23775
rect -17677 -23825 -17421 -23809
rect -12314 -23785 -11764 -23773
rect -12314 -23819 -12302 -23785
rect -11776 -23819 -11764 -23785
rect -12314 -23831 -11764 -23819
rect -17677 -23871 -17421 -23855
rect -17677 -23905 -17665 -23871
rect -17433 -23905 -17421 -23871
rect -17677 -23917 -17421 -23905
rect -24396 -24027 -24182 -24011
rect -24396 -24061 -24384 -24027
rect -24194 -24061 -24182 -24027
rect 7138 -23961 7200 -23949
rect -24396 -24073 -24182 -24061
rect 7138 -24259 7150 -23961
rect 7184 -24259 7200 -23961
rect 7138 -24271 7200 -24259
rect 7230 -23961 7296 -23949
rect 7230 -24259 7246 -23961
rect 7280 -24259 7296 -23961
rect 7230 -24271 7296 -24259
rect 7326 -23961 7392 -23949
rect 7326 -24259 7342 -23961
rect 7376 -24259 7392 -23961
rect 7326 -24271 7392 -24259
rect 7422 -23961 7488 -23949
rect 7422 -24259 7438 -23961
rect 7472 -24259 7488 -23961
rect 7422 -24271 7488 -24259
rect 7518 -23961 7584 -23949
rect 7518 -24259 7534 -23961
rect 7568 -24259 7584 -23961
rect 7518 -24271 7584 -24259
rect 7614 -23961 7680 -23949
rect 7614 -24259 7630 -23961
rect 7664 -24259 7680 -23961
rect 7614 -24271 7680 -24259
rect 7710 -23961 7776 -23949
rect 7710 -24259 7726 -23961
rect 7760 -24259 7776 -23961
rect 7710 -24271 7776 -24259
rect 7806 -23961 7872 -23949
rect 7806 -24259 7822 -23961
rect 7856 -24259 7872 -23961
rect 7806 -24271 7872 -24259
rect 7902 -23961 7964 -23949
rect 7902 -24259 7918 -23961
rect 7952 -24259 7964 -23961
rect 7902 -24271 7964 -24259
rect 8086 -23961 8148 -23949
rect 8086 -24259 8098 -23961
rect 8132 -24259 8148 -23961
rect 8086 -24271 8148 -24259
rect 8178 -23961 8244 -23949
rect 8178 -24259 8194 -23961
rect 8228 -24259 8244 -23961
rect 8178 -24271 8244 -24259
rect 8274 -23961 8340 -23949
rect 8274 -24259 8290 -23961
rect 8324 -24259 8340 -23961
rect 8274 -24271 8340 -24259
rect 8370 -23961 8436 -23949
rect 8370 -24259 8386 -23961
rect 8420 -24259 8436 -23961
rect 8370 -24271 8436 -24259
rect 8466 -23961 8532 -23949
rect 8466 -24259 8482 -23961
rect 8516 -24259 8532 -23961
rect 8466 -24271 8532 -24259
rect 8562 -23961 8628 -23949
rect 8562 -24259 8578 -23961
rect 8612 -24259 8628 -23961
rect 8562 -24271 8628 -24259
rect 8658 -23961 8724 -23949
rect 8658 -24259 8674 -23961
rect 8708 -24259 8724 -23961
rect 8658 -24271 8724 -24259
rect 8754 -23961 8820 -23949
rect 8754 -24259 8770 -23961
rect 8804 -24259 8820 -23961
rect 8754 -24271 8820 -24259
rect 8850 -23961 8912 -23949
rect 8850 -24259 8866 -23961
rect 8900 -24259 8912 -23961
rect 8850 -24271 8912 -24259
rect 9022 -23961 9084 -23949
rect 9022 -24259 9034 -23961
rect 9068 -24259 9084 -23961
rect 9022 -24271 9084 -24259
rect 9114 -23961 9180 -23949
rect 9114 -24259 9130 -23961
rect 9164 -24259 9180 -23961
rect 9114 -24271 9180 -24259
rect 9210 -23961 9276 -23949
rect 9210 -24259 9226 -23961
rect 9260 -24259 9276 -23961
rect 9210 -24271 9276 -24259
rect 9306 -23961 9372 -23949
rect 9306 -24259 9322 -23961
rect 9356 -24259 9372 -23961
rect 9306 -24271 9372 -24259
rect 9402 -23961 9468 -23949
rect 9402 -24259 9418 -23961
rect 9452 -24259 9468 -23961
rect 9402 -24271 9468 -24259
rect 9498 -23961 9564 -23949
rect 9498 -24259 9514 -23961
rect 9548 -24259 9564 -23961
rect 9498 -24271 9564 -24259
rect 9594 -23961 9660 -23949
rect 9594 -24259 9610 -23961
rect 9644 -24259 9660 -23961
rect 9594 -24271 9660 -24259
rect 9690 -23961 9756 -23949
rect 9690 -24259 9706 -23961
rect 9740 -24259 9756 -23961
rect 9690 -24271 9756 -24259
rect 9786 -23961 9848 -23949
rect 9786 -24259 9802 -23961
rect 9836 -24259 9848 -23961
rect 9786 -24271 9848 -24259
rect 9953 -23961 10015 -23949
rect 9953 -24259 9965 -23961
rect 9999 -24259 10015 -23961
rect 9953 -24271 10015 -24259
rect 10045 -23961 10111 -23949
rect 10045 -24259 10061 -23961
rect 10095 -24259 10111 -23961
rect 10045 -24271 10111 -24259
rect 10141 -23961 10207 -23949
rect 10141 -24259 10157 -23961
rect 10191 -24259 10207 -23961
rect 10141 -24271 10207 -24259
rect 10237 -23961 10303 -23949
rect 10237 -24259 10253 -23961
rect 10287 -24259 10303 -23961
rect 10237 -24271 10303 -24259
rect 10333 -23961 10399 -23949
rect 10333 -24259 10349 -23961
rect 10383 -24259 10399 -23961
rect 10333 -24271 10399 -24259
rect 10429 -23961 10495 -23949
rect 10429 -24259 10445 -23961
rect 10479 -24259 10495 -23961
rect 10429 -24271 10495 -24259
rect 10525 -23961 10591 -23949
rect 10525 -24259 10541 -23961
rect 10575 -24259 10591 -23961
rect 10525 -24271 10591 -24259
rect 10621 -23961 10687 -23949
rect 10621 -24259 10637 -23961
rect 10671 -24259 10687 -23961
rect 10621 -24271 10687 -24259
rect 10717 -23961 10779 -23949
rect 10717 -24259 10733 -23961
rect 10767 -24259 10779 -23961
rect 10717 -24271 10779 -24259
rect 10880 -23961 10942 -23949
rect 10880 -24259 10892 -23961
rect 10926 -24259 10942 -23961
rect 10880 -24271 10942 -24259
rect 10972 -23961 11038 -23949
rect 10972 -24259 10988 -23961
rect 11022 -24259 11038 -23961
rect 10972 -24271 11038 -24259
rect 11068 -23961 11134 -23949
rect 11068 -24259 11084 -23961
rect 11118 -24259 11134 -23961
rect 11068 -24271 11134 -24259
rect 11164 -23961 11230 -23949
rect 11164 -24259 11180 -23961
rect 11214 -24259 11230 -23961
rect 11164 -24271 11230 -24259
rect 11260 -23961 11326 -23949
rect 11260 -24259 11276 -23961
rect 11310 -24259 11326 -23961
rect 11260 -24271 11326 -24259
rect 11356 -23961 11422 -23949
rect 11356 -24259 11372 -23961
rect 11406 -24259 11422 -23961
rect 11356 -24271 11422 -24259
rect 11452 -23961 11518 -23949
rect 11452 -24259 11468 -23961
rect 11502 -24259 11518 -23961
rect 11452 -24271 11518 -24259
rect 11548 -23961 11614 -23949
rect 11548 -24259 11564 -23961
rect 11598 -24259 11614 -23961
rect 11548 -24271 11614 -24259
rect 11644 -23961 11706 -23949
rect 11644 -24259 11660 -23961
rect 11694 -24259 11706 -23961
rect 11644 -24271 11706 -24259
rect -17677 -24311 -17421 -24299
rect -17677 -24345 -17665 -24311
rect -17433 -24345 -17421 -24311
rect -17677 -24361 -17421 -24345
rect -17677 -24407 -17421 -24391
rect -17677 -24441 -17665 -24407
rect -17433 -24441 -17421 -24407
rect -17677 -24457 -17421 -24441
rect -17677 -24503 -17421 -24487
rect -17677 -24537 -17665 -24503
rect -17433 -24537 -17421 -24503
rect -17677 -24553 -17421 -24537
rect -17677 -24599 -17421 -24583
rect -17677 -24633 -17665 -24599
rect -17433 -24633 -17421 -24599
rect -17677 -24649 -17421 -24633
rect -17677 -24695 -17421 -24679
rect -17677 -24729 -17665 -24695
rect -17433 -24729 -17421 -24695
rect -17677 -24745 -17421 -24729
rect -17677 -24791 -17421 -24775
rect -17677 -24825 -17665 -24791
rect -17433 -24825 -17421 -24791
rect -17677 -24841 -17421 -24825
rect -17677 -24887 -17421 -24871
rect -17677 -24921 -17665 -24887
rect -17433 -24921 -17421 -24887
rect -17677 -24937 -17421 -24921
rect -17677 -24983 -17421 -24967
rect -17677 -25017 -17665 -24983
rect -17433 -25017 -17421 -24983
rect -17677 -25033 -17421 -25017
rect -17677 -25079 -17421 -25063
rect -17677 -25113 -17665 -25079
rect -17433 -25113 -17421 -25079
rect -17677 -25129 -17421 -25113
rect -17677 -25175 -17421 -25159
rect -17677 -25209 -17665 -25175
rect -17433 -25209 -17421 -25175
rect -17677 -25225 -17421 -25209
rect -12314 -25225 -11764 -25213
rect -17677 -25271 -17421 -25255
rect -12314 -25259 -12302 -25225
rect -11776 -25259 -11764 -25225
rect -12314 -25271 -11764 -25259
rect -17677 -25305 -17665 -25271
rect -17433 -25305 -17421 -25271
rect -17677 -25317 -17421 -25305
rect -12314 -25313 -11764 -25301
rect -12314 -25347 -12302 -25313
rect -11776 -25347 -11764 -25313
rect -12314 -25363 -11764 -25347
rect -12314 -25409 -11764 -25393
rect -12314 -25443 -12302 -25409
rect -11776 -25443 -11764 -25409
rect -12314 -25459 -11764 -25443
rect -12314 -25505 -11764 -25489
rect -12314 -25539 -12302 -25505
rect -11776 -25539 -11764 -25505
rect -12314 -25555 -11764 -25539
rect -12314 -25601 -11764 -25585
rect -12314 -25635 -12302 -25601
rect -11776 -25635 -11764 -25601
rect -12314 -25651 -11764 -25635
rect -12314 -25697 -11764 -25681
rect -12314 -25731 -12302 -25697
rect -11776 -25731 -11764 -25697
rect -12314 -25747 -11764 -25731
rect -12314 -25793 -11764 -25777
rect -12314 -25827 -12302 -25793
rect -11776 -25827 -11764 -25793
rect -12314 -25843 -11764 -25827
rect -12314 -25889 -11764 -25873
rect -12314 -25923 -12302 -25889
rect -11776 -25923 -11764 -25889
rect -12314 -25939 -11764 -25923
rect -12314 -25985 -11764 -25969
rect -12314 -26019 -12302 -25985
rect -11776 -26019 -11764 -25985
rect -12314 -26035 -11764 -26019
rect -12314 -26081 -11764 -26065
rect -12314 -26115 -12302 -26081
rect -11776 -26115 -11764 -26081
rect -12314 -26131 -11764 -26115
rect -12314 -26177 -11764 -26161
rect -12314 -26211 -12302 -26177
rect -11776 -26211 -11764 -26177
rect -12314 -26227 -11764 -26211
rect -12314 -26273 -11764 -26257
rect -12314 -26307 -12302 -26273
rect -11776 -26307 -11764 -26273
rect -12314 -26323 -11764 -26307
rect -12314 -26369 -11764 -26353
rect -12314 -26403 -12302 -26369
rect -11776 -26403 -11764 -26369
rect -12314 -26419 -11764 -26403
rect -12314 -26465 -11764 -26449
rect -12314 -26499 -12302 -26465
rect -11776 -26499 -11764 -26465
rect -12314 -26511 -11764 -26499
rect 11773 -25171 11835 -25159
rect 11773 -25403 11785 -25171
rect 11819 -25403 11835 -25171
rect 11773 -25415 11835 -25403
rect 11865 -25171 11931 -25159
rect 11865 -25403 11881 -25171
rect 11915 -25403 11931 -25171
rect 11865 -25415 11931 -25403
rect 11961 -25171 12027 -25159
rect 11961 -25403 11977 -25171
rect 12011 -25403 12027 -25171
rect 11961 -25415 12027 -25403
rect 12057 -25171 12123 -25159
rect 12057 -25403 12073 -25171
rect 12107 -25403 12123 -25171
rect 12057 -25415 12123 -25403
rect 12153 -25171 12219 -25159
rect 12153 -25403 12169 -25171
rect 12203 -25403 12219 -25171
rect 12153 -25415 12219 -25403
rect 12249 -25171 12315 -25159
rect 12249 -25403 12265 -25171
rect 12299 -25403 12315 -25171
rect 12249 -25415 12315 -25403
rect 12345 -25171 12411 -25159
rect 12345 -25403 12361 -25171
rect 12395 -25403 12411 -25171
rect 12345 -25415 12411 -25403
rect 12441 -25171 12507 -25159
rect 12441 -25403 12457 -25171
rect 12491 -25403 12507 -25171
rect 12441 -25415 12507 -25403
rect 12537 -25171 12603 -25159
rect 12537 -25403 12553 -25171
rect 12587 -25403 12603 -25171
rect 12537 -25415 12603 -25403
rect 12633 -25171 12699 -25159
rect 12633 -25403 12649 -25171
rect 12683 -25403 12699 -25171
rect 12633 -25415 12699 -25403
rect 12729 -25171 12791 -25159
rect 12729 -25403 12745 -25171
rect 12779 -25403 12791 -25171
rect 12923 -25275 13137 -25263
rect 12729 -25415 12791 -25403
rect -12314 -26553 -11764 -26541
rect -12314 -26587 -12302 -26553
rect -11776 -26587 -11764 -26553
rect -12314 -26599 -11764 -26587
rect 12923 -25309 12935 -25275
rect 13125 -25309 13137 -25275
rect 12923 -25325 13137 -25309
rect 12923 -25371 13137 -25355
rect 12923 -25405 12935 -25371
rect 13129 -25405 13137 -25371
rect 12923 -25421 13137 -25405
rect 12923 -25467 13137 -25451
rect 12923 -25501 12935 -25467
rect 13125 -25501 13137 -25467
rect 12923 -25517 13137 -25501
rect 12923 -25563 13137 -25547
rect 12923 -25597 12935 -25563
rect 13129 -25597 13137 -25563
rect 12923 -25609 13137 -25597
rect 7138 -26825 7200 -26813
rect 7138 -27123 7150 -26825
rect 7184 -27123 7200 -26825
rect 7138 -27135 7200 -27123
rect 7230 -26825 7296 -26813
rect 7230 -27123 7246 -26825
rect 7280 -27123 7296 -26825
rect 7230 -27135 7296 -27123
rect 7326 -26825 7392 -26813
rect 7326 -27123 7342 -26825
rect 7376 -27123 7392 -26825
rect 7326 -27135 7392 -27123
rect 7422 -26825 7488 -26813
rect 7422 -27123 7438 -26825
rect 7472 -27123 7488 -26825
rect 7422 -27135 7488 -27123
rect 7518 -26825 7584 -26813
rect 7518 -27123 7534 -26825
rect 7568 -27123 7584 -26825
rect 7518 -27135 7584 -27123
rect 7614 -26825 7680 -26813
rect 7614 -27123 7630 -26825
rect 7664 -27123 7680 -26825
rect 7614 -27135 7680 -27123
rect 7710 -26825 7776 -26813
rect 7710 -27123 7726 -26825
rect 7760 -27123 7776 -26825
rect 7710 -27135 7776 -27123
rect 7806 -26825 7872 -26813
rect 7806 -27123 7822 -26825
rect 7856 -27123 7872 -26825
rect 7806 -27135 7872 -27123
rect 7902 -26825 7964 -26813
rect 7902 -27123 7918 -26825
rect 7952 -27123 7964 -26825
rect 7902 -27135 7964 -27123
rect 8086 -26825 8148 -26813
rect 8086 -27123 8098 -26825
rect 8132 -27123 8148 -26825
rect 8086 -27135 8148 -27123
rect 8178 -26825 8244 -26813
rect 8178 -27123 8194 -26825
rect 8228 -27123 8244 -26825
rect 8178 -27135 8244 -27123
rect 8274 -26825 8340 -26813
rect 8274 -27123 8290 -26825
rect 8324 -27123 8340 -26825
rect 8274 -27135 8340 -27123
rect 8370 -26825 8436 -26813
rect 8370 -27123 8386 -26825
rect 8420 -27123 8436 -26825
rect 8370 -27135 8436 -27123
rect 8466 -26825 8532 -26813
rect 8466 -27123 8482 -26825
rect 8516 -27123 8532 -26825
rect 8466 -27135 8532 -27123
rect 8562 -26825 8628 -26813
rect 8562 -27123 8578 -26825
rect 8612 -27123 8628 -26825
rect 8562 -27135 8628 -27123
rect 8658 -26825 8724 -26813
rect 8658 -27123 8674 -26825
rect 8708 -27123 8724 -26825
rect 8658 -27135 8724 -27123
rect 8754 -26825 8820 -26813
rect 8754 -27123 8770 -26825
rect 8804 -27123 8820 -26825
rect 8754 -27135 8820 -27123
rect 8850 -26825 8912 -26813
rect 8850 -27123 8866 -26825
rect 8900 -27123 8912 -26825
rect 8850 -27135 8912 -27123
rect 9022 -26825 9084 -26813
rect 9022 -27123 9034 -26825
rect 9068 -27123 9084 -26825
rect 9022 -27135 9084 -27123
rect 9114 -26825 9180 -26813
rect 9114 -27123 9130 -26825
rect 9164 -27123 9180 -26825
rect 9114 -27135 9180 -27123
rect 9210 -26825 9276 -26813
rect 9210 -27123 9226 -26825
rect 9260 -27123 9276 -26825
rect 9210 -27135 9276 -27123
rect 9306 -26825 9372 -26813
rect 9306 -27123 9322 -26825
rect 9356 -27123 9372 -26825
rect 9306 -27135 9372 -27123
rect 9402 -26825 9468 -26813
rect 9402 -27123 9418 -26825
rect 9452 -27123 9468 -26825
rect 9402 -27135 9468 -27123
rect 9498 -26825 9564 -26813
rect 9498 -27123 9514 -26825
rect 9548 -27123 9564 -26825
rect 9498 -27135 9564 -27123
rect 9594 -26825 9660 -26813
rect 9594 -27123 9610 -26825
rect 9644 -27123 9660 -26825
rect 9594 -27135 9660 -27123
rect 9690 -26825 9756 -26813
rect 9690 -27123 9706 -26825
rect 9740 -27123 9756 -26825
rect 9690 -27135 9756 -27123
rect 9786 -26825 9848 -26813
rect 9786 -27123 9802 -26825
rect 9836 -27123 9848 -26825
rect 9786 -27135 9848 -27123
rect 9953 -26824 10015 -26812
rect 9953 -27122 9965 -26824
rect 9999 -27122 10015 -26824
rect 9953 -27134 10015 -27122
rect 10045 -26824 10111 -26812
rect 10045 -27122 10061 -26824
rect 10095 -27122 10111 -26824
rect 10045 -27134 10111 -27122
rect 10141 -26824 10207 -26812
rect 10141 -27122 10157 -26824
rect 10191 -27122 10207 -26824
rect 10141 -27134 10207 -27122
rect 10237 -26824 10303 -26812
rect 10237 -27122 10253 -26824
rect 10287 -27122 10303 -26824
rect 10237 -27134 10303 -27122
rect 10333 -26824 10399 -26812
rect 10333 -27122 10349 -26824
rect 10383 -27122 10399 -26824
rect 10333 -27134 10399 -27122
rect 10429 -26824 10495 -26812
rect 10429 -27122 10445 -26824
rect 10479 -27122 10495 -26824
rect 10429 -27134 10495 -27122
rect 10525 -26824 10591 -26812
rect 10525 -27122 10541 -26824
rect 10575 -27122 10591 -26824
rect 10525 -27134 10591 -27122
rect 10621 -26824 10687 -26812
rect 10621 -27122 10637 -26824
rect 10671 -27122 10687 -26824
rect 10621 -27134 10687 -27122
rect 10717 -26824 10779 -26812
rect 10717 -27122 10733 -26824
rect 10767 -27122 10779 -26824
rect 10717 -27134 10779 -27122
rect 10880 -26825 10942 -26813
rect 10880 -27123 10892 -26825
rect 10926 -27123 10942 -26825
rect 10880 -27135 10942 -27123
rect 10972 -26825 11038 -26813
rect 10972 -27123 10988 -26825
rect 11022 -27123 11038 -26825
rect 10972 -27135 11038 -27123
rect 11068 -26825 11134 -26813
rect 11068 -27123 11084 -26825
rect 11118 -27123 11134 -26825
rect 11068 -27135 11134 -27123
rect 11164 -26825 11230 -26813
rect 11164 -27123 11180 -26825
rect 11214 -27123 11230 -26825
rect 11164 -27135 11230 -27123
rect 11260 -26825 11326 -26813
rect 11260 -27123 11276 -26825
rect 11310 -27123 11326 -26825
rect 11260 -27135 11326 -27123
rect 11356 -26825 11422 -26813
rect 11356 -27123 11372 -26825
rect 11406 -27123 11422 -26825
rect 11356 -27135 11422 -27123
rect 11452 -26825 11518 -26813
rect 11452 -27123 11468 -26825
rect 11502 -27123 11518 -26825
rect 11452 -27135 11518 -27123
rect 11548 -26825 11614 -26813
rect 11548 -27123 11564 -26825
rect 11598 -27123 11614 -26825
rect 11548 -27135 11614 -27123
rect 11644 -26825 11706 -26813
rect 11644 -27123 11660 -26825
rect 11694 -27123 11706 -26825
rect 11644 -27135 11706 -27123
rect 5658 -27785 5872 -27773
rect -12314 -27858 -11764 -27846
rect -12314 -27892 -12302 -27858
rect -11776 -27892 -11764 -27858
rect -12314 -27904 -11764 -27892
rect -12314 -27946 -11764 -27934
rect -12314 -27980 -12302 -27946
rect -11776 -27980 -11764 -27946
rect -12314 -27996 -11764 -27980
rect -12314 -28042 -11764 -28026
rect -12314 -28076 -12302 -28042
rect -11776 -28076 -11764 -28042
rect -12314 -28092 -11764 -28076
rect -12314 -28138 -11764 -28122
rect -12314 -28172 -12302 -28138
rect -11776 -28172 -11764 -28138
rect -12314 -28188 -11764 -28172
rect -12314 -28234 -11764 -28218
rect -12314 -28268 -12302 -28234
rect -11776 -28268 -11764 -28234
rect -12314 -28284 -11764 -28268
rect -12314 -28330 -11764 -28314
rect -12314 -28364 -12302 -28330
rect -11776 -28364 -11764 -28330
rect -12314 -28380 -11764 -28364
rect -12314 -28426 -11764 -28410
rect -12314 -28460 -12302 -28426
rect -11776 -28460 -11764 -28426
rect -12314 -28476 -11764 -28460
rect -12314 -28522 -11764 -28506
rect -12314 -28556 -12302 -28522
rect -11776 -28556 -11764 -28522
rect -12314 -28572 -11764 -28556
rect -12314 -28618 -11764 -28602
rect -12314 -28652 -12302 -28618
rect -11776 -28652 -11764 -28618
rect -12314 -28668 -11764 -28652
rect -12314 -28714 -11764 -28698
rect -12314 -28748 -12302 -28714
rect -11776 -28748 -11764 -28714
rect -12314 -28764 -11764 -28748
rect -12314 -28810 -11764 -28794
rect -12314 -28844 -12302 -28810
rect -11776 -28844 -11764 -28810
rect -12314 -28860 -11764 -28844
rect -12314 -28906 -11764 -28890
rect -12314 -28940 -12302 -28906
rect -11776 -28940 -11764 -28906
rect -12314 -28956 -11764 -28940
rect -12314 -29002 -11764 -28986
rect -12314 -29036 -12302 -29002
rect -11776 -29036 -11764 -29002
rect -12314 -29052 -11764 -29036
rect -12314 -29098 -11764 -29082
rect -12314 -29132 -12302 -29098
rect -11776 -29132 -11764 -29098
rect -12314 -29144 -11764 -29132
rect 5658 -27819 5670 -27785
rect 5860 -27819 5872 -27785
rect 6098 -27785 6312 -27773
rect 5658 -27835 5872 -27819
rect 5658 -27881 5872 -27865
rect 5658 -27915 5670 -27881
rect 5864 -27915 5872 -27881
rect 5658 -27931 5872 -27915
rect 5658 -27977 5872 -27961
rect 5658 -28011 5670 -27977
rect 5860 -28011 5872 -27977
rect 5658 -28027 5872 -28011
rect 5658 -28073 5872 -28057
rect 5658 -28107 5670 -28073
rect 5864 -28107 5872 -28073
rect 6098 -27819 6110 -27785
rect 6300 -27819 6312 -27785
rect 6538 -27785 6752 -27773
rect 6098 -27835 6312 -27819
rect 6098 -27881 6312 -27865
rect 6098 -27915 6110 -27881
rect 6304 -27915 6312 -27881
rect 6098 -27931 6312 -27915
rect 6098 -27977 6312 -27961
rect 6098 -28011 6110 -27977
rect 6300 -28011 6312 -27977
rect 6098 -28027 6312 -28011
rect 6098 -28073 6312 -28057
rect 5658 -28119 5872 -28107
rect 6098 -28107 6110 -28073
rect 6304 -28107 6312 -28073
rect 6538 -27819 6550 -27785
rect 6740 -27819 6752 -27785
rect 6538 -27835 6752 -27819
rect 6538 -27881 6752 -27865
rect 6538 -27915 6550 -27881
rect 6744 -27915 6752 -27881
rect 6538 -27931 6752 -27915
rect 6538 -27977 6752 -27961
rect 6538 -28011 6550 -27977
rect 6740 -28011 6752 -27977
rect 6538 -28027 6752 -28011
rect 6538 -28073 6752 -28057
rect 6098 -28119 6312 -28107
rect 6538 -28107 6550 -28073
rect 6744 -28107 6752 -28073
rect 6538 -28119 6752 -28107
rect 7138 -28489 7200 -28477
rect 7138 -28787 7150 -28489
rect 7184 -28787 7200 -28489
rect 7138 -28799 7200 -28787
rect 7230 -28489 7296 -28477
rect 7230 -28787 7246 -28489
rect 7280 -28787 7296 -28489
rect 7230 -28799 7296 -28787
rect 7326 -28489 7392 -28477
rect 7326 -28787 7342 -28489
rect 7376 -28787 7392 -28489
rect 7326 -28799 7392 -28787
rect 7422 -28489 7488 -28477
rect 7422 -28787 7438 -28489
rect 7472 -28787 7488 -28489
rect 7422 -28799 7488 -28787
rect 7518 -28489 7584 -28477
rect 7518 -28787 7534 -28489
rect 7568 -28787 7584 -28489
rect 7518 -28799 7584 -28787
rect 7614 -28489 7680 -28477
rect 7614 -28787 7630 -28489
rect 7664 -28787 7680 -28489
rect 7614 -28799 7680 -28787
rect 7710 -28489 7776 -28477
rect 7710 -28787 7726 -28489
rect 7760 -28787 7776 -28489
rect 7710 -28799 7776 -28787
rect 7806 -28489 7872 -28477
rect 7806 -28787 7822 -28489
rect 7856 -28787 7872 -28489
rect 7806 -28799 7872 -28787
rect 7902 -28489 7964 -28477
rect 7902 -28787 7918 -28489
rect 7952 -28787 7964 -28489
rect 7902 -28799 7964 -28787
rect 8086 -28489 8148 -28477
rect 8086 -28787 8098 -28489
rect 8132 -28787 8148 -28489
rect 8086 -28799 8148 -28787
rect 8178 -28489 8244 -28477
rect 8178 -28787 8194 -28489
rect 8228 -28787 8244 -28489
rect 8178 -28799 8244 -28787
rect 8274 -28489 8340 -28477
rect 8274 -28787 8290 -28489
rect 8324 -28787 8340 -28489
rect 8274 -28799 8340 -28787
rect 8370 -28489 8436 -28477
rect 8370 -28787 8386 -28489
rect 8420 -28787 8436 -28489
rect 8370 -28799 8436 -28787
rect 8466 -28489 8532 -28477
rect 8466 -28787 8482 -28489
rect 8516 -28787 8532 -28489
rect 8466 -28799 8532 -28787
rect 8562 -28489 8628 -28477
rect 8562 -28787 8578 -28489
rect 8612 -28787 8628 -28489
rect 8562 -28799 8628 -28787
rect 8658 -28489 8724 -28477
rect 8658 -28787 8674 -28489
rect 8708 -28787 8724 -28489
rect 8658 -28799 8724 -28787
rect 8754 -28489 8820 -28477
rect 8754 -28787 8770 -28489
rect 8804 -28787 8820 -28489
rect 8754 -28799 8820 -28787
rect 8850 -28489 8912 -28477
rect 8850 -28787 8866 -28489
rect 8900 -28787 8912 -28489
rect 8850 -28799 8912 -28787
rect 9022 -28489 9084 -28477
rect 9022 -28787 9034 -28489
rect 9068 -28787 9084 -28489
rect 9022 -28799 9084 -28787
rect 9114 -28489 9180 -28477
rect 9114 -28787 9130 -28489
rect 9164 -28787 9180 -28489
rect 9114 -28799 9180 -28787
rect 9210 -28489 9276 -28477
rect 9210 -28787 9226 -28489
rect 9260 -28787 9276 -28489
rect 9210 -28799 9276 -28787
rect 9306 -28489 9372 -28477
rect 9306 -28787 9322 -28489
rect 9356 -28787 9372 -28489
rect 9306 -28799 9372 -28787
rect 9402 -28489 9468 -28477
rect 9402 -28787 9418 -28489
rect 9452 -28787 9468 -28489
rect 9402 -28799 9468 -28787
rect 9498 -28489 9564 -28477
rect 9498 -28787 9514 -28489
rect 9548 -28787 9564 -28489
rect 9498 -28799 9564 -28787
rect 9594 -28489 9660 -28477
rect 9594 -28787 9610 -28489
rect 9644 -28787 9660 -28489
rect 9594 -28799 9660 -28787
rect 9690 -28489 9756 -28477
rect 9690 -28787 9706 -28489
rect 9740 -28787 9756 -28489
rect 9690 -28799 9756 -28787
rect 9786 -28489 9848 -28477
rect 9786 -28787 9802 -28489
rect 9836 -28787 9848 -28489
rect 9786 -28799 9848 -28787
rect 9953 -28489 10015 -28477
rect 9953 -28787 9965 -28489
rect 9999 -28787 10015 -28489
rect 9953 -28799 10015 -28787
rect 10045 -28489 10111 -28477
rect 10045 -28787 10061 -28489
rect 10095 -28787 10111 -28489
rect 10045 -28799 10111 -28787
rect 10141 -28489 10207 -28477
rect 10141 -28787 10157 -28489
rect 10191 -28787 10207 -28489
rect 10141 -28799 10207 -28787
rect 10237 -28489 10303 -28477
rect 10237 -28787 10253 -28489
rect 10287 -28787 10303 -28489
rect 10237 -28799 10303 -28787
rect 10333 -28489 10399 -28477
rect 10333 -28787 10349 -28489
rect 10383 -28787 10399 -28489
rect 10333 -28799 10399 -28787
rect 10429 -28489 10495 -28477
rect 10429 -28787 10445 -28489
rect 10479 -28787 10495 -28489
rect 10429 -28799 10495 -28787
rect 10525 -28489 10591 -28477
rect 10525 -28787 10541 -28489
rect 10575 -28787 10591 -28489
rect 10525 -28799 10591 -28787
rect 10621 -28489 10687 -28477
rect 10621 -28787 10637 -28489
rect 10671 -28787 10687 -28489
rect 10621 -28799 10687 -28787
rect 10717 -28489 10779 -28477
rect 10717 -28787 10733 -28489
rect 10767 -28787 10779 -28489
rect 10717 -28799 10779 -28787
rect 10880 -28489 10942 -28477
rect 10880 -28787 10892 -28489
rect 10926 -28787 10942 -28489
rect 10880 -28799 10942 -28787
rect 10972 -28489 11038 -28477
rect 10972 -28787 10988 -28489
rect 11022 -28787 11038 -28489
rect 10972 -28799 11038 -28787
rect 11068 -28489 11134 -28477
rect 11068 -28787 11084 -28489
rect 11118 -28787 11134 -28489
rect 11068 -28799 11134 -28787
rect 11164 -28489 11230 -28477
rect 11164 -28787 11180 -28489
rect 11214 -28787 11230 -28489
rect 11164 -28799 11230 -28787
rect 11260 -28489 11326 -28477
rect 11260 -28787 11276 -28489
rect 11310 -28787 11326 -28489
rect 11260 -28799 11326 -28787
rect 11356 -28489 11422 -28477
rect 11356 -28787 11372 -28489
rect 11406 -28787 11422 -28489
rect 11356 -28799 11422 -28787
rect 11452 -28489 11518 -28477
rect 11452 -28787 11468 -28489
rect 11502 -28787 11518 -28489
rect 11452 -28799 11518 -28787
rect 11548 -28489 11614 -28477
rect 11548 -28787 11564 -28489
rect 11598 -28787 11614 -28489
rect 11548 -28799 11614 -28787
rect 11644 -28489 11706 -28477
rect 11644 -28787 11660 -28489
rect 11694 -28787 11706 -28489
rect 11644 -28799 11706 -28787
rect -12314 -29186 -11764 -29174
rect -12314 -29220 -12302 -29186
rect -11776 -29220 -11764 -29186
rect -12314 -29232 -11764 -29220
rect 11773 -29699 11835 -29687
rect 11773 -29931 11785 -29699
rect 11819 -29931 11835 -29699
rect 11773 -29943 11835 -29931
rect 11865 -29699 11931 -29687
rect 11865 -29931 11881 -29699
rect 11915 -29931 11931 -29699
rect 11865 -29943 11931 -29931
rect 11961 -29699 12027 -29687
rect 11961 -29931 11977 -29699
rect 12011 -29931 12027 -29699
rect 11961 -29943 12027 -29931
rect 12057 -29699 12123 -29687
rect 12057 -29931 12073 -29699
rect 12107 -29931 12123 -29699
rect 12057 -29943 12123 -29931
rect 12153 -29699 12219 -29687
rect 12153 -29931 12169 -29699
rect 12203 -29931 12219 -29699
rect 12153 -29943 12219 -29931
rect 12249 -29699 12315 -29687
rect 12249 -29931 12265 -29699
rect 12299 -29931 12315 -29699
rect 12249 -29943 12315 -29931
rect 12345 -29699 12411 -29687
rect 12345 -29931 12361 -29699
rect 12395 -29931 12411 -29699
rect 12345 -29943 12411 -29931
rect 12441 -29699 12507 -29687
rect 12441 -29931 12457 -29699
rect 12491 -29931 12507 -29699
rect 12441 -29943 12507 -29931
rect 12537 -29699 12603 -29687
rect 12537 -29931 12553 -29699
rect 12587 -29931 12603 -29699
rect 12537 -29943 12603 -29931
rect 12633 -29699 12699 -29687
rect 12633 -29931 12649 -29699
rect 12683 -29931 12699 -29699
rect 12633 -29943 12699 -29931
rect 12729 -29699 12791 -29687
rect 12729 -29931 12745 -29699
rect 12779 -29931 12791 -29699
rect 12923 -29803 13137 -29791
rect 12729 -29943 12791 -29931
rect -12314 -30467 -11764 -30455
rect -12314 -30501 -12302 -30467
rect -11776 -30501 -11764 -30467
rect -12314 -30513 -11764 -30501
rect -12314 -30555 -11764 -30543
rect -12314 -30589 -12302 -30555
rect -11776 -30589 -11764 -30555
rect -12314 -30605 -11764 -30589
rect -12314 -30651 -11764 -30635
rect -12314 -30685 -12302 -30651
rect -11776 -30685 -11764 -30651
rect -12314 -30701 -11764 -30685
rect -12314 -30747 -11764 -30731
rect -12314 -30781 -12302 -30747
rect -11776 -30781 -11764 -30747
rect -12314 -30797 -11764 -30781
rect -12314 -30843 -11764 -30827
rect -12314 -30877 -12302 -30843
rect -11776 -30877 -11764 -30843
rect -12314 -30893 -11764 -30877
rect -12314 -30939 -11764 -30923
rect -12314 -30973 -12302 -30939
rect -11776 -30973 -11764 -30939
rect -12314 -30989 -11764 -30973
rect -12314 -31035 -11764 -31019
rect -12314 -31069 -12302 -31035
rect -11776 -31069 -11764 -31035
rect -12314 -31085 -11764 -31069
rect -12314 -31131 -11764 -31115
rect -12314 -31165 -12302 -31131
rect -11776 -31165 -11764 -31131
rect -12314 -31181 -11764 -31165
rect -12314 -31227 -11764 -31211
rect -12314 -31261 -12302 -31227
rect -11776 -31261 -11764 -31227
rect -12314 -31277 -11764 -31261
rect -12314 -31323 -11764 -31307
rect -12314 -31357 -12302 -31323
rect -11776 -31357 -11764 -31323
rect -12314 -31373 -11764 -31357
rect -12314 -31419 -11764 -31403
rect -12314 -31453 -12302 -31419
rect -11776 -31453 -11764 -31419
rect -12314 -31469 -11764 -31453
rect -12314 -31515 -11764 -31499
rect -12314 -31549 -12302 -31515
rect -11776 -31549 -11764 -31515
rect -12314 -31565 -11764 -31549
rect -12314 -31611 -11764 -31595
rect -12314 -31645 -12302 -31611
rect -11776 -31645 -11764 -31611
rect -12314 -31661 -11764 -31645
rect -12314 -31707 -11764 -31691
rect -12314 -31741 -12302 -31707
rect -11776 -31741 -11764 -31707
rect -12314 -31753 -11764 -31741
rect 12923 -29837 12935 -29803
rect 13125 -29837 13137 -29803
rect 12923 -29853 13137 -29837
rect 12923 -29899 13137 -29883
rect 12923 -29933 12935 -29899
rect 13129 -29933 13137 -29899
rect 12923 -29949 13137 -29933
rect 12923 -29995 13137 -29979
rect 12923 -30029 12935 -29995
rect 13125 -30029 13137 -29995
rect 12923 -30045 13137 -30029
rect 12923 -30091 13137 -30075
rect 12923 -30125 12935 -30091
rect 13129 -30125 13137 -30091
rect 12923 -30137 13137 -30125
rect 7138 -31353 7200 -31341
rect 7138 -31651 7150 -31353
rect 7184 -31651 7200 -31353
rect 7138 -31663 7200 -31651
rect 7230 -31353 7296 -31341
rect 7230 -31651 7246 -31353
rect 7280 -31651 7296 -31353
rect 7230 -31663 7296 -31651
rect 7326 -31353 7392 -31341
rect 7326 -31651 7342 -31353
rect 7376 -31651 7392 -31353
rect 7326 -31663 7392 -31651
rect 7422 -31353 7488 -31341
rect 7422 -31651 7438 -31353
rect 7472 -31651 7488 -31353
rect 7422 -31663 7488 -31651
rect 7518 -31353 7584 -31341
rect 7518 -31651 7534 -31353
rect 7568 -31651 7584 -31353
rect 7518 -31663 7584 -31651
rect 7614 -31353 7680 -31341
rect 7614 -31651 7630 -31353
rect 7664 -31651 7680 -31353
rect 7614 -31663 7680 -31651
rect 7710 -31353 7776 -31341
rect 7710 -31651 7726 -31353
rect 7760 -31651 7776 -31353
rect 7710 -31663 7776 -31651
rect 7806 -31353 7872 -31341
rect 7806 -31651 7822 -31353
rect 7856 -31651 7872 -31353
rect 7806 -31663 7872 -31651
rect 7902 -31353 7964 -31341
rect 7902 -31651 7918 -31353
rect 7952 -31651 7964 -31353
rect 7902 -31663 7964 -31651
rect 8086 -31353 8148 -31341
rect 8086 -31651 8098 -31353
rect 8132 -31651 8148 -31353
rect 8086 -31663 8148 -31651
rect 8178 -31353 8244 -31341
rect 8178 -31651 8194 -31353
rect 8228 -31651 8244 -31353
rect 8178 -31663 8244 -31651
rect 8274 -31353 8340 -31341
rect 8274 -31651 8290 -31353
rect 8324 -31651 8340 -31353
rect 8274 -31663 8340 -31651
rect 8370 -31353 8436 -31341
rect 8370 -31651 8386 -31353
rect 8420 -31651 8436 -31353
rect 8370 -31663 8436 -31651
rect 8466 -31353 8532 -31341
rect 8466 -31651 8482 -31353
rect 8516 -31651 8532 -31353
rect 8466 -31663 8532 -31651
rect 8562 -31353 8628 -31341
rect 8562 -31651 8578 -31353
rect 8612 -31651 8628 -31353
rect 8562 -31663 8628 -31651
rect 8658 -31353 8724 -31341
rect 8658 -31651 8674 -31353
rect 8708 -31651 8724 -31353
rect 8658 -31663 8724 -31651
rect 8754 -31353 8820 -31341
rect 8754 -31651 8770 -31353
rect 8804 -31651 8820 -31353
rect 8754 -31663 8820 -31651
rect 8850 -31353 8912 -31341
rect 8850 -31651 8866 -31353
rect 8900 -31651 8912 -31353
rect 8850 -31663 8912 -31651
rect 9022 -31353 9084 -31341
rect 9022 -31651 9034 -31353
rect 9068 -31651 9084 -31353
rect 9022 -31663 9084 -31651
rect 9114 -31353 9180 -31341
rect 9114 -31651 9130 -31353
rect 9164 -31651 9180 -31353
rect 9114 -31663 9180 -31651
rect 9210 -31353 9276 -31341
rect 9210 -31651 9226 -31353
rect 9260 -31651 9276 -31353
rect 9210 -31663 9276 -31651
rect 9306 -31353 9372 -31341
rect 9306 -31651 9322 -31353
rect 9356 -31651 9372 -31353
rect 9306 -31663 9372 -31651
rect 9402 -31353 9468 -31341
rect 9402 -31651 9418 -31353
rect 9452 -31651 9468 -31353
rect 9402 -31663 9468 -31651
rect 9498 -31353 9564 -31341
rect 9498 -31651 9514 -31353
rect 9548 -31651 9564 -31353
rect 9498 -31663 9564 -31651
rect 9594 -31353 9660 -31341
rect 9594 -31651 9610 -31353
rect 9644 -31651 9660 -31353
rect 9594 -31663 9660 -31651
rect 9690 -31353 9756 -31341
rect 9690 -31651 9706 -31353
rect 9740 -31651 9756 -31353
rect 9690 -31663 9756 -31651
rect 9786 -31353 9848 -31341
rect 9786 -31651 9802 -31353
rect 9836 -31651 9848 -31353
rect 9786 -31663 9848 -31651
rect 9953 -31352 10015 -31340
rect 9953 -31650 9965 -31352
rect 9999 -31650 10015 -31352
rect 9953 -31662 10015 -31650
rect 10045 -31352 10111 -31340
rect 10045 -31650 10061 -31352
rect 10095 -31650 10111 -31352
rect 10045 -31662 10111 -31650
rect 10141 -31352 10207 -31340
rect 10141 -31650 10157 -31352
rect 10191 -31650 10207 -31352
rect 10141 -31662 10207 -31650
rect 10237 -31352 10303 -31340
rect 10237 -31650 10253 -31352
rect 10287 -31650 10303 -31352
rect 10237 -31662 10303 -31650
rect 10333 -31352 10399 -31340
rect 10333 -31650 10349 -31352
rect 10383 -31650 10399 -31352
rect 10333 -31662 10399 -31650
rect 10429 -31352 10495 -31340
rect 10429 -31650 10445 -31352
rect 10479 -31650 10495 -31352
rect 10429 -31662 10495 -31650
rect 10525 -31352 10591 -31340
rect 10525 -31650 10541 -31352
rect 10575 -31650 10591 -31352
rect 10525 -31662 10591 -31650
rect 10621 -31352 10687 -31340
rect 10621 -31650 10637 -31352
rect 10671 -31650 10687 -31352
rect 10621 -31662 10687 -31650
rect 10717 -31352 10779 -31340
rect 10717 -31650 10733 -31352
rect 10767 -31650 10779 -31352
rect 10717 -31662 10779 -31650
rect 10880 -31353 10942 -31341
rect 10880 -31651 10892 -31353
rect 10926 -31651 10942 -31353
rect 10880 -31663 10942 -31651
rect 10972 -31353 11038 -31341
rect 10972 -31651 10988 -31353
rect 11022 -31651 11038 -31353
rect 10972 -31663 11038 -31651
rect 11068 -31353 11134 -31341
rect 11068 -31651 11084 -31353
rect 11118 -31651 11134 -31353
rect 11068 -31663 11134 -31651
rect 11164 -31353 11230 -31341
rect 11164 -31651 11180 -31353
rect 11214 -31651 11230 -31353
rect 11164 -31663 11230 -31651
rect 11260 -31353 11326 -31341
rect 11260 -31651 11276 -31353
rect 11310 -31651 11326 -31353
rect 11260 -31663 11326 -31651
rect 11356 -31353 11422 -31341
rect 11356 -31651 11372 -31353
rect 11406 -31651 11422 -31353
rect 11356 -31663 11422 -31651
rect 11452 -31353 11518 -31341
rect 11452 -31651 11468 -31353
rect 11502 -31651 11518 -31353
rect 11452 -31663 11518 -31651
rect 11548 -31353 11614 -31341
rect 11548 -31651 11564 -31353
rect 11598 -31651 11614 -31353
rect 11548 -31663 11614 -31651
rect 11644 -31353 11706 -31341
rect 11644 -31651 11660 -31353
rect 11694 -31651 11706 -31353
rect 11644 -31663 11706 -31651
rect -12314 -31795 -11764 -31783
rect -12314 -31829 -12302 -31795
rect -11776 -31829 -11764 -31795
rect -12314 -31841 -11764 -31829
rect 5658 -32313 5872 -32301
rect 5658 -32347 5670 -32313
rect 5860 -32347 5872 -32313
rect 6098 -32313 6312 -32301
rect 5658 -32363 5872 -32347
rect 5658 -32409 5872 -32393
rect 5658 -32443 5670 -32409
rect 5864 -32443 5872 -32409
rect 5658 -32459 5872 -32443
rect 5658 -32505 5872 -32489
rect 5658 -32539 5670 -32505
rect 5860 -32539 5872 -32505
rect 5658 -32555 5872 -32539
rect 5658 -32601 5872 -32585
rect 5658 -32635 5670 -32601
rect 5864 -32635 5872 -32601
rect 6098 -32347 6110 -32313
rect 6300 -32347 6312 -32313
rect 6538 -32313 6752 -32301
rect 6098 -32363 6312 -32347
rect 6098 -32409 6312 -32393
rect 6098 -32443 6110 -32409
rect 6304 -32443 6312 -32409
rect 6098 -32459 6312 -32443
rect 6098 -32505 6312 -32489
rect 6098 -32539 6110 -32505
rect 6300 -32539 6312 -32505
rect 6098 -32555 6312 -32539
rect 6098 -32601 6312 -32585
rect 5658 -32647 5872 -32635
rect 6098 -32635 6110 -32601
rect 6304 -32635 6312 -32601
rect 6538 -32347 6550 -32313
rect 6740 -32347 6752 -32313
rect 6538 -32363 6752 -32347
rect 6538 -32409 6752 -32393
rect 6538 -32443 6550 -32409
rect 6744 -32443 6752 -32409
rect 6538 -32459 6752 -32443
rect 6538 -32505 6752 -32489
rect 6538 -32539 6550 -32505
rect 6740 -32539 6752 -32505
rect 6538 -32555 6752 -32539
rect 6538 -32601 6752 -32585
rect 6098 -32647 6312 -32635
rect 6538 -32635 6550 -32601
rect 6744 -32635 6752 -32601
rect 6538 -32647 6752 -32635
rect 7138 -33017 7200 -33005
rect -12316 -33087 -11766 -33075
rect -12316 -33121 -12304 -33087
rect -11778 -33121 -11766 -33087
rect -12316 -33133 -11766 -33121
rect -12316 -33175 -11766 -33163
rect -12316 -33209 -12304 -33175
rect -11778 -33209 -11766 -33175
rect -12316 -33225 -11766 -33209
rect -12316 -33271 -11766 -33255
rect -12316 -33305 -12304 -33271
rect -11778 -33305 -11766 -33271
rect -12316 -33321 -11766 -33305
rect -12316 -33367 -11766 -33351
rect -12316 -33401 -12304 -33367
rect -11778 -33401 -11766 -33367
rect -12316 -33417 -11766 -33401
rect -12316 -33463 -11766 -33447
rect -12316 -33497 -12304 -33463
rect -11778 -33497 -11766 -33463
rect -12316 -33513 -11766 -33497
rect -12316 -33559 -11766 -33543
rect -12316 -33593 -12304 -33559
rect -11778 -33593 -11766 -33559
rect -12316 -33609 -11766 -33593
rect -12316 -33655 -11766 -33639
rect -12316 -33689 -12304 -33655
rect -11778 -33689 -11766 -33655
rect -12316 -33705 -11766 -33689
rect -12316 -33751 -11766 -33735
rect -12316 -33785 -12304 -33751
rect -11778 -33785 -11766 -33751
rect -12316 -33801 -11766 -33785
rect -12316 -33847 -11766 -33831
rect -12316 -33881 -12304 -33847
rect -11778 -33881 -11766 -33847
rect -12316 -33897 -11766 -33881
rect -12316 -33943 -11766 -33927
rect -12316 -33977 -12304 -33943
rect -11778 -33977 -11766 -33943
rect -12316 -33993 -11766 -33977
rect -12316 -34039 -11766 -34023
rect -12316 -34073 -12304 -34039
rect -11778 -34073 -11766 -34039
rect -12316 -34089 -11766 -34073
rect -12316 -34135 -11766 -34119
rect -12316 -34169 -12304 -34135
rect -11778 -34169 -11766 -34135
rect -12316 -34185 -11766 -34169
rect -12316 -34231 -11766 -34215
rect -12316 -34265 -12304 -34231
rect -11778 -34265 -11766 -34231
rect -12316 -34281 -11766 -34265
rect -12316 -34327 -11766 -34311
rect -12316 -34361 -12304 -34327
rect -11778 -34361 -11766 -34327
rect -12316 -34373 -11766 -34361
rect 7138 -33315 7150 -33017
rect 7184 -33315 7200 -33017
rect 7138 -33327 7200 -33315
rect 7230 -33017 7296 -33005
rect 7230 -33315 7246 -33017
rect 7280 -33315 7296 -33017
rect 7230 -33327 7296 -33315
rect 7326 -33017 7392 -33005
rect 7326 -33315 7342 -33017
rect 7376 -33315 7392 -33017
rect 7326 -33327 7392 -33315
rect 7422 -33017 7488 -33005
rect 7422 -33315 7438 -33017
rect 7472 -33315 7488 -33017
rect 7422 -33327 7488 -33315
rect 7518 -33017 7584 -33005
rect 7518 -33315 7534 -33017
rect 7568 -33315 7584 -33017
rect 7518 -33327 7584 -33315
rect 7614 -33017 7680 -33005
rect 7614 -33315 7630 -33017
rect 7664 -33315 7680 -33017
rect 7614 -33327 7680 -33315
rect 7710 -33017 7776 -33005
rect 7710 -33315 7726 -33017
rect 7760 -33315 7776 -33017
rect 7710 -33327 7776 -33315
rect 7806 -33017 7872 -33005
rect 7806 -33315 7822 -33017
rect 7856 -33315 7872 -33017
rect 7806 -33327 7872 -33315
rect 7902 -33017 7964 -33005
rect 7902 -33315 7918 -33017
rect 7952 -33315 7964 -33017
rect 7902 -33327 7964 -33315
rect 8086 -33017 8148 -33005
rect 8086 -33315 8098 -33017
rect 8132 -33315 8148 -33017
rect 8086 -33327 8148 -33315
rect 8178 -33017 8244 -33005
rect 8178 -33315 8194 -33017
rect 8228 -33315 8244 -33017
rect 8178 -33327 8244 -33315
rect 8274 -33017 8340 -33005
rect 8274 -33315 8290 -33017
rect 8324 -33315 8340 -33017
rect 8274 -33327 8340 -33315
rect 8370 -33017 8436 -33005
rect 8370 -33315 8386 -33017
rect 8420 -33315 8436 -33017
rect 8370 -33327 8436 -33315
rect 8466 -33017 8532 -33005
rect 8466 -33315 8482 -33017
rect 8516 -33315 8532 -33017
rect 8466 -33327 8532 -33315
rect 8562 -33017 8628 -33005
rect 8562 -33315 8578 -33017
rect 8612 -33315 8628 -33017
rect 8562 -33327 8628 -33315
rect 8658 -33017 8724 -33005
rect 8658 -33315 8674 -33017
rect 8708 -33315 8724 -33017
rect 8658 -33327 8724 -33315
rect 8754 -33017 8820 -33005
rect 8754 -33315 8770 -33017
rect 8804 -33315 8820 -33017
rect 8754 -33327 8820 -33315
rect 8850 -33017 8912 -33005
rect 8850 -33315 8866 -33017
rect 8900 -33315 8912 -33017
rect 8850 -33327 8912 -33315
rect 9022 -33017 9084 -33005
rect 9022 -33315 9034 -33017
rect 9068 -33315 9084 -33017
rect 9022 -33327 9084 -33315
rect 9114 -33017 9180 -33005
rect 9114 -33315 9130 -33017
rect 9164 -33315 9180 -33017
rect 9114 -33327 9180 -33315
rect 9210 -33017 9276 -33005
rect 9210 -33315 9226 -33017
rect 9260 -33315 9276 -33017
rect 9210 -33327 9276 -33315
rect 9306 -33017 9372 -33005
rect 9306 -33315 9322 -33017
rect 9356 -33315 9372 -33017
rect 9306 -33327 9372 -33315
rect 9402 -33017 9468 -33005
rect 9402 -33315 9418 -33017
rect 9452 -33315 9468 -33017
rect 9402 -33327 9468 -33315
rect 9498 -33017 9564 -33005
rect 9498 -33315 9514 -33017
rect 9548 -33315 9564 -33017
rect 9498 -33327 9564 -33315
rect 9594 -33017 9660 -33005
rect 9594 -33315 9610 -33017
rect 9644 -33315 9660 -33017
rect 9594 -33327 9660 -33315
rect 9690 -33017 9756 -33005
rect 9690 -33315 9706 -33017
rect 9740 -33315 9756 -33017
rect 9690 -33327 9756 -33315
rect 9786 -33017 9848 -33005
rect 9786 -33315 9802 -33017
rect 9836 -33315 9848 -33017
rect 9786 -33327 9848 -33315
rect 9953 -33017 10015 -33005
rect 9953 -33315 9965 -33017
rect 9999 -33315 10015 -33017
rect 9953 -33327 10015 -33315
rect 10045 -33017 10111 -33005
rect 10045 -33315 10061 -33017
rect 10095 -33315 10111 -33017
rect 10045 -33327 10111 -33315
rect 10141 -33017 10207 -33005
rect 10141 -33315 10157 -33017
rect 10191 -33315 10207 -33017
rect 10141 -33327 10207 -33315
rect 10237 -33017 10303 -33005
rect 10237 -33315 10253 -33017
rect 10287 -33315 10303 -33017
rect 10237 -33327 10303 -33315
rect 10333 -33017 10399 -33005
rect 10333 -33315 10349 -33017
rect 10383 -33315 10399 -33017
rect 10333 -33327 10399 -33315
rect 10429 -33017 10495 -33005
rect 10429 -33315 10445 -33017
rect 10479 -33315 10495 -33017
rect 10429 -33327 10495 -33315
rect 10525 -33017 10591 -33005
rect 10525 -33315 10541 -33017
rect 10575 -33315 10591 -33017
rect 10525 -33327 10591 -33315
rect 10621 -33017 10687 -33005
rect 10621 -33315 10637 -33017
rect 10671 -33315 10687 -33017
rect 10621 -33327 10687 -33315
rect 10717 -33017 10779 -33005
rect 10717 -33315 10733 -33017
rect 10767 -33315 10779 -33017
rect 10717 -33327 10779 -33315
rect 10880 -33017 10942 -33005
rect 10880 -33315 10892 -33017
rect 10926 -33315 10942 -33017
rect 10880 -33327 10942 -33315
rect 10972 -33017 11038 -33005
rect 10972 -33315 10988 -33017
rect 11022 -33315 11038 -33017
rect 10972 -33327 11038 -33315
rect 11068 -33017 11134 -33005
rect 11068 -33315 11084 -33017
rect 11118 -33315 11134 -33017
rect 11068 -33327 11134 -33315
rect 11164 -33017 11230 -33005
rect 11164 -33315 11180 -33017
rect 11214 -33315 11230 -33017
rect 11164 -33327 11230 -33315
rect 11260 -33017 11326 -33005
rect 11260 -33315 11276 -33017
rect 11310 -33315 11326 -33017
rect 11260 -33327 11326 -33315
rect 11356 -33017 11422 -33005
rect 11356 -33315 11372 -33017
rect 11406 -33315 11422 -33017
rect 11356 -33327 11422 -33315
rect 11452 -33017 11518 -33005
rect 11452 -33315 11468 -33017
rect 11502 -33315 11518 -33017
rect 11452 -33327 11518 -33315
rect 11548 -33017 11614 -33005
rect 11548 -33315 11564 -33017
rect 11598 -33315 11614 -33017
rect 11548 -33327 11614 -33315
rect 11644 -33017 11706 -33005
rect 11644 -33315 11660 -33017
rect 11694 -33315 11706 -33017
rect 11644 -33327 11706 -33315
rect -12316 -34415 -11766 -34403
rect -12316 -34449 -12304 -34415
rect -11778 -34449 -11766 -34415
rect -12316 -34461 -11766 -34449
rect 11773 -34227 11835 -34215
rect 11773 -34459 11785 -34227
rect 11819 -34459 11835 -34227
rect 11773 -34471 11835 -34459
rect 11865 -34227 11931 -34215
rect 11865 -34459 11881 -34227
rect 11915 -34459 11931 -34227
rect 11865 -34471 11931 -34459
rect 11961 -34227 12027 -34215
rect 11961 -34459 11977 -34227
rect 12011 -34459 12027 -34227
rect 11961 -34471 12027 -34459
rect 12057 -34227 12123 -34215
rect 12057 -34459 12073 -34227
rect 12107 -34459 12123 -34227
rect 12057 -34471 12123 -34459
rect 12153 -34227 12219 -34215
rect 12153 -34459 12169 -34227
rect 12203 -34459 12219 -34227
rect 12153 -34471 12219 -34459
rect 12249 -34227 12315 -34215
rect 12249 -34459 12265 -34227
rect 12299 -34459 12315 -34227
rect 12249 -34471 12315 -34459
rect 12345 -34227 12411 -34215
rect 12345 -34459 12361 -34227
rect 12395 -34459 12411 -34227
rect 12345 -34471 12411 -34459
rect 12441 -34227 12507 -34215
rect 12441 -34459 12457 -34227
rect 12491 -34459 12507 -34227
rect 12441 -34471 12507 -34459
rect 12537 -34227 12603 -34215
rect 12537 -34459 12553 -34227
rect 12587 -34459 12603 -34227
rect 12537 -34471 12603 -34459
rect 12633 -34227 12699 -34215
rect 12633 -34459 12649 -34227
rect 12683 -34459 12699 -34227
rect 12633 -34471 12699 -34459
rect 12729 -34227 12791 -34215
rect 12729 -34459 12745 -34227
rect 12779 -34459 12791 -34227
rect 12923 -34331 13137 -34319
rect 12729 -34471 12791 -34459
rect 12923 -34365 12935 -34331
rect 13125 -34365 13137 -34331
rect 12923 -34381 13137 -34365
rect 12923 -34427 13137 -34411
rect 12923 -34461 12935 -34427
rect 13129 -34461 13137 -34427
rect 12923 -34477 13137 -34461
rect 12923 -34523 13137 -34507
rect 12923 -34557 12935 -34523
rect 13125 -34557 13137 -34523
rect 12923 -34573 13137 -34557
rect 12923 -34619 13137 -34603
rect 12923 -34653 12935 -34619
rect 13129 -34653 13137 -34619
rect 12923 -34665 13137 -34653
rect 7138 -35881 7200 -35869
rect 7138 -36179 7150 -35881
rect 7184 -36179 7200 -35881
rect 7138 -36191 7200 -36179
rect 7230 -35881 7296 -35869
rect 7230 -36179 7246 -35881
rect 7280 -36179 7296 -35881
rect 7230 -36191 7296 -36179
rect 7326 -35881 7392 -35869
rect 7326 -36179 7342 -35881
rect 7376 -36179 7392 -35881
rect 7326 -36191 7392 -36179
rect 7422 -35881 7488 -35869
rect 7422 -36179 7438 -35881
rect 7472 -36179 7488 -35881
rect 7422 -36191 7488 -36179
rect 7518 -35881 7584 -35869
rect 7518 -36179 7534 -35881
rect 7568 -36179 7584 -35881
rect 7518 -36191 7584 -36179
rect 7614 -35881 7680 -35869
rect 7614 -36179 7630 -35881
rect 7664 -36179 7680 -35881
rect 7614 -36191 7680 -36179
rect 7710 -35881 7776 -35869
rect 7710 -36179 7726 -35881
rect 7760 -36179 7776 -35881
rect 7710 -36191 7776 -36179
rect 7806 -35881 7872 -35869
rect 7806 -36179 7822 -35881
rect 7856 -36179 7872 -35881
rect 7806 -36191 7872 -36179
rect 7902 -35881 7964 -35869
rect 7902 -36179 7918 -35881
rect 7952 -36179 7964 -35881
rect 7902 -36191 7964 -36179
rect 8086 -35881 8148 -35869
rect 8086 -36179 8098 -35881
rect 8132 -36179 8148 -35881
rect 8086 -36191 8148 -36179
rect 8178 -35881 8244 -35869
rect 8178 -36179 8194 -35881
rect 8228 -36179 8244 -35881
rect 8178 -36191 8244 -36179
rect 8274 -35881 8340 -35869
rect 8274 -36179 8290 -35881
rect 8324 -36179 8340 -35881
rect 8274 -36191 8340 -36179
rect 8370 -35881 8436 -35869
rect 8370 -36179 8386 -35881
rect 8420 -36179 8436 -35881
rect 8370 -36191 8436 -36179
rect 8466 -35881 8532 -35869
rect 8466 -36179 8482 -35881
rect 8516 -36179 8532 -35881
rect 8466 -36191 8532 -36179
rect 8562 -35881 8628 -35869
rect 8562 -36179 8578 -35881
rect 8612 -36179 8628 -35881
rect 8562 -36191 8628 -36179
rect 8658 -35881 8724 -35869
rect 8658 -36179 8674 -35881
rect 8708 -36179 8724 -35881
rect 8658 -36191 8724 -36179
rect 8754 -35881 8820 -35869
rect 8754 -36179 8770 -35881
rect 8804 -36179 8820 -35881
rect 8754 -36191 8820 -36179
rect 8850 -35881 8912 -35869
rect 8850 -36179 8866 -35881
rect 8900 -36179 8912 -35881
rect 8850 -36191 8912 -36179
rect 9022 -35881 9084 -35869
rect 9022 -36179 9034 -35881
rect 9068 -36179 9084 -35881
rect 9022 -36191 9084 -36179
rect 9114 -35881 9180 -35869
rect 9114 -36179 9130 -35881
rect 9164 -36179 9180 -35881
rect 9114 -36191 9180 -36179
rect 9210 -35881 9276 -35869
rect 9210 -36179 9226 -35881
rect 9260 -36179 9276 -35881
rect 9210 -36191 9276 -36179
rect 9306 -35881 9372 -35869
rect 9306 -36179 9322 -35881
rect 9356 -36179 9372 -35881
rect 9306 -36191 9372 -36179
rect 9402 -35881 9468 -35869
rect 9402 -36179 9418 -35881
rect 9452 -36179 9468 -35881
rect 9402 -36191 9468 -36179
rect 9498 -35881 9564 -35869
rect 9498 -36179 9514 -35881
rect 9548 -36179 9564 -35881
rect 9498 -36191 9564 -36179
rect 9594 -35881 9660 -35869
rect 9594 -36179 9610 -35881
rect 9644 -36179 9660 -35881
rect 9594 -36191 9660 -36179
rect 9690 -35881 9756 -35869
rect 9690 -36179 9706 -35881
rect 9740 -36179 9756 -35881
rect 9690 -36191 9756 -36179
rect 9786 -35881 9848 -35869
rect 9786 -36179 9802 -35881
rect 9836 -36179 9848 -35881
rect 9786 -36191 9848 -36179
rect 9953 -35880 10015 -35868
rect 9953 -36178 9965 -35880
rect 9999 -36178 10015 -35880
rect 9953 -36190 10015 -36178
rect 10045 -35880 10111 -35868
rect 10045 -36178 10061 -35880
rect 10095 -36178 10111 -35880
rect 10045 -36190 10111 -36178
rect 10141 -35880 10207 -35868
rect 10141 -36178 10157 -35880
rect 10191 -36178 10207 -35880
rect 10141 -36190 10207 -36178
rect 10237 -35880 10303 -35868
rect 10237 -36178 10253 -35880
rect 10287 -36178 10303 -35880
rect 10237 -36190 10303 -36178
rect 10333 -35880 10399 -35868
rect 10333 -36178 10349 -35880
rect 10383 -36178 10399 -35880
rect 10333 -36190 10399 -36178
rect 10429 -35880 10495 -35868
rect 10429 -36178 10445 -35880
rect 10479 -36178 10495 -35880
rect 10429 -36190 10495 -36178
rect 10525 -35880 10591 -35868
rect 10525 -36178 10541 -35880
rect 10575 -36178 10591 -35880
rect 10525 -36190 10591 -36178
rect 10621 -35880 10687 -35868
rect 10621 -36178 10637 -35880
rect 10671 -36178 10687 -35880
rect 10621 -36190 10687 -36178
rect 10717 -35880 10779 -35868
rect 10717 -36178 10733 -35880
rect 10767 -36178 10779 -35880
rect 10717 -36190 10779 -36178
rect 10880 -35881 10942 -35869
rect 10880 -36179 10892 -35881
rect 10926 -36179 10942 -35881
rect 10880 -36191 10942 -36179
rect 10972 -35881 11038 -35869
rect 10972 -36179 10988 -35881
rect 11022 -36179 11038 -35881
rect 10972 -36191 11038 -36179
rect 11068 -35881 11134 -35869
rect 11068 -36179 11084 -35881
rect 11118 -36179 11134 -35881
rect 11068 -36191 11134 -36179
rect 11164 -35881 11230 -35869
rect 11164 -36179 11180 -35881
rect 11214 -36179 11230 -35881
rect 11164 -36191 11230 -36179
rect 11260 -35881 11326 -35869
rect 11260 -36179 11276 -35881
rect 11310 -36179 11326 -35881
rect 11260 -36191 11326 -36179
rect 11356 -35881 11422 -35869
rect 11356 -36179 11372 -35881
rect 11406 -36179 11422 -35881
rect 11356 -36191 11422 -36179
rect 11452 -35881 11518 -35869
rect 11452 -36179 11468 -35881
rect 11502 -36179 11518 -35881
rect 11452 -36191 11518 -36179
rect 11548 -35881 11614 -35869
rect 11548 -36179 11564 -35881
rect 11598 -36179 11614 -35881
rect 11548 -36191 11614 -36179
rect 11644 -35881 11706 -35869
rect 11644 -36179 11660 -35881
rect 11694 -36179 11706 -35881
rect 13124 -35727 13186 -35715
rect 13124 -35921 13136 -35727
rect 13170 -35921 13186 -35727
rect 13124 -35929 13186 -35921
rect 13216 -35727 13282 -35715
rect 13216 -35917 13232 -35727
rect 13266 -35917 13282 -35727
rect 13216 -35929 13282 -35917
rect 13312 -35727 13378 -35715
rect 13312 -35921 13328 -35727
rect 13362 -35921 13378 -35727
rect 13312 -35929 13378 -35921
rect 13408 -35727 13470 -35715
rect 13408 -35917 13424 -35727
rect 13458 -35917 13470 -35727
rect 13408 -35929 13470 -35917
rect 11644 -36191 11706 -36179
rect 13124 -36106 13186 -36094
rect 13124 -36300 13136 -36106
rect 13170 -36300 13186 -36106
rect 13124 -36308 13186 -36300
rect 13216 -36106 13282 -36094
rect 13216 -36296 13232 -36106
rect 13266 -36296 13282 -36106
rect 13216 -36308 13282 -36296
rect 13312 -36106 13378 -36094
rect 13312 -36300 13328 -36106
rect 13362 -36300 13378 -36106
rect 13312 -36308 13378 -36300
rect 13408 -36106 13470 -36094
rect 13408 -36296 13424 -36106
rect 13458 -36296 13470 -36106
rect 13408 -36308 13470 -36296
<< ndiffc >>
rect 1719 4926 1753 5032
rect 1807 4926 1841 5032
rect 1903 4926 1937 5032
rect 1999 4926 2033 5032
rect 2095 4926 2129 5032
rect 2191 4926 2225 5032
rect 2287 4926 2321 5032
rect 2383 4926 2417 5032
rect 2479 4926 2513 5032
rect 2575 4926 2609 5032
rect 2671 4926 2705 5032
rect 2767 4926 2801 5032
rect 2863 4926 2897 5032
rect 2959 4926 2993 5032
rect 3047 4926 3081 5032
rect 3325 4926 3359 5032
rect 3413 4926 3447 5032
rect 3509 4926 3543 5032
rect 3605 4926 3639 5032
rect 3701 4926 3735 5032
rect 3797 4926 3831 5032
rect 3893 4926 3927 5032
rect 3989 4926 4023 5032
rect 4085 4926 4119 5032
rect 4181 4926 4215 5032
rect 4277 4926 4311 5032
rect 4373 4926 4407 5032
rect 4469 4926 4503 5032
rect 4565 4926 4599 5032
rect 4653 4926 4687 5032
rect 5029 4924 5063 5030
rect 5117 4924 5151 5030
rect 5213 4924 5247 5030
rect 5309 4924 5343 5030
rect 5405 4924 5439 5030
rect 5501 4924 5535 5030
rect 5597 4924 5631 5030
rect 5693 4924 5727 5030
rect 5789 4924 5823 5030
rect 5885 4924 5919 5030
rect 5981 4924 6015 5030
rect 6077 4924 6111 5030
rect 6173 4924 6207 5030
rect 6269 4924 6303 5030
rect 6357 4924 6391 5030
rect 7185 5051 7561 5085
rect 7821 4975 7997 5009
rect 7185 4859 7561 4893
rect 7821 4887 7997 4921
rect 5670 3427 5846 3461
rect 5670 3339 5846 3373
rect 6110 3427 6286 3461
rect 6110 3339 6286 3373
rect 6550 3427 6726 3461
rect 6550 3339 6726 3373
rect -24118 3202 -24084 3308
rect -24030 3202 -23996 3308
rect -23934 3202 -23900 3308
rect -23838 3202 -23804 3308
rect -23742 3202 -23708 3308
rect -23646 3202 -23612 3308
rect -23550 3202 -23516 3308
rect -23454 3202 -23420 3308
rect -23358 3202 -23324 3308
rect -23262 3202 -23228 3308
rect -23166 3202 -23132 3308
rect -23070 3202 -23036 3308
rect -22974 3202 -22940 3308
rect -22878 3202 -22844 3308
rect -22790 3202 -22756 3308
rect -20827 3202 -20793 3308
rect -20739 3202 -20705 3308
rect -20643 3202 -20609 3308
rect -20547 3202 -20513 3308
rect -20451 3202 -20417 3308
rect -20355 3202 -20321 3308
rect -20259 3202 -20225 3308
rect -20163 3202 -20129 3308
rect -20067 3202 -20033 3308
rect -19971 3202 -19937 3308
rect -19875 3202 -19841 3308
rect -19779 3202 -19745 3308
rect -19683 3202 -19649 3308
rect -19587 3202 -19553 3308
rect -19499 3202 -19465 3308
rect -17536 3202 -17502 3308
rect -17448 3202 -17414 3308
rect -17352 3202 -17318 3308
rect -17256 3202 -17222 3308
rect -17160 3202 -17126 3308
rect -17064 3202 -17030 3308
rect -16968 3202 -16934 3308
rect -16872 3202 -16838 3308
rect -16776 3202 -16742 3308
rect -16680 3202 -16646 3308
rect -16584 3202 -16550 3308
rect -16488 3202 -16454 3308
rect -16392 3202 -16358 3308
rect -16296 3202 -16262 3308
rect -16208 3202 -16174 3308
rect -14245 3202 -14211 3308
rect -14157 3202 -14123 3308
rect -14061 3202 -14027 3308
rect -13965 3202 -13931 3308
rect -13869 3202 -13835 3308
rect -13773 3202 -13739 3308
rect -13677 3202 -13643 3308
rect -13581 3202 -13547 3308
rect -13485 3202 -13451 3308
rect -13389 3202 -13355 3308
rect -13293 3202 -13259 3308
rect -13197 3202 -13163 3308
rect -13101 3202 -13067 3308
rect -13005 3202 -12971 3308
rect -12917 3202 -12883 3308
rect -10954 3202 -10920 3308
rect -10866 3202 -10832 3308
rect -10770 3202 -10736 3308
rect -10674 3202 -10640 3308
rect -10578 3202 -10544 3308
rect -10482 3202 -10448 3308
rect -10386 3202 -10352 3308
rect -10290 3202 -10256 3308
rect -10194 3202 -10160 3308
rect -10098 3202 -10064 3308
rect -10002 3202 -9968 3308
rect -9906 3202 -9872 3308
rect -9810 3202 -9776 3308
rect -9714 3202 -9680 3308
rect -9626 3202 -9592 3308
rect -7664 3202 -7630 3308
rect -7576 3202 -7542 3308
rect -7480 3202 -7446 3308
rect -7384 3202 -7350 3308
rect -7288 3202 -7254 3308
rect -7192 3202 -7158 3308
rect -7096 3202 -7062 3308
rect -7000 3202 -6966 3308
rect -6904 3202 -6870 3308
rect -6808 3202 -6774 3308
rect -6712 3202 -6678 3308
rect -6616 3202 -6582 3308
rect -6520 3202 -6486 3308
rect -6424 3202 -6390 3308
rect -6336 3202 -6302 3308
rect -4373 3202 -4339 3308
rect -4285 3202 -4251 3308
rect -4189 3202 -4155 3308
rect -4093 3202 -4059 3308
rect -3997 3202 -3963 3308
rect -3901 3202 -3867 3308
rect -3805 3202 -3771 3308
rect -3709 3202 -3675 3308
rect -3613 3202 -3579 3308
rect -3517 3202 -3483 3308
rect -3421 3202 -3387 3308
rect -3325 3202 -3291 3308
rect -3229 3202 -3195 3308
rect -3133 3202 -3099 3308
rect -3045 3202 -3011 3308
rect -1082 3202 -1048 3308
rect -994 3202 -960 3308
rect -898 3202 -864 3308
rect -802 3202 -768 3308
rect -706 3202 -672 3308
rect -610 3202 -576 3308
rect -514 3202 -480 3308
rect -418 3202 -384 3308
rect -322 3202 -288 3308
rect -226 3202 -192 3308
rect -130 3202 -96 3308
rect -34 3202 0 3308
rect 62 3202 96 3308
rect 158 3202 192 3308
rect 246 3202 280 3308
rect 7372 1702 7406 2478
rect 7756 1702 7790 2478
rect 8320 1702 8354 2478
rect 8704 1702 8738 2478
rect 9256 1702 9290 2478
rect 9640 1702 9674 2478
rect 10187 1702 10221 2478
rect 10571 1702 10605 2478
rect 11114 1702 11148 2478
rect 11498 1702 11532 2478
rect -24792 1418 -24758 1524
rect -24704 1418 -24670 1524
rect -24608 1418 -24574 1524
rect -24512 1418 -24478 1524
rect -24416 1418 -24382 1524
rect -24320 1418 -24286 1524
rect -24224 1418 -24190 1524
rect -24128 1418 -24094 1524
rect -24032 1418 -23998 1524
rect -23936 1418 -23902 1524
rect -23840 1418 -23806 1524
rect -23744 1418 -23710 1524
rect -23648 1418 -23614 1524
rect -23552 1418 -23518 1524
rect -23464 1418 -23430 1524
rect -23233 1418 -23199 1524
rect -23145 1418 -23111 1524
rect -23049 1418 -23015 1524
rect -22953 1418 -22919 1524
rect -22857 1418 -22823 1524
rect -22761 1418 -22727 1524
rect -22665 1418 -22631 1524
rect -22569 1418 -22535 1524
rect -22473 1418 -22439 1524
rect -22377 1418 -22343 1524
rect -22281 1418 -22247 1524
rect -22185 1418 -22151 1524
rect -22089 1418 -22055 1524
rect -21993 1418 -21959 1524
rect -21905 1418 -21871 1524
rect -21501 1418 -21467 1524
rect -21413 1418 -21379 1524
rect -21317 1418 -21283 1524
rect -21221 1418 -21187 1524
rect -21125 1418 -21091 1524
rect -21029 1418 -20995 1524
rect -20933 1418 -20899 1524
rect -20837 1418 -20803 1524
rect -20741 1418 -20707 1524
rect -20645 1418 -20611 1524
rect -20549 1418 -20515 1524
rect -20453 1418 -20419 1524
rect -20357 1418 -20323 1524
rect -20261 1418 -20227 1524
rect -20173 1418 -20139 1524
rect -19942 1418 -19908 1524
rect -19854 1418 -19820 1524
rect -19758 1418 -19724 1524
rect -19662 1418 -19628 1524
rect -19566 1418 -19532 1524
rect -19470 1418 -19436 1524
rect -19374 1418 -19340 1524
rect -19278 1418 -19244 1524
rect -19182 1418 -19148 1524
rect -19086 1418 -19052 1524
rect -18990 1418 -18956 1524
rect -18894 1418 -18860 1524
rect -18798 1418 -18764 1524
rect -18702 1418 -18668 1524
rect -18614 1418 -18580 1524
rect -18210 1418 -18176 1524
rect -18122 1418 -18088 1524
rect -18026 1418 -17992 1524
rect -17930 1418 -17896 1524
rect -17834 1418 -17800 1524
rect -17738 1418 -17704 1524
rect -17642 1418 -17608 1524
rect -17546 1418 -17512 1524
rect -17450 1418 -17416 1524
rect -17354 1418 -17320 1524
rect -17258 1418 -17224 1524
rect -17162 1418 -17128 1524
rect -17066 1418 -17032 1524
rect -16970 1418 -16936 1524
rect -16882 1418 -16848 1524
rect -16651 1418 -16617 1524
rect -16563 1418 -16529 1524
rect -16467 1418 -16433 1524
rect -16371 1418 -16337 1524
rect -16275 1418 -16241 1524
rect -16179 1418 -16145 1524
rect -16083 1418 -16049 1524
rect -15987 1418 -15953 1524
rect -15891 1418 -15857 1524
rect -15795 1418 -15761 1524
rect -15699 1418 -15665 1524
rect -15603 1418 -15569 1524
rect -15507 1418 -15473 1524
rect -15411 1418 -15377 1524
rect -15323 1418 -15289 1524
rect -14919 1418 -14885 1524
rect -14831 1418 -14797 1524
rect -14735 1418 -14701 1524
rect -14639 1418 -14605 1524
rect -14543 1418 -14509 1524
rect -14447 1418 -14413 1524
rect -14351 1418 -14317 1524
rect -14255 1418 -14221 1524
rect -14159 1418 -14125 1524
rect -14063 1418 -14029 1524
rect -13967 1418 -13933 1524
rect -13871 1418 -13837 1524
rect -13775 1418 -13741 1524
rect -13679 1418 -13645 1524
rect -13591 1418 -13557 1524
rect -13360 1418 -13326 1524
rect -13272 1418 -13238 1524
rect -13176 1418 -13142 1524
rect -13080 1418 -13046 1524
rect -12984 1418 -12950 1524
rect -12888 1418 -12854 1524
rect -12792 1418 -12758 1524
rect -12696 1418 -12662 1524
rect -12600 1418 -12566 1524
rect -12504 1418 -12470 1524
rect -12408 1418 -12374 1524
rect -12312 1418 -12278 1524
rect -12216 1418 -12182 1524
rect -12120 1418 -12086 1524
rect -12032 1418 -11998 1524
rect -11628 1418 -11594 1524
rect -11540 1418 -11506 1524
rect -11444 1418 -11410 1524
rect -11348 1418 -11314 1524
rect -11252 1418 -11218 1524
rect -11156 1418 -11122 1524
rect -11060 1418 -11026 1524
rect -10964 1418 -10930 1524
rect -10868 1418 -10834 1524
rect -10772 1418 -10738 1524
rect -10676 1418 -10642 1524
rect -10580 1418 -10546 1524
rect -10484 1418 -10450 1524
rect -10388 1418 -10354 1524
rect -10300 1418 -10266 1524
rect -10069 1418 -10035 1524
rect -9981 1418 -9947 1524
rect -9885 1418 -9851 1524
rect -9789 1418 -9755 1524
rect -9693 1418 -9659 1524
rect -9597 1418 -9563 1524
rect -9501 1418 -9467 1524
rect -9405 1418 -9371 1524
rect -9309 1418 -9275 1524
rect -9213 1418 -9179 1524
rect -9117 1418 -9083 1524
rect -9021 1418 -8987 1524
rect -8925 1418 -8891 1524
rect -8829 1418 -8795 1524
rect -8741 1418 -8707 1524
rect -8338 1418 -8304 1524
rect -8250 1418 -8216 1524
rect -8154 1418 -8120 1524
rect -8058 1418 -8024 1524
rect -7962 1418 -7928 1524
rect -7866 1418 -7832 1524
rect -7770 1418 -7736 1524
rect -7674 1418 -7640 1524
rect -7578 1418 -7544 1524
rect -7482 1418 -7448 1524
rect -7386 1418 -7352 1524
rect -7290 1418 -7256 1524
rect -7194 1418 -7160 1524
rect -7098 1418 -7064 1524
rect -7010 1418 -6976 1524
rect -6779 1418 -6745 1524
rect -6691 1418 -6657 1524
rect -6595 1418 -6561 1524
rect -6499 1418 -6465 1524
rect -6403 1418 -6369 1524
rect -6307 1418 -6273 1524
rect -6211 1418 -6177 1524
rect -6115 1418 -6081 1524
rect -6019 1418 -5985 1524
rect -5923 1418 -5889 1524
rect -5827 1418 -5793 1524
rect -5731 1418 -5697 1524
rect -5635 1418 -5601 1524
rect -5539 1418 -5505 1524
rect -5451 1418 -5417 1524
rect -5047 1418 -5013 1524
rect -4959 1418 -4925 1524
rect -4863 1418 -4829 1524
rect -4767 1418 -4733 1524
rect -4671 1418 -4637 1524
rect -4575 1418 -4541 1524
rect -4479 1418 -4445 1524
rect -4383 1418 -4349 1524
rect -4287 1418 -4253 1524
rect -4191 1418 -4157 1524
rect -4095 1418 -4061 1524
rect -3999 1418 -3965 1524
rect -3903 1418 -3869 1524
rect -3807 1418 -3773 1524
rect -3719 1418 -3685 1524
rect -3488 1418 -3454 1524
rect -3400 1418 -3366 1524
rect -3304 1418 -3270 1524
rect -3208 1418 -3174 1524
rect -3112 1418 -3078 1524
rect -3016 1418 -2982 1524
rect -2920 1418 -2886 1524
rect -2824 1418 -2790 1524
rect -2728 1418 -2694 1524
rect -2632 1418 -2598 1524
rect -2536 1418 -2502 1524
rect -2440 1418 -2406 1524
rect -2344 1418 -2310 1524
rect -2248 1418 -2214 1524
rect -2160 1418 -2126 1524
rect -1756 1418 -1722 1524
rect -1668 1418 -1634 1524
rect -1572 1418 -1538 1524
rect -1476 1418 -1442 1524
rect -1380 1418 -1346 1524
rect -1284 1418 -1250 1524
rect -1188 1418 -1154 1524
rect -1092 1418 -1058 1524
rect -996 1418 -962 1524
rect -900 1418 -866 1524
rect -804 1418 -770 1524
rect -708 1418 -674 1524
rect -612 1418 -578 1524
rect -516 1418 -482 1524
rect -428 1418 -394 1524
rect -197 1418 -163 1524
rect -109 1418 -75 1524
rect -13 1418 21 1524
rect 83 1418 117 1524
rect 179 1418 213 1524
rect 275 1418 309 1524
rect 371 1418 405 1524
rect 467 1418 501 1524
rect 563 1418 597 1524
rect 659 1418 693 1524
rect 755 1418 789 1524
rect 851 1418 885 1524
rect 947 1418 981 1524
rect 1043 1418 1077 1524
rect 1131 1418 1165 1524
rect 7372 774 7406 1550
rect 7756 774 7790 1550
rect 8320 774 8354 1550
rect 8704 774 8738 1550
rect 9256 774 9290 1550
rect 9640 774 9674 1550
rect 10187 775 10221 1551
rect 10571 775 10605 1551
rect -24351 485 -23975 519
rect -23242 485 -22866 519
rect -22360 485 -21984 519
rect -21060 485 -20684 519
rect -19951 485 -19575 519
rect -19069 485 -18693 519
rect -17769 485 -17393 519
rect -16660 485 -16284 519
rect -15778 485 -15402 519
rect -14478 485 -14102 519
rect -13369 485 -12993 519
rect -12487 485 -12111 519
rect -11187 485 -10811 519
rect -10078 485 -9702 519
rect -9196 485 -8820 519
rect -7897 485 -7521 519
rect -6788 485 -6412 519
rect -5906 485 -5530 519
rect -4606 485 -4230 519
rect -3497 485 -3121 519
rect -2615 485 -2239 519
rect -1315 485 -939 519
rect -206 485 170 519
rect 676 485 1052 519
rect 11114 774 11148 1550
rect 11498 774 11532 1550
rect 12169 1332 12203 1508
rect 12265 1332 12299 1508
rect 12361 1332 12395 1508
rect 12935 1409 13111 1443
rect 12935 1321 13111 1355
rect -24351 293 -23975 327
rect -23242 293 -22866 327
rect -22360 293 -21984 327
rect -21060 293 -20684 327
rect -19951 293 -19575 327
rect -19069 293 -18693 327
rect -17769 293 -17393 327
rect -16660 293 -16284 327
rect -15778 293 -15402 327
rect -14478 293 -14102 327
rect -13369 293 -12993 327
rect -12487 293 -12111 327
rect -11187 293 -10811 327
rect -10078 293 -9702 327
rect -9196 293 -8820 327
rect -7897 293 -7521 327
rect -6788 293 -6412 327
rect -5906 293 -5530 327
rect -4606 293 -4230 327
rect -3497 293 -3121 327
rect -2615 293 -2239 327
rect -1315 293 -939 327
rect -206 293 170 327
rect 676 293 1052 327
rect 5670 -1101 5846 -1067
rect 5670 -1189 5846 -1155
rect 6110 -1101 6286 -1067
rect 6110 -1189 6286 -1155
rect 6550 -1101 6726 -1067
rect 6550 -1189 6726 -1155
rect -24201 -2803 -23825 -2769
rect -23616 -2803 -23440 -2769
rect -23616 -2891 -23440 -2857
rect -22164 -2803 -21788 -2769
rect -21596 -2803 -21420 -2769
rect -21596 -2891 -21420 -2857
rect -20434 -2803 -20058 -2769
rect -19855 -2803 -19679 -2769
rect -19855 -2891 -19679 -2857
rect -18674 -2803 -18298 -2769
rect -18076 -2803 -17900 -2769
rect 7372 -2826 7406 -2050
rect 7756 -2826 7790 -2050
rect 8320 -2826 8354 -2050
rect 8704 -2826 8738 -2050
rect 9256 -2826 9290 -2050
rect 9640 -2826 9674 -2050
rect 10187 -2826 10221 -2050
rect 10571 -2826 10605 -2050
rect 11114 -2826 11148 -2050
rect 11498 -2826 11532 -2050
rect -18076 -2891 -17900 -2857
rect -24201 -2995 -23825 -2961
rect -22164 -2995 -21788 -2961
rect -20434 -2995 -20058 -2961
rect -18674 -2995 -18298 -2961
rect 7372 -3754 7406 -2978
rect 7756 -3754 7790 -2978
rect 8320 -3754 8354 -2978
rect 8704 -3754 8738 -2978
rect 9256 -3754 9290 -2978
rect 9640 -3754 9674 -2978
rect 10187 -3753 10221 -2977
rect 10571 -3753 10605 -2977
rect -24150 -4615 -23774 -4581
rect -23572 -4615 -23396 -4581
rect -23572 -4703 -23396 -4669
rect 11114 -3754 11148 -2978
rect 11498 -3754 11532 -2978
rect 12169 -3196 12203 -3020
rect 12265 -3196 12299 -3020
rect 12361 -3196 12395 -3020
rect 12935 -3119 13111 -3085
rect 12935 -3207 13111 -3173
rect -22414 -4615 -22038 -4581
rect -21834 -4615 -21658 -4581
rect -21834 -4703 -21658 -4669
rect -24150 -4807 -23774 -4773
rect -22414 -4807 -22038 -4773
rect -20725 -5142 -20691 -5036
rect -20637 -5142 -20603 -5036
rect -20541 -5142 -20507 -5036
rect -20445 -5142 -20411 -5036
rect -20349 -5142 -20315 -5036
rect -20253 -5142 -20219 -5036
rect -20157 -5142 -20123 -5036
rect -20061 -5142 -20027 -5036
rect -19965 -5142 -19931 -5036
rect -19869 -5142 -19835 -5036
rect -19773 -5142 -19739 -5036
rect -19677 -5142 -19643 -5036
rect -19581 -5142 -19547 -5036
rect -19485 -5142 -19451 -5036
rect -19397 -5142 -19363 -5036
rect -19166 -5142 -19132 -5036
rect -19078 -5142 -19044 -5036
rect -18982 -5142 -18948 -5036
rect -18886 -5142 -18852 -5036
rect -18790 -5142 -18756 -5036
rect -18694 -5142 -18660 -5036
rect -18598 -5142 -18564 -5036
rect -18502 -5142 -18468 -5036
rect -18406 -5142 -18372 -5036
rect -18310 -5142 -18276 -5036
rect -18214 -5142 -18180 -5036
rect -18118 -5142 -18084 -5036
rect -18022 -5142 -17988 -5036
rect -17926 -5142 -17892 -5036
rect -17838 -5142 -17804 -5036
rect -17434 -5142 -17400 -5036
rect -17346 -5142 -17312 -5036
rect -17250 -5142 -17216 -5036
rect -17154 -5142 -17120 -5036
rect -17058 -5142 -17024 -5036
rect -16962 -5142 -16928 -5036
rect -16866 -5142 -16832 -5036
rect -16770 -5142 -16736 -5036
rect -16674 -5142 -16640 -5036
rect -16578 -5142 -16544 -5036
rect -16482 -5142 -16448 -5036
rect -16386 -5142 -16352 -5036
rect -16290 -5142 -16256 -5036
rect -16194 -5142 -16160 -5036
rect -16106 -5142 -16072 -5036
rect -15875 -5142 -15841 -5036
rect -15787 -5142 -15753 -5036
rect -15691 -5142 -15657 -5036
rect -15595 -5142 -15561 -5036
rect -15499 -5142 -15465 -5036
rect -15403 -5142 -15369 -5036
rect -15307 -5142 -15273 -5036
rect -15211 -5142 -15177 -5036
rect -15115 -5142 -15081 -5036
rect -15019 -5142 -14985 -5036
rect -14923 -5142 -14889 -5036
rect -14827 -5142 -14793 -5036
rect -14731 -5142 -14697 -5036
rect -14635 -5142 -14601 -5036
rect -14547 -5142 -14513 -5036
rect -14143 -5142 -14109 -5036
rect -14055 -5142 -14021 -5036
rect -13959 -5142 -13925 -5036
rect -13863 -5142 -13829 -5036
rect -13767 -5142 -13733 -5036
rect -13671 -5142 -13637 -5036
rect -13575 -5142 -13541 -5036
rect -13479 -5142 -13445 -5036
rect -13383 -5142 -13349 -5036
rect -13287 -5142 -13253 -5036
rect -13191 -5142 -13157 -5036
rect -13095 -5142 -13061 -5036
rect -12999 -5142 -12965 -5036
rect -12903 -5142 -12869 -5036
rect -12815 -5142 -12781 -5036
rect -12584 -5142 -12550 -5036
rect -12496 -5142 -12462 -5036
rect -12400 -5142 -12366 -5036
rect -12304 -5142 -12270 -5036
rect -12208 -5142 -12174 -5036
rect -12112 -5142 -12078 -5036
rect -12016 -5142 -11982 -5036
rect -11920 -5142 -11886 -5036
rect -11824 -5142 -11790 -5036
rect -11728 -5142 -11694 -5036
rect -11632 -5142 -11598 -5036
rect -11536 -5142 -11502 -5036
rect -11440 -5142 -11406 -5036
rect -11344 -5142 -11310 -5036
rect -11256 -5142 -11222 -5036
rect -10852 -5142 -10818 -5036
rect -10764 -5142 -10730 -5036
rect -10668 -5142 -10634 -5036
rect -10572 -5142 -10538 -5036
rect -10476 -5142 -10442 -5036
rect -10380 -5142 -10346 -5036
rect -10284 -5142 -10250 -5036
rect -10188 -5142 -10154 -5036
rect -10092 -5142 -10058 -5036
rect -9996 -5142 -9962 -5036
rect -9900 -5142 -9866 -5036
rect -9804 -5142 -9770 -5036
rect -9708 -5142 -9674 -5036
rect -9612 -5142 -9578 -5036
rect -9524 -5142 -9490 -5036
rect -9293 -5142 -9259 -5036
rect -9205 -5142 -9171 -5036
rect -9109 -5142 -9075 -5036
rect -9013 -5142 -8979 -5036
rect -8917 -5142 -8883 -5036
rect -8821 -5142 -8787 -5036
rect -8725 -5142 -8691 -5036
rect -8629 -5142 -8595 -5036
rect -8533 -5142 -8499 -5036
rect -8437 -5142 -8403 -5036
rect -8341 -5142 -8307 -5036
rect -8245 -5142 -8211 -5036
rect -8149 -5142 -8115 -5036
rect -8053 -5142 -8019 -5036
rect -7965 -5142 -7931 -5036
rect 5670 -5529 5846 -5495
rect 5670 -5617 5846 -5583
rect 6110 -5529 6286 -5495
rect 6110 -5617 6286 -5583
rect 6550 -5529 6726 -5495
rect 6550 -5617 6726 -5583
rect -24150 -5907 -23774 -5873
rect -23574 -5907 -23398 -5873
rect -23574 -5995 -23398 -5961
rect -22414 -5907 -22038 -5873
rect -21840 -5907 -21664 -5873
rect -21840 -5995 -21664 -5961
rect -24150 -6099 -23774 -6065
rect -22414 -6099 -22038 -6065
rect -20284 -6075 -19908 -6041
rect -19175 -6075 -18799 -6041
rect -18293 -6075 -17917 -6041
rect -16993 -6075 -16617 -6041
rect -15884 -6075 -15508 -6041
rect -15002 -6075 -14626 -6041
rect -13702 -6075 -13326 -6041
rect -12593 -6075 -12217 -6041
rect -11711 -6075 -11335 -6041
rect -10411 -6075 -10035 -6041
rect -9302 -6075 -8926 -6041
rect -8420 -6075 -8044 -6041
rect -20284 -6267 -19908 -6233
rect -19175 -6267 -18799 -6233
rect -18293 -6267 -17917 -6233
rect -16993 -6267 -16617 -6233
rect -15884 -6267 -15508 -6233
rect -15002 -6267 -14626 -6233
rect -13702 -6267 -13326 -6233
rect -12593 -6267 -12217 -6233
rect -11711 -6267 -11335 -6233
rect -10411 -6267 -10035 -6233
rect -9302 -6267 -8926 -6233
rect -8420 -6267 -8044 -6233
rect -24150 -7880 -23774 -7846
rect -23572 -7880 -23396 -7846
rect -23572 -7968 -23396 -7934
rect 7372 -7254 7406 -6478
rect 7756 -7254 7790 -6478
rect 8320 -7254 8354 -6478
rect 8704 -7254 8738 -6478
rect 9256 -7254 9290 -6478
rect 9640 -7254 9674 -6478
rect 10187 -7254 10221 -6478
rect 10571 -7254 10605 -6478
rect 11114 -7254 11148 -6478
rect 11498 -7254 11532 -6478
rect -22413 -7880 -22037 -7846
rect -21838 -7880 -21662 -7846
rect -21838 -7968 -21662 -7934
rect -24150 -8072 -23774 -8038
rect -22413 -8072 -22037 -8038
rect 7372 -8182 7406 -7406
rect 7756 -8182 7790 -7406
rect 8320 -8182 8354 -7406
rect 8704 -8182 8738 -7406
rect 9256 -8182 9290 -7406
rect 9640 -8182 9674 -7406
rect 10187 -8181 10221 -7405
rect 10571 -8181 10605 -7405
rect -20725 -8407 -20691 -8301
rect -20637 -8407 -20603 -8301
rect -20541 -8407 -20507 -8301
rect -20445 -8407 -20411 -8301
rect -20349 -8407 -20315 -8301
rect -20253 -8407 -20219 -8301
rect -20157 -8407 -20123 -8301
rect -20061 -8407 -20027 -8301
rect -19965 -8407 -19931 -8301
rect -19869 -8407 -19835 -8301
rect -19773 -8407 -19739 -8301
rect -19677 -8407 -19643 -8301
rect -19581 -8407 -19547 -8301
rect -19485 -8407 -19451 -8301
rect -19397 -8407 -19363 -8301
rect -19166 -8407 -19132 -8301
rect -19078 -8407 -19044 -8301
rect -18982 -8407 -18948 -8301
rect -18886 -8407 -18852 -8301
rect -18790 -8407 -18756 -8301
rect -18694 -8407 -18660 -8301
rect -18598 -8407 -18564 -8301
rect -18502 -8407 -18468 -8301
rect -18406 -8407 -18372 -8301
rect -18310 -8407 -18276 -8301
rect -18214 -8407 -18180 -8301
rect -18118 -8407 -18084 -8301
rect -18022 -8407 -17988 -8301
rect -17926 -8407 -17892 -8301
rect -17838 -8407 -17804 -8301
rect -17434 -8407 -17400 -8301
rect -17346 -8407 -17312 -8301
rect -17250 -8407 -17216 -8301
rect -17154 -8407 -17120 -8301
rect -17058 -8407 -17024 -8301
rect -16962 -8407 -16928 -8301
rect -16866 -8407 -16832 -8301
rect -16770 -8407 -16736 -8301
rect -16674 -8407 -16640 -8301
rect -16578 -8407 -16544 -8301
rect -16482 -8407 -16448 -8301
rect -16386 -8407 -16352 -8301
rect -16290 -8407 -16256 -8301
rect -16194 -8407 -16160 -8301
rect -16106 -8407 -16072 -8301
rect -15875 -8407 -15841 -8301
rect -15787 -8407 -15753 -8301
rect -15691 -8407 -15657 -8301
rect -15595 -8407 -15561 -8301
rect -15499 -8407 -15465 -8301
rect -15403 -8407 -15369 -8301
rect -15307 -8407 -15273 -8301
rect -15211 -8407 -15177 -8301
rect -15115 -8407 -15081 -8301
rect -15019 -8407 -14985 -8301
rect -14923 -8407 -14889 -8301
rect -14827 -8407 -14793 -8301
rect -14731 -8407 -14697 -8301
rect -14635 -8407 -14601 -8301
rect -14547 -8407 -14513 -8301
rect -14143 -8407 -14109 -8301
rect -14055 -8407 -14021 -8301
rect -13959 -8407 -13925 -8301
rect -13863 -8407 -13829 -8301
rect -13767 -8407 -13733 -8301
rect -13671 -8407 -13637 -8301
rect -13575 -8407 -13541 -8301
rect -13479 -8407 -13445 -8301
rect -13383 -8407 -13349 -8301
rect -13287 -8407 -13253 -8301
rect -13191 -8407 -13157 -8301
rect -13095 -8407 -13061 -8301
rect -12999 -8407 -12965 -8301
rect -12903 -8407 -12869 -8301
rect -12815 -8407 -12781 -8301
rect -12584 -8407 -12550 -8301
rect -12496 -8407 -12462 -8301
rect -12400 -8407 -12366 -8301
rect -12304 -8407 -12270 -8301
rect -12208 -8407 -12174 -8301
rect -12112 -8407 -12078 -8301
rect -12016 -8407 -11982 -8301
rect -11920 -8407 -11886 -8301
rect -11824 -8407 -11790 -8301
rect -11728 -8407 -11694 -8301
rect -11632 -8407 -11598 -8301
rect -11536 -8407 -11502 -8301
rect -11440 -8407 -11406 -8301
rect -11344 -8407 -11310 -8301
rect -11256 -8407 -11222 -8301
rect -10852 -8407 -10818 -8301
rect -10764 -8407 -10730 -8301
rect -10668 -8407 -10634 -8301
rect -10572 -8407 -10538 -8301
rect -10476 -8407 -10442 -8301
rect -10380 -8407 -10346 -8301
rect -10284 -8407 -10250 -8301
rect -10188 -8407 -10154 -8301
rect -10092 -8407 -10058 -8301
rect -9996 -8407 -9962 -8301
rect -9900 -8407 -9866 -8301
rect -9804 -8407 -9770 -8301
rect -9708 -8407 -9674 -8301
rect -9612 -8407 -9578 -8301
rect -9524 -8407 -9490 -8301
rect -9293 -8407 -9259 -8301
rect -9205 -8407 -9171 -8301
rect -9109 -8407 -9075 -8301
rect -9013 -8407 -8979 -8301
rect -8917 -8407 -8883 -8301
rect -8821 -8407 -8787 -8301
rect -8725 -8407 -8691 -8301
rect -8629 -8407 -8595 -8301
rect -8533 -8407 -8499 -8301
rect -8437 -8407 -8403 -8301
rect -8341 -8407 -8307 -8301
rect -8245 -8407 -8211 -8301
rect -8149 -8407 -8115 -8301
rect -8053 -8407 -8019 -8301
rect -7965 -8407 -7931 -8301
rect 11114 -8182 11148 -7406
rect 11498 -8182 11532 -7406
rect 12169 -7624 12203 -7448
rect 12265 -7624 12299 -7448
rect 12361 -7624 12395 -7448
rect 12935 -7547 13111 -7513
rect 12935 -7635 13111 -7601
rect -24150 -9172 -23774 -9138
rect -23571 -9172 -23395 -9138
rect -23571 -9260 -23395 -9226
rect -22414 -9172 -22038 -9138
rect -21834 -9172 -21658 -9138
rect -21834 -9260 -21658 -9226
rect -24150 -9364 -23774 -9330
rect -22414 -9364 -22038 -9330
rect -20284 -9340 -19908 -9306
rect -19175 -9340 -18799 -9306
rect -18293 -9340 -17917 -9306
rect -16993 -9340 -16617 -9306
rect -15884 -9340 -15508 -9306
rect -15002 -9340 -14626 -9306
rect -13702 -9340 -13326 -9306
rect -12593 -9340 -12217 -9306
rect -11711 -9340 -11335 -9306
rect -10411 -9340 -10035 -9306
rect -9302 -9340 -8926 -9306
rect -8420 -9340 -8044 -9306
rect -20284 -9532 -19908 -9498
rect -19175 -9532 -18799 -9498
rect -18293 -9532 -17917 -9498
rect -16993 -9532 -16617 -9498
rect -15884 -9532 -15508 -9498
rect -15002 -9532 -14626 -9498
rect -13702 -9532 -13326 -9498
rect -12593 -9532 -12217 -9498
rect -11711 -9532 -11335 -9498
rect -10411 -9532 -10035 -9498
rect -9302 -9532 -8926 -9498
rect -8420 -9532 -8044 -9498
rect 5670 -10157 5846 -10123
rect 5670 -10245 5846 -10211
rect 6110 -10157 6286 -10123
rect 6110 -10245 6286 -10211
rect 6550 -10157 6726 -10123
rect 6550 -10245 6726 -10211
rect -24150 -11144 -23774 -11110
rect -23571 -11144 -23395 -11110
rect -23571 -11232 -23395 -11198
rect -22413 -11144 -22037 -11110
rect -21838 -11144 -21662 -11110
rect -21838 -11232 -21662 -11198
rect -24150 -11336 -23774 -11302
rect -22413 -11336 -22037 -11302
rect -20725 -11671 -20691 -11565
rect -20637 -11671 -20603 -11565
rect -20541 -11671 -20507 -11565
rect -20445 -11671 -20411 -11565
rect -20349 -11671 -20315 -11565
rect -20253 -11671 -20219 -11565
rect -20157 -11671 -20123 -11565
rect -20061 -11671 -20027 -11565
rect -19965 -11671 -19931 -11565
rect -19869 -11671 -19835 -11565
rect -19773 -11671 -19739 -11565
rect -19677 -11671 -19643 -11565
rect -19581 -11671 -19547 -11565
rect -19485 -11671 -19451 -11565
rect -19397 -11671 -19363 -11565
rect -19166 -11671 -19132 -11565
rect -19078 -11671 -19044 -11565
rect -18982 -11671 -18948 -11565
rect -18886 -11671 -18852 -11565
rect -18790 -11671 -18756 -11565
rect -18694 -11671 -18660 -11565
rect -18598 -11671 -18564 -11565
rect -18502 -11671 -18468 -11565
rect -18406 -11671 -18372 -11565
rect -18310 -11671 -18276 -11565
rect -18214 -11671 -18180 -11565
rect -18118 -11671 -18084 -11565
rect -18022 -11671 -17988 -11565
rect -17926 -11671 -17892 -11565
rect -17838 -11671 -17804 -11565
rect -17434 -11671 -17400 -11565
rect -17346 -11671 -17312 -11565
rect -17250 -11671 -17216 -11565
rect -17154 -11671 -17120 -11565
rect -17058 -11671 -17024 -11565
rect -16962 -11671 -16928 -11565
rect -16866 -11671 -16832 -11565
rect -16770 -11671 -16736 -11565
rect -16674 -11671 -16640 -11565
rect -16578 -11671 -16544 -11565
rect -16482 -11671 -16448 -11565
rect -16386 -11671 -16352 -11565
rect -16290 -11671 -16256 -11565
rect -16194 -11671 -16160 -11565
rect -16106 -11671 -16072 -11565
rect -15875 -11671 -15841 -11565
rect -15787 -11671 -15753 -11565
rect -15691 -11671 -15657 -11565
rect -15595 -11671 -15561 -11565
rect -15499 -11671 -15465 -11565
rect -15403 -11671 -15369 -11565
rect -15307 -11671 -15273 -11565
rect -15211 -11671 -15177 -11565
rect -15115 -11671 -15081 -11565
rect -15019 -11671 -14985 -11565
rect -14923 -11671 -14889 -11565
rect -14827 -11671 -14793 -11565
rect -14731 -11671 -14697 -11565
rect -14635 -11671 -14601 -11565
rect -14547 -11671 -14513 -11565
rect -14143 -11671 -14109 -11565
rect -14055 -11671 -14021 -11565
rect -13959 -11671 -13925 -11565
rect -13863 -11671 -13829 -11565
rect -13767 -11671 -13733 -11565
rect -13671 -11671 -13637 -11565
rect -13575 -11671 -13541 -11565
rect -13479 -11671 -13445 -11565
rect -13383 -11671 -13349 -11565
rect -13287 -11671 -13253 -11565
rect -13191 -11671 -13157 -11565
rect -13095 -11671 -13061 -11565
rect -12999 -11671 -12965 -11565
rect -12903 -11671 -12869 -11565
rect -12815 -11671 -12781 -11565
rect -12584 -11671 -12550 -11565
rect -12496 -11671 -12462 -11565
rect -12400 -11671 -12366 -11565
rect -12304 -11671 -12270 -11565
rect -12208 -11671 -12174 -11565
rect -12112 -11671 -12078 -11565
rect -12016 -11671 -11982 -11565
rect -11920 -11671 -11886 -11565
rect -11824 -11671 -11790 -11565
rect -11728 -11671 -11694 -11565
rect -11632 -11671 -11598 -11565
rect -11536 -11671 -11502 -11565
rect -11440 -11671 -11406 -11565
rect -11344 -11671 -11310 -11565
rect -11256 -11671 -11222 -11565
rect -10852 -11671 -10818 -11565
rect -10764 -11671 -10730 -11565
rect -10668 -11671 -10634 -11565
rect -10572 -11671 -10538 -11565
rect -10476 -11671 -10442 -11565
rect -10380 -11671 -10346 -11565
rect -10284 -11671 -10250 -11565
rect -10188 -11671 -10154 -11565
rect -10092 -11671 -10058 -11565
rect -9996 -11671 -9962 -11565
rect -9900 -11671 -9866 -11565
rect -9804 -11671 -9770 -11565
rect -9708 -11671 -9674 -11565
rect -9612 -11671 -9578 -11565
rect -9524 -11671 -9490 -11565
rect -9293 -11671 -9259 -11565
rect -9205 -11671 -9171 -11565
rect -9109 -11671 -9075 -11565
rect -9013 -11671 -8979 -11565
rect -8917 -11671 -8883 -11565
rect -8821 -11671 -8787 -11565
rect -8725 -11671 -8691 -11565
rect -8629 -11671 -8595 -11565
rect -8533 -11671 -8499 -11565
rect -8437 -11671 -8403 -11565
rect -8341 -11671 -8307 -11565
rect -8245 -11671 -8211 -11565
rect -8149 -11671 -8115 -11565
rect -8053 -11671 -8019 -11565
rect -7965 -11671 -7931 -11565
rect 7372 -11882 7406 -11106
rect 7756 -11882 7790 -11106
rect 8320 -11882 8354 -11106
rect 8704 -11882 8738 -11106
rect 9256 -11882 9290 -11106
rect 9640 -11882 9674 -11106
rect 10187 -11882 10221 -11106
rect 10571 -11882 10605 -11106
rect 11114 -11882 11148 -11106
rect 11498 -11882 11532 -11106
rect -24150 -12436 -23774 -12402
rect -23571 -12436 -23395 -12402
rect -23571 -12524 -23395 -12490
rect -22413 -12436 -22037 -12402
rect -21842 -12436 -21666 -12402
rect -21842 -12524 -21666 -12490
rect -24150 -12628 -23774 -12594
rect -22413 -12628 -22037 -12594
rect -20284 -12604 -19908 -12570
rect -19175 -12604 -18799 -12570
rect -18293 -12604 -17917 -12570
rect -16993 -12604 -16617 -12570
rect -15884 -12604 -15508 -12570
rect -15002 -12604 -14626 -12570
rect -13702 -12604 -13326 -12570
rect -12593 -12604 -12217 -12570
rect -11711 -12604 -11335 -12570
rect -10411 -12604 -10035 -12570
rect -9302 -12604 -8926 -12570
rect -8420 -12604 -8044 -12570
rect -20284 -12796 -19908 -12762
rect -19175 -12796 -18799 -12762
rect -18293 -12796 -17917 -12762
rect -16993 -12796 -16617 -12762
rect -15884 -12796 -15508 -12762
rect -15002 -12796 -14626 -12762
rect -13702 -12796 -13326 -12762
rect -12593 -12796 -12217 -12762
rect -11711 -12796 -11335 -12762
rect -10411 -12796 -10035 -12762
rect -9302 -12796 -8926 -12762
rect -8420 -12796 -8044 -12762
rect 7372 -12810 7406 -12034
rect 7756 -12810 7790 -12034
rect 8320 -12810 8354 -12034
rect 8704 -12810 8738 -12034
rect 9256 -12810 9290 -12034
rect 9640 -12810 9674 -12034
rect 10187 -12809 10221 -12033
rect 10571 -12809 10605 -12033
rect 11114 -12810 11148 -12034
rect 11498 -12810 11532 -12034
rect 12169 -12252 12203 -12076
rect 12265 -12252 12299 -12076
rect 12361 -12252 12395 -12076
rect 12935 -12175 13111 -12141
rect 12935 -12263 13111 -12229
rect -1650 -14020 -1616 -13844
rect -1562 -14020 -1528 -13844
rect -11264 -14139 -11158 -14105
rect -24093 -15304 -24059 -14928
rect -23901 -15304 -23867 -14928
rect -17176 -14929 -17000 -14895
rect -17176 -15025 -17000 -14991
rect -17176 -15121 -17000 -15087
rect -11264 -14227 -11158 -14193
rect -11264 -14323 -11158 -14289
rect -11264 -14419 -11158 -14385
rect -11264 -14515 -11158 -14481
rect -11264 -14611 -11158 -14577
rect -11264 -14707 -11158 -14673
rect -11264 -14803 -11158 -14769
rect -11264 -14899 -11158 -14865
rect -11264 -14995 -11158 -14961
rect -11264 -15091 -11158 -15057
rect -11264 -15187 -11158 -15153
rect -11264 -15283 -11158 -15249
rect -11264 -15379 -11158 -15345
rect -4366 -14391 -4332 -14215
rect -4278 -14391 -4244 -14215
rect -1650 -14399 -1616 -14223
rect -1562 -14399 -1528 -14223
rect -4366 -14831 -4332 -14655
rect -4278 -14831 -4244 -14655
rect -1650 -14839 -1616 -14663
rect -1562 -14839 -1528 -14663
rect 5670 -14685 5846 -14651
rect 5670 -14773 5846 -14739
rect 6110 -14685 6286 -14651
rect 6110 -14773 6286 -14739
rect 6550 -14685 6726 -14651
rect 6550 -14773 6726 -14739
rect -4366 -15210 -4332 -15034
rect -4278 -15210 -4244 -15034
rect -1650 -15218 -1616 -15042
rect -1562 -15218 -1528 -15042
rect -11264 -15467 -11158 -15433
rect -7717 -15548 -7683 -15372
rect -7629 -15548 -7595 -15372
rect -4366 -15650 -4332 -15474
rect -4278 -15650 -4244 -15474
rect -1650 -15658 -1616 -15482
rect -1562 -15658 -1528 -15482
rect -7716 -16048 -7682 -15872
rect -7628 -16048 -7594 -15872
rect -4366 -16029 -4332 -15853
rect -4278 -16029 -4244 -15853
rect -24092 -16489 -24058 -16113
rect -23900 -16489 -23866 -16113
rect -1650 -16037 -1616 -15861
rect -1562 -16037 -1528 -15861
rect -17176 -16329 -17000 -16295
rect -17176 -16425 -17000 -16391
rect -17176 -16521 -17000 -16487
rect -7717 -16528 -7683 -16352
rect -7629 -16528 -7595 -16352
rect -4366 -16469 -4332 -16293
rect -4278 -16469 -4244 -16293
rect -1650 -16477 -1616 -16301
rect -1562 -16477 -1528 -16301
rect 7372 -16410 7406 -15634
rect 7756 -16410 7790 -15634
rect 8320 -16410 8354 -15634
rect 8704 -16410 8738 -15634
rect 9256 -16410 9290 -15634
rect 9640 -16410 9674 -15634
rect 10187 -16410 10221 -15634
rect 10571 -16410 10605 -15634
rect 11114 -16410 11148 -15634
rect 11498 -16410 11532 -15634
rect -11262 -16955 -11156 -16921
rect -24087 -17702 -24053 -17326
rect -23895 -17702 -23861 -17326
rect -17176 -17729 -17000 -17695
rect -17176 -17825 -17000 -17791
rect -21156 -18236 -21122 -18060
rect -21068 -18236 -21034 -18060
rect -17176 -17921 -17000 -17887
rect -15565 -18107 -15531 -17931
rect -15477 -18107 -15443 -17931
rect -11262 -17043 -11156 -17009
rect -11262 -17139 -11156 -17105
rect -11262 -17235 -11156 -17201
rect -11262 -17331 -11156 -17297
rect -11262 -17427 -11156 -17393
rect -11262 -17523 -11156 -17489
rect -11262 -17619 -11156 -17585
rect -11262 -17715 -11156 -17681
rect -11262 -17811 -11156 -17777
rect -11262 -17907 -11156 -17873
rect -11262 -18003 -11156 -17969
rect -11262 -18099 -11156 -18065
rect -11262 -18195 -11156 -18161
rect -7717 -17028 -7683 -16852
rect -7629 -17028 -7595 -16852
rect -4366 -16848 -4332 -16672
rect -4278 -16848 -4244 -16672
rect -1650 -16856 -1616 -16680
rect -1562 -16856 -1528 -16680
rect -4366 -17288 -4332 -17112
rect -4278 -17288 -4244 -17112
rect -7717 -17508 -7683 -17332
rect -7629 -17508 -7595 -17332
rect -1650 -17296 -1616 -17120
rect -1562 -17296 -1528 -17120
rect 7372 -17338 7406 -16562
rect 7756 -17338 7790 -16562
rect 8320 -17338 8354 -16562
rect 8704 -17338 8738 -16562
rect 9256 -17338 9290 -16562
rect 9640 -17338 9674 -16562
rect 10187 -17337 10221 -16561
rect 10571 -17337 10605 -16561
rect -4366 -17667 -4332 -17491
rect -4278 -17667 -4244 -17491
rect -1650 -17675 -1616 -17499
rect -1562 -17675 -1528 -17499
rect -7717 -17968 -7683 -17792
rect -7629 -17968 -7595 -17792
rect 11114 -17338 11148 -16562
rect 11498 -17338 11532 -16562
rect 12169 -16780 12203 -16604
rect 12265 -16780 12299 -16604
rect 12361 -16780 12395 -16604
rect 12935 -16703 13111 -16669
rect 12935 -16791 13111 -16757
rect 16159 -17237 16193 -17061
rect 16255 -17237 16289 -17061
rect 16351 -17237 16385 -17061
rect 16447 -17237 16481 -17061
rect 16543 -17237 16577 -17061
rect -4366 -18107 -4332 -17931
rect -4278 -18107 -4244 -17931
rect -1650 -18115 -1616 -17939
rect -1562 -18115 -1528 -17939
rect -11262 -18283 -11156 -18249
rect -24072 -18821 -24038 -18445
rect -23880 -18821 -23846 -18445
rect -21155 -18736 -21121 -18560
rect -21067 -18736 -21033 -18560
rect -15564 -18607 -15530 -18431
rect -15476 -18607 -15442 -18431
rect -7731 -18428 -7697 -18252
rect -7643 -18428 -7609 -18252
rect -4366 -18486 -4332 -18310
rect -4278 -18486 -4244 -18310
rect -1650 -18494 -1616 -18318
rect -1562 -18494 -1528 -18318
rect -21156 -19216 -21122 -19040
rect -21068 -19216 -21034 -19040
rect -17176 -19129 -17000 -19095
rect -15565 -19087 -15531 -18911
rect -15477 -19087 -15443 -18911
rect -7729 -18908 -7695 -18732
rect -7641 -18908 -7607 -18732
rect -4366 -18926 -4332 -18750
rect -4278 -18926 -4244 -18750
rect -1650 -18934 -1616 -18758
rect -1562 -18934 -1528 -18758
rect -17176 -19225 -17000 -19191
rect -24070 -20015 -24036 -19639
rect -23878 -20015 -23844 -19639
rect -21156 -19716 -21122 -19540
rect -21068 -19716 -21034 -19540
rect -17176 -19321 -17000 -19287
rect -4366 -19305 -4332 -19129
rect -4278 -19305 -4244 -19129
rect -1650 -19313 -1616 -19137
rect -1562 -19313 -1528 -19137
rect 5670 -19213 5846 -19179
rect 5670 -19301 5846 -19267
rect 6110 -19213 6286 -19179
rect 6110 -19301 6286 -19267
rect 6550 -19213 6726 -19179
rect 6550 -19301 6726 -19267
rect -15565 -19587 -15531 -19411
rect -15477 -19587 -15443 -19411
rect -4366 -19745 -4332 -19569
rect -4278 -19745 -4244 -19569
rect -1650 -19753 -1616 -19577
rect -1562 -19753 -1528 -19577
rect 17540 -18665 17916 -18631
rect 18108 -18743 18284 -18709
rect 17540 -18857 17916 -18823
rect 18108 -18831 18284 -18797
rect -21156 -20196 -21122 -20020
rect -21068 -20196 -21034 -20020
rect -15565 -20067 -15531 -19891
rect -15477 -20067 -15443 -19891
rect -11262 -19912 -11156 -19878
rect -21156 -20656 -21122 -20480
rect -21068 -20656 -21034 -20480
rect -17176 -20529 -17000 -20495
rect -17176 -20625 -17000 -20591
rect -24039 -21215 -24005 -20839
rect -23847 -21215 -23813 -20839
rect -21170 -21116 -21136 -20940
rect -21082 -21116 -21048 -20940
rect -17176 -20721 -17000 -20687
rect -15565 -20527 -15531 -20351
rect -15477 -20527 -15443 -20351
rect -15579 -20987 -15545 -20811
rect -15491 -20987 -15457 -20811
rect -11262 -20000 -11156 -19966
rect -11262 -20096 -11156 -20062
rect -11262 -20192 -11156 -20158
rect -11262 -20288 -11156 -20254
rect -11262 -20384 -11156 -20350
rect -11262 -20480 -11156 -20446
rect -11262 -20576 -11156 -20542
rect -11262 -20672 -11156 -20638
rect -11262 -20768 -11156 -20734
rect -11262 -20864 -11156 -20830
rect -11262 -20960 -11156 -20926
rect -11262 -21056 -11156 -21022
rect -11262 -21152 -11156 -21118
rect -4366 -20124 -4332 -19948
rect -4278 -20124 -4244 -19948
rect -1650 -20132 -1616 -19956
rect -1562 -20132 -1528 -19956
rect 16159 -20111 16193 -19935
rect 16255 -20111 16289 -19935
rect 16351 -20111 16385 -19935
rect 16447 -20111 16481 -19935
rect 16543 -20111 16577 -19935
rect -4366 -20564 -4332 -20388
rect -4278 -20564 -4244 -20388
rect -1650 -20572 -1616 -20396
rect -1562 -20572 -1528 -20396
rect -4366 -20943 -4332 -20767
rect -4278 -20943 -4244 -20767
rect 7372 -20938 7406 -20162
rect 7756 -20938 7790 -20162
rect 8320 -20938 8354 -20162
rect 8704 -20938 8738 -20162
rect 9256 -20938 9290 -20162
rect 9640 -20938 9674 -20162
rect 10187 -20938 10221 -20162
rect 10571 -20938 10605 -20162
rect 11114 -20938 11148 -20162
rect 11498 -20938 11532 -20162
rect -21168 -21596 -21134 -21420
rect -21080 -21596 -21046 -21420
rect -15577 -21467 -15543 -21291
rect -15489 -21467 -15455 -21291
rect -11262 -21240 -11156 -21206
rect 7372 -21866 7406 -21090
rect 7756 -21866 7790 -21090
rect 8320 -21866 8354 -21090
rect 8704 -21866 8738 -21090
rect 9256 -21866 9290 -21090
rect 9640 -21866 9674 -21090
rect 10187 -21865 10221 -21089
rect 10571 -21865 10605 -21089
rect -17176 -21929 -17000 -21895
rect -17176 -22025 -17000 -21991
rect -24040 -22518 -24006 -22142
rect -23848 -22518 -23814 -22142
rect -17176 -22121 -17000 -22087
rect 11114 -21866 11148 -21090
rect 11498 -21866 11532 -21090
rect 12169 -21308 12203 -21132
rect 12265 -21308 12299 -21132
rect 12361 -21308 12395 -21132
rect 12935 -21231 13111 -21197
rect 12935 -21319 13111 -21285
rect -11262 -22491 -11156 -22457
rect -17176 -23329 -17000 -23295
rect -24040 -23827 -24006 -23451
rect -23848 -23827 -23814 -23451
rect -17176 -23425 -17000 -23391
rect -17176 -23521 -17000 -23487
rect -11262 -22579 -11156 -22545
rect -11262 -22675 -11156 -22641
rect -11262 -22771 -11156 -22737
rect -11262 -22867 -11156 -22833
rect -11262 -22963 -11156 -22929
rect -11262 -23059 -11156 -23025
rect -11262 -23155 -11156 -23121
rect -11262 -23251 -11156 -23217
rect -11262 -23347 -11156 -23313
rect -11262 -23443 -11156 -23409
rect -11262 -23539 -11156 -23505
rect -11262 -23635 -11156 -23601
rect -11262 -23731 -11156 -23697
rect -11262 -23819 -11156 -23785
rect 5670 -23741 5846 -23707
rect 5670 -23829 5846 -23795
rect 6110 -23741 6286 -23707
rect 6110 -23829 6286 -23795
rect 6550 -23741 6726 -23707
rect 6550 -23829 6726 -23795
rect -17176 -24729 -17000 -24695
rect -17176 -24825 -17000 -24791
rect -17176 -24921 -17000 -24887
rect -11262 -25259 -11156 -25225
rect -11262 -25347 -11156 -25313
rect -11262 -25443 -11156 -25409
rect -11262 -25539 -11156 -25505
rect -11262 -25635 -11156 -25601
rect -11262 -25731 -11156 -25697
rect -11262 -25827 -11156 -25793
rect -11262 -25923 -11156 -25889
rect -11262 -26019 -11156 -25985
rect -11262 -26115 -11156 -26081
rect -11262 -26211 -11156 -26177
rect -11262 -26307 -11156 -26273
rect -11262 -26403 -11156 -26369
rect -11262 -26499 -11156 -26465
rect 7372 -25466 7406 -24690
rect 7756 -25466 7790 -24690
rect 8320 -25466 8354 -24690
rect 8704 -25466 8738 -24690
rect 9256 -25466 9290 -24690
rect 9640 -25466 9674 -24690
rect 10187 -25466 10221 -24690
rect 10571 -25466 10605 -24690
rect 11114 -25466 11148 -24690
rect 11498 -25466 11532 -24690
rect 7372 -26394 7406 -25618
rect 7756 -26394 7790 -25618
rect 8320 -26394 8354 -25618
rect 8704 -26394 8738 -25618
rect 9256 -26394 9290 -25618
rect 9640 -26394 9674 -25618
rect 10187 -26393 10221 -25617
rect 10571 -26393 10605 -25617
rect -11262 -26587 -11156 -26553
rect 11114 -26394 11148 -25618
rect 11498 -26394 11532 -25618
rect 12169 -25836 12203 -25660
rect 12265 -25836 12299 -25660
rect 12361 -25836 12395 -25660
rect 12935 -25759 13111 -25725
rect 12935 -25847 13111 -25813
rect -11262 -27892 -11156 -27858
rect -11262 -27980 -11156 -27946
rect -11262 -28076 -11156 -28042
rect -11262 -28172 -11156 -28138
rect -11262 -28268 -11156 -28234
rect -11262 -28364 -11156 -28330
rect -11262 -28460 -11156 -28426
rect -11262 -28556 -11156 -28522
rect -11262 -28652 -11156 -28618
rect -11262 -28748 -11156 -28714
rect -11262 -28844 -11156 -28810
rect -11262 -28940 -11156 -28906
rect -11262 -29036 -11156 -29002
rect -11262 -29132 -11156 -29098
rect 5670 -28269 5846 -28235
rect 5670 -28357 5846 -28323
rect 6110 -28269 6286 -28235
rect 6110 -28357 6286 -28323
rect 6550 -28269 6726 -28235
rect 6550 -28357 6726 -28323
rect -11262 -29220 -11156 -29186
rect 7372 -29994 7406 -29218
rect 7756 -29994 7790 -29218
rect 8320 -29994 8354 -29218
rect 8704 -29994 8738 -29218
rect 9256 -29994 9290 -29218
rect 9640 -29994 9674 -29218
rect 10187 -29994 10221 -29218
rect 10571 -29994 10605 -29218
rect 11114 -29994 11148 -29218
rect 11498 -29994 11532 -29218
rect -11262 -30501 -11156 -30467
rect -11262 -30589 -11156 -30555
rect -11262 -30685 -11156 -30651
rect -11262 -30781 -11156 -30747
rect -11262 -30877 -11156 -30843
rect -11262 -30973 -11156 -30939
rect -11262 -31069 -11156 -31035
rect -11262 -31165 -11156 -31131
rect -11262 -31261 -11156 -31227
rect -11262 -31357 -11156 -31323
rect -11262 -31453 -11156 -31419
rect -11262 -31549 -11156 -31515
rect -11262 -31645 -11156 -31611
rect -11262 -31741 -11156 -31707
rect 7372 -30922 7406 -30146
rect 7756 -30922 7790 -30146
rect 8320 -30922 8354 -30146
rect 8704 -30922 8738 -30146
rect 9256 -30922 9290 -30146
rect 9640 -30922 9674 -30146
rect 10187 -30921 10221 -30145
rect 10571 -30921 10605 -30145
rect 11114 -30922 11148 -30146
rect 11498 -30922 11532 -30146
rect 12169 -30364 12203 -30188
rect 12265 -30364 12299 -30188
rect 12361 -30364 12395 -30188
rect 12935 -30287 13111 -30253
rect 12935 -30375 13111 -30341
rect -11262 -31829 -11156 -31795
rect 5670 -32797 5846 -32763
rect 5670 -32885 5846 -32851
rect 6110 -32797 6286 -32763
rect 6110 -32885 6286 -32851
rect 6550 -32797 6726 -32763
rect 6550 -32885 6726 -32851
rect -11264 -33121 -11158 -33087
rect -11264 -33209 -11158 -33175
rect -11264 -33305 -11158 -33271
rect -11264 -33401 -11158 -33367
rect -11264 -33497 -11158 -33463
rect -11264 -33593 -11158 -33559
rect -11264 -33689 -11158 -33655
rect -11264 -33785 -11158 -33751
rect -11264 -33881 -11158 -33847
rect -11264 -33977 -11158 -33943
rect -11264 -34073 -11158 -34039
rect -11264 -34169 -11158 -34135
rect -11264 -34265 -11158 -34231
rect -11264 -34361 -11158 -34327
rect -11264 -34449 -11158 -34415
rect 7372 -34522 7406 -33746
rect 7756 -34522 7790 -33746
rect 8320 -34522 8354 -33746
rect 8704 -34522 8738 -33746
rect 9256 -34522 9290 -33746
rect 9640 -34522 9674 -33746
rect 10187 -34522 10221 -33746
rect 10571 -34522 10605 -33746
rect 11114 -34522 11148 -33746
rect 11498 -34522 11532 -33746
rect 7372 -35450 7406 -34674
rect 7756 -35450 7790 -34674
rect 8320 -35450 8354 -34674
rect 8704 -35450 8738 -34674
rect 9256 -35450 9290 -34674
rect 9640 -35450 9674 -34674
rect 10187 -35449 10221 -34673
rect 10571 -35449 10605 -34673
rect 11114 -35450 11148 -34674
rect 11498 -35450 11532 -34674
rect 12169 -34892 12203 -34716
rect 12265 -34892 12299 -34716
rect 12361 -34892 12395 -34716
rect 12935 -34815 13111 -34781
rect 12935 -34903 13111 -34869
rect 12886 -35903 12920 -35727
rect 12974 -35903 13008 -35727
rect 12886 -36282 12920 -36106
rect 12974 -36282 13008 -36106
<< pdiffc >>
rect 1719 5546 1753 6072
rect 1807 5546 1841 6072
rect 1903 5546 1937 6072
rect 1999 5546 2033 6072
rect 2095 5546 2129 6072
rect 2191 5546 2225 6072
rect 2287 5546 2321 6072
rect 2383 5546 2417 6072
rect 2479 5546 2513 6072
rect 2575 5546 2609 6072
rect 2671 5546 2705 6072
rect 2767 5546 2801 6072
rect 2863 5546 2897 6072
rect 2959 5546 2993 6072
rect 3047 5546 3081 6072
rect 3325 5546 3359 6072
rect 3413 5546 3447 6072
rect 3509 5546 3543 6072
rect 3605 5546 3639 6072
rect 3701 5546 3735 6072
rect 3797 5546 3831 6072
rect 3893 5546 3927 6072
rect 3989 5546 4023 6072
rect 4085 5546 4119 6072
rect 4181 5546 4215 6072
rect 4277 5546 4311 6072
rect 4373 5546 4407 6072
rect 4469 5546 4503 6072
rect 4565 5546 4599 6072
rect 4653 5546 4687 6072
rect 5029 5544 5063 6070
rect 5117 5544 5151 6070
rect 5213 5544 5247 6070
rect 5309 5544 5343 6070
rect 5405 5544 5439 6070
rect 5501 5544 5535 6070
rect 5597 5544 5631 6070
rect 5693 5544 5727 6070
rect 5789 5544 5823 6070
rect 5885 5544 5919 6070
rect 5981 5544 6015 6070
rect 6077 5544 6111 6070
rect 6173 5544 6207 6070
rect 6269 5544 6303 6070
rect 6357 5544 6391 6070
rect 6951 5239 6985 5429
rect 7047 5239 7081 5429
rect 7143 5239 7177 5429
rect 7239 5239 7273 5429
rect 7335 5239 7369 5429
rect 7431 5239 7465 5429
rect 7527 5239 7561 5429
rect 7821 5425 8011 5459
rect 7821 5329 8015 5363
rect 7821 5233 8011 5267
rect 7821 5137 8015 5171
rect -24118 3822 -24084 4348
rect -24030 3822 -23996 4348
rect -23934 3822 -23900 4348
rect -23838 3822 -23804 4348
rect -23742 3822 -23708 4348
rect -23646 3822 -23612 4348
rect -23550 3822 -23516 4348
rect -23454 3822 -23420 4348
rect -23358 3822 -23324 4348
rect -23262 3822 -23228 4348
rect -23166 3822 -23132 4348
rect -23070 3822 -23036 4348
rect -22974 3822 -22940 4348
rect -22878 3822 -22844 4348
rect -22790 3822 -22756 4348
rect -20827 3822 -20793 4348
rect -20739 3822 -20705 4348
rect -20643 3822 -20609 4348
rect -20547 3822 -20513 4348
rect -20451 3822 -20417 4348
rect -20355 3822 -20321 4348
rect -20259 3822 -20225 4348
rect -20163 3822 -20129 4348
rect -20067 3822 -20033 4348
rect -19971 3822 -19937 4348
rect -19875 3822 -19841 4348
rect -19779 3822 -19745 4348
rect -19683 3822 -19649 4348
rect -19587 3822 -19553 4348
rect -19499 3822 -19465 4348
rect -17536 3822 -17502 4348
rect -17448 3822 -17414 4348
rect -17352 3822 -17318 4348
rect -17256 3822 -17222 4348
rect -17160 3822 -17126 4348
rect -17064 3822 -17030 4348
rect -16968 3822 -16934 4348
rect -16872 3822 -16838 4348
rect -16776 3822 -16742 4348
rect -16680 3822 -16646 4348
rect -16584 3822 -16550 4348
rect -16488 3822 -16454 4348
rect -16392 3822 -16358 4348
rect -16296 3822 -16262 4348
rect -16208 3822 -16174 4348
rect -14245 3822 -14211 4348
rect -14157 3822 -14123 4348
rect -14061 3822 -14027 4348
rect -13965 3822 -13931 4348
rect -13869 3822 -13835 4348
rect -13773 3822 -13739 4348
rect -13677 3822 -13643 4348
rect -13581 3822 -13547 4348
rect -13485 3822 -13451 4348
rect -13389 3822 -13355 4348
rect -13293 3822 -13259 4348
rect -13197 3822 -13163 4348
rect -13101 3822 -13067 4348
rect -13005 3822 -12971 4348
rect -12917 3822 -12883 4348
rect -10954 3822 -10920 4348
rect -10866 3822 -10832 4348
rect -10770 3822 -10736 4348
rect -10674 3822 -10640 4348
rect -10578 3822 -10544 4348
rect -10482 3822 -10448 4348
rect -10386 3822 -10352 4348
rect -10290 3822 -10256 4348
rect -10194 3822 -10160 4348
rect -10098 3822 -10064 4348
rect -10002 3822 -9968 4348
rect -9906 3822 -9872 4348
rect -9810 3822 -9776 4348
rect -9714 3822 -9680 4348
rect -9626 3822 -9592 4348
rect -7664 3822 -7630 4348
rect -7576 3822 -7542 4348
rect -7480 3822 -7446 4348
rect -7384 3822 -7350 4348
rect -7288 3822 -7254 4348
rect -7192 3822 -7158 4348
rect -7096 3822 -7062 4348
rect -7000 3822 -6966 4348
rect -6904 3822 -6870 4348
rect -6808 3822 -6774 4348
rect -6712 3822 -6678 4348
rect -6616 3822 -6582 4348
rect -6520 3822 -6486 4348
rect -6424 3822 -6390 4348
rect -6336 3822 -6302 4348
rect -4373 3822 -4339 4348
rect -4285 3822 -4251 4348
rect -4189 3822 -4155 4348
rect -4093 3822 -4059 4348
rect -3997 3822 -3963 4348
rect -3901 3822 -3867 4348
rect -3805 3822 -3771 4348
rect -3709 3822 -3675 4348
rect -3613 3822 -3579 4348
rect -3517 3822 -3483 4348
rect -3421 3822 -3387 4348
rect -3325 3822 -3291 4348
rect -3229 3822 -3195 4348
rect -3133 3822 -3099 4348
rect -3045 3822 -3011 4348
rect -1082 3822 -1048 4348
rect -994 3822 -960 4348
rect -898 3822 -864 4348
rect -802 3822 -768 4348
rect -706 3822 -672 4348
rect -610 3822 -576 4348
rect -514 3822 -480 4348
rect -418 3822 -384 4348
rect -322 3822 -288 4348
rect -226 3822 -192 4348
rect -130 3822 -96 4348
rect -34 3822 0 4348
rect 62 3822 96 4348
rect 158 3822 192 4348
rect 246 3822 280 4348
rect 5670 3877 5860 3911
rect 5670 3781 5864 3815
rect 5670 3685 5860 3719
rect 5670 3589 5864 3623
rect 6110 3877 6300 3911
rect 6110 3781 6304 3815
rect 6110 3685 6300 3719
rect 6110 3589 6304 3623
rect 6550 3877 6740 3911
rect 6550 3781 6744 3815
rect 6550 3685 6740 3719
rect 6550 3589 6744 3623
rect 7150 2909 7184 3207
rect 7246 2909 7280 3207
rect 7342 2909 7376 3207
rect 7438 2909 7472 3207
rect 7534 2909 7568 3207
rect 7630 2909 7664 3207
rect 7726 2909 7760 3207
rect 7822 2909 7856 3207
rect 7918 2909 7952 3207
rect 8098 2909 8132 3207
rect 8194 2909 8228 3207
rect 8290 2909 8324 3207
rect 8386 2909 8420 3207
rect 8482 2909 8516 3207
rect 8578 2909 8612 3207
rect 8674 2909 8708 3207
rect 8770 2909 8804 3207
rect 8866 2909 8900 3207
rect 9034 2909 9068 3207
rect 9130 2909 9164 3207
rect 9226 2909 9260 3207
rect 9322 2909 9356 3207
rect 9418 2909 9452 3207
rect 9514 2909 9548 3207
rect 9610 2909 9644 3207
rect 9706 2909 9740 3207
rect 9802 2909 9836 3207
rect 9965 2909 9999 3207
rect 10061 2909 10095 3207
rect 10157 2909 10191 3207
rect 10253 2909 10287 3207
rect 10349 2909 10383 3207
rect 10445 2909 10479 3207
rect 10541 2909 10575 3207
rect 10637 2909 10671 3207
rect 10733 2909 10767 3207
rect 10892 2909 10926 3207
rect 10988 2909 11022 3207
rect 11084 2909 11118 3207
rect 11180 2909 11214 3207
rect 11276 2909 11310 3207
rect 11372 2909 11406 3207
rect 11468 2909 11502 3207
rect 11564 2909 11598 3207
rect 11660 2909 11694 3207
rect -24792 2038 -24758 2564
rect -24704 2038 -24670 2564
rect -24608 2038 -24574 2564
rect -24512 2038 -24478 2564
rect -24416 2038 -24382 2564
rect -24320 2038 -24286 2564
rect -24224 2038 -24190 2564
rect -24128 2038 -24094 2564
rect -24032 2038 -23998 2564
rect -23936 2038 -23902 2564
rect -23840 2038 -23806 2564
rect -23744 2038 -23710 2564
rect -23648 2038 -23614 2564
rect -23552 2038 -23518 2564
rect -23464 2038 -23430 2564
rect -23233 2038 -23199 2564
rect -23145 2038 -23111 2564
rect -23049 2038 -23015 2564
rect -22953 2038 -22919 2564
rect -22857 2038 -22823 2564
rect -22761 2038 -22727 2564
rect -22665 2038 -22631 2564
rect -22569 2038 -22535 2564
rect -22473 2038 -22439 2564
rect -22377 2038 -22343 2564
rect -22281 2038 -22247 2564
rect -22185 2038 -22151 2564
rect -22089 2038 -22055 2564
rect -21993 2038 -21959 2564
rect -21905 2038 -21871 2564
rect -21501 2038 -21467 2564
rect -21413 2038 -21379 2564
rect -21317 2038 -21283 2564
rect -21221 2038 -21187 2564
rect -21125 2038 -21091 2564
rect -21029 2038 -20995 2564
rect -20933 2038 -20899 2564
rect -20837 2038 -20803 2564
rect -20741 2038 -20707 2564
rect -20645 2038 -20611 2564
rect -20549 2038 -20515 2564
rect -20453 2038 -20419 2564
rect -20357 2038 -20323 2564
rect -20261 2038 -20227 2564
rect -20173 2038 -20139 2564
rect -19942 2038 -19908 2564
rect -19854 2038 -19820 2564
rect -19758 2038 -19724 2564
rect -19662 2038 -19628 2564
rect -19566 2038 -19532 2564
rect -19470 2038 -19436 2564
rect -19374 2038 -19340 2564
rect -19278 2038 -19244 2564
rect -19182 2038 -19148 2564
rect -19086 2038 -19052 2564
rect -18990 2038 -18956 2564
rect -18894 2038 -18860 2564
rect -18798 2038 -18764 2564
rect -18702 2038 -18668 2564
rect -18614 2038 -18580 2564
rect -18210 2038 -18176 2564
rect -18122 2038 -18088 2564
rect -18026 2038 -17992 2564
rect -17930 2038 -17896 2564
rect -17834 2038 -17800 2564
rect -17738 2038 -17704 2564
rect -17642 2038 -17608 2564
rect -17546 2038 -17512 2564
rect -17450 2038 -17416 2564
rect -17354 2038 -17320 2564
rect -17258 2038 -17224 2564
rect -17162 2038 -17128 2564
rect -17066 2038 -17032 2564
rect -16970 2038 -16936 2564
rect -16882 2038 -16848 2564
rect -16651 2038 -16617 2564
rect -16563 2038 -16529 2564
rect -16467 2038 -16433 2564
rect -16371 2038 -16337 2564
rect -16275 2038 -16241 2564
rect -16179 2038 -16145 2564
rect -16083 2038 -16049 2564
rect -15987 2038 -15953 2564
rect -15891 2038 -15857 2564
rect -15795 2038 -15761 2564
rect -15699 2038 -15665 2564
rect -15603 2038 -15569 2564
rect -15507 2038 -15473 2564
rect -15411 2038 -15377 2564
rect -15323 2038 -15289 2564
rect -14919 2038 -14885 2564
rect -14831 2038 -14797 2564
rect -14735 2038 -14701 2564
rect -14639 2038 -14605 2564
rect -14543 2038 -14509 2564
rect -14447 2038 -14413 2564
rect -14351 2038 -14317 2564
rect -14255 2038 -14221 2564
rect -14159 2038 -14125 2564
rect -14063 2038 -14029 2564
rect -13967 2038 -13933 2564
rect -13871 2038 -13837 2564
rect -13775 2038 -13741 2564
rect -13679 2038 -13645 2564
rect -13591 2038 -13557 2564
rect -13360 2038 -13326 2564
rect -13272 2038 -13238 2564
rect -13176 2038 -13142 2564
rect -13080 2038 -13046 2564
rect -12984 2038 -12950 2564
rect -12888 2038 -12854 2564
rect -12792 2038 -12758 2564
rect -12696 2038 -12662 2564
rect -12600 2038 -12566 2564
rect -12504 2038 -12470 2564
rect -12408 2038 -12374 2564
rect -12312 2038 -12278 2564
rect -12216 2038 -12182 2564
rect -12120 2038 -12086 2564
rect -12032 2038 -11998 2564
rect -11628 2038 -11594 2564
rect -11540 2038 -11506 2564
rect -11444 2038 -11410 2564
rect -11348 2038 -11314 2564
rect -11252 2038 -11218 2564
rect -11156 2038 -11122 2564
rect -11060 2038 -11026 2564
rect -10964 2038 -10930 2564
rect -10868 2038 -10834 2564
rect -10772 2038 -10738 2564
rect -10676 2038 -10642 2564
rect -10580 2038 -10546 2564
rect -10484 2038 -10450 2564
rect -10388 2038 -10354 2564
rect -10300 2038 -10266 2564
rect -10069 2038 -10035 2564
rect -9981 2038 -9947 2564
rect -9885 2038 -9851 2564
rect -9789 2038 -9755 2564
rect -9693 2038 -9659 2564
rect -9597 2038 -9563 2564
rect -9501 2038 -9467 2564
rect -9405 2038 -9371 2564
rect -9309 2038 -9275 2564
rect -9213 2038 -9179 2564
rect -9117 2038 -9083 2564
rect -9021 2038 -8987 2564
rect -8925 2038 -8891 2564
rect -8829 2038 -8795 2564
rect -8741 2038 -8707 2564
rect -8338 2038 -8304 2564
rect -8250 2038 -8216 2564
rect -8154 2038 -8120 2564
rect -8058 2038 -8024 2564
rect -7962 2038 -7928 2564
rect -7866 2038 -7832 2564
rect -7770 2038 -7736 2564
rect -7674 2038 -7640 2564
rect -7578 2038 -7544 2564
rect -7482 2038 -7448 2564
rect -7386 2038 -7352 2564
rect -7290 2038 -7256 2564
rect -7194 2038 -7160 2564
rect -7098 2038 -7064 2564
rect -7010 2038 -6976 2564
rect -6779 2038 -6745 2564
rect -6691 2038 -6657 2564
rect -6595 2038 -6561 2564
rect -6499 2038 -6465 2564
rect -6403 2038 -6369 2564
rect -6307 2038 -6273 2564
rect -6211 2038 -6177 2564
rect -6115 2038 -6081 2564
rect -6019 2038 -5985 2564
rect -5923 2038 -5889 2564
rect -5827 2038 -5793 2564
rect -5731 2038 -5697 2564
rect -5635 2038 -5601 2564
rect -5539 2038 -5505 2564
rect -5451 2038 -5417 2564
rect -5047 2038 -5013 2564
rect -4959 2038 -4925 2564
rect -4863 2038 -4829 2564
rect -4767 2038 -4733 2564
rect -4671 2038 -4637 2564
rect -4575 2038 -4541 2564
rect -4479 2038 -4445 2564
rect -4383 2038 -4349 2564
rect -4287 2038 -4253 2564
rect -4191 2038 -4157 2564
rect -4095 2038 -4061 2564
rect -3999 2038 -3965 2564
rect -3903 2038 -3869 2564
rect -3807 2038 -3773 2564
rect -3719 2038 -3685 2564
rect -3488 2038 -3454 2564
rect -3400 2038 -3366 2564
rect -3304 2038 -3270 2564
rect -3208 2038 -3174 2564
rect -3112 2038 -3078 2564
rect -3016 2038 -2982 2564
rect -2920 2038 -2886 2564
rect -2824 2038 -2790 2564
rect -2728 2038 -2694 2564
rect -2632 2038 -2598 2564
rect -2536 2038 -2502 2564
rect -2440 2038 -2406 2564
rect -2344 2038 -2310 2564
rect -2248 2038 -2214 2564
rect -2160 2038 -2126 2564
rect -1756 2038 -1722 2564
rect -1668 2038 -1634 2564
rect -1572 2038 -1538 2564
rect -1476 2038 -1442 2564
rect -1380 2038 -1346 2564
rect -1284 2038 -1250 2564
rect -1188 2038 -1154 2564
rect -1092 2038 -1058 2564
rect -996 2038 -962 2564
rect -900 2038 -866 2564
rect -804 2038 -770 2564
rect -708 2038 -674 2564
rect -612 2038 -578 2564
rect -516 2038 -482 2564
rect -428 2038 -394 2564
rect -197 2038 -163 2564
rect -109 2038 -75 2564
rect -13 2038 21 2564
rect 83 2038 117 2564
rect 179 2038 213 2564
rect 275 2038 309 2564
rect 371 2038 405 2564
rect 467 2038 501 2564
rect 563 2038 597 2564
rect 659 2038 693 2564
rect 755 2038 789 2564
rect 851 2038 885 2564
rect 947 2038 981 2564
rect 1043 2038 1077 2564
rect 1131 2038 1165 2564
rect 11785 1765 11819 1997
rect 11881 1765 11915 1997
rect 11977 1765 12011 1997
rect 12073 1765 12107 1997
rect 12169 1765 12203 1997
rect 12265 1765 12299 1997
rect 12361 1765 12395 1997
rect 12457 1765 12491 1997
rect 12553 1765 12587 1997
rect 12649 1765 12683 1997
rect 12745 1765 12779 1997
rect -24585 673 -24551 863
rect -24489 673 -24455 863
rect -24393 673 -24359 863
rect -24297 673 -24263 863
rect -24201 673 -24167 863
rect -24105 673 -24071 863
rect -24009 673 -23975 863
rect -23476 673 -23442 863
rect -23380 673 -23346 863
rect -23284 673 -23250 863
rect -23188 673 -23154 863
rect -23092 673 -23058 863
rect -22996 673 -22962 863
rect -22900 673 -22866 863
rect -22594 673 -22560 863
rect -22498 673 -22464 863
rect -22402 673 -22368 863
rect -22306 673 -22272 863
rect -22210 673 -22176 863
rect -22114 673 -22080 863
rect -22018 673 -21984 863
rect -21294 673 -21260 863
rect -21198 673 -21164 863
rect -21102 673 -21068 863
rect -21006 673 -20972 863
rect -20910 673 -20876 863
rect -20814 673 -20780 863
rect -20718 673 -20684 863
rect -20185 673 -20151 863
rect -20089 673 -20055 863
rect -19993 673 -19959 863
rect -19897 673 -19863 863
rect -19801 673 -19767 863
rect -19705 673 -19671 863
rect -19609 673 -19575 863
rect -19303 673 -19269 863
rect -19207 673 -19173 863
rect -19111 673 -19077 863
rect -19015 673 -18981 863
rect -18919 673 -18885 863
rect -18823 673 -18789 863
rect -18727 673 -18693 863
rect -18003 673 -17969 863
rect -17907 673 -17873 863
rect -17811 673 -17777 863
rect -17715 673 -17681 863
rect -17619 673 -17585 863
rect -17523 673 -17489 863
rect -17427 673 -17393 863
rect -16894 673 -16860 863
rect -16798 673 -16764 863
rect -16702 673 -16668 863
rect -16606 673 -16572 863
rect -16510 673 -16476 863
rect -16414 673 -16380 863
rect -16318 673 -16284 863
rect -16012 673 -15978 863
rect -15916 673 -15882 863
rect -15820 673 -15786 863
rect -15724 673 -15690 863
rect -15628 673 -15594 863
rect -15532 673 -15498 863
rect -15436 673 -15402 863
rect -14712 673 -14678 863
rect -14616 673 -14582 863
rect -14520 673 -14486 863
rect -14424 673 -14390 863
rect -14328 673 -14294 863
rect -14232 673 -14198 863
rect -14136 673 -14102 863
rect -13603 673 -13569 863
rect -13507 673 -13473 863
rect -13411 673 -13377 863
rect -13315 673 -13281 863
rect -13219 673 -13185 863
rect -13123 673 -13089 863
rect -13027 673 -12993 863
rect -12721 673 -12687 863
rect -12625 673 -12591 863
rect -12529 673 -12495 863
rect -12433 673 -12399 863
rect -12337 673 -12303 863
rect -12241 673 -12207 863
rect -12145 673 -12111 863
rect -11421 673 -11387 863
rect -11325 673 -11291 863
rect -11229 673 -11195 863
rect -11133 673 -11099 863
rect -11037 673 -11003 863
rect -10941 673 -10907 863
rect -10845 673 -10811 863
rect -10312 673 -10278 863
rect -10216 673 -10182 863
rect -10120 673 -10086 863
rect -10024 673 -9990 863
rect -9928 673 -9894 863
rect -9832 673 -9798 863
rect -9736 673 -9702 863
rect -9430 673 -9396 863
rect -9334 673 -9300 863
rect -9238 673 -9204 863
rect -9142 673 -9108 863
rect -9046 673 -9012 863
rect -8950 673 -8916 863
rect -8854 673 -8820 863
rect -8131 673 -8097 863
rect -8035 673 -8001 863
rect -7939 673 -7905 863
rect -7843 673 -7809 863
rect -7747 673 -7713 863
rect -7651 673 -7617 863
rect -7555 673 -7521 863
rect -7022 673 -6988 863
rect -6926 673 -6892 863
rect -6830 673 -6796 863
rect -6734 673 -6700 863
rect -6638 673 -6604 863
rect -6542 673 -6508 863
rect -6446 673 -6412 863
rect -6140 673 -6106 863
rect -6044 673 -6010 863
rect -5948 673 -5914 863
rect -5852 673 -5818 863
rect -5756 673 -5722 863
rect -5660 673 -5626 863
rect -5564 673 -5530 863
rect -4840 673 -4806 863
rect -4744 673 -4710 863
rect -4648 673 -4614 863
rect -4552 673 -4518 863
rect -4456 673 -4422 863
rect -4360 673 -4326 863
rect -4264 673 -4230 863
rect -3731 673 -3697 863
rect -3635 673 -3601 863
rect -3539 673 -3505 863
rect -3443 673 -3409 863
rect -3347 673 -3313 863
rect -3251 673 -3217 863
rect -3155 673 -3121 863
rect -2849 673 -2815 863
rect -2753 673 -2719 863
rect -2657 673 -2623 863
rect -2561 673 -2527 863
rect -2465 673 -2431 863
rect -2369 673 -2335 863
rect -2273 673 -2239 863
rect -1549 673 -1515 863
rect -1453 673 -1419 863
rect -1357 673 -1323 863
rect -1261 673 -1227 863
rect -1165 673 -1131 863
rect -1069 673 -1035 863
rect -973 673 -939 863
rect -440 673 -406 863
rect -344 673 -310 863
rect -248 673 -214 863
rect -152 673 -118 863
rect -56 673 -22 863
rect 40 673 74 863
rect 136 673 170 863
rect 442 673 476 863
rect 538 673 572 863
rect 634 673 668 863
rect 730 673 764 863
rect 826 673 860 863
rect 922 673 956 863
rect 1018 673 1052 863
rect 12935 1859 13125 1893
rect 12935 1763 13129 1797
rect 12935 1667 13125 1701
rect 12935 1571 13129 1605
rect 7150 45 7184 343
rect 7246 45 7280 343
rect 7342 45 7376 343
rect 7438 45 7472 343
rect 7534 45 7568 343
rect 7630 45 7664 343
rect 7726 45 7760 343
rect 7822 45 7856 343
rect 7918 45 7952 343
rect 8098 45 8132 343
rect 8194 45 8228 343
rect 8290 45 8324 343
rect 8386 45 8420 343
rect 8482 45 8516 343
rect 8578 45 8612 343
rect 8674 45 8708 343
rect 8770 45 8804 343
rect 8866 45 8900 343
rect 9034 45 9068 343
rect 9130 45 9164 343
rect 9226 45 9260 343
rect 9322 45 9356 343
rect 9418 45 9452 343
rect 9514 45 9548 343
rect 9610 45 9644 343
rect 9706 45 9740 343
rect 9802 45 9836 343
rect 9965 46 9999 344
rect 10061 46 10095 344
rect 10157 46 10191 344
rect 10253 46 10287 344
rect 10349 46 10383 344
rect 10445 46 10479 344
rect 10541 46 10575 344
rect 10637 46 10671 344
rect 10733 46 10767 344
rect 10892 45 10926 343
rect 10988 45 11022 343
rect 11084 45 11118 343
rect 11180 45 11214 343
rect 11276 45 11310 343
rect 11372 45 11406 343
rect 11468 45 11502 343
rect 11564 45 11598 343
rect 11660 45 11694 343
rect 5670 -651 5860 -617
rect 5670 -747 5864 -713
rect 5670 -843 5860 -809
rect 5670 -939 5864 -905
rect 6110 -651 6300 -617
rect 6110 -747 6304 -713
rect 6110 -843 6300 -809
rect 6110 -939 6304 -905
rect 6550 -651 6740 -617
rect 6550 -747 6744 -713
rect 6550 -843 6740 -809
rect 6550 -939 6744 -905
rect 7150 -1619 7184 -1321
rect 7246 -1619 7280 -1321
rect 7342 -1619 7376 -1321
rect 7438 -1619 7472 -1321
rect 7534 -1619 7568 -1321
rect 7630 -1619 7664 -1321
rect 7726 -1619 7760 -1321
rect 7822 -1619 7856 -1321
rect 7918 -1619 7952 -1321
rect 8098 -1619 8132 -1321
rect 8194 -1619 8228 -1321
rect 8290 -1619 8324 -1321
rect 8386 -1619 8420 -1321
rect 8482 -1619 8516 -1321
rect 8578 -1619 8612 -1321
rect 8674 -1619 8708 -1321
rect 8770 -1619 8804 -1321
rect 8866 -1619 8900 -1321
rect 9034 -1619 9068 -1321
rect 9130 -1619 9164 -1321
rect 9226 -1619 9260 -1321
rect 9322 -1619 9356 -1321
rect 9418 -1619 9452 -1321
rect 9514 -1619 9548 -1321
rect 9610 -1619 9644 -1321
rect 9706 -1619 9740 -1321
rect 9802 -1619 9836 -1321
rect 9965 -1619 9999 -1321
rect 10061 -1619 10095 -1321
rect 10157 -1619 10191 -1321
rect 10253 -1619 10287 -1321
rect 10349 -1619 10383 -1321
rect 10445 -1619 10479 -1321
rect 10541 -1619 10575 -1321
rect 10637 -1619 10671 -1321
rect 10733 -1619 10767 -1321
rect 10892 -1619 10926 -1321
rect 10988 -1619 11022 -1321
rect 11084 -1619 11118 -1321
rect 11180 -1619 11214 -1321
rect 11276 -1619 11310 -1321
rect 11372 -1619 11406 -1321
rect 11468 -1619 11502 -1321
rect 11564 -1619 11598 -1321
rect 11660 -1619 11694 -1321
rect -24435 -2615 -24401 -2425
rect -24339 -2615 -24305 -2425
rect -24243 -2615 -24209 -2425
rect -24147 -2615 -24113 -2425
rect -24051 -2615 -24017 -2425
rect -23955 -2615 -23921 -2425
rect -23859 -2615 -23825 -2425
rect -23616 -2353 -23426 -2319
rect -23616 -2449 -23422 -2415
rect -23616 -2545 -23426 -2511
rect -23616 -2641 -23422 -2607
rect -22398 -2615 -22364 -2425
rect -22302 -2615 -22268 -2425
rect -22206 -2615 -22172 -2425
rect -22110 -2615 -22076 -2425
rect -22014 -2615 -21980 -2425
rect -21918 -2615 -21884 -2425
rect -21822 -2615 -21788 -2425
rect -21596 -2353 -21406 -2319
rect -21596 -2449 -21402 -2415
rect -21596 -2545 -21406 -2511
rect -21596 -2641 -21402 -2607
rect -20668 -2615 -20634 -2425
rect -20572 -2615 -20538 -2425
rect -20476 -2615 -20442 -2425
rect -20380 -2615 -20346 -2425
rect -20284 -2615 -20250 -2425
rect -20188 -2615 -20154 -2425
rect -20092 -2615 -20058 -2425
rect -19855 -2353 -19665 -2319
rect -19855 -2449 -19661 -2415
rect -19855 -2545 -19665 -2511
rect -19855 -2641 -19661 -2607
rect -18908 -2615 -18874 -2425
rect -18812 -2615 -18778 -2425
rect -18716 -2615 -18682 -2425
rect -18620 -2615 -18586 -2425
rect -18524 -2615 -18490 -2425
rect -18428 -2615 -18394 -2425
rect -18332 -2615 -18298 -2425
rect -18076 -2353 -17886 -2319
rect -18076 -2449 -17882 -2415
rect -18076 -2545 -17886 -2511
rect -18076 -2641 -17882 -2607
rect 11785 -2763 11819 -2531
rect 11881 -2763 11915 -2531
rect 11977 -2763 12011 -2531
rect 12073 -2763 12107 -2531
rect 12169 -2763 12203 -2531
rect 12265 -2763 12299 -2531
rect 12361 -2763 12395 -2531
rect 12457 -2763 12491 -2531
rect 12553 -2763 12587 -2531
rect 12649 -2763 12683 -2531
rect 12745 -2763 12779 -2531
rect -24384 -4427 -24350 -4237
rect -24288 -4427 -24254 -4237
rect -24192 -4427 -24158 -4237
rect -24096 -4427 -24062 -4237
rect -24000 -4427 -23966 -4237
rect -23904 -4427 -23870 -4237
rect -23808 -4427 -23774 -4237
rect -23572 -4165 -23382 -4131
rect -23572 -4261 -23378 -4227
rect -23572 -4357 -23382 -4323
rect -23572 -4453 -23378 -4419
rect -22648 -4427 -22614 -4237
rect -22552 -4427 -22518 -4237
rect -22456 -4427 -22422 -4237
rect -22360 -4427 -22326 -4237
rect -22264 -4427 -22230 -4237
rect -22168 -4427 -22134 -4237
rect -22072 -4427 -22038 -4237
rect -21834 -4165 -21644 -4131
rect -21834 -4261 -21640 -4227
rect -21834 -4357 -21644 -4323
rect -21834 -4453 -21640 -4419
rect -20725 -4522 -20691 -3996
rect -20637 -4522 -20603 -3996
rect -20541 -4522 -20507 -3996
rect -20445 -4522 -20411 -3996
rect -20349 -4522 -20315 -3996
rect -20253 -4522 -20219 -3996
rect -20157 -4522 -20123 -3996
rect -20061 -4522 -20027 -3996
rect -19965 -4522 -19931 -3996
rect -19869 -4522 -19835 -3996
rect -19773 -4522 -19739 -3996
rect -19677 -4522 -19643 -3996
rect -19581 -4522 -19547 -3996
rect -19485 -4522 -19451 -3996
rect -19397 -4522 -19363 -3996
rect -19166 -4522 -19132 -3996
rect -19078 -4522 -19044 -3996
rect -18982 -4522 -18948 -3996
rect -18886 -4522 -18852 -3996
rect -18790 -4522 -18756 -3996
rect -18694 -4522 -18660 -3996
rect -18598 -4522 -18564 -3996
rect -18502 -4522 -18468 -3996
rect -18406 -4522 -18372 -3996
rect -18310 -4522 -18276 -3996
rect -18214 -4522 -18180 -3996
rect -18118 -4522 -18084 -3996
rect -18022 -4522 -17988 -3996
rect -17926 -4522 -17892 -3996
rect -17838 -4522 -17804 -3996
rect -17434 -4522 -17400 -3996
rect -17346 -4522 -17312 -3996
rect -17250 -4522 -17216 -3996
rect -17154 -4522 -17120 -3996
rect -17058 -4522 -17024 -3996
rect -16962 -4522 -16928 -3996
rect -16866 -4522 -16832 -3996
rect -16770 -4522 -16736 -3996
rect -16674 -4522 -16640 -3996
rect -16578 -4522 -16544 -3996
rect -16482 -4522 -16448 -3996
rect -16386 -4522 -16352 -3996
rect -16290 -4522 -16256 -3996
rect -16194 -4522 -16160 -3996
rect -16106 -4522 -16072 -3996
rect -15875 -4522 -15841 -3996
rect -15787 -4522 -15753 -3996
rect -15691 -4522 -15657 -3996
rect -15595 -4522 -15561 -3996
rect -15499 -4522 -15465 -3996
rect -15403 -4522 -15369 -3996
rect -15307 -4522 -15273 -3996
rect -15211 -4522 -15177 -3996
rect -15115 -4522 -15081 -3996
rect -15019 -4522 -14985 -3996
rect -14923 -4522 -14889 -3996
rect -14827 -4522 -14793 -3996
rect -14731 -4522 -14697 -3996
rect -14635 -4522 -14601 -3996
rect -14547 -4522 -14513 -3996
rect -14143 -4522 -14109 -3996
rect -14055 -4522 -14021 -3996
rect -13959 -4522 -13925 -3996
rect -13863 -4522 -13829 -3996
rect -13767 -4522 -13733 -3996
rect -13671 -4522 -13637 -3996
rect -13575 -4522 -13541 -3996
rect -13479 -4522 -13445 -3996
rect -13383 -4522 -13349 -3996
rect -13287 -4522 -13253 -3996
rect -13191 -4522 -13157 -3996
rect -13095 -4522 -13061 -3996
rect -12999 -4522 -12965 -3996
rect -12903 -4522 -12869 -3996
rect -12815 -4522 -12781 -3996
rect -12584 -4522 -12550 -3996
rect -12496 -4522 -12462 -3996
rect -12400 -4522 -12366 -3996
rect -12304 -4522 -12270 -3996
rect -12208 -4522 -12174 -3996
rect -12112 -4522 -12078 -3996
rect -12016 -4522 -11982 -3996
rect -11920 -4522 -11886 -3996
rect -11824 -4522 -11790 -3996
rect -11728 -4522 -11694 -3996
rect -11632 -4522 -11598 -3996
rect -11536 -4522 -11502 -3996
rect -11440 -4522 -11406 -3996
rect -11344 -4522 -11310 -3996
rect -11256 -4522 -11222 -3996
rect -10852 -4522 -10818 -3996
rect -10764 -4522 -10730 -3996
rect -10668 -4522 -10634 -3996
rect -10572 -4522 -10538 -3996
rect -10476 -4522 -10442 -3996
rect -10380 -4522 -10346 -3996
rect -10284 -4522 -10250 -3996
rect -10188 -4522 -10154 -3996
rect -10092 -4522 -10058 -3996
rect -9996 -4522 -9962 -3996
rect -9900 -4522 -9866 -3996
rect -9804 -4522 -9770 -3996
rect -9708 -4522 -9674 -3996
rect -9612 -4522 -9578 -3996
rect -9524 -4522 -9490 -3996
rect -9293 -4522 -9259 -3996
rect -9205 -4522 -9171 -3996
rect -9109 -4522 -9075 -3996
rect -9013 -4522 -8979 -3996
rect -8917 -4522 -8883 -3996
rect -8821 -4522 -8787 -3996
rect -8725 -4522 -8691 -3996
rect -8629 -4522 -8595 -3996
rect -8533 -4522 -8499 -3996
rect -8437 -4522 -8403 -3996
rect -8341 -4522 -8307 -3996
rect -8245 -4522 -8211 -3996
rect -8149 -4522 -8115 -3996
rect -8053 -4522 -8019 -3996
rect -7965 -4522 -7931 -3996
rect 12935 -2669 13125 -2635
rect 12935 -2765 13129 -2731
rect 12935 -2861 13125 -2827
rect 12935 -2957 13129 -2923
rect 7150 -4483 7184 -4185
rect 7246 -4483 7280 -4185
rect 7342 -4483 7376 -4185
rect 7438 -4483 7472 -4185
rect 7534 -4483 7568 -4185
rect 7630 -4483 7664 -4185
rect 7726 -4483 7760 -4185
rect 7822 -4483 7856 -4185
rect 7918 -4483 7952 -4185
rect 8098 -4483 8132 -4185
rect 8194 -4483 8228 -4185
rect 8290 -4483 8324 -4185
rect 8386 -4483 8420 -4185
rect 8482 -4483 8516 -4185
rect 8578 -4483 8612 -4185
rect 8674 -4483 8708 -4185
rect 8770 -4483 8804 -4185
rect 8866 -4483 8900 -4185
rect 9034 -4483 9068 -4185
rect 9130 -4483 9164 -4185
rect 9226 -4483 9260 -4185
rect 9322 -4483 9356 -4185
rect 9418 -4483 9452 -4185
rect 9514 -4483 9548 -4185
rect 9610 -4483 9644 -4185
rect 9706 -4483 9740 -4185
rect 9802 -4483 9836 -4185
rect 9965 -4482 9999 -4184
rect 10061 -4482 10095 -4184
rect 10157 -4482 10191 -4184
rect 10253 -4482 10287 -4184
rect 10349 -4482 10383 -4184
rect 10445 -4482 10479 -4184
rect 10541 -4482 10575 -4184
rect 10637 -4482 10671 -4184
rect 10733 -4482 10767 -4184
rect 10892 -4483 10926 -4185
rect 10988 -4483 11022 -4185
rect 11084 -4483 11118 -4185
rect 11180 -4483 11214 -4185
rect 11276 -4483 11310 -4185
rect 11372 -4483 11406 -4185
rect 11468 -4483 11502 -4185
rect 11564 -4483 11598 -4185
rect 11660 -4483 11694 -4185
rect 5670 -5079 5860 -5045
rect 5670 -5175 5864 -5141
rect 5670 -5271 5860 -5237
rect 5670 -5367 5864 -5333
rect 6110 -5079 6300 -5045
rect 6110 -5175 6304 -5141
rect 6110 -5271 6300 -5237
rect 6110 -5367 6304 -5333
rect 6550 -5079 6740 -5045
rect 6550 -5175 6744 -5141
rect 6550 -5271 6740 -5237
rect 6550 -5367 6744 -5333
rect -24384 -5719 -24350 -5529
rect -24288 -5719 -24254 -5529
rect -24192 -5719 -24158 -5529
rect -24096 -5719 -24062 -5529
rect -24000 -5719 -23966 -5529
rect -23904 -5719 -23870 -5529
rect -23808 -5719 -23774 -5529
rect -23574 -5457 -23384 -5423
rect -23574 -5553 -23380 -5519
rect -23574 -5649 -23384 -5615
rect -23574 -5745 -23380 -5711
rect -22648 -5719 -22614 -5529
rect -22552 -5719 -22518 -5529
rect -22456 -5719 -22422 -5529
rect -22360 -5719 -22326 -5529
rect -22264 -5719 -22230 -5529
rect -22168 -5719 -22134 -5529
rect -22072 -5719 -22038 -5529
rect -21840 -5457 -21650 -5423
rect -21840 -5553 -21646 -5519
rect -21840 -5649 -21650 -5615
rect -21840 -5745 -21646 -5711
rect -20518 -5887 -20484 -5697
rect -20422 -5887 -20388 -5697
rect -20326 -5887 -20292 -5697
rect -20230 -5887 -20196 -5697
rect -20134 -5887 -20100 -5697
rect -20038 -5887 -20004 -5697
rect -19942 -5887 -19908 -5697
rect -19409 -5887 -19375 -5697
rect -19313 -5887 -19279 -5697
rect -19217 -5887 -19183 -5697
rect -19121 -5887 -19087 -5697
rect -19025 -5887 -18991 -5697
rect -18929 -5887 -18895 -5697
rect -18833 -5887 -18799 -5697
rect -18527 -5887 -18493 -5697
rect -18431 -5887 -18397 -5697
rect -18335 -5887 -18301 -5697
rect -18239 -5887 -18205 -5697
rect -18143 -5887 -18109 -5697
rect -18047 -5887 -18013 -5697
rect -17951 -5887 -17917 -5697
rect -17227 -5887 -17193 -5697
rect -17131 -5887 -17097 -5697
rect -17035 -5887 -17001 -5697
rect -16939 -5887 -16905 -5697
rect -16843 -5887 -16809 -5697
rect -16747 -5887 -16713 -5697
rect -16651 -5887 -16617 -5697
rect -16118 -5887 -16084 -5697
rect -16022 -5887 -15988 -5697
rect -15926 -5887 -15892 -5697
rect -15830 -5887 -15796 -5697
rect -15734 -5887 -15700 -5697
rect -15638 -5887 -15604 -5697
rect -15542 -5887 -15508 -5697
rect -15236 -5887 -15202 -5697
rect -15140 -5887 -15106 -5697
rect -15044 -5887 -15010 -5697
rect -14948 -5887 -14914 -5697
rect -14852 -5887 -14818 -5697
rect -14756 -5887 -14722 -5697
rect -14660 -5887 -14626 -5697
rect -13936 -5887 -13902 -5697
rect -13840 -5887 -13806 -5697
rect -13744 -5887 -13710 -5697
rect -13648 -5887 -13614 -5697
rect -13552 -5887 -13518 -5697
rect -13456 -5887 -13422 -5697
rect -13360 -5887 -13326 -5697
rect -12827 -5887 -12793 -5697
rect -12731 -5887 -12697 -5697
rect -12635 -5887 -12601 -5697
rect -12539 -5887 -12505 -5697
rect -12443 -5887 -12409 -5697
rect -12347 -5887 -12313 -5697
rect -12251 -5887 -12217 -5697
rect -11945 -5887 -11911 -5697
rect -11849 -5887 -11815 -5697
rect -11753 -5887 -11719 -5697
rect -11657 -5887 -11623 -5697
rect -11561 -5887 -11527 -5697
rect -11465 -5887 -11431 -5697
rect -11369 -5887 -11335 -5697
rect -10645 -5887 -10611 -5697
rect -10549 -5887 -10515 -5697
rect -10453 -5887 -10419 -5697
rect -10357 -5887 -10323 -5697
rect -10261 -5887 -10227 -5697
rect -10165 -5887 -10131 -5697
rect -10069 -5887 -10035 -5697
rect -9536 -5887 -9502 -5697
rect -9440 -5887 -9406 -5697
rect -9344 -5887 -9310 -5697
rect -9248 -5887 -9214 -5697
rect -9152 -5887 -9118 -5697
rect -9056 -5887 -9022 -5697
rect -8960 -5887 -8926 -5697
rect -8654 -5887 -8620 -5697
rect -8558 -5887 -8524 -5697
rect -8462 -5887 -8428 -5697
rect -8366 -5887 -8332 -5697
rect -8270 -5887 -8236 -5697
rect -8174 -5887 -8140 -5697
rect -8078 -5887 -8044 -5697
rect 7150 -6047 7184 -5749
rect 7246 -6047 7280 -5749
rect 7342 -6047 7376 -5749
rect 7438 -6047 7472 -5749
rect 7534 -6047 7568 -5749
rect 7630 -6047 7664 -5749
rect 7726 -6047 7760 -5749
rect 7822 -6047 7856 -5749
rect 7918 -6047 7952 -5749
rect 8098 -6047 8132 -5749
rect 8194 -6047 8228 -5749
rect 8290 -6047 8324 -5749
rect 8386 -6047 8420 -5749
rect 8482 -6047 8516 -5749
rect 8578 -6047 8612 -5749
rect 8674 -6047 8708 -5749
rect 8770 -6047 8804 -5749
rect 8866 -6047 8900 -5749
rect 9034 -6047 9068 -5749
rect 9130 -6047 9164 -5749
rect 9226 -6047 9260 -5749
rect 9322 -6047 9356 -5749
rect 9418 -6047 9452 -5749
rect 9514 -6047 9548 -5749
rect 9610 -6047 9644 -5749
rect 9706 -6047 9740 -5749
rect 9802 -6047 9836 -5749
rect 9965 -6047 9999 -5749
rect 10061 -6047 10095 -5749
rect 10157 -6047 10191 -5749
rect 10253 -6047 10287 -5749
rect 10349 -6047 10383 -5749
rect 10445 -6047 10479 -5749
rect 10541 -6047 10575 -5749
rect 10637 -6047 10671 -5749
rect 10733 -6047 10767 -5749
rect 10892 -6047 10926 -5749
rect 10988 -6047 11022 -5749
rect 11084 -6047 11118 -5749
rect 11180 -6047 11214 -5749
rect 11276 -6047 11310 -5749
rect 11372 -6047 11406 -5749
rect 11468 -6047 11502 -5749
rect 11564 -6047 11598 -5749
rect 11660 -6047 11694 -5749
rect -24384 -7692 -24350 -7502
rect -24288 -7692 -24254 -7502
rect -24192 -7692 -24158 -7502
rect -24096 -7692 -24062 -7502
rect -24000 -7692 -23966 -7502
rect -23904 -7692 -23870 -7502
rect -23808 -7692 -23774 -7502
rect -23572 -7430 -23382 -7396
rect -23572 -7526 -23378 -7492
rect -23572 -7622 -23382 -7588
rect -23572 -7718 -23378 -7684
rect -22647 -7692 -22613 -7502
rect -22551 -7692 -22517 -7502
rect -22455 -7692 -22421 -7502
rect -22359 -7692 -22325 -7502
rect -22263 -7692 -22229 -7502
rect -22167 -7692 -22133 -7502
rect -22071 -7692 -22037 -7502
rect -21838 -7430 -21648 -7396
rect -21838 -7526 -21644 -7492
rect -21838 -7622 -21648 -7588
rect -21838 -7718 -21644 -7684
rect -20725 -7787 -20691 -7261
rect -20637 -7787 -20603 -7261
rect -20541 -7787 -20507 -7261
rect -20445 -7787 -20411 -7261
rect -20349 -7787 -20315 -7261
rect -20253 -7787 -20219 -7261
rect -20157 -7787 -20123 -7261
rect -20061 -7787 -20027 -7261
rect -19965 -7787 -19931 -7261
rect -19869 -7787 -19835 -7261
rect -19773 -7787 -19739 -7261
rect -19677 -7787 -19643 -7261
rect -19581 -7787 -19547 -7261
rect -19485 -7787 -19451 -7261
rect -19397 -7787 -19363 -7261
rect -19166 -7787 -19132 -7261
rect -19078 -7787 -19044 -7261
rect -18982 -7787 -18948 -7261
rect -18886 -7787 -18852 -7261
rect -18790 -7787 -18756 -7261
rect -18694 -7787 -18660 -7261
rect -18598 -7787 -18564 -7261
rect -18502 -7787 -18468 -7261
rect -18406 -7787 -18372 -7261
rect -18310 -7787 -18276 -7261
rect -18214 -7787 -18180 -7261
rect -18118 -7787 -18084 -7261
rect -18022 -7787 -17988 -7261
rect -17926 -7787 -17892 -7261
rect -17838 -7787 -17804 -7261
rect -17434 -7787 -17400 -7261
rect -17346 -7787 -17312 -7261
rect -17250 -7787 -17216 -7261
rect -17154 -7787 -17120 -7261
rect -17058 -7787 -17024 -7261
rect -16962 -7787 -16928 -7261
rect -16866 -7787 -16832 -7261
rect -16770 -7787 -16736 -7261
rect -16674 -7787 -16640 -7261
rect -16578 -7787 -16544 -7261
rect -16482 -7787 -16448 -7261
rect -16386 -7787 -16352 -7261
rect -16290 -7787 -16256 -7261
rect -16194 -7787 -16160 -7261
rect -16106 -7787 -16072 -7261
rect -15875 -7787 -15841 -7261
rect -15787 -7787 -15753 -7261
rect -15691 -7787 -15657 -7261
rect -15595 -7787 -15561 -7261
rect -15499 -7787 -15465 -7261
rect -15403 -7787 -15369 -7261
rect -15307 -7787 -15273 -7261
rect -15211 -7787 -15177 -7261
rect -15115 -7787 -15081 -7261
rect -15019 -7787 -14985 -7261
rect -14923 -7787 -14889 -7261
rect -14827 -7787 -14793 -7261
rect -14731 -7787 -14697 -7261
rect -14635 -7787 -14601 -7261
rect -14547 -7787 -14513 -7261
rect -14143 -7787 -14109 -7261
rect -14055 -7787 -14021 -7261
rect -13959 -7787 -13925 -7261
rect -13863 -7787 -13829 -7261
rect -13767 -7787 -13733 -7261
rect -13671 -7787 -13637 -7261
rect -13575 -7787 -13541 -7261
rect -13479 -7787 -13445 -7261
rect -13383 -7787 -13349 -7261
rect -13287 -7787 -13253 -7261
rect -13191 -7787 -13157 -7261
rect -13095 -7787 -13061 -7261
rect -12999 -7787 -12965 -7261
rect -12903 -7787 -12869 -7261
rect -12815 -7787 -12781 -7261
rect -12584 -7787 -12550 -7261
rect -12496 -7787 -12462 -7261
rect -12400 -7787 -12366 -7261
rect -12304 -7787 -12270 -7261
rect -12208 -7787 -12174 -7261
rect -12112 -7787 -12078 -7261
rect -12016 -7787 -11982 -7261
rect -11920 -7787 -11886 -7261
rect -11824 -7787 -11790 -7261
rect -11728 -7787 -11694 -7261
rect -11632 -7787 -11598 -7261
rect -11536 -7787 -11502 -7261
rect -11440 -7787 -11406 -7261
rect -11344 -7787 -11310 -7261
rect -11256 -7787 -11222 -7261
rect -10852 -7787 -10818 -7261
rect -10764 -7787 -10730 -7261
rect -10668 -7787 -10634 -7261
rect -10572 -7787 -10538 -7261
rect -10476 -7787 -10442 -7261
rect -10380 -7787 -10346 -7261
rect -10284 -7787 -10250 -7261
rect -10188 -7787 -10154 -7261
rect -10092 -7787 -10058 -7261
rect -9996 -7787 -9962 -7261
rect -9900 -7787 -9866 -7261
rect -9804 -7787 -9770 -7261
rect -9708 -7787 -9674 -7261
rect -9612 -7787 -9578 -7261
rect -9524 -7787 -9490 -7261
rect -9293 -7787 -9259 -7261
rect -9205 -7787 -9171 -7261
rect -9109 -7787 -9075 -7261
rect -9013 -7787 -8979 -7261
rect -8917 -7787 -8883 -7261
rect -8821 -7787 -8787 -7261
rect -8725 -7787 -8691 -7261
rect -8629 -7787 -8595 -7261
rect -8533 -7787 -8499 -7261
rect -8437 -7787 -8403 -7261
rect -8341 -7787 -8307 -7261
rect -8245 -7787 -8211 -7261
rect -8149 -7787 -8115 -7261
rect -8053 -7787 -8019 -7261
rect -7965 -7787 -7931 -7261
rect 11785 -7191 11819 -6959
rect 11881 -7191 11915 -6959
rect 11977 -7191 12011 -6959
rect 12073 -7191 12107 -6959
rect 12169 -7191 12203 -6959
rect 12265 -7191 12299 -6959
rect 12361 -7191 12395 -6959
rect 12457 -7191 12491 -6959
rect 12553 -7191 12587 -6959
rect 12649 -7191 12683 -6959
rect 12745 -7191 12779 -6959
rect 12935 -7097 13125 -7063
rect 12935 -7193 13129 -7159
rect 12935 -7289 13125 -7255
rect 12935 -7385 13129 -7351
rect -24384 -8984 -24350 -8794
rect -24288 -8984 -24254 -8794
rect -24192 -8984 -24158 -8794
rect -24096 -8984 -24062 -8794
rect -24000 -8984 -23966 -8794
rect -23904 -8984 -23870 -8794
rect -23808 -8984 -23774 -8794
rect -23571 -8722 -23381 -8688
rect -23571 -8818 -23377 -8784
rect -23571 -8914 -23381 -8880
rect -23571 -9010 -23377 -8976
rect -22648 -8984 -22614 -8794
rect -22552 -8984 -22518 -8794
rect -22456 -8984 -22422 -8794
rect -22360 -8984 -22326 -8794
rect -22264 -8984 -22230 -8794
rect -22168 -8984 -22134 -8794
rect -22072 -8984 -22038 -8794
rect -21834 -8722 -21644 -8688
rect -21834 -8818 -21640 -8784
rect -21834 -8914 -21644 -8880
rect 7150 -8911 7184 -8613
rect 7246 -8911 7280 -8613
rect 7342 -8911 7376 -8613
rect 7438 -8911 7472 -8613
rect 7534 -8911 7568 -8613
rect 7630 -8911 7664 -8613
rect 7726 -8911 7760 -8613
rect 7822 -8911 7856 -8613
rect 7918 -8911 7952 -8613
rect 8098 -8911 8132 -8613
rect 8194 -8911 8228 -8613
rect 8290 -8911 8324 -8613
rect 8386 -8911 8420 -8613
rect 8482 -8911 8516 -8613
rect 8578 -8911 8612 -8613
rect 8674 -8911 8708 -8613
rect 8770 -8911 8804 -8613
rect 8866 -8911 8900 -8613
rect 9034 -8911 9068 -8613
rect 9130 -8911 9164 -8613
rect 9226 -8911 9260 -8613
rect 9322 -8911 9356 -8613
rect 9418 -8911 9452 -8613
rect 9514 -8911 9548 -8613
rect 9610 -8911 9644 -8613
rect 9706 -8911 9740 -8613
rect 9802 -8911 9836 -8613
rect 9965 -8910 9999 -8612
rect 10061 -8910 10095 -8612
rect 10157 -8910 10191 -8612
rect 10253 -8910 10287 -8612
rect 10349 -8910 10383 -8612
rect 10445 -8910 10479 -8612
rect 10541 -8910 10575 -8612
rect 10637 -8910 10671 -8612
rect 10733 -8910 10767 -8612
rect 10892 -8911 10926 -8613
rect 10988 -8911 11022 -8613
rect 11084 -8911 11118 -8613
rect 11180 -8911 11214 -8613
rect 11276 -8911 11310 -8613
rect 11372 -8911 11406 -8613
rect 11468 -8911 11502 -8613
rect 11564 -8911 11598 -8613
rect 11660 -8911 11694 -8613
rect -21834 -9010 -21640 -8976
rect -20518 -9152 -20484 -8962
rect -20422 -9152 -20388 -8962
rect -20326 -9152 -20292 -8962
rect -20230 -9152 -20196 -8962
rect -20134 -9152 -20100 -8962
rect -20038 -9152 -20004 -8962
rect -19942 -9152 -19908 -8962
rect -19409 -9152 -19375 -8962
rect -19313 -9152 -19279 -8962
rect -19217 -9152 -19183 -8962
rect -19121 -9152 -19087 -8962
rect -19025 -9152 -18991 -8962
rect -18929 -9152 -18895 -8962
rect -18833 -9152 -18799 -8962
rect -18527 -9152 -18493 -8962
rect -18431 -9152 -18397 -8962
rect -18335 -9152 -18301 -8962
rect -18239 -9152 -18205 -8962
rect -18143 -9152 -18109 -8962
rect -18047 -9152 -18013 -8962
rect -17951 -9152 -17917 -8962
rect -17227 -9152 -17193 -8962
rect -17131 -9152 -17097 -8962
rect -17035 -9152 -17001 -8962
rect -16939 -9152 -16905 -8962
rect -16843 -9152 -16809 -8962
rect -16747 -9152 -16713 -8962
rect -16651 -9152 -16617 -8962
rect -16118 -9152 -16084 -8962
rect -16022 -9152 -15988 -8962
rect -15926 -9152 -15892 -8962
rect -15830 -9152 -15796 -8962
rect -15734 -9152 -15700 -8962
rect -15638 -9152 -15604 -8962
rect -15542 -9152 -15508 -8962
rect -15236 -9152 -15202 -8962
rect -15140 -9152 -15106 -8962
rect -15044 -9152 -15010 -8962
rect -14948 -9152 -14914 -8962
rect -14852 -9152 -14818 -8962
rect -14756 -9152 -14722 -8962
rect -14660 -9152 -14626 -8962
rect -13936 -9152 -13902 -8962
rect -13840 -9152 -13806 -8962
rect -13744 -9152 -13710 -8962
rect -13648 -9152 -13614 -8962
rect -13552 -9152 -13518 -8962
rect -13456 -9152 -13422 -8962
rect -13360 -9152 -13326 -8962
rect -12827 -9152 -12793 -8962
rect -12731 -9152 -12697 -8962
rect -12635 -9152 -12601 -8962
rect -12539 -9152 -12505 -8962
rect -12443 -9152 -12409 -8962
rect -12347 -9152 -12313 -8962
rect -12251 -9152 -12217 -8962
rect -11945 -9152 -11911 -8962
rect -11849 -9152 -11815 -8962
rect -11753 -9152 -11719 -8962
rect -11657 -9152 -11623 -8962
rect -11561 -9152 -11527 -8962
rect -11465 -9152 -11431 -8962
rect -11369 -9152 -11335 -8962
rect -10645 -9152 -10611 -8962
rect -10549 -9152 -10515 -8962
rect -10453 -9152 -10419 -8962
rect -10357 -9152 -10323 -8962
rect -10261 -9152 -10227 -8962
rect -10165 -9152 -10131 -8962
rect -10069 -9152 -10035 -8962
rect -9536 -9152 -9502 -8962
rect -9440 -9152 -9406 -8962
rect -9344 -9152 -9310 -8962
rect -9248 -9152 -9214 -8962
rect -9152 -9152 -9118 -8962
rect -9056 -9152 -9022 -8962
rect -8960 -9152 -8926 -8962
rect -8654 -9152 -8620 -8962
rect -8558 -9152 -8524 -8962
rect -8462 -9152 -8428 -8962
rect -8366 -9152 -8332 -8962
rect -8270 -9152 -8236 -8962
rect -8174 -9152 -8140 -8962
rect -8078 -9152 -8044 -8962
rect 5670 -9707 5860 -9673
rect 5670 -9803 5864 -9769
rect 5670 -9899 5860 -9865
rect 5670 -9995 5864 -9961
rect 6110 -9707 6300 -9673
rect 6110 -9803 6304 -9769
rect 6110 -9899 6300 -9865
rect 6110 -9995 6304 -9961
rect 6550 -9707 6740 -9673
rect 6550 -9803 6744 -9769
rect 6550 -9899 6740 -9865
rect 6550 -9995 6744 -9961
rect -24384 -10956 -24350 -10766
rect -24288 -10956 -24254 -10766
rect -24192 -10956 -24158 -10766
rect -24096 -10956 -24062 -10766
rect -24000 -10956 -23966 -10766
rect -23904 -10956 -23870 -10766
rect -23808 -10956 -23774 -10766
rect -23571 -10694 -23381 -10660
rect -23571 -10790 -23377 -10756
rect -23571 -10886 -23381 -10852
rect -23571 -10982 -23377 -10948
rect -22647 -10956 -22613 -10766
rect -22551 -10956 -22517 -10766
rect -22455 -10956 -22421 -10766
rect -22359 -10956 -22325 -10766
rect -22263 -10956 -22229 -10766
rect -22167 -10956 -22133 -10766
rect -22071 -10956 -22037 -10766
rect -21838 -10694 -21648 -10660
rect -21838 -10790 -21644 -10756
rect -21838 -10886 -21648 -10852
rect -21838 -10982 -21644 -10948
rect -20725 -11051 -20691 -10525
rect -20637 -11051 -20603 -10525
rect -20541 -11051 -20507 -10525
rect -20445 -11051 -20411 -10525
rect -20349 -11051 -20315 -10525
rect -20253 -11051 -20219 -10525
rect -20157 -11051 -20123 -10525
rect -20061 -11051 -20027 -10525
rect -19965 -11051 -19931 -10525
rect -19869 -11051 -19835 -10525
rect -19773 -11051 -19739 -10525
rect -19677 -11051 -19643 -10525
rect -19581 -11051 -19547 -10525
rect -19485 -11051 -19451 -10525
rect -19397 -11051 -19363 -10525
rect -19166 -11051 -19132 -10525
rect -19078 -11051 -19044 -10525
rect -18982 -11051 -18948 -10525
rect -18886 -11051 -18852 -10525
rect -18790 -11051 -18756 -10525
rect -18694 -11051 -18660 -10525
rect -18598 -11051 -18564 -10525
rect -18502 -11051 -18468 -10525
rect -18406 -11051 -18372 -10525
rect -18310 -11051 -18276 -10525
rect -18214 -11051 -18180 -10525
rect -18118 -11051 -18084 -10525
rect -18022 -11051 -17988 -10525
rect -17926 -11051 -17892 -10525
rect -17838 -11051 -17804 -10525
rect -17434 -11051 -17400 -10525
rect -17346 -11051 -17312 -10525
rect -17250 -11051 -17216 -10525
rect -17154 -11051 -17120 -10525
rect -17058 -11051 -17024 -10525
rect -16962 -11051 -16928 -10525
rect -16866 -11051 -16832 -10525
rect -16770 -11051 -16736 -10525
rect -16674 -11051 -16640 -10525
rect -16578 -11051 -16544 -10525
rect -16482 -11051 -16448 -10525
rect -16386 -11051 -16352 -10525
rect -16290 -11051 -16256 -10525
rect -16194 -11051 -16160 -10525
rect -16106 -11051 -16072 -10525
rect -15875 -11051 -15841 -10525
rect -15787 -11051 -15753 -10525
rect -15691 -11051 -15657 -10525
rect -15595 -11051 -15561 -10525
rect -15499 -11051 -15465 -10525
rect -15403 -11051 -15369 -10525
rect -15307 -11051 -15273 -10525
rect -15211 -11051 -15177 -10525
rect -15115 -11051 -15081 -10525
rect -15019 -11051 -14985 -10525
rect -14923 -11051 -14889 -10525
rect -14827 -11051 -14793 -10525
rect -14731 -11051 -14697 -10525
rect -14635 -11051 -14601 -10525
rect -14547 -11051 -14513 -10525
rect -14143 -11051 -14109 -10525
rect -14055 -11051 -14021 -10525
rect -13959 -11051 -13925 -10525
rect -13863 -11051 -13829 -10525
rect -13767 -11051 -13733 -10525
rect -13671 -11051 -13637 -10525
rect -13575 -11051 -13541 -10525
rect -13479 -11051 -13445 -10525
rect -13383 -11051 -13349 -10525
rect -13287 -11051 -13253 -10525
rect -13191 -11051 -13157 -10525
rect -13095 -11051 -13061 -10525
rect -12999 -11051 -12965 -10525
rect -12903 -11051 -12869 -10525
rect -12815 -11051 -12781 -10525
rect -12584 -11051 -12550 -10525
rect -12496 -11051 -12462 -10525
rect -12400 -11051 -12366 -10525
rect -12304 -11051 -12270 -10525
rect -12208 -11051 -12174 -10525
rect -12112 -11051 -12078 -10525
rect -12016 -11051 -11982 -10525
rect -11920 -11051 -11886 -10525
rect -11824 -11051 -11790 -10525
rect -11728 -11051 -11694 -10525
rect -11632 -11051 -11598 -10525
rect -11536 -11051 -11502 -10525
rect -11440 -11051 -11406 -10525
rect -11344 -11051 -11310 -10525
rect -11256 -11051 -11222 -10525
rect -10852 -11051 -10818 -10525
rect -10764 -11051 -10730 -10525
rect -10668 -11051 -10634 -10525
rect -10572 -11051 -10538 -10525
rect -10476 -11051 -10442 -10525
rect -10380 -11051 -10346 -10525
rect -10284 -11051 -10250 -10525
rect -10188 -11051 -10154 -10525
rect -10092 -11051 -10058 -10525
rect -9996 -11051 -9962 -10525
rect -9900 -11051 -9866 -10525
rect -9804 -11051 -9770 -10525
rect -9708 -11051 -9674 -10525
rect -9612 -11051 -9578 -10525
rect -9524 -11051 -9490 -10525
rect -9293 -11051 -9259 -10525
rect -9205 -11051 -9171 -10525
rect -9109 -11051 -9075 -10525
rect -9013 -11051 -8979 -10525
rect -8917 -11051 -8883 -10525
rect -8821 -11051 -8787 -10525
rect -8725 -11051 -8691 -10525
rect -8629 -11051 -8595 -10525
rect -8533 -11051 -8499 -10525
rect -8437 -11051 -8403 -10525
rect -8341 -11051 -8307 -10525
rect -8245 -11051 -8211 -10525
rect -8149 -11051 -8115 -10525
rect -8053 -11051 -8019 -10525
rect -7965 -11051 -7931 -10525
rect 7150 -10675 7184 -10377
rect 7246 -10675 7280 -10377
rect 7342 -10675 7376 -10377
rect 7438 -10675 7472 -10377
rect 7534 -10675 7568 -10377
rect 7630 -10675 7664 -10377
rect 7726 -10675 7760 -10377
rect 7822 -10675 7856 -10377
rect 7918 -10675 7952 -10377
rect 8098 -10675 8132 -10377
rect 8194 -10675 8228 -10377
rect 8290 -10675 8324 -10377
rect 8386 -10675 8420 -10377
rect 8482 -10675 8516 -10377
rect 8578 -10675 8612 -10377
rect 8674 -10675 8708 -10377
rect 8770 -10675 8804 -10377
rect 8866 -10675 8900 -10377
rect 9034 -10675 9068 -10377
rect 9130 -10675 9164 -10377
rect 9226 -10675 9260 -10377
rect 9322 -10675 9356 -10377
rect 9418 -10675 9452 -10377
rect 9514 -10675 9548 -10377
rect 9610 -10675 9644 -10377
rect 9706 -10675 9740 -10377
rect 9802 -10675 9836 -10377
rect 9965 -10675 9999 -10377
rect 10061 -10675 10095 -10377
rect 10157 -10675 10191 -10377
rect 10253 -10675 10287 -10377
rect 10349 -10675 10383 -10377
rect 10445 -10675 10479 -10377
rect 10541 -10675 10575 -10377
rect 10637 -10675 10671 -10377
rect 10733 -10675 10767 -10377
rect 10892 -10675 10926 -10377
rect 10988 -10675 11022 -10377
rect 11084 -10675 11118 -10377
rect 11180 -10675 11214 -10377
rect 11276 -10675 11310 -10377
rect 11372 -10675 11406 -10377
rect 11468 -10675 11502 -10377
rect 11564 -10675 11598 -10377
rect 11660 -10675 11694 -10377
rect 11785 -11819 11819 -11587
rect 11881 -11819 11915 -11587
rect 11977 -11819 12011 -11587
rect 12073 -11819 12107 -11587
rect 12169 -11819 12203 -11587
rect 12265 -11819 12299 -11587
rect 12361 -11819 12395 -11587
rect 12457 -11819 12491 -11587
rect 12553 -11819 12587 -11587
rect 12649 -11819 12683 -11587
rect 12745 -11819 12779 -11587
rect -24384 -12248 -24350 -12058
rect -24288 -12248 -24254 -12058
rect -24192 -12248 -24158 -12058
rect -24096 -12248 -24062 -12058
rect -24000 -12248 -23966 -12058
rect -23904 -12248 -23870 -12058
rect -23808 -12248 -23774 -12058
rect -23571 -11986 -23381 -11952
rect -23571 -12082 -23377 -12048
rect -23571 -12178 -23381 -12144
rect -23571 -12274 -23377 -12240
rect -22647 -12248 -22613 -12058
rect -22551 -12248 -22517 -12058
rect -22455 -12248 -22421 -12058
rect -22359 -12248 -22325 -12058
rect -22263 -12248 -22229 -12058
rect -22167 -12248 -22133 -12058
rect -22071 -12248 -22037 -12058
rect -21842 -11986 -21652 -11952
rect -21842 -12082 -21648 -12048
rect -21842 -12178 -21652 -12144
rect -21842 -12274 -21648 -12240
rect -20518 -12416 -20484 -12226
rect -20422 -12416 -20388 -12226
rect -20326 -12416 -20292 -12226
rect -20230 -12416 -20196 -12226
rect -20134 -12416 -20100 -12226
rect -20038 -12416 -20004 -12226
rect -19942 -12416 -19908 -12226
rect -19409 -12416 -19375 -12226
rect -19313 -12416 -19279 -12226
rect -19217 -12416 -19183 -12226
rect -19121 -12416 -19087 -12226
rect -19025 -12416 -18991 -12226
rect -18929 -12416 -18895 -12226
rect -18833 -12416 -18799 -12226
rect -18527 -12416 -18493 -12226
rect -18431 -12416 -18397 -12226
rect -18335 -12416 -18301 -12226
rect -18239 -12416 -18205 -12226
rect -18143 -12416 -18109 -12226
rect -18047 -12416 -18013 -12226
rect -17951 -12416 -17917 -12226
rect -17227 -12416 -17193 -12226
rect -17131 -12416 -17097 -12226
rect -17035 -12416 -17001 -12226
rect -16939 -12416 -16905 -12226
rect -16843 -12416 -16809 -12226
rect -16747 -12416 -16713 -12226
rect -16651 -12416 -16617 -12226
rect -16118 -12416 -16084 -12226
rect -16022 -12416 -15988 -12226
rect -15926 -12416 -15892 -12226
rect -15830 -12416 -15796 -12226
rect -15734 -12416 -15700 -12226
rect -15638 -12416 -15604 -12226
rect -15542 -12416 -15508 -12226
rect -15236 -12416 -15202 -12226
rect -15140 -12416 -15106 -12226
rect -15044 -12416 -15010 -12226
rect -14948 -12416 -14914 -12226
rect -14852 -12416 -14818 -12226
rect -14756 -12416 -14722 -12226
rect -14660 -12416 -14626 -12226
rect -13936 -12416 -13902 -12226
rect -13840 -12416 -13806 -12226
rect -13744 -12416 -13710 -12226
rect -13648 -12416 -13614 -12226
rect -13552 -12416 -13518 -12226
rect -13456 -12416 -13422 -12226
rect -13360 -12416 -13326 -12226
rect -12827 -12416 -12793 -12226
rect -12731 -12416 -12697 -12226
rect -12635 -12416 -12601 -12226
rect -12539 -12416 -12505 -12226
rect -12443 -12416 -12409 -12226
rect -12347 -12416 -12313 -12226
rect -12251 -12416 -12217 -12226
rect -11945 -12416 -11911 -12226
rect -11849 -12416 -11815 -12226
rect -11753 -12416 -11719 -12226
rect -11657 -12416 -11623 -12226
rect -11561 -12416 -11527 -12226
rect -11465 -12416 -11431 -12226
rect -11369 -12416 -11335 -12226
rect -10645 -12416 -10611 -12226
rect -10549 -12416 -10515 -12226
rect -10453 -12416 -10419 -12226
rect -10357 -12416 -10323 -12226
rect -10261 -12416 -10227 -12226
rect -10165 -12416 -10131 -12226
rect -10069 -12416 -10035 -12226
rect -9536 -12416 -9502 -12226
rect -9440 -12416 -9406 -12226
rect -9344 -12416 -9310 -12226
rect -9248 -12416 -9214 -12226
rect -9152 -12416 -9118 -12226
rect -9056 -12416 -9022 -12226
rect -8960 -12416 -8926 -12226
rect -8654 -12416 -8620 -12226
rect -8558 -12416 -8524 -12226
rect -8462 -12416 -8428 -12226
rect -8366 -12416 -8332 -12226
rect -8270 -12416 -8236 -12226
rect -8174 -12416 -8140 -12226
rect -8078 -12416 -8044 -12226
rect 12935 -11725 13125 -11691
rect 12935 -11821 13129 -11787
rect 12935 -11917 13125 -11883
rect 12935 -12013 13129 -11979
rect 7150 -13539 7184 -13241
rect 7246 -13539 7280 -13241
rect 7342 -13539 7376 -13241
rect 7438 -13539 7472 -13241
rect 7534 -13539 7568 -13241
rect 7630 -13539 7664 -13241
rect 7726 -13539 7760 -13241
rect 7822 -13539 7856 -13241
rect 7918 -13539 7952 -13241
rect 8098 -13539 8132 -13241
rect 8194 -13539 8228 -13241
rect 8290 -13539 8324 -13241
rect 8386 -13539 8420 -13241
rect 8482 -13539 8516 -13241
rect 8578 -13539 8612 -13241
rect 8674 -13539 8708 -13241
rect 8770 -13539 8804 -13241
rect 8866 -13539 8900 -13241
rect 9034 -13539 9068 -13241
rect 9130 -13539 9164 -13241
rect 9226 -13539 9260 -13241
rect 9322 -13539 9356 -13241
rect 9418 -13539 9452 -13241
rect 9514 -13539 9548 -13241
rect 9610 -13539 9644 -13241
rect 9706 -13539 9740 -13241
rect 9802 -13539 9836 -13241
rect 9965 -13538 9999 -13240
rect 10061 -13538 10095 -13240
rect 10157 -13538 10191 -13240
rect 10253 -13538 10287 -13240
rect 10349 -13538 10383 -13240
rect 10445 -13538 10479 -13240
rect 10541 -13538 10575 -13240
rect 10637 -13538 10671 -13240
rect 10733 -13538 10767 -13240
rect 10892 -13539 10926 -13241
rect 10988 -13539 11022 -13241
rect 11084 -13539 11118 -13241
rect 11180 -13539 11214 -13241
rect 11276 -13539 11310 -13241
rect 11372 -13539 11406 -13241
rect 11468 -13539 11502 -13241
rect 11564 -13539 11598 -13241
rect 11660 -13539 11694 -13241
rect -2100 -14020 -2066 -13830
rect -2004 -14020 -1970 -13826
rect -1908 -14020 -1874 -13830
rect -1812 -14020 -1778 -13826
rect -12304 -14139 -11778 -14105
rect -17665 -14545 -17433 -14511
rect -17665 -14641 -17433 -14607
rect -17665 -14737 -17433 -14703
rect -17665 -14833 -17433 -14799
rect -24437 -14962 -24247 -14928
rect -24437 -15058 -24247 -15024
rect -24437 -15154 -24247 -15120
rect -24437 -15250 -24247 -15216
rect -24437 -15346 -24247 -15312
rect -17665 -14929 -17433 -14895
rect -17665 -15025 -17433 -14991
rect -24437 -15442 -24247 -15408
rect -17665 -15121 -17433 -15087
rect -17665 -15217 -17433 -15183
rect -17665 -15313 -17433 -15279
rect -17665 -15409 -17433 -15375
rect -12304 -14227 -11778 -14193
rect -12304 -14323 -11778 -14289
rect -12304 -14419 -11778 -14385
rect -12304 -14515 -11778 -14481
rect -12304 -14611 -11778 -14577
rect -12304 -14707 -11778 -14673
rect -12304 -14803 -11778 -14769
rect -12304 -14899 -11778 -14865
rect -12304 -14995 -11778 -14961
rect -12304 -15091 -11778 -15057
rect -12304 -15187 -11778 -15153
rect -12304 -15283 -11778 -15249
rect -12304 -15379 -11778 -15345
rect -4816 -14405 -4782 -14215
rect -4720 -14409 -4686 -14215
rect -4624 -14405 -4590 -14215
rect -4528 -14409 -4494 -14215
rect -2100 -14399 -2066 -14209
rect -2004 -14399 -1970 -14205
rect -1908 -14399 -1874 -14209
rect -1812 -14399 -1778 -14205
rect 5670 -14235 5860 -14201
rect 5670 -14331 5864 -14297
rect 5670 -14427 5860 -14393
rect 5670 -14523 5864 -14489
rect 6110 -14235 6300 -14201
rect 6110 -14331 6304 -14297
rect 6110 -14427 6300 -14393
rect 6110 -14523 6304 -14489
rect 6550 -14235 6740 -14201
rect 6550 -14331 6744 -14297
rect 6550 -14427 6740 -14393
rect 6550 -14523 6744 -14489
rect -4816 -14845 -4782 -14655
rect -4720 -14849 -4686 -14655
rect -4624 -14845 -4590 -14655
rect -4528 -14849 -4494 -14655
rect -2100 -14839 -2066 -14649
rect -2004 -14839 -1970 -14645
rect -1908 -14839 -1874 -14649
rect -1812 -14839 -1778 -14645
rect -4816 -15224 -4782 -15034
rect -4720 -15228 -4686 -15034
rect -4624 -15224 -4590 -15034
rect -4528 -15228 -4494 -15034
rect -2100 -15218 -2066 -15028
rect -2004 -15218 -1970 -15024
rect -1908 -15218 -1874 -15028
rect -1812 -15218 -1778 -15024
rect 7150 -15203 7184 -14905
rect 7246 -15203 7280 -14905
rect 7342 -15203 7376 -14905
rect 7438 -15203 7472 -14905
rect 7534 -15203 7568 -14905
rect 7630 -15203 7664 -14905
rect 7726 -15203 7760 -14905
rect 7822 -15203 7856 -14905
rect 7918 -15203 7952 -14905
rect 8098 -15203 8132 -14905
rect 8194 -15203 8228 -14905
rect 8290 -15203 8324 -14905
rect 8386 -15203 8420 -14905
rect 8482 -15203 8516 -14905
rect 8578 -15203 8612 -14905
rect 8674 -15203 8708 -14905
rect 8770 -15203 8804 -14905
rect 8866 -15203 8900 -14905
rect 9034 -15203 9068 -14905
rect 9130 -15203 9164 -14905
rect 9226 -15203 9260 -14905
rect 9322 -15203 9356 -14905
rect 9418 -15203 9452 -14905
rect 9514 -15203 9548 -14905
rect 9610 -15203 9644 -14905
rect 9706 -15203 9740 -14905
rect 9802 -15203 9836 -14905
rect 9965 -15203 9999 -14905
rect 10061 -15203 10095 -14905
rect 10157 -15203 10191 -14905
rect 10253 -15203 10287 -14905
rect 10349 -15203 10383 -14905
rect 10445 -15203 10479 -14905
rect 10541 -15203 10575 -14905
rect 10637 -15203 10671 -14905
rect 10733 -15203 10767 -14905
rect 10892 -15203 10926 -14905
rect 10988 -15203 11022 -14905
rect 11084 -15203 11118 -14905
rect 11180 -15203 11214 -14905
rect 11276 -15203 11310 -14905
rect 11372 -15203 11406 -14905
rect 11468 -15203 11502 -14905
rect 11564 -15203 11598 -14905
rect 11660 -15203 11694 -14905
rect -24437 -15538 -24247 -15504
rect -17665 -15505 -17433 -15471
rect -12304 -15467 -11778 -15433
rect -8167 -15548 -8133 -15358
rect -8071 -15548 -8037 -15354
rect -7975 -15548 -7941 -15358
rect -7879 -15548 -7845 -15354
rect -4816 -15664 -4782 -15474
rect -4720 -15668 -4686 -15474
rect -4624 -15664 -4590 -15474
rect -4528 -15668 -4494 -15474
rect -2100 -15658 -2066 -15468
rect -2004 -15658 -1970 -15464
rect -1908 -15658 -1874 -15468
rect -1812 -15658 -1778 -15464
rect -17665 -15945 -17433 -15911
rect -17665 -16041 -17433 -16007
rect -8166 -16048 -8132 -15858
rect -8070 -16048 -8036 -15854
rect -7974 -16048 -7940 -15858
rect -7878 -16048 -7844 -15854
rect -4816 -16043 -4782 -15853
rect -4720 -16047 -4686 -15853
rect -4624 -16043 -4590 -15853
rect -4528 -16047 -4494 -15853
rect -24436 -16147 -24246 -16113
rect -24436 -16243 -24246 -16209
rect -24436 -16339 -24246 -16305
rect -24436 -16435 -24246 -16401
rect -24436 -16531 -24246 -16497
rect -17665 -16137 -17433 -16103
rect -2100 -16037 -2066 -15847
rect -2004 -16037 -1970 -15843
rect -1908 -16037 -1874 -15847
rect -1812 -16037 -1778 -15843
rect -17665 -16233 -17433 -16199
rect -17665 -16329 -17433 -16295
rect -17665 -16425 -17433 -16391
rect -24436 -16627 -24246 -16593
rect -24436 -16723 -24246 -16689
rect -17665 -16521 -17433 -16487
rect -8167 -16528 -8133 -16338
rect -8071 -16528 -8037 -16334
rect -7975 -16528 -7941 -16338
rect -7879 -16528 -7845 -16334
rect -4816 -16483 -4782 -16293
rect -4720 -16487 -4686 -16293
rect -4624 -16483 -4590 -16293
rect -4528 -16487 -4494 -16293
rect -2100 -16477 -2066 -16287
rect -2004 -16477 -1970 -16283
rect -1908 -16477 -1874 -16287
rect -1812 -16477 -1778 -16283
rect 11785 -16347 11819 -16115
rect 11881 -16347 11915 -16115
rect 11977 -16347 12011 -16115
rect 12073 -16347 12107 -16115
rect 12169 -16347 12203 -16115
rect 12265 -16347 12299 -16115
rect 12361 -16347 12395 -16115
rect 12457 -16347 12491 -16115
rect 12553 -16347 12587 -16115
rect 12649 -16347 12683 -16115
rect 12745 -16347 12779 -16115
rect -17665 -16617 -17433 -16583
rect -17665 -16713 -17433 -16679
rect -17665 -16809 -17433 -16775
rect -17665 -16905 -17433 -16871
rect -12302 -16955 -11776 -16921
rect -24431 -17360 -24241 -17326
rect -24431 -17456 -24241 -17422
rect -24431 -17552 -24241 -17518
rect -24431 -17648 -24241 -17614
rect -24431 -17744 -24241 -17710
rect -17665 -17345 -17433 -17311
rect -17665 -17441 -17433 -17407
rect -17665 -17537 -17433 -17503
rect -17665 -17633 -17433 -17599
rect -24431 -17840 -24241 -17806
rect -17665 -17729 -17433 -17695
rect -17665 -17825 -17433 -17791
rect -24431 -17936 -24241 -17902
rect -21606 -18236 -21572 -18046
rect -21510 -18236 -21476 -18042
rect -21414 -18236 -21380 -18046
rect -21318 -18236 -21284 -18042
rect -17665 -17921 -17433 -17887
rect -17665 -18017 -17433 -17983
rect -17665 -18113 -17433 -18079
rect -16015 -18107 -15981 -17917
rect -15919 -18107 -15885 -17913
rect -15823 -18107 -15789 -17917
rect -15727 -18107 -15693 -17913
rect -17665 -18209 -17433 -18175
rect -12302 -17043 -11776 -17009
rect -12302 -17139 -11776 -17105
rect -12302 -17235 -11776 -17201
rect -12302 -17331 -11776 -17297
rect -12302 -17427 -11776 -17393
rect -12302 -17523 -11776 -17489
rect -12302 -17619 -11776 -17585
rect -12302 -17715 -11776 -17681
rect -12302 -17811 -11776 -17777
rect -12302 -17907 -11776 -17873
rect -12302 -18003 -11776 -17969
rect -12302 -18099 -11776 -18065
rect -12302 -18195 -11776 -18161
rect -8167 -17028 -8133 -16838
rect -8071 -17028 -8037 -16834
rect -7975 -17028 -7941 -16838
rect -7879 -17028 -7845 -16834
rect -4816 -16862 -4782 -16672
rect -4720 -16866 -4686 -16672
rect -4624 -16862 -4590 -16672
rect -4528 -16866 -4494 -16672
rect -2100 -16856 -2066 -16666
rect -2004 -16856 -1970 -16662
rect -1908 -16856 -1874 -16666
rect -1812 -16856 -1778 -16662
rect -8167 -17508 -8133 -17318
rect -8071 -17508 -8037 -17314
rect -7975 -17508 -7941 -17318
rect -7879 -17508 -7845 -17314
rect -4816 -17302 -4782 -17112
rect -4720 -17306 -4686 -17112
rect -4624 -17302 -4590 -17112
rect -4528 -17306 -4494 -17112
rect -2100 -17296 -2066 -17106
rect -2004 -17296 -1970 -17102
rect -1908 -17296 -1874 -17106
rect -1812 -17296 -1778 -17102
rect -4816 -17681 -4782 -17491
rect -4720 -17685 -4686 -17491
rect -4624 -17681 -4590 -17491
rect -4528 -17685 -4494 -17491
rect -2100 -17675 -2066 -17485
rect -2004 -17675 -1970 -17481
rect -1908 -17675 -1874 -17485
rect -1812 -17675 -1778 -17481
rect -8167 -17968 -8133 -17778
rect -8071 -17968 -8037 -17774
rect -7975 -17968 -7941 -17778
rect -7879 -17968 -7845 -17774
rect 12935 -16253 13125 -16219
rect 12935 -16349 13129 -16315
rect 12935 -16445 13125 -16411
rect 12935 -16541 13129 -16507
rect -4816 -18121 -4782 -17931
rect -4720 -18125 -4686 -17931
rect -4624 -18121 -4590 -17931
rect -4528 -18125 -4494 -17931
rect -2100 -18115 -2066 -17925
rect -2004 -18115 -1970 -17921
rect -1908 -18115 -1874 -17925
rect -1812 -18115 -1778 -17921
rect 7150 -18067 7184 -17769
rect 7246 -18067 7280 -17769
rect 7342 -18067 7376 -17769
rect 7438 -18067 7472 -17769
rect 7534 -18067 7568 -17769
rect 7630 -18067 7664 -17769
rect 7726 -18067 7760 -17769
rect 7822 -18067 7856 -17769
rect 7918 -18067 7952 -17769
rect 8098 -18067 8132 -17769
rect 8194 -18067 8228 -17769
rect 8290 -18067 8324 -17769
rect 8386 -18067 8420 -17769
rect 8482 -18067 8516 -17769
rect 8578 -18067 8612 -17769
rect 8674 -18067 8708 -17769
rect 8770 -18067 8804 -17769
rect 8866 -18067 8900 -17769
rect 9034 -18067 9068 -17769
rect 9130 -18067 9164 -17769
rect 9226 -18067 9260 -17769
rect 9322 -18067 9356 -17769
rect 9418 -18067 9452 -17769
rect 9514 -18067 9548 -17769
rect 9610 -18067 9644 -17769
rect 9706 -18067 9740 -17769
rect 9802 -18067 9836 -17769
rect 9965 -18066 9999 -17768
rect 10061 -18066 10095 -17768
rect 10157 -18066 10191 -17768
rect 10253 -18066 10287 -17768
rect 10349 -18066 10383 -17768
rect 10445 -18066 10479 -17768
rect 10541 -18066 10575 -17768
rect 10637 -18066 10671 -17768
rect 10733 -18066 10767 -17768
rect 10892 -18067 10926 -17769
rect 10988 -18067 11022 -17769
rect 11084 -18067 11118 -17769
rect 11180 -18067 11214 -17769
rect 11276 -18067 11310 -17769
rect 11372 -18067 11406 -17769
rect 11468 -18067 11502 -17769
rect 11564 -18067 11598 -17769
rect 11660 -18067 11694 -17769
rect -17665 -18305 -17433 -18271
rect -12302 -18283 -11776 -18249
rect -24416 -18479 -24226 -18445
rect -24416 -18575 -24226 -18541
rect -24416 -18671 -24226 -18637
rect -24416 -18767 -24226 -18733
rect -24416 -18863 -24226 -18829
rect -21605 -18736 -21571 -18546
rect -21509 -18736 -21475 -18542
rect -21413 -18736 -21379 -18546
rect -21317 -18736 -21283 -18542
rect -16014 -18607 -15980 -18417
rect -15918 -18607 -15884 -18413
rect -15822 -18607 -15788 -18417
rect -15726 -18607 -15692 -18413
rect -8181 -18428 -8147 -18238
rect -8085 -18428 -8051 -18234
rect -7989 -18428 -7955 -18238
rect -7893 -18428 -7859 -18234
rect -4816 -18500 -4782 -18310
rect -4720 -18504 -4686 -18310
rect -4624 -18500 -4590 -18310
rect -4528 -18504 -4494 -18310
rect -2100 -18494 -2066 -18304
rect -2004 -18494 -1970 -18300
rect -1908 -18494 -1874 -18304
rect -1812 -18494 -1778 -18300
rect 15775 -18511 15809 -17679
rect 15871 -18511 15905 -17679
rect 15967 -18511 16001 -17679
rect 16063 -18511 16097 -17679
rect 16159 -18511 16193 -17679
rect 16255 -18511 16289 -17679
rect 16351 -18511 16385 -17679
rect 16447 -18511 16481 -17679
rect 16543 -18511 16577 -17679
rect 16639 -18511 16673 -17679
rect 16735 -18511 16769 -17679
rect 16831 -18511 16865 -17679
rect 16927 -18511 16961 -17679
rect 17306 -18477 17340 -18287
rect 17402 -18477 17436 -18287
rect 17498 -18477 17532 -18287
rect 17594 -18477 17628 -18287
rect 17690 -18477 17724 -18287
rect 17786 -18477 17820 -18287
rect 17882 -18477 17916 -18287
rect -17665 -18745 -17433 -18711
rect -24416 -18959 -24226 -18925
rect -17665 -18841 -17433 -18807
rect -17665 -18937 -17433 -18903
rect -24416 -19055 -24226 -19021
rect -21606 -19216 -21572 -19026
rect -21510 -19216 -21476 -19022
rect -21414 -19216 -21380 -19026
rect -21318 -19216 -21284 -19022
rect -17665 -19033 -17433 -18999
rect -17665 -19129 -17433 -19095
rect -17665 -19225 -17433 -19191
rect -16015 -19087 -15981 -18897
rect -15919 -19087 -15885 -18893
rect -15823 -19087 -15789 -18897
rect -15727 -19087 -15693 -18893
rect -8179 -18908 -8145 -18718
rect -8083 -18908 -8049 -18714
rect -7987 -18908 -7953 -18718
rect -7891 -18908 -7857 -18714
rect 18108 -18293 18298 -18259
rect 18108 -18389 18302 -18355
rect 18108 -18485 18298 -18451
rect 18108 -18581 18302 -18547
rect -4816 -18940 -4782 -18750
rect -4720 -18944 -4686 -18750
rect -4624 -18940 -4590 -18750
rect -4528 -18944 -4494 -18750
rect -2100 -18934 -2066 -18744
rect -2004 -18934 -1970 -18740
rect -1908 -18934 -1874 -18744
rect -1812 -18934 -1778 -18740
rect 5670 -18763 5860 -18729
rect 5670 -18859 5864 -18825
rect 5670 -18955 5860 -18921
rect 5670 -19051 5864 -19017
rect 6110 -18763 6300 -18729
rect 6110 -18859 6304 -18825
rect 6110 -18955 6300 -18921
rect 6110 -19051 6304 -19017
rect 6550 -18763 6740 -18729
rect 6550 -18859 6744 -18825
rect 6550 -18955 6740 -18921
rect 6550 -19051 6744 -19017
rect -24414 -19673 -24224 -19639
rect -24414 -19769 -24224 -19735
rect -24414 -19865 -24224 -19831
rect -24414 -19961 -24224 -19927
rect -24414 -20057 -24224 -20023
rect -21606 -19716 -21572 -19526
rect -21510 -19716 -21476 -19522
rect -21414 -19716 -21380 -19526
rect -21318 -19716 -21284 -19522
rect -17665 -19321 -17433 -19287
rect -4816 -19319 -4782 -19129
rect -4720 -19323 -4686 -19129
rect -4624 -19319 -4590 -19129
rect -4528 -19323 -4494 -19129
rect -2100 -19313 -2066 -19123
rect -2004 -19313 -1970 -19119
rect -1908 -19313 -1874 -19123
rect -1812 -19313 -1778 -19119
rect -17665 -19417 -17433 -19383
rect -17665 -19513 -17433 -19479
rect -17665 -19609 -17433 -19575
rect -16015 -19587 -15981 -19397
rect -15919 -19587 -15885 -19393
rect -15823 -19587 -15789 -19397
rect -15727 -19587 -15693 -19393
rect -17665 -19705 -17433 -19671
rect -4816 -19759 -4782 -19569
rect -4720 -19763 -4686 -19569
rect -4624 -19759 -4590 -19569
rect -4528 -19763 -4494 -19569
rect -2100 -19753 -2066 -19563
rect -2004 -19753 -1970 -19559
rect -1908 -19753 -1874 -19563
rect -1812 -19753 -1778 -19559
rect 7150 -19731 7184 -19433
rect 7246 -19731 7280 -19433
rect 7342 -19731 7376 -19433
rect 7438 -19731 7472 -19433
rect 7534 -19731 7568 -19433
rect 7630 -19731 7664 -19433
rect 7726 -19731 7760 -19433
rect 7822 -19731 7856 -19433
rect 7918 -19731 7952 -19433
rect 8098 -19731 8132 -19433
rect 8194 -19731 8228 -19433
rect 8290 -19731 8324 -19433
rect 8386 -19731 8420 -19433
rect 8482 -19731 8516 -19433
rect 8578 -19731 8612 -19433
rect 8674 -19731 8708 -19433
rect 8770 -19731 8804 -19433
rect 8866 -19731 8900 -19433
rect 9034 -19731 9068 -19433
rect 9130 -19731 9164 -19433
rect 9226 -19731 9260 -19433
rect 9322 -19731 9356 -19433
rect 9418 -19731 9452 -19433
rect 9514 -19731 9548 -19433
rect 9610 -19731 9644 -19433
rect 9706 -19731 9740 -19433
rect 9802 -19731 9836 -19433
rect 9965 -19731 9999 -19433
rect 10061 -19731 10095 -19433
rect 10157 -19731 10191 -19433
rect 10253 -19731 10287 -19433
rect 10349 -19731 10383 -19433
rect 10445 -19731 10479 -19433
rect 10541 -19731 10575 -19433
rect 10637 -19731 10671 -19433
rect 10733 -19731 10767 -19433
rect 10892 -19731 10926 -19433
rect 10988 -19731 11022 -19433
rect 11084 -19731 11118 -19433
rect 11180 -19731 11214 -19433
rect 11276 -19731 11310 -19433
rect 11372 -19731 11406 -19433
rect 11468 -19731 11502 -19433
rect 11564 -19731 11598 -19433
rect 11660 -19731 11694 -19433
rect 15775 -19493 15809 -18661
rect 15871 -19493 15905 -18661
rect 15967 -19493 16001 -18661
rect 16063 -19493 16097 -18661
rect 16159 -19493 16193 -18661
rect 16255 -19493 16289 -18661
rect 16351 -19493 16385 -18661
rect 16447 -19493 16481 -18661
rect 16543 -19493 16577 -18661
rect 16639 -19493 16673 -18661
rect 16735 -19493 16769 -18661
rect 16831 -19493 16865 -18661
rect 16927 -19493 16961 -18661
rect -24414 -20153 -24224 -20119
rect -21606 -20196 -21572 -20006
rect -21510 -20196 -21476 -20002
rect -21414 -20196 -21380 -20006
rect -21318 -20196 -21284 -20002
rect -16015 -20067 -15981 -19877
rect -15919 -20067 -15885 -19873
rect -15823 -20067 -15789 -19877
rect -15727 -20067 -15693 -19873
rect -12302 -19912 -11776 -19878
rect -17665 -20145 -17433 -20111
rect -24414 -20249 -24224 -20215
rect -17665 -20241 -17433 -20207
rect -17665 -20337 -17433 -20303
rect -17665 -20433 -17433 -20399
rect -21606 -20656 -21572 -20466
rect -21510 -20656 -21476 -20462
rect -21414 -20656 -21380 -20466
rect -21318 -20656 -21284 -20462
rect -17665 -20529 -17433 -20495
rect -17665 -20625 -17433 -20591
rect -24383 -20873 -24193 -20839
rect -24383 -20969 -24193 -20935
rect -24383 -21065 -24193 -21031
rect -24383 -21161 -24193 -21127
rect -24383 -21257 -24193 -21223
rect -21620 -21116 -21586 -20926
rect -21524 -21116 -21490 -20922
rect -21428 -21116 -21394 -20926
rect -21332 -21116 -21298 -20922
rect -17665 -20721 -17433 -20687
rect -16015 -20527 -15981 -20337
rect -15919 -20527 -15885 -20333
rect -15823 -20527 -15789 -20337
rect -15727 -20527 -15693 -20333
rect -17665 -20817 -17433 -20783
rect -17665 -20913 -17433 -20879
rect -17665 -21009 -17433 -20975
rect -16029 -20987 -15995 -20797
rect -15933 -20987 -15899 -20793
rect -15837 -20987 -15803 -20797
rect -15741 -20987 -15707 -20793
rect -17665 -21105 -17433 -21071
rect -12302 -20000 -11776 -19966
rect -12302 -20096 -11776 -20062
rect -12302 -20192 -11776 -20158
rect -12302 -20288 -11776 -20254
rect -12302 -20384 -11776 -20350
rect -12302 -20480 -11776 -20446
rect -12302 -20576 -11776 -20542
rect -12302 -20672 -11776 -20638
rect -12302 -20768 -11776 -20734
rect -12302 -20864 -11776 -20830
rect -12302 -20960 -11776 -20926
rect -12302 -21056 -11776 -21022
rect -12302 -21152 -11776 -21118
rect -4816 -20138 -4782 -19948
rect -4720 -20142 -4686 -19948
rect -4624 -20138 -4590 -19948
rect -4528 -20142 -4494 -19948
rect -2100 -20132 -2066 -19942
rect -2004 -20132 -1970 -19938
rect -1908 -20132 -1874 -19942
rect -1812 -20132 -1778 -19938
rect -4816 -20578 -4782 -20388
rect -4720 -20582 -4686 -20388
rect -4624 -20578 -4590 -20388
rect -4528 -20582 -4494 -20388
rect -2100 -20572 -2066 -20382
rect -2004 -20572 -1970 -20378
rect -1908 -20572 -1874 -20382
rect -1812 -20572 -1778 -20378
rect -4816 -20957 -4782 -20767
rect -4720 -20961 -4686 -20767
rect -4624 -20957 -4590 -20767
rect -4528 -20961 -4494 -20767
rect 11785 -20875 11819 -20643
rect 11881 -20875 11915 -20643
rect 11977 -20875 12011 -20643
rect 12073 -20875 12107 -20643
rect 12169 -20875 12203 -20643
rect 12265 -20875 12299 -20643
rect 12361 -20875 12395 -20643
rect 12457 -20875 12491 -20643
rect 12553 -20875 12587 -20643
rect 12649 -20875 12683 -20643
rect 12745 -20875 12779 -20643
rect -24383 -21353 -24193 -21319
rect -12302 -21240 -11776 -21206
rect -24383 -21449 -24193 -21415
rect -21618 -21596 -21584 -21406
rect -21522 -21596 -21488 -21402
rect -21426 -21596 -21392 -21406
rect -21330 -21596 -21296 -21402
rect -16027 -21467 -15993 -21277
rect -15931 -21467 -15897 -21273
rect -15835 -21467 -15801 -21277
rect -15739 -21467 -15705 -21273
rect -17665 -21545 -17433 -21511
rect -17665 -21641 -17433 -21607
rect -17665 -21737 -17433 -21703
rect -17665 -21833 -17433 -21799
rect -17665 -21929 -17433 -21895
rect -17665 -22025 -17433 -21991
rect -24384 -22176 -24194 -22142
rect -24384 -22272 -24194 -22238
rect -24384 -22368 -24194 -22334
rect -24384 -22464 -24194 -22430
rect -24384 -22560 -24194 -22526
rect -17665 -22121 -17433 -22087
rect -17665 -22217 -17433 -22183
rect 12935 -20781 13125 -20747
rect 12935 -20877 13129 -20843
rect 12935 -20973 13125 -20939
rect 12935 -21069 13129 -21035
rect -17665 -22313 -17433 -22279
rect -17665 -22409 -17433 -22375
rect -17665 -22505 -17433 -22471
rect -12302 -22491 -11776 -22457
rect -24384 -22656 -24194 -22622
rect -24384 -22752 -24194 -22718
rect -17665 -22945 -17433 -22911
rect -17665 -23041 -17433 -23007
rect -17665 -23137 -17433 -23103
rect -17665 -23233 -17433 -23199
rect -17665 -23329 -17433 -23295
rect -17665 -23425 -17433 -23391
rect -24384 -23485 -24194 -23451
rect -24384 -23581 -24194 -23547
rect -24384 -23677 -24194 -23643
rect -24384 -23773 -24194 -23739
rect -24384 -23869 -24194 -23835
rect -24384 -23965 -24194 -23931
rect -17665 -23521 -17433 -23487
rect -17665 -23617 -17433 -23583
rect -17665 -23713 -17433 -23679
rect -12302 -22579 -11776 -22545
rect -12302 -22675 -11776 -22641
rect -12302 -22771 -11776 -22737
rect -12302 -22867 -11776 -22833
rect -12302 -22963 -11776 -22929
rect -12302 -23059 -11776 -23025
rect -12302 -23155 -11776 -23121
rect -12302 -23251 -11776 -23217
rect -12302 -23347 -11776 -23313
rect -12302 -23443 -11776 -23409
rect -12302 -23539 -11776 -23505
rect -12302 -23635 -11776 -23601
rect -12302 -23731 -11776 -23697
rect 7150 -22595 7184 -22297
rect 7246 -22595 7280 -22297
rect 7342 -22595 7376 -22297
rect 7438 -22595 7472 -22297
rect 7534 -22595 7568 -22297
rect 7630 -22595 7664 -22297
rect 7726 -22595 7760 -22297
rect 7822 -22595 7856 -22297
rect 7918 -22595 7952 -22297
rect 8098 -22595 8132 -22297
rect 8194 -22595 8228 -22297
rect 8290 -22595 8324 -22297
rect 8386 -22595 8420 -22297
rect 8482 -22595 8516 -22297
rect 8578 -22595 8612 -22297
rect 8674 -22595 8708 -22297
rect 8770 -22595 8804 -22297
rect 8866 -22595 8900 -22297
rect 9034 -22595 9068 -22297
rect 9130 -22595 9164 -22297
rect 9226 -22595 9260 -22297
rect 9322 -22595 9356 -22297
rect 9418 -22595 9452 -22297
rect 9514 -22595 9548 -22297
rect 9610 -22595 9644 -22297
rect 9706 -22595 9740 -22297
rect 9802 -22595 9836 -22297
rect 9965 -22594 9999 -22296
rect 10061 -22594 10095 -22296
rect 10157 -22594 10191 -22296
rect 10253 -22594 10287 -22296
rect 10349 -22594 10383 -22296
rect 10445 -22594 10479 -22296
rect 10541 -22594 10575 -22296
rect 10637 -22594 10671 -22296
rect 10733 -22594 10767 -22296
rect 10892 -22595 10926 -22297
rect 10988 -22595 11022 -22297
rect 11084 -22595 11118 -22297
rect 11180 -22595 11214 -22297
rect 11276 -22595 11310 -22297
rect 11372 -22595 11406 -22297
rect 11468 -22595 11502 -22297
rect 11564 -22595 11598 -22297
rect 11660 -22595 11694 -22297
rect 5670 -23291 5860 -23257
rect 5670 -23387 5864 -23353
rect 5670 -23483 5860 -23449
rect 5670 -23579 5864 -23545
rect 6110 -23291 6300 -23257
rect 6110 -23387 6304 -23353
rect 6110 -23483 6300 -23449
rect 6110 -23579 6304 -23545
rect 6550 -23291 6740 -23257
rect 6550 -23387 6744 -23353
rect 6550 -23483 6740 -23449
rect 6550 -23579 6744 -23545
rect -17665 -23809 -17433 -23775
rect -12302 -23819 -11776 -23785
rect -17665 -23905 -17433 -23871
rect -24384 -24061 -24194 -24027
rect 7150 -24259 7184 -23961
rect 7246 -24259 7280 -23961
rect 7342 -24259 7376 -23961
rect 7438 -24259 7472 -23961
rect 7534 -24259 7568 -23961
rect 7630 -24259 7664 -23961
rect 7726 -24259 7760 -23961
rect 7822 -24259 7856 -23961
rect 7918 -24259 7952 -23961
rect 8098 -24259 8132 -23961
rect 8194 -24259 8228 -23961
rect 8290 -24259 8324 -23961
rect 8386 -24259 8420 -23961
rect 8482 -24259 8516 -23961
rect 8578 -24259 8612 -23961
rect 8674 -24259 8708 -23961
rect 8770 -24259 8804 -23961
rect 8866 -24259 8900 -23961
rect 9034 -24259 9068 -23961
rect 9130 -24259 9164 -23961
rect 9226 -24259 9260 -23961
rect 9322 -24259 9356 -23961
rect 9418 -24259 9452 -23961
rect 9514 -24259 9548 -23961
rect 9610 -24259 9644 -23961
rect 9706 -24259 9740 -23961
rect 9802 -24259 9836 -23961
rect 9965 -24259 9999 -23961
rect 10061 -24259 10095 -23961
rect 10157 -24259 10191 -23961
rect 10253 -24259 10287 -23961
rect 10349 -24259 10383 -23961
rect 10445 -24259 10479 -23961
rect 10541 -24259 10575 -23961
rect 10637 -24259 10671 -23961
rect 10733 -24259 10767 -23961
rect 10892 -24259 10926 -23961
rect 10988 -24259 11022 -23961
rect 11084 -24259 11118 -23961
rect 11180 -24259 11214 -23961
rect 11276 -24259 11310 -23961
rect 11372 -24259 11406 -23961
rect 11468 -24259 11502 -23961
rect 11564 -24259 11598 -23961
rect 11660 -24259 11694 -23961
rect -17665 -24345 -17433 -24311
rect -17665 -24441 -17433 -24407
rect -17665 -24537 -17433 -24503
rect -17665 -24633 -17433 -24599
rect -17665 -24729 -17433 -24695
rect -17665 -24825 -17433 -24791
rect -17665 -24921 -17433 -24887
rect -17665 -25017 -17433 -24983
rect -17665 -25113 -17433 -25079
rect -17665 -25209 -17433 -25175
rect -12302 -25259 -11776 -25225
rect -17665 -25305 -17433 -25271
rect -12302 -25347 -11776 -25313
rect -12302 -25443 -11776 -25409
rect -12302 -25539 -11776 -25505
rect -12302 -25635 -11776 -25601
rect -12302 -25731 -11776 -25697
rect -12302 -25827 -11776 -25793
rect -12302 -25923 -11776 -25889
rect -12302 -26019 -11776 -25985
rect -12302 -26115 -11776 -26081
rect -12302 -26211 -11776 -26177
rect -12302 -26307 -11776 -26273
rect -12302 -26403 -11776 -26369
rect -12302 -26499 -11776 -26465
rect 11785 -25403 11819 -25171
rect 11881 -25403 11915 -25171
rect 11977 -25403 12011 -25171
rect 12073 -25403 12107 -25171
rect 12169 -25403 12203 -25171
rect 12265 -25403 12299 -25171
rect 12361 -25403 12395 -25171
rect 12457 -25403 12491 -25171
rect 12553 -25403 12587 -25171
rect 12649 -25403 12683 -25171
rect 12745 -25403 12779 -25171
rect -12302 -26587 -11776 -26553
rect 12935 -25309 13125 -25275
rect 12935 -25405 13129 -25371
rect 12935 -25501 13125 -25467
rect 12935 -25597 13129 -25563
rect 7150 -27123 7184 -26825
rect 7246 -27123 7280 -26825
rect 7342 -27123 7376 -26825
rect 7438 -27123 7472 -26825
rect 7534 -27123 7568 -26825
rect 7630 -27123 7664 -26825
rect 7726 -27123 7760 -26825
rect 7822 -27123 7856 -26825
rect 7918 -27123 7952 -26825
rect 8098 -27123 8132 -26825
rect 8194 -27123 8228 -26825
rect 8290 -27123 8324 -26825
rect 8386 -27123 8420 -26825
rect 8482 -27123 8516 -26825
rect 8578 -27123 8612 -26825
rect 8674 -27123 8708 -26825
rect 8770 -27123 8804 -26825
rect 8866 -27123 8900 -26825
rect 9034 -27123 9068 -26825
rect 9130 -27123 9164 -26825
rect 9226 -27123 9260 -26825
rect 9322 -27123 9356 -26825
rect 9418 -27123 9452 -26825
rect 9514 -27123 9548 -26825
rect 9610 -27123 9644 -26825
rect 9706 -27123 9740 -26825
rect 9802 -27123 9836 -26825
rect 9965 -27122 9999 -26824
rect 10061 -27122 10095 -26824
rect 10157 -27122 10191 -26824
rect 10253 -27122 10287 -26824
rect 10349 -27122 10383 -26824
rect 10445 -27122 10479 -26824
rect 10541 -27122 10575 -26824
rect 10637 -27122 10671 -26824
rect 10733 -27122 10767 -26824
rect 10892 -27123 10926 -26825
rect 10988 -27123 11022 -26825
rect 11084 -27123 11118 -26825
rect 11180 -27123 11214 -26825
rect 11276 -27123 11310 -26825
rect 11372 -27123 11406 -26825
rect 11468 -27123 11502 -26825
rect 11564 -27123 11598 -26825
rect 11660 -27123 11694 -26825
rect -12302 -27892 -11776 -27858
rect -12302 -27980 -11776 -27946
rect -12302 -28076 -11776 -28042
rect -12302 -28172 -11776 -28138
rect -12302 -28268 -11776 -28234
rect -12302 -28364 -11776 -28330
rect -12302 -28460 -11776 -28426
rect -12302 -28556 -11776 -28522
rect -12302 -28652 -11776 -28618
rect -12302 -28748 -11776 -28714
rect -12302 -28844 -11776 -28810
rect -12302 -28940 -11776 -28906
rect -12302 -29036 -11776 -29002
rect -12302 -29132 -11776 -29098
rect 5670 -27819 5860 -27785
rect 5670 -27915 5864 -27881
rect 5670 -28011 5860 -27977
rect 5670 -28107 5864 -28073
rect 6110 -27819 6300 -27785
rect 6110 -27915 6304 -27881
rect 6110 -28011 6300 -27977
rect 6110 -28107 6304 -28073
rect 6550 -27819 6740 -27785
rect 6550 -27915 6744 -27881
rect 6550 -28011 6740 -27977
rect 6550 -28107 6744 -28073
rect 7150 -28787 7184 -28489
rect 7246 -28787 7280 -28489
rect 7342 -28787 7376 -28489
rect 7438 -28787 7472 -28489
rect 7534 -28787 7568 -28489
rect 7630 -28787 7664 -28489
rect 7726 -28787 7760 -28489
rect 7822 -28787 7856 -28489
rect 7918 -28787 7952 -28489
rect 8098 -28787 8132 -28489
rect 8194 -28787 8228 -28489
rect 8290 -28787 8324 -28489
rect 8386 -28787 8420 -28489
rect 8482 -28787 8516 -28489
rect 8578 -28787 8612 -28489
rect 8674 -28787 8708 -28489
rect 8770 -28787 8804 -28489
rect 8866 -28787 8900 -28489
rect 9034 -28787 9068 -28489
rect 9130 -28787 9164 -28489
rect 9226 -28787 9260 -28489
rect 9322 -28787 9356 -28489
rect 9418 -28787 9452 -28489
rect 9514 -28787 9548 -28489
rect 9610 -28787 9644 -28489
rect 9706 -28787 9740 -28489
rect 9802 -28787 9836 -28489
rect 9965 -28787 9999 -28489
rect 10061 -28787 10095 -28489
rect 10157 -28787 10191 -28489
rect 10253 -28787 10287 -28489
rect 10349 -28787 10383 -28489
rect 10445 -28787 10479 -28489
rect 10541 -28787 10575 -28489
rect 10637 -28787 10671 -28489
rect 10733 -28787 10767 -28489
rect 10892 -28787 10926 -28489
rect 10988 -28787 11022 -28489
rect 11084 -28787 11118 -28489
rect 11180 -28787 11214 -28489
rect 11276 -28787 11310 -28489
rect 11372 -28787 11406 -28489
rect 11468 -28787 11502 -28489
rect 11564 -28787 11598 -28489
rect 11660 -28787 11694 -28489
rect -12302 -29220 -11776 -29186
rect 11785 -29931 11819 -29699
rect 11881 -29931 11915 -29699
rect 11977 -29931 12011 -29699
rect 12073 -29931 12107 -29699
rect 12169 -29931 12203 -29699
rect 12265 -29931 12299 -29699
rect 12361 -29931 12395 -29699
rect 12457 -29931 12491 -29699
rect 12553 -29931 12587 -29699
rect 12649 -29931 12683 -29699
rect 12745 -29931 12779 -29699
rect -12302 -30501 -11776 -30467
rect -12302 -30589 -11776 -30555
rect -12302 -30685 -11776 -30651
rect -12302 -30781 -11776 -30747
rect -12302 -30877 -11776 -30843
rect -12302 -30973 -11776 -30939
rect -12302 -31069 -11776 -31035
rect -12302 -31165 -11776 -31131
rect -12302 -31261 -11776 -31227
rect -12302 -31357 -11776 -31323
rect -12302 -31453 -11776 -31419
rect -12302 -31549 -11776 -31515
rect -12302 -31645 -11776 -31611
rect -12302 -31741 -11776 -31707
rect 12935 -29837 13125 -29803
rect 12935 -29933 13129 -29899
rect 12935 -30029 13125 -29995
rect 12935 -30125 13129 -30091
rect 7150 -31651 7184 -31353
rect 7246 -31651 7280 -31353
rect 7342 -31651 7376 -31353
rect 7438 -31651 7472 -31353
rect 7534 -31651 7568 -31353
rect 7630 -31651 7664 -31353
rect 7726 -31651 7760 -31353
rect 7822 -31651 7856 -31353
rect 7918 -31651 7952 -31353
rect 8098 -31651 8132 -31353
rect 8194 -31651 8228 -31353
rect 8290 -31651 8324 -31353
rect 8386 -31651 8420 -31353
rect 8482 -31651 8516 -31353
rect 8578 -31651 8612 -31353
rect 8674 -31651 8708 -31353
rect 8770 -31651 8804 -31353
rect 8866 -31651 8900 -31353
rect 9034 -31651 9068 -31353
rect 9130 -31651 9164 -31353
rect 9226 -31651 9260 -31353
rect 9322 -31651 9356 -31353
rect 9418 -31651 9452 -31353
rect 9514 -31651 9548 -31353
rect 9610 -31651 9644 -31353
rect 9706 -31651 9740 -31353
rect 9802 -31651 9836 -31353
rect 9965 -31650 9999 -31352
rect 10061 -31650 10095 -31352
rect 10157 -31650 10191 -31352
rect 10253 -31650 10287 -31352
rect 10349 -31650 10383 -31352
rect 10445 -31650 10479 -31352
rect 10541 -31650 10575 -31352
rect 10637 -31650 10671 -31352
rect 10733 -31650 10767 -31352
rect 10892 -31651 10926 -31353
rect 10988 -31651 11022 -31353
rect 11084 -31651 11118 -31353
rect 11180 -31651 11214 -31353
rect 11276 -31651 11310 -31353
rect 11372 -31651 11406 -31353
rect 11468 -31651 11502 -31353
rect 11564 -31651 11598 -31353
rect 11660 -31651 11694 -31353
rect -12302 -31829 -11776 -31795
rect 5670 -32347 5860 -32313
rect 5670 -32443 5864 -32409
rect 5670 -32539 5860 -32505
rect 5670 -32635 5864 -32601
rect 6110 -32347 6300 -32313
rect 6110 -32443 6304 -32409
rect 6110 -32539 6300 -32505
rect 6110 -32635 6304 -32601
rect 6550 -32347 6740 -32313
rect 6550 -32443 6744 -32409
rect 6550 -32539 6740 -32505
rect 6550 -32635 6744 -32601
rect -12304 -33121 -11778 -33087
rect -12304 -33209 -11778 -33175
rect -12304 -33305 -11778 -33271
rect -12304 -33401 -11778 -33367
rect -12304 -33497 -11778 -33463
rect -12304 -33593 -11778 -33559
rect -12304 -33689 -11778 -33655
rect -12304 -33785 -11778 -33751
rect -12304 -33881 -11778 -33847
rect -12304 -33977 -11778 -33943
rect -12304 -34073 -11778 -34039
rect -12304 -34169 -11778 -34135
rect -12304 -34265 -11778 -34231
rect -12304 -34361 -11778 -34327
rect 7150 -33315 7184 -33017
rect 7246 -33315 7280 -33017
rect 7342 -33315 7376 -33017
rect 7438 -33315 7472 -33017
rect 7534 -33315 7568 -33017
rect 7630 -33315 7664 -33017
rect 7726 -33315 7760 -33017
rect 7822 -33315 7856 -33017
rect 7918 -33315 7952 -33017
rect 8098 -33315 8132 -33017
rect 8194 -33315 8228 -33017
rect 8290 -33315 8324 -33017
rect 8386 -33315 8420 -33017
rect 8482 -33315 8516 -33017
rect 8578 -33315 8612 -33017
rect 8674 -33315 8708 -33017
rect 8770 -33315 8804 -33017
rect 8866 -33315 8900 -33017
rect 9034 -33315 9068 -33017
rect 9130 -33315 9164 -33017
rect 9226 -33315 9260 -33017
rect 9322 -33315 9356 -33017
rect 9418 -33315 9452 -33017
rect 9514 -33315 9548 -33017
rect 9610 -33315 9644 -33017
rect 9706 -33315 9740 -33017
rect 9802 -33315 9836 -33017
rect 9965 -33315 9999 -33017
rect 10061 -33315 10095 -33017
rect 10157 -33315 10191 -33017
rect 10253 -33315 10287 -33017
rect 10349 -33315 10383 -33017
rect 10445 -33315 10479 -33017
rect 10541 -33315 10575 -33017
rect 10637 -33315 10671 -33017
rect 10733 -33315 10767 -33017
rect 10892 -33315 10926 -33017
rect 10988 -33315 11022 -33017
rect 11084 -33315 11118 -33017
rect 11180 -33315 11214 -33017
rect 11276 -33315 11310 -33017
rect 11372 -33315 11406 -33017
rect 11468 -33315 11502 -33017
rect 11564 -33315 11598 -33017
rect 11660 -33315 11694 -33017
rect -12304 -34449 -11778 -34415
rect 11785 -34459 11819 -34227
rect 11881 -34459 11915 -34227
rect 11977 -34459 12011 -34227
rect 12073 -34459 12107 -34227
rect 12169 -34459 12203 -34227
rect 12265 -34459 12299 -34227
rect 12361 -34459 12395 -34227
rect 12457 -34459 12491 -34227
rect 12553 -34459 12587 -34227
rect 12649 -34459 12683 -34227
rect 12745 -34459 12779 -34227
rect 12935 -34365 13125 -34331
rect 12935 -34461 13129 -34427
rect 12935 -34557 13125 -34523
rect 12935 -34653 13129 -34619
rect 7150 -36179 7184 -35881
rect 7246 -36179 7280 -35881
rect 7342 -36179 7376 -35881
rect 7438 -36179 7472 -35881
rect 7534 -36179 7568 -35881
rect 7630 -36179 7664 -35881
rect 7726 -36179 7760 -35881
rect 7822 -36179 7856 -35881
rect 7918 -36179 7952 -35881
rect 8098 -36179 8132 -35881
rect 8194 -36179 8228 -35881
rect 8290 -36179 8324 -35881
rect 8386 -36179 8420 -35881
rect 8482 -36179 8516 -35881
rect 8578 -36179 8612 -35881
rect 8674 -36179 8708 -35881
rect 8770 -36179 8804 -35881
rect 8866 -36179 8900 -35881
rect 9034 -36179 9068 -35881
rect 9130 -36179 9164 -35881
rect 9226 -36179 9260 -35881
rect 9322 -36179 9356 -35881
rect 9418 -36179 9452 -35881
rect 9514 -36179 9548 -35881
rect 9610 -36179 9644 -35881
rect 9706 -36179 9740 -35881
rect 9802 -36179 9836 -35881
rect 9965 -36178 9999 -35880
rect 10061 -36178 10095 -35880
rect 10157 -36178 10191 -35880
rect 10253 -36178 10287 -35880
rect 10349 -36178 10383 -35880
rect 10445 -36178 10479 -35880
rect 10541 -36178 10575 -35880
rect 10637 -36178 10671 -35880
rect 10733 -36178 10767 -35880
rect 10892 -36179 10926 -35881
rect 10988 -36179 11022 -35881
rect 11084 -36179 11118 -35881
rect 11180 -36179 11214 -35881
rect 11276 -36179 11310 -35881
rect 11372 -36179 11406 -35881
rect 11468 -36179 11502 -35881
rect 11564 -36179 11598 -35881
rect 11660 -36179 11694 -35881
rect 13136 -35921 13170 -35727
rect 13232 -35917 13266 -35727
rect 13328 -35921 13362 -35727
rect 13424 -35917 13458 -35727
rect 13136 -36300 13170 -36106
rect 13232 -36296 13266 -36106
rect 13328 -36300 13362 -36106
rect 13424 -36296 13458 -36106
<< psubdiff >>
rect 1800 4838 3002 4860
rect 1800 4792 1841 4838
rect 2964 4792 3002 4838
rect 1800 4769 3002 4792
rect 3406 4838 4608 4860
rect 3406 4792 3447 4838
rect 4570 4792 4608 4838
rect 3406 4769 4608 4792
rect 5110 4836 6312 4858
rect 5110 4790 5151 4836
rect 6274 4790 6312 4836
rect 5110 4767 6312 4790
rect 7173 4821 7573 4847
rect 7173 4787 7200 4821
rect 7535 4787 7573 4821
rect 7173 4776 7573 4787
rect 7809 4819 8009 4821
rect 7809 4785 7840 4819
rect 7972 4785 8009 4819
rect 7809 4778 8009 4785
rect 5658 3271 5858 3273
rect 5658 3237 5689 3271
rect 5821 3237 5858 3271
rect 5658 3230 5858 3237
rect 6098 3271 6298 3273
rect 6098 3237 6129 3271
rect 6261 3237 6298 3271
rect 6098 3230 6298 3237
rect 6538 3271 6738 3273
rect 6538 3237 6569 3271
rect 6701 3237 6738 3271
rect 6538 3230 6738 3237
rect -24039 3114 -22837 3136
rect -24039 3068 -24001 3114
rect -22878 3068 -22837 3114
rect -24039 3045 -22837 3068
rect -20748 3114 -19546 3136
rect -20748 3068 -20710 3114
rect -19587 3068 -19546 3114
rect -20748 3045 -19546 3068
rect -17457 3114 -16255 3136
rect -17457 3068 -17419 3114
rect -16296 3068 -16255 3114
rect -17457 3045 -16255 3068
rect -14166 3114 -12964 3136
rect -14166 3068 -14128 3114
rect -13005 3068 -12964 3114
rect -14166 3045 -12964 3068
rect -10875 3114 -9673 3136
rect -10875 3068 -10837 3114
rect -9714 3068 -9673 3114
rect -10875 3045 -9673 3068
rect -7585 3114 -6383 3136
rect -7585 3068 -7547 3114
rect -6424 3068 -6383 3114
rect -7585 3045 -6383 3068
rect -4294 3114 -3092 3136
rect -4294 3068 -4256 3114
rect -3133 3068 -3092 3114
rect -4294 3045 -3092 3068
rect -1003 3114 199 3136
rect -1003 3068 -965 3114
rect 158 3068 199 3114
rect -1003 3045 199 3068
rect 7298 2466 7360 2490
rect 7332 2118 7360 2466
rect 7298 2066 7360 2118
rect 7332 1715 7360 2066
rect 7298 1690 7360 1715
rect 8246 2466 8308 2490
rect 8280 2118 8308 2466
rect 8246 2066 8308 2118
rect 8280 1715 8308 2066
rect 8246 1690 8308 1715
rect 9182 2466 9244 2490
rect 9216 2118 9244 2466
rect 9182 2066 9244 2118
rect 9216 1715 9244 2066
rect 9182 1690 9244 1715
rect 10113 2466 10175 2490
rect 10147 2118 10175 2466
rect 10113 2066 10175 2118
rect 10147 1715 10175 2066
rect 10113 1690 10175 1715
rect 11040 2466 11102 2490
rect 11074 2118 11102 2466
rect 11040 2066 11102 2118
rect 11074 1715 11102 2066
rect 11040 1690 11102 1715
rect 7298 1537 7360 1562
rect -24711 1330 -23509 1352
rect -24711 1284 -24670 1330
rect -23547 1284 -23509 1330
rect -24711 1261 -23509 1284
rect -23152 1330 -21950 1352
rect -23152 1284 -23111 1330
rect -21988 1284 -21950 1330
rect -23152 1261 -21950 1284
rect -21420 1330 -20218 1352
rect -21420 1284 -21379 1330
rect -20256 1284 -20218 1330
rect -21420 1261 -20218 1284
rect -19861 1330 -18659 1352
rect -19861 1284 -19820 1330
rect -18697 1284 -18659 1330
rect -19861 1261 -18659 1284
rect -18129 1330 -16927 1352
rect -18129 1284 -18088 1330
rect -16965 1284 -16927 1330
rect -18129 1261 -16927 1284
rect -16570 1330 -15368 1352
rect -16570 1284 -16529 1330
rect -15406 1284 -15368 1330
rect -16570 1261 -15368 1284
rect -14838 1330 -13636 1352
rect -14838 1284 -14797 1330
rect -13674 1284 -13636 1330
rect -14838 1261 -13636 1284
rect -13279 1330 -12077 1352
rect -13279 1284 -13238 1330
rect -12115 1284 -12077 1330
rect -13279 1261 -12077 1284
rect -11547 1330 -10345 1352
rect -11547 1284 -11506 1330
rect -10383 1284 -10345 1330
rect -11547 1261 -10345 1284
rect -9988 1330 -8786 1352
rect -9988 1284 -9947 1330
rect -8824 1284 -8786 1330
rect -9988 1261 -8786 1284
rect -8257 1330 -7055 1352
rect -8257 1284 -8216 1330
rect -7093 1284 -7055 1330
rect -8257 1261 -7055 1284
rect -6698 1330 -5496 1352
rect -6698 1284 -6657 1330
rect -5534 1284 -5496 1330
rect -6698 1261 -5496 1284
rect -4966 1330 -3764 1352
rect -4966 1284 -4925 1330
rect -3802 1284 -3764 1330
rect -4966 1261 -3764 1284
rect -3407 1330 -2205 1352
rect -3407 1284 -3366 1330
rect -2243 1284 -2205 1330
rect -3407 1261 -2205 1284
rect -1675 1330 -473 1352
rect -1675 1284 -1634 1330
rect -511 1284 -473 1330
rect -1675 1261 -473 1284
rect -116 1330 1086 1352
rect -116 1284 -75 1330
rect 1048 1284 1086 1330
rect -116 1261 1086 1284
rect 7332 1186 7360 1537
rect 7298 1134 7360 1186
rect 7332 786 7360 1134
rect 7298 762 7360 786
rect 8246 1537 8308 1562
rect 8280 1186 8308 1537
rect 8246 1134 8308 1186
rect 8280 786 8308 1134
rect 8246 762 8308 786
rect 9182 1537 9244 1562
rect 9216 1186 9244 1537
rect 9182 1134 9244 1186
rect 9216 786 9244 1134
rect 9182 762 9244 786
rect 10113 1538 10175 1563
rect 10147 1187 10175 1538
rect 10113 1135 10175 1187
rect 10147 787 10175 1135
rect 10113 763 10175 787
rect 11040 1537 11102 1562
rect 11074 1186 11102 1537
rect 11040 1134 11102 1186
rect 11074 786 11102 1134
rect 11040 762 11102 786
rect 12157 1249 12407 1266
rect 12157 1188 12183 1249
rect 12382 1188 12407 1249
rect 12923 1253 13123 1255
rect 12923 1219 12954 1253
rect 13086 1219 13123 1253
rect 12923 1212 13123 1219
rect 12157 1170 12407 1188
rect -24363 255 -23963 281
rect -24363 221 -24336 255
rect -24001 221 -23963 255
rect -24363 210 -23963 221
rect -23254 255 -22854 281
rect -23254 221 -23227 255
rect -22892 221 -22854 255
rect -23254 210 -22854 221
rect -22372 255 -21972 281
rect -22372 221 -22345 255
rect -22010 221 -21972 255
rect -22372 210 -21972 221
rect -21072 255 -20672 281
rect -21072 221 -21045 255
rect -20710 221 -20672 255
rect -21072 210 -20672 221
rect -19963 255 -19563 281
rect -19963 221 -19936 255
rect -19601 221 -19563 255
rect -19963 210 -19563 221
rect -19081 255 -18681 281
rect -19081 221 -19054 255
rect -18719 221 -18681 255
rect -19081 210 -18681 221
rect -17781 255 -17381 281
rect -17781 221 -17754 255
rect -17419 221 -17381 255
rect -17781 210 -17381 221
rect -16672 255 -16272 281
rect -16672 221 -16645 255
rect -16310 221 -16272 255
rect -16672 210 -16272 221
rect -15790 255 -15390 281
rect -15790 221 -15763 255
rect -15428 221 -15390 255
rect -15790 210 -15390 221
rect -14490 255 -14090 281
rect -14490 221 -14463 255
rect -14128 221 -14090 255
rect -14490 210 -14090 221
rect -13381 255 -12981 281
rect -13381 221 -13354 255
rect -13019 221 -12981 255
rect -13381 210 -12981 221
rect -12499 255 -12099 281
rect -12499 221 -12472 255
rect -12137 221 -12099 255
rect -12499 210 -12099 221
rect -11199 255 -10799 281
rect -11199 221 -11172 255
rect -10837 221 -10799 255
rect -11199 210 -10799 221
rect -10090 255 -9690 281
rect -10090 221 -10063 255
rect -9728 221 -9690 255
rect -10090 210 -9690 221
rect -9208 255 -8808 281
rect -9208 221 -9181 255
rect -8846 221 -8808 255
rect -9208 210 -8808 221
rect -7909 255 -7509 281
rect -7909 221 -7882 255
rect -7547 221 -7509 255
rect -7909 210 -7509 221
rect -6800 255 -6400 281
rect -6800 221 -6773 255
rect -6438 221 -6400 255
rect -6800 210 -6400 221
rect -5918 255 -5518 281
rect -5918 221 -5891 255
rect -5556 221 -5518 255
rect -5918 210 -5518 221
rect -4618 255 -4218 281
rect -4618 221 -4591 255
rect -4256 221 -4218 255
rect -4618 210 -4218 221
rect -3509 255 -3109 281
rect -3509 221 -3482 255
rect -3147 221 -3109 255
rect -3509 210 -3109 221
rect -2627 255 -2227 281
rect -2627 221 -2600 255
rect -2265 221 -2227 255
rect -2627 210 -2227 221
rect -1327 255 -927 281
rect -1327 221 -1300 255
rect -965 221 -927 255
rect -1327 210 -927 221
rect -218 255 182 281
rect -218 221 -191 255
rect 144 221 182 255
rect -218 210 182 221
rect 664 255 1064 281
rect 664 221 691 255
rect 1026 221 1064 255
rect 664 210 1064 221
rect 5658 -1257 5858 -1255
rect 5658 -1291 5689 -1257
rect 5821 -1291 5858 -1257
rect 5658 -1298 5858 -1291
rect 6098 -1257 6298 -1255
rect 6098 -1291 6129 -1257
rect 6261 -1291 6298 -1257
rect 6098 -1298 6298 -1291
rect 6538 -1257 6738 -1255
rect 6538 -1291 6569 -1257
rect 6701 -1291 6738 -1257
rect 6538 -1298 6738 -1291
rect 7298 -2062 7360 -2038
rect 7332 -2410 7360 -2062
rect 7298 -2462 7360 -2410
rect 7332 -2813 7360 -2462
rect 7298 -2838 7360 -2813
rect 8246 -2062 8308 -2038
rect 8280 -2410 8308 -2062
rect 8246 -2462 8308 -2410
rect 8280 -2813 8308 -2462
rect 8246 -2838 8308 -2813
rect 9182 -2062 9244 -2038
rect 9216 -2410 9244 -2062
rect 9182 -2462 9244 -2410
rect 9216 -2813 9244 -2462
rect 9182 -2838 9244 -2813
rect 10113 -2062 10175 -2038
rect 10147 -2410 10175 -2062
rect 10113 -2462 10175 -2410
rect 10147 -2813 10175 -2462
rect 10113 -2838 10175 -2813
rect 11040 -2062 11102 -2038
rect 11074 -2410 11102 -2062
rect 11040 -2462 11102 -2410
rect 11074 -2813 11102 -2462
rect 11040 -2838 11102 -2813
rect -23628 -2959 -23428 -2957
rect -23628 -2993 -23597 -2959
rect -23465 -2993 -23428 -2959
rect -23628 -3000 -23428 -2993
rect -24213 -3033 -23813 -3007
rect -24213 -3067 -24186 -3033
rect -23851 -3067 -23813 -3033
rect -24213 -3078 -23813 -3067
rect -21608 -2959 -21408 -2957
rect -21608 -2993 -21577 -2959
rect -21445 -2993 -21408 -2959
rect -21608 -3000 -21408 -2993
rect -22176 -3033 -21776 -3007
rect -22176 -3067 -22149 -3033
rect -21814 -3067 -21776 -3033
rect -22176 -3078 -21776 -3067
rect -19867 -2959 -19667 -2957
rect -19867 -2993 -19836 -2959
rect -19704 -2993 -19667 -2959
rect -19867 -3000 -19667 -2993
rect -20446 -3033 -20046 -3007
rect -20446 -3067 -20419 -3033
rect -20084 -3067 -20046 -3033
rect -20446 -3078 -20046 -3067
rect -18088 -2959 -17888 -2957
rect -18088 -2993 -18057 -2959
rect -17925 -2993 -17888 -2959
rect -18088 -3000 -17888 -2993
rect 7298 -2991 7360 -2966
rect -18686 -3033 -18286 -3007
rect -18686 -3067 -18659 -3033
rect -18324 -3067 -18286 -3033
rect -18686 -3078 -18286 -3067
rect 7332 -3342 7360 -2991
rect 7298 -3394 7360 -3342
rect 7332 -3742 7360 -3394
rect 7298 -3766 7360 -3742
rect 8246 -2991 8308 -2966
rect 8280 -3342 8308 -2991
rect 8246 -3394 8308 -3342
rect 8280 -3742 8308 -3394
rect 8246 -3766 8308 -3742
rect 9182 -2991 9244 -2966
rect 9216 -3342 9244 -2991
rect 9182 -3394 9244 -3342
rect 9216 -3742 9244 -3394
rect 9182 -3766 9244 -3742
rect 10113 -2990 10175 -2965
rect 10147 -3341 10175 -2990
rect 10113 -3393 10175 -3341
rect 10147 -3741 10175 -3393
rect 10113 -3765 10175 -3741
rect 11040 -2991 11102 -2966
rect 11074 -3342 11102 -2991
rect 11040 -3394 11102 -3342
rect 11074 -3742 11102 -3394
rect 11040 -3766 11102 -3742
rect 12157 -3279 12407 -3262
rect 12157 -3340 12183 -3279
rect 12382 -3340 12407 -3279
rect 12923 -3275 13123 -3273
rect 12923 -3309 12954 -3275
rect 13086 -3309 13123 -3275
rect 12923 -3316 13123 -3309
rect 12157 -3358 12407 -3340
rect -23584 -4771 -23384 -4769
rect -23584 -4805 -23553 -4771
rect -23421 -4805 -23384 -4771
rect -23584 -4812 -23384 -4805
rect -24162 -4845 -23762 -4819
rect -24162 -4879 -24135 -4845
rect -23800 -4879 -23762 -4845
rect -24162 -4890 -23762 -4879
rect -21846 -4771 -21646 -4769
rect -21846 -4805 -21815 -4771
rect -21683 -4805 -21646 -4771
rect -21846 -4812 -21646 -4805
rect -22426 -4845 -22026 -4819
rect -22426 -4879 -22399 -4845
rect -22064 -4879 -22026 -4845
rect -22426 -4890 -22026 -4879
rect -20644 -5230 -19442 -5208
rect -20644 -5276 -20603 -5230
rect -19480 -5276 -19442 -5230
rect -20644 -5299 -19442 -5276
rect -19085 -5230 -17883 -5208
rect -19085 -5276 -19044 -5230
rect -17921 -5276 -17883 -5230
rect -19085 -5299 -17883 -5276
rect -17353 -5230 -16151 -5208
rect -17353 -5276 -17312 -5230
rect -16189 -5276 -16151 -5230
rect -17353 -5299 -16151 -5276
rect -15794 -5230 -14592 -5208
rect -15794 -5276 -15753 -5230
rect -14630 -5276 -14592 -5230
rect -15794 -5299 -14592 -5276
rect -14062 -5230 -12860 -5208
rect -14062 -5276 -14021 -5230
rect -12898 -5276 -12860 -5230
rect -14062 -5299 -12860 -5276
rect -12503 -5230 -11301 -5208
rect -12503 -5276 -12462 -5230
rect -11339 -5276 -11301 -5230
rect -12503 -5299 -11301 -5276
rect -10771 -5230 -9569 -5208
rect -10771 -5276 -10730 -5230
rect -9607 -5276 -9569 -5230
rect -10771 -5299 -9569 -5276
rect -9212 -5230 -8010 -5208
rect -9212 -5276 -9171 -5230
rect -8048 -5276 -8010 -5230
rect -9212 -5299 -8010 -5276
rect 5658 -5685 5858 -5683
rect 5658 -5719 5689 -5685
rect 5821 -5719 5858 -5685
rect 5658 -5726 5858 -5719
rect 6098 -5685 6298 -5683
rect 6098 -5719 6129 -5685
rect 6261 -5719 6298 -5685
rect 6098 -5726 6298 -5719
rect 6538 -5685 6738 -5683
rect 6538 -5719 6569 -5685
rect 6701 -5719 6738 -5685
rect 6538 -5726 6738 -5719
rect -23586 -6063 -23386 -6061
rect -23586 -6097 -23555 -6063
rect -23423 -6097 -23386 -6063
rect -23586 -6104 -23386 -6097
rect -24162 -6137 -23762 -6111
rect -24162 -6171 -24135 -6137
rect -23800 -6171 -23762 -6137
rect -24162 -6182 -23762 -6171
rect -21852 -6063 -21652 -6061
rect -21852 -6097 -21821 -6063
rect -21689 -6097 -21652 -6063
rect -21852 -6104 -21652 -6097
rect -22426 -6137 -22026 -6111
rect -22426 -6171 -22399 -6137
rect -22064 -6171 -22026 -6137
rect -22426 -6182 -22026 -6171
rect -20296 -6305 -19896 -6279
rect -20296 -6339 -20269 -6305
rect -19934 -6339 -19896 -6305
rect -20296 -6350 -19896 -6339
rect -19187 -6305 -18787 -6279
rect -19187 -6339 -19160 -6305
rect -18825 -6339 -18787 -6305
rect -19187 -6350 -18787 -6339
rect -18305 -6305 -17905 -6279
rect -18305 -6339 -18278 -6305
rect -17943 -6339 -17905 -6305
rect -18305 -6350 -17905 -6339
rect -17005 -6305 -16605 -6279
rect -17005 -6339 -16978 -6305
rect -16643 -6339 -16605 -6305
rect -17005 -6350 -16605 -6339
rect -15896 -6305 -15496 -6279
rect -15896 -6339 -15869 -6305
rect -15534 -6339 -15496 -6305
rect -15896 -6350 -15496 -6339
rect -15014 -6305 -14614 -6279
rect -15014 -6339 -14987 -6305
rect -14652 -6339 -14614 -6305
rect -15014 -6350 -14614 -6339
rect -13714 -6305 -13314 -6279
rect -13714 -6339 -13687 -6305
rect -13352 -6339 -13314 -6305
rect -13714 -6350 -13314 -6339
rect -12605 -6305 -12205 -6279
rect -12605 -6339 -12578 -6305
rect -12243 -6339 -12205 -6305
rect -12605 -6350 -12205 -6339
rect -11723 -6305 -11323 -6279
rect -11723 -6339 -11696 -6305
rect -11361 -6339 -11323 -6305
rect -11723 -6350 -11323 -6339
rect -10423 -6305 -10023 -6279
rect -10423 -6339 -10396 -6305
rect -10061 -6339 -10023 -6305
rect -10423 -6350 -10023 -6339
rect -9314 -6305 -8914 -6279
rect -9314 -6339 -9287 -6305
rect -8952 -6339 -8914 -6305
rect -9314 -6350 -8914 -6339
rect -8432 -6305 -8032 -6279
rect -8432 -6339 -8405 -6305
rect -8070 -6339 -8032 -6305
rect -8432 -6350 -8032 -6339
rect 7298 -6490 7360 -6466
rect 7332 -6838 7360 -6490
rect 7298 -6890 7360 -6838
rect 7332 -7241 7360 -6890
rect 7298 -7266 7360 -7241
rect 8246 -6490 8308 -6466
rect 8280 -6838 8308 -6490
rect 8246 -6890 8308 -6838
rect 8280 -7241 8308 -6890
rect 8246 -7266 8308 -7241
rect 9182 -6490 9244 -6466
rect 9216 -6838 9244 -6490
rect 9182 -6890 9244 -6838
rect 9216 -7241 9244 -6890
rect 9182 -7266 9244 -7241
rect 10113 -6490 10175 -6466
rect 10147 -6838 10175 -6490
rect 10113 -6890 10175 -6838
rect 10147 -7241 10175 -6890
rect 10113 -7266 10175 -7241
rect 11040 -6490 11102 -6466
rect 11074 -6838 11102 -6490
rect 11040 -6890 11102 -6838
rect 11074 -7241 11102 -6890
rect 11040 -7266 11102 -7241
rect 7298 -7419 7360 -7394
rect 7332 -7770 7360 -7419
rect -23584 -8036 -23384 -8034
rect -23584 -8070 -23553 -8036
rect -23421 -8070 -23384 -8036
rect -23584 -8077 -23384 -8070
rect -24162 -8110 -23762 -8084
rect -24162 -8144 -24135 -8110
rect -23800 -8144 -23762 -8110
rect -24162 -8155 -23762 -8144
rect -21850 -8036 -21650 -8034
rect -21850 -8070 -21819 -8036
rect -21687 -8070 -21650 -8036
rect -21850 -8077 -21650 -8070
rect -22425 -8110 -22025 -8084
rect -22425 -8144 -22398 -8110
rect -22063 -8144 -22025 -8110
rect -22425 -8155 -22025 -8144
rect 7298 -7822 7360 -7770
rect 7332 -8170 7360 -7822
rect 7298 -8194 7360 -8170
rect 8246 -7419 8308 -7394
rect 8280 -7770 8308 -7419
rect 8246 -7822 8308 -7770
rect 8280 -8170 8308 -7822
rect 8246 -8194 8308 -8170
rect 9182 -7419 9244 -7394
rect 9216 -7770 9244 -7419
rect 9182 -7822 9244 -7770
rect 9216 -8170 9244 -7822
rect 9182 -8194 9244 -8170
rect 10113 -7418 10175 -7393
rect 10147 -7769 10175 -7418
rect 10113 -7821 10175 -7769
rect 10147 -8169 10175 -7821
rect 10113 -8193 10175 -8169
rect 11040 -7419 11102 -7394
rect 11074 -7770 11102 -7419
rect 11040 -7822 11102 -7770
rect 11074 -8170 11102 -7822
rect -20644 -8495 -19442 -8473
rect -20644 -8541 -20603 -8495
rect -19480 -8541 -19442 -8495
rect -20644 -8564 -19442 -8541
rect -19085 -8495 -17883 -8473
rect -19085 -8541 -19044 -8495
rect -17921 -8541 -17883 -8495
rect -19085 -8564 -17883 -8541
rect -17353 -8495 -16151 -8473
rect -17353 -8541 -17312 -8495
rect -16189 -8541 -16151 -8495
rect -17353 -8564 -16151 -8541
rect -15794 -8495 -14592 -8473
rect -15794 -8541 -15753 -8495
rect -14630 -8541 -14592 -8495
rect -15794 -8564 -14592 -8541
rect -14062 -8495 -12860 -8473
rect -14062 -8541 -14021 -8495
rect -12898 -8541 -12860 -8495
rect -14062 -8564 -12860 -8541
rect -12503 -8495 -11301 -8473
rect -12503 -8541 -12462 -8495
rect -11339 -8541 -11301 -8495
rect -12503 -8564 -11301 -8541
rect -10771 -8495 -9569 -8473
rect -10771 -8541 -10730 -8495
rect -9607 -8541 -9569 -8495
rect -10771 -8564 -9569 -8541
rect -9212 -8495 -8010 -8473
rect -9212 -8541 -9171 -8495
rect -8048 -8541 -8010 -8495
rect -9212 -8564 -8010 -8541
rect 11040 -8194 11102 -8170
rect 12157 -7707 12407 -7690
rect 12157 -7768 12183 -7707
rect 12382 -7768 12407 -7707
rect 12923 -7703 13123 -7701
rect 12923 -7737 12954 -7703
rect 13086 -7737 13123 -7703
rect 12923 -7744 13123 -7737
rect 12157 -7786 12407 -7768
rect -23583 -9328 -23383 -9326
rect -23583 -9362 -23552 -9328
rect -23420 -9362 -23383 -9328
rect -23583 -9369 -23383 -9362
rect -24162 -9402 -23762 -9376
rect -24162 -9436 -24135 -9402
rect -23800 -9436 -23762 -9402
rect -24162 -9447 -23762 -9436
rect -21846 -9328 -21646 -9326
rect -21846 -9362 -21815 -9328
rect -21683 -9362 -21646 -9328
rect -21846 -9369 -21646 -9362
rect -22426 -9402 -22026 -9376
rect -22426 -9436 -22399 -9402
rect -22064 -9436 -22026 -9402
rect -22426 -9447 -22026 -9436
rect -20296 -9570 -19896 -9544
rect -20296 -9604 -20269 -9570
rect -19934 -9604 -19896 -9570
rect -20296 -9615 -19896 -9604
rect -19187 -9570 -18787 -9544
rect -19187 -9604 -19160 -9570
rect -18825 -9604 -18787 -9570
rect -19187 -9615 -18787 -9604
rect -18305 -9570 -17905 -9544
rect -18305 -9604 -18278 -9570
rect -17943 -9604 -17905 -9570
rect -18305 -9615 -17905 -9604
rect -17005 -9570 -16605 -9544
rect -17005 -9604 -16978 -9570
rect -16643 -9604 -16605 -9570
rect -17005 -9615 -16605 -9604
rect -15896 -9570 -15496 -9544
rect -15896 -9604 -15869 -9570
rect -15534 -9604 -15496 -9570
rect -15896 -9615 -15496 -9604
rect -15014 -9570 -14614 -9544
rect -15014 -9604 -14987 -9570
rect -14652 -9604 -14614 -9570
rect -15014 -9615 -14614 -9604
rect -13714 -9570 -13314 -9544
rect -13714 -9604 -13687 -9570
rect -13352 -9604 -13314 -9570
rect -13714 -9615 -13314 -9604
rect -12605 -9570 -12205 -9544
rect -12605 -9604 -12578 -9570
rect -12243 -9604 -12205 -9570
rect -12605 -9615 -12205 -9604
rect -11723 -9570 -11323 -9544
rect -11723 -9604 -11696 -9570
rect -11361 -9604 -11323 -9570
rect -11723 -9615 -11323 -9604
rect -10423 -9570 -10023 -9544
rect -10423 -9604 -10396 -9570
rect -10061 -9604 -10023 -9570
rect -10423 -9615 -10023 -9604
rect -9314 -9570 -8914 -9544
rect -9314 -9604 -9287 -9570
rect -8952 -9604 -8914 -9570
rect -9314 -9615 -8914 -9604
rect -8432 -9570 -8032 -9544
rect -8432 -9604 -8405 -9570
rect -8070 -9604 -8032 -9570
rect -8432 -9615 -8032 -9604
rect 5658 -10313 5858 -10311
rect 5658 -10347 5689 -10313
rect 5821 -10347 5858 -10313
rect 5658 -10354 5858 -10347
rect 6098 -10313 6298 -10311
rect 6098 -10347 6129 -10313
rect 6261 -10347 6298 -10313
rect 6098 -10354 6298 -10347
rect 6538 -10313 6738 -10311
rect 6538 -10347 6569 -10313
rect 6701 -10347 6738 -10313
rect 6538 -10354 6738 -10347
rect -23583 -11300 -23383 -11298
rect -23583 -11334 -23552 -11300
rect -23420 -11334 -23383 -11300
rect -23583 -11341 -23383 -11334
rect -24162 -11374 -23762 -11348
rect -24162 -11408 -24135 -11374
rect -23800 -11408 -23762 -11374
rect -24162 -11419 -23762 -11408
rect -21850 -11300 -21650 -11298
rect -21850 -11334 -21819 -11300
rect -21687 -11334 -21650 -11300
rect -21850 -11341 -21650 -11334
rect -22425 -11374 -22025 -11348
rect -22425 -11408 -22398 -11374
rect -22063 -11408 -22025 -11374
rect -22425 -11419 -22025 -11408
rect 7298 -11118 7360 -11094
rect 7332 -11466 7360 -11118
rect 7298 -11518 7360 -11466
rect -20644 -11759 -19442 -11737
rect -20644 -11805 -20603 -11759
rect -19480 -11805 -19442 -11759
rect -20644 -11828 -19442 -11805
rect -19085 -11759 -17883 -11737
rect -19085 -11805 -19044 -11759
rect -17921 -11805 -17883 -11759
rect -19085 -11828 -17883 -11805
rect -17353 -11759 -16151 -11737
rect -17353 -11805 -17312 -11759
rect -16189 -11805 -16151 -11759
rect -17353 -11828 -16151 -11805
rect -15794 -11759 -14592 -11737
rect -15794 -11805 -15753 -11759
rect -14630 -11805 -14592 -11759
rect -15794 -11828 -14592 -11805
rect -14062 -11759 -12860 -11737
rect -14062 -11805 -14021 -11759
rect -12898 -11805 -12860 -11759
rect -14062 -11828 -12860 -11805
rect -12503 -11759 -11301 -11737
rect -12503 -11805 -12462 -11759
rect -11339 -11805 -11301 -11759
rect -12503 -11828 -11301 -11805
rect -10771 -11759 -9569 -11737
rect -10771 -11805 -10730 -11759
rect -9607 -11805 -9569 -11759
rect -10771 -11828 -9569 -11805
rect -9212 -11759 -8010 -11737
rect -9212 -11805 -9171 -11759
rect -8048 -11805 -8010 -11759
rect -9212 -11828 -8010 -11805
rect 7332 -11869 7360 -11518
rect 7298 -11894 7360 -11869
rect 8246 -11118 8308 -11094
rect 8280 -11466 8308 -11118
rect 8246 -11518 8308 -11466
rect 8280 -11869 8308 -11518
rect 8246 -11894 8308 -11869
rect 9182 -11118 9244 -11094
rect 9216 -11466 9244 -11118
rect 9182 -11518 9244 -11466
rect 9216 -11869 9244 -11518
rect 9182 -11894 9244 -11869
rect 10113 -11118 10175 -11094
rect 10147 -11466 10175 -11118
rect 10113 -11518 10175 -11466
rect 10147 -11869 10175 -11518
rect 10113 -11894 10175 -11869
rect 11040 -11118 11102 -11094
rect 11074 -11466 11102 -11118
rect 11040 -11518 11102 -11466
rect 11074 -11869 11102 -11518
rect 11040 -11894 11102 -11869
rect 7298 -12047 7360 -12022
rect 7332 -12398 7360 -12047
rect 7298 -12450 7360 -12398
rect -23583 -12592 -23383 -12590
rect -23583 -12626 -23552 -12592
rect -23420 -12626 -23383 -12592
rect -23583 -12633 -23383 -12626
rect -24162 -12666 -23762 -12640
rect -24162 -12700 -24135 -12666
rect -23800 -12700 -23762 -12666
rect -24162 -12711 -23762 -12700
rect -21854 -12592 -21654 -12590
rect -21854 -12626 -21823 -12592
rect -21691 -12626 -21654 -12592
rect -21854 -12633 -21654 -12626
rect -22425 -12666 -22025 -12640
rect -22425 -12700 -22398 -12666
rect -22063 -12700 -22025 -12666
rect -22425 -12711 -22025 -12700
rect -20296 -12834 -19896 -12808
rect -20296 -12868 -20269 -12834
rect -19934 -12868 -19896 -12834
rect -20296 -12879 -19896 -12868
rect -19187 -12834 -18787 -12808
rect -19187 -12868 -19160 -12834
rect -18825 -12868 -18787 -12834
rect -19187 -12879 -18787 -12868
rect -18305 -12834 -17905 -12808
rect -18305 -12868 -18278 -12834
rect -17943 -12868 -17905 -12834
rect -18305 -12879 -17905 -12868
rect -17005 -12834 -16605 -12808
rect -17005 -12868 -16978 -12834
rect -16643 -12868 -16605 -12834
rect -17005 -12879 -16605 -12868
rect -15896 -12834 -15496 -12808
rect -15896 -12868 -15869 -12834
rect -15534 -12868 -15496 -12834
rect -15896 -12879 -15496 -12868
rect -15014 -12834 -14614 -12808
rect -15014 -12868 -14987 -12834
rect -14652 -12868 -14614 -12834
rect -15014 -12879 -14614 -12868
rect -13714 -12834 -13314 -12808
rect -13714 -12868 -13687 -12834
rect -13352 -12868 -13314 -12834
rect -13714 -12879 -13314 -12868
rect -12605 -12834 -12205 -12808
rect -12605 -12868 -12578 -12834
rect -12243 -12868 -12205 -12834
rect -12605 -12879 -12205 -12868
rect -11723 -12834 -11323 -12808
rect -11723 -12868 -11696 -12834
rect -11361 -12868 -11323 -12834
rect -11723 -12879 -11323 -12868
rect -10423 -12834 -10023 -12808
rect -10423 -12868 -10396 -12834
rect -10061 -12868 -10023 -12834
rect -10423 -12879 -10023 -12868
rect -9314 -12834 -8914 -12808
rect -9314 -12868 -9287 -12834
rect -8952 -12868 -8914 -12834
rect -9314 -12879 -8914 -12868
rect -8432 -12834 -8032 -12808
rect 7332 -12798 7360 -12450
rect 7298 -12822 7360 -12798
rect 8246 -12047 8308 -12022
rect 8280 -12398 8308 -12047
rect 8246 -12450 8308 -12398
rect 8280 -12798 8308 -12450
rect 8246 -12822 8308 -12798
rect 9182 -12047 9244 -12022
rect 9216 -12398 9244 -12047
rect 9182 -12450 9244 -12398
rect 9216 -12798 9244 -12450
rect 9182 -12822 9244 -12798
rect 10113 -12046 10175 -12021
rect 10147 -12397 10175 -12046
rect 10113 -12449 10175 -12397
rect 10147 -12797 10175 -12449
rect 10113 -12821 10175 -12797
rect 11040 -12047 11102 -12022
rect 11074 -12398 11102 -12047
rect 11040 -12450 11102 -12398
rect 11074 -12798 11102 -12450
rect -8432 -12868 -8405 -12834
rect -8070 -12868 -8032 -12834
rect -8432 -12879 -8032 -12868
rect 11040 -12822 11102 -12798
rect 12157 -12335 12407 -12318
rect 12157 -12396 12183 -12335
rect 12382 -12396 12407 -12335
rect 12923 -12331 13123 -12329
rect 12923 -12365 12954 -12331
rect 13086 -12365 13123 -12331
rect 12923 -12372 13123 -12365
rect 12157 -12414 12407 -12396
rect -1462 -13869 -1419 -13832
rect -1462 -14001 -1460 -13869
rect -1426 -14001 -1419 -13869
rect -1462 -14032 -1419 -14001
rect -23855 -14954 -23784 -14916
rect -23855 -15289 -23829 -14954
rect -23795 -15289 -23784 -14954
rect -16934 -14908 -16838 -14883
rect -23855 -15316 -23784 -15289
rect -16934 -15107 -16917 -14908
rect -16856 -15107 -16838 -14908
rect -16934 -15133 -16838 -15107
rect -11092 -14222 -11001 -14184
rect -11092 -15345 -11070 -14222
rect -11024 -15345 -11001 -14222
rect -4178 -14234 -4135 -14203
rect -4178 -14366 -4176 -14234
rect -4142 -14366 -4135 -14234
rect -4178 -14403 -4135 -14366
rect -1462 -14248 -1419 -14211
rect -1462 -14380 -1460 -14248
rect -1426 -14380 -1419 -14248
rect -1462 -14411 -1419 -14380
rect -4178 -14674 -4135 -14643
rect -4178 -14806 -4176 -14674
rect -4142 -14806 -4135 -14674
rect -4178 -14843 -4135 -14806
rect -1462 -14688 -1419 -14651
rect -1462 -14820 -1460 -14688
rect -1426 -14820 -1419 -14688
rect -1462 -14851 -1419 -14820
rect 5658 -14841 5858 -14839
rect 5658 -14875 5689 -14841
rect 5821 -14875 5858 -14841
rect 5658 -14882 5858 -14875
rect 6098 -14841 6298 -14839
rect 6098 -14875 6129 -14841
rect 6261 -14875 6298 -14841
rect 6098 -14882 6298 -14875
rect 6538 -14841 6738 -14839
rect 6538 -14875 6569 -14841
rect 6701 -14875 6738 -14841
rect 6538 -14882 6738 -14875
rect -4178 -15053 -4135 -15022
rect -4178 -15185 -4176 -15053
rect -4142 -15185 -4135 -15053
rect -4178 -15222 -4135 -15185
rect -1462 -15067 -1419 -15030
rect -1462 -15199 -1460 -15067
rect -1426 -15199 -1419 -15067
rect -1462 -15230 -1419 -15199
rect -11092 -15386 -11001 -15345
rect -7529 -15397 -7486 -15360
rect -7529 -15529 -7527 -15397
rect -7493 -15529 -7486 -15397
rect -7529 -15560 -7486 -15529
rect -4178 -15493 -4135 -15462
rect -4178 -15625 -4176 -15493
rect -4142 -15625 -4135 -15493
rect -4178 -15662 -4135 -15625
rect -1462 -15507 -1419 -15470
rect -1462 -15639 -1460 -15507
rect -1426 -15639 -1419 -15507
rect -1462 -15670 -1419 -15639
rect 7298 -15646 7360 -15622
rect -7528 -15897 -7485 -15860
rect -7528 -16029 -7526 -15897
rect -7492 -16029 -7485 -15897
rect -7528 -16060 -7485 -16029
rect -4178 -15872 -4135 -15841
rect -4178 -16004 -4176 -15872
rect -4142 -16004 -4135 -15872
rect -4178 -16041 -4135 -16004
rect -23854 -16139 -23783 -16101
rect -23854 -16474 -23828 -16139
rect -23794 -16474 -23783 -16139
rect -1462 -15886 -1419 -15849
rect -1462 -16018 -1460 -15886
rect -1426 -16018 -1419 -15886
rect -1462 -16049 -1419 -16018
rect 7332 -15994 7360 -15646
rect 7298 -16046 7360 -15994
rect -16934 -16308 -16838 -16283
rect -23854 -16501 -23783 -16474
rect -16934 -16507 -16917 -16308
rect -16856 -16507 -16838 -16308
rect -16934 -16533 -16838 -16507
rect -7529 -16377 -7486 -16340
rect -7529 -16509 -7527 -16377
rect -7493 -16509 -7486 -16377
rect -4178 -16312 -4135 -16281
rect -4178 -16444 -4176 -16312
rect -4142 -16444 -4135 -16312
rect -4178 -16481 -4135 -16444
rect -7529 -16540 -7486 -16509
rect -1462 -16326 -1419 -16289
rect -1462 -16458 -1460 -16326
rect -1426 -16458 -1419 -16326
rect 7332 -16397 7360 -16046
rect 7298 -16422 7360 -16397
rect 8246 -15646 8308 -15622
rect 8280 -15994 8308 -15646
rect 8246 -16046 8308 -15994
rect 8280 -16397 8308 -16046
rect 8246 -16422 8308 -16397
rect 9182 -15646 9244 -15622
rect 9216 -15994 9244 -15646
rect 9182 -16046 9244 -15994
rect 9216 -16397 9244 -16046
rect 9182 -16422 9244 -16397
rect 10113 -15646 10175 -15622
rect 10147 -15994 10175 -15646
rect 10113 -16046 10175 -15994
rect 10147 -16397 10175 -16046
rect 10113 -16422 10175 -16397
rect 11040 -15646 11102 -15622
rect 11074 -15994 11102 -15646
rect 11040 -16046 11102 -15994
rect 11074 -16397 11102 -16046
rect 11040 -16422 11102 -16397
rect -1462 -16489 -1419 -16458
rect 7298 -16575 7360 -16550
rect -23849 -17352 -23778 -17314
rect -23849 -17687 -23823 -17352
rect -23789 -17687 -23778 -17352
rect -23849 -17714 -23778 -17687
rect -16934 -17708 -16838 -17683
rect -20968 -18085 -20925 -18048
rect -20968 -18217 -20966 -18085
rect -20932 -18217 -20925 -18085
rect -20968 -18248 -20925 -18217
rect -16934 -17907 -16917 -17708
rect -16856 -17907 -16838 -17708
rect -16934 -17933 -16838 -17907
rect -15377 -17956 -15334 -17919
rect -15377 -18088 -15375 -17956
rect -15341 -18088 -15334 -17956
rect -15377 -18119 -15334 -18088
rect -11090 -17038 -10999 -17000
rect -11090 -18161 -11068 -17038
rect -11022 -18161 -10999 -17038
rect -7529 -16877 -7486 -16840
rect -4178 -16691 -4135 -16660
rect -4178 -16823 -4176 -16691
rect -4142 -16823 -4135 -16691
rect -4178 -16860 -4135 -16823
rect -7529 -17009 -7527 -16877
rect -7493 -17009 -7486 -16877
rect -1462 -16705 -1419 -16668
rect -1462 -16837 -1460 -16705
rect -1426 -16837 -1419 -16705
rect -1462 -16868 -1419 -16837
rect 7332 -16926 7360 -16575
rect 7298 -16978 7360 -16926
rect -7529 -17040 -7486 -17009
rect -4178 -17131 -4135 -17100
rect -4178 -17263 -4176 -17131
rect -4142 -17263 -4135 -17131
rect -4178 -17300 -4135 -17263
rect -7529 -17357 -7486 -17320
rect -1462 -17145 -1419 -17108
rect -1462 -17277 -1460 -17145
rect -1426 -17277 -1419 -17145
rect -1462 -17308 -1419 -17277
rect 7332 -17326 7360 -16978
rect -7529 -17489 -7527 -17357
rect -7493 -17489 -7486 -17357
rect 7298 -17350 7360 -17326
rect 8246 -16575 8308 -16550
rect 8280 -16926 8308 -16575
rect 8246 -16978 8308 -16926
rect 8280 -17326 8308 -16978
rect 8246 -17350 8308 -17326
rect 9182 -16575 9244 -16550
rect 9216 -16926 9244 -16575
rect 9182 -16978 9244 -16926
rect 9216 -17326 9244 -16978
rect 9182 -17350 9244 -17326
rect 10113 -16574 10175 -16549
rect 10147 -16925 10175 -16574
rect 10113 -16977 10175 -16925
rect 10147 -17325 10175 -16977
rect 10113 -17349 10175 -17325
rect 11040 -16575 11102 -16550
rect 11074 -16926 11102 -16575
rect 11040 -16978 11102 -16926
rect 11074 -17326 11102 -16978
rect -7529 -17520 -7486 -17489
rect -4178 -17510 -4135 -17479
rect -4178 -17642 -4176 -17510
rect -4142 -17642 -4135 -17510
rect -4178 -17679 -4135 -17642
rect -1462 -17524 -1419 -17487
rect -1462 -17656 -1460 -17524
rect -1426 -17656 -1419 -17524
rect -1462 -17687 -1419 -17656
rect -7529 -17817 -7486 -17780
rect 11040 -17350 11102 -17326
rect 16147 -16814 16589 -16738
rect 12157 -16863 12407 -16846
rect 12157 -16924 12183 -16863
rect 12382 -16924 12407 -16863
rect 12923 -16859 13123 -16857
rect 12923 -16893 12954 -16859
rect 13086 -16893 13123 -16859
rect 12923 -16900 13123 -16893
rect 12157 -16942 12407 -16924
rect 16147 -16927 16211 -16814
rect 16541 -16927 16589 -16814
rect 16147 -16995 16589 -16927
rect -7529 -17949 -7527 -17817
rect -7493 -17949 -7486 -17817
rect -7529 -17980 -7486 -17949
rect -4178 -17950 -4135 -17919
rect -4178 -18082 -4176 -17950
rect -4142 -18082 -4135 -17950
rect -4178 -18119 -4135 -18082
rect -1462 -17964 -1419 -17927
rect -1462 -18096 -1460 -17964
rect -1426 -18096 -1419 -17964
rect -1462 -18127 -1419 -18096
rect -11090 -18202 -10999 -18161
rect -23834 -18471 -23763 -18433
rect -23834 -18806 -23808 -18471
rect -23774 -18806 -23763 -18471
rect -20967 -18585 -20924 -18548
rect -20967 -18717 -20965 -18585
rect -20931 -18717 -20924 -18585
rect -15376 -18456 -15333 -18419
rect -15376 -18588 -15374 -18456
rect -15340 -18588 -15333 -18456
rect -7543 -18277 -7500 -18240
rect -7543 -18409 -7541 -18277
rect -7507 -18409 -7500 -18277
rect -7543 -18440 -7500 -18409
rect -4178 -18329 -4135 -18298
rect -4178 -18461 -4176 -18329
rect -4142 -18461 -4135 -18329
rect -4178 -18498 -4135 -18461
rect -1462 -18343 -1419 -18306
rect -1462 -18475 -1460 -18343
rect -1426 -18475 -1419 -18343
rect -1462 -18506 -1419 -18475
rect -15376 -18619 -15333 -18588
rect -20967 -18748 -20924 -18717
rect -23834 -18833 -23763 -18806
rect -20968 -19065 -20925 -19028
rect -20968 -19197 -20966 -19065
rect -20932 -19197 -20925 -19065
rect -20968 -19228 -20925 -19197
rect -16934 -19108 -16838 -19083
rect -15377 -18936 -15334 -18899
rect -7541 -18757 -7498 -18720
rect -7541 -18889 -7539 -18757
rect -7505 -18889 -7498 -18757
rect -7541 -18920 -7498 -18889
rect -15377 -19068 -15375 -18936
rect -15341 -19068 -15334 -18936
rect -4178 -18769 -4135 -18738
rect -4178 -18901 -4176 -18769
rect -4142 -18901 -4135 -18769
rect -4178 -18938 -4135 -18901
rect -1462 -18783 -1419 -18746
rect -1462 -18915 -1460 -18783
rect -1426 -18915 -1419 -18783
rect -1462 -18946 -1419 -18915
rect -15377 -19099 -15334 -19068
rect -23832 -19665 -23761 -19627
rect -23832 -20000 -23806 -19665
rect -23772 -20000 -23761 -19665
rect -20968 -19565 -20925 -19528
rect -20968 -19697 -20966 -19565
rect -20932 -19697 -20925 -19565
rect -20968 -19728 -20925 -19697
rect -16934 -19307 -16917 -19108
rect -16856 -19307 -16838 -19108
rect -16934 -19333 -16838 -19307
rect -4178 -19148 -4135 -19117
rect -4178 -19280 -4176 -19148
rect -4142 -19280 -4135 -19148
rect -4178 -19317 -4135 -19280
rect -1462 -19162 -1419 -19125
rect -1462 -19294 -1460 -19162
rect -1426 -19294 -1419 -19162
rect -1462 -19325 -1419 -19294
rect -15377 -19436 -15334 -19399
rect 5658 -19369 5858 -19367
rect 5658 -19403 5689 -19369
rect 5821 -19403 5858 -19369
rect 5658 -19410 5858 -19403
rect 6098 -19369 6298 -19367
rect 6098 -19403 6129 -19369
rect 6261 -19403 6298 -19369
rect 6098 -19410 6298 -19403
rect 6538 -19369 6738 -19367
rect 6538 -19403 6569 -19369
rect 6701 -19403 6738 -19369
rect 6538 -19410 6738 -19403
rect -15377 -19568 -15375 -19436
rect -15341 -19568 -15334 -19436
rect -15377 -19599 -15334 -19568
rect -4178 -19588 -4135 -19557
rect -4178 -19720 -4176 -19588
rect -4142 -19720 -4135 -19588
rect -4178 -19757 -4135 -19720
rect -1462 -19602 -1419 -19565
rect -1462 -19734 -1460 -19602
rect -1426 -19734 -1419 -19602
rect -1462 -19765 -1419 -19734
rect 17528 -18895 17928 -18869
rect 17528 -18929 17555 -18895
rect 17890 -18929 17928 -18895
rect 17528 -18940 17928 -18929
rect 18096 -18899 18296 -18897
rect 18096 -18933 18127 -18899
rect 18259 -18933 18296 -18899
rect 18096 -18940 18296 -18933
rect -23832 -20027 -23761 -20000
rect -20968 -20045 -20925 -20008
rect -20968 -20177 -20966 -20045
rect -20932 -20177 -20925 -20045
rect -15377 -19916 -15334 -19879
rect -15377 -20048 -15375 -19916
rect -15341 -20048 -15334 -19916
rect -15377 -20079 -15334 -20048
rect -20968 -20208 -20925 -20177
rect -20968 -20505 -20925 -20468
rect -20968 -20637 -20966 -20505
rect -20932 -20637 -20925 -20505
rect -20968 -20668 -20925 -20637
rect -16934 -20508 -16838 -20483
rect -23801 -20865 -23730 -20827
rect -23801 -21200 -23775 -20865
rect -23741 -21200 -23730 -20865
rect -20982 -20965 -20939 -20928
rect -20982 -21097 -20980 -20965
rect -20946 -21097 -20939 -20965
rect -20982 -21128 -20939 -21097
rect -16934 -20707 -16917 -20508
rect -16856 -20707 -16838 -20508
rect -15377 -20376 -15334 -20339
rect -15377 -20508 -15375 -20376
rect -15341 -20508 -15334 -20376
rect -15377 -20539 -15334 -20508
rect -16934 -20733 -16838 -20707
rect -15391 -20836 -15348 -20799
rect -15391 -20968 -15389 -20836
rect -15355 -20968 -15348 -20836
rect -15391 -20999 -15348 -20968
rect -11090 -19995 -10999 -19957
rect -23801 -21227 -23730 -21200
rect -11090 -21118 -11068 -19995
rect -11022 -21118 -10999 -19995
rect -4178 -19967 -4135 -19936
rect -4178 -20099 -4176 -19967
rect -4142 -20099 -4135 -19967
rect -4178 -20136 -4135 -20099
rect -1462 -19981 -1419 -19944
rect -1462 -20113 -1460 -19981
rect -1426 -20113 -1419 -19981
rect -1462 -20144 -1419 -20113
rect 7298 -20174 7360 -20150
rect -4178 -20407 -4135 -20376
rect -4178 -20539 -4176 -20407
rect -4142 -20539 -4135 -20407
rect -4178 -20576 -4135 -20539
rect -1462 -20421 -1419 -20384
rect -1462 -20553 -1460 -20421
rect -1426 -20553 -1419 -20421
rect -1462 -20584 -1419 -20553
rect 7332 -20522 7360 -20174
rect 7298 -20574 7360 -20522
rect -4178 -20786 -4135 -20755
rect -4178 -20918 -4176 -20786
rect -4142 -20918 -4135 -20786
rect -4178 -20955 -4135 -20918
rect 7332 -20925 7360 -20574
rect 7298 -20950 7360 -20925
rect 8246 -20174 8308 -20150
rect 8280 -20522 8308 -20174
rect 8246 -20574 8308 -20522
rect 8280 -20925 8308 -20574
rect 8246 -20950 8308 -20925
rect 9182 -20174 9244 -20150
rect 9216 -20522 9244 -20174
rect 9182 -20574 9244 -20522
rect 9216 -20925 9244 -20574
rect 9182 -20950 9244 -20925
rect 10113 -20174 10175 -20150
rect 10147 -20522 10175 -20174
rect 10113 -20574 10175 -20522
rect 10147 -20925 10175 -20574
rect 10113 -20950 10175 -20925
rect 11040 -20174 11102 -20150
rect 11074 -20522 11102 -20174
rect 11040 -20574 11102 -20522
rect 11074 -20925 11102 -20574
rect 11040 -20950 11102 -20925
rect 16147 -20245 16589 -20177
rect 16147 -20358 16211 -20245
rect 16541 -20358 16589 -20245
rect 16147 -20434 16589 -20358
rect -11090 -21159 -10999 -21118
rect 7298 -21103 7360 -21078
rect -20980 -21445 -20937 -21408
rect -20980 -21577 -20978 -21445
rect -20944 -21577 -20937 -21445
rect -15389 -21316 -15346 -21279
rect -15389 -21448 -15387 -21316
rect -15353 -21448 -15346 -21316
rect -15389 -21479 -15346 -21448
rect 7332 -21454 7360 -21103
rect 7298 -21506 7360 -21454
rect -20980 -21608 -20937 -21577
rect 7332 -21854 7360 -21506
rect 7298 -21878 7360 -21854
rect 8246 -21103 8308 -21078
rect 8280 -21454 8308 -21103
rect 8246 -21506 8308 -21454
rect 8280 -21854 8308 -21506
rect 8246 -21878 8308 -21854
rect 9182 -21103 9244 -21078
rect 9216 -21454 9244 -21103
rect 9182 -21506 9244 -21454
rect 9216 -21854 9244 -21506
rect 9182 -21878 9244 -21854
rect 10113 -21102 10175 -21077
rect 10147 -21453 10175 -21102
rect 10113 -21505 10175 -21453
rect 10147 -21853 10175 -21505
rect 10113 -21877 10175 -21853
rect 11040 -21103 11102 -21078
rect 11074 -21454 11102 -21103
rect 11040 -21506 11102 -21454
rect 11074 -21854 11102 -21506
rect -16934 -21908 -16838 -21883
rect -23802 -22168 -23731 -22130
rect -23802 -22503 -23776 -22168
rect -23742 -22503 -23731 -22168
rect -23802 -22530 -23731 -22503
rect -16934 -22107 -16917 -21908
rect -16856 -22107 -16838 -21908
rect -16934 -22133 -16838 -22107
rect 11040 -21878 11102 -21854
rect 12157 -21391 12407 -21374
rect 12157 -21452 12183 -21391
rect 12382 -21452 12407 -21391
rect 12923 -21387 13123 -21385
rect 12923 -21421 12954 -21387
rect 13086 -21421 13123 -21387
rect 12923 -21428 13123 -21421
rect 12157 -21470 12407 -21452
rect -16934 -23308 -16838 -23283
rect -23802 -23477 -23731 -23439
rect -23802 -23812 -23776 -23477
rect -23742 -23812 -23731 -23477
rect -23802 -23839 -23731 -23812
rect -16934 -23507 -16917 -23308
rect -16856 -23507 -16838 -23308
rect -16934 -23533 -16838 -23507
rect -11090 -22574 -10999 -22536
rect -11090 -23697 -11068 -22574
rect -11022 -23697 -10999 -22574
rect -11090 -23738 -10999 -23697
rect 5658 -23897 5858 -23895
rect 5658 -23931 5689 -23897
rect 5821 -23931 5858 -23897
rect 5658 -23938 5858 -23931
rect 6098 -23897 6298 -23895
rect 6098 -23931 6129 -23897
rect 6261 -23931 6298 -23897
rect 6098 -23938 6298 -23931
rect 6538 -23897 6738 -23895
rect 6538 -23931 6569 -23897
rect 6701 -23931 6738 -23897
rect 6538 -23938 6738 -23931
rect -16934 -24708 -16838 -24683
rect -16934 -24907 -16917 -24708
rect -16856 -24907 -16838 -24708
rect -16934 -24933 -16838 -24907
rect 7298 -24702 7360 -24678
rect 7332 -25050 7360 -24702
rect 7298 -25102 7360 -25050
rect -11090 -25342 -10999 -25304
rect -11090 -26465 -11068 -25342
rect -11022 -26465 -10999 -25342
rect 7332 -25453 7360 -25102
rect 7298 -25478 7360 -25453
rect 8246 -24702 8308 -24678
rect 8280 -25050 8308 -24702
rect 8246 -25102 8308 -25050
rect 8280 -25453 8308 -25102
rect 8246 -25478 8308 -25453
rect 9182 -24702 9244 -24678
rect 9216 -25050 9244 -24702
rect 9182 -25102 9244 -25050
rect 9216 -25453 9244 -25102
rect 9182 -25478 9244 -25453
rect 10113 -24702 10175 -24678
rect 10147 -25050 10175 -24702
rect 10113 -25102 10175 -25050
rect 10147 -25453 10175 -25102
rect 10113 -25478 10175 -25453
rect 11040 -24702 11102 -24678
rect 11074 -25050 11102 -24702
rect 11040 -25102 11102 -25050
rect 11074 -25453 11102 -25102
rect 11040 -25478 11102 -25453
rect 7298 -25631 7360 -25606
rect 7332 -25982 7360 -25631
rect 7298 -26034 7360 -25982
rect 7332 -26382 7360 -26034
rect 7298 -26406 7360 -26382
rect 8246 -25631 8308 -25606
rect 8280 -25982 8308 -25631
rect 8246 -26034 8308 -25982
rect 8280 -26382 8308 -26034
rect 8246 -26406 8308 -26382
rect 9182 -25631 9244 -25606
rect 9216 -25982 9244 -25631
rect 9182 -26034 9244 -25982
rect 9216 -26382 9244 -26034
rect 9182 -26406 9244 -26382
rect 10113 -25630 10175 -25605
rect 10147 -25981 10175 -25630
rect 10113 -26033 10175 -25981
rect 10147 -26381 10175 -26033
rect 10113 -26405 10175 -26381
rect 11040 -25631 11102 -25606
rect 11074 -25982 11102 -25631
rect 11040 -26034 11102 -25982
rect 11074 -26382 11102 -26034
rect -11090 -26506 -10999 -26465
rect 11040 -26406 11102 -26382
rect 12157 -25919 12407 -25902
rect 12157 -25980 12183 -25919
rect 12382 -25980 12407 -25919
rect 12923 -25915 13123 -25913
rect 12923 -25949 12954 -25915
rect 13086 -25949 13123 -25915
rect 12923 -25956 13123 -25949
rect 12157 -25998 12407 -25980
rect -11090 -27975 -10999 -27937
rect -11090 -29098 -11068 -27975
rect -11022 -29098 -10999 -27975
rect 5658 -28425 5858 -28423
rect 5658 -28459 5689 -28425
rect 5821 -28459 5858 -28425
rect 5658 -28466 5858 -28459
rect 6098 -28425 6298 -28423
rect 6098 -28459 6129 -28425
rect 6261 -28459 6298 -28425
rect 6098 -28466 6298 -28459
rect 6538 -28425 6738 -28423
rect 6538 -28459 6569 -28425
rect 6701 -28459 6738 -28425
rect 6538 -28466 6738 -28459
rect -11090 -29139 -10999 -29098
rect 7298 -29230 7360 -29206
rect 7332 -29578 7360 -29230
rect 7298 -29630 7360 -29578
rect 7332 -29981 7360 -29630
rect 7298 -30006 7360 -29981
rect 8246 -29230 8308 -29206
rect 8280 -29578 8308 -29230
rect 8246 -29630 8308 -29578
rect 8280 -29981 8308 -29630
rect 8246 -30006 8308 -29981
rect 9182 -29230 9244 -29206
rect 9216 -29578 9244 -29230
rect 9182 -29630 9244 -29578
rect 9216 -29981 9244 -29630
rect 9182 -30006 9244 -29981
rect 10113 -29230 10175 -29206
rect 10147 -29578 10175 -29230
rect 10113 -29630 10175 -29578
rect 10147 -29981 10175 -29630
rect 10113 -30006 10175 -29981
rect 11040 -29230 11102 -29206
rect 11074 -29578 11102 -29230
rect 11040 -29630 11102 -29578
rect 11074 -29981 11102 -29630
rect 11040 -30006 11102 -29981
rect 7298 -30159 7360 -30134
rect 7332 -30510 7360 -30159
rect -11090 -30584 -10999 -30546
rect -11090 -31707 -11068 -30584
rect -11022 -31707 -10999 -30584
rect 7298 -30562 7360 -30510
rect 7332 -30910 7360 -30562
rect 7298 -30934 7360 -30910
rect 8246 -30159 8308 -30134
rect 8280 -30510 8308 -30159
rect 8246 -30562 8308 -30510
rect 8280 -30910 8308 -30562
rect 8246 -30934 8308 -30910
rect 9182 -30159 9244 -30134
rect 9216 -30510 9244 -30159
rect 9182 -30562 9244 -30510
rect 9216 -30910 9244 -30562
rect 9182 -30934 9244 -30910
rect 10113 -30158 10175 -30133
rect 10147 -30509 10175 -30158
rect 10113 -30561 10175 -30509
rect 10147 -30909 10175 -30561
rect 10113 -30933 10175 -30909
rect 11040 -30159 11102 -30134
rect 11074 -30510 11102 -30159
rect 11040 -30562 11102 -30510
rect 11074 -30910 11102 -30562
rect 11040 -30934 11102 -30910
rect 12157 -30447 12407 -30430
rect 12157 -30508 12183 -30447
rect 12382 -30508 12407 -30447
rect 12923 -30443 13123 -30441
rect 12923 -30477 12954 -30443
rect 13086 -30477 13123 -30443
rect 12923 -30484 13123 -30477
rect 12157 -30526 12407 -30508
rect -11090 -31748 -10999 -31707
rect 5658 -32953 5858 -32951
rect 5658 -32987 5689 -32953
rect 5821 -32987 5858 -32953
rect 5658 -32994 5858 -32987
rect 6098 -32953 6298 -32951
rect 6098 -32987 6129 -32953
rect 6261 -32987 6298 -32953
rect 6098 -32994 6298 -32987
rect 6538 -32953 6738 -32951
rect 6538 -32987 6569 -32953
rect 6701 -32987 6738 -32953
rect 6538 -32994 6738 -32987
rect -11092 -33204 -11001 -33166
rect -11092 -34327 -11070 -33204
rect -11024 -34327 -11001 -33204
rect -11092 -34368 -11001 -34327
rect 7298 -33758 7360 -33734
rect 7332 -34106 7360 -33758
rect 7298 -34158 7360 -34106
rect 7332 -34509 7360 -34158
rect 7298 -34534 7360 -34509
rect 8246 -33758 8308 -33734
rect 8280 -34106 8308 -33758
rect 8246 -34158 8308 -34106
rect 8280 -34509 8308 -34158
rect 8246 -34534 8308 -34509
rect 9182 -33758 9244 -33734
rect 9216 -34106 9244 -33758
rect 9182 -34158 9244 -34106
rect 9216 -34509 9244 -34158
rect 9182 -34534 9244 -34509
rect 10113 -33758 10175 -33734
rect 10147 -34106 10175 -33758
rect 10113 -34158 10175 -34106
rect 10147 -34509 10175 -34158
rect 10113 -34534 10175 -34509
rect 11040 -33758 11102 -33734
rect 11074 -34106 11102 -33758
rect 11040 -34158 11102 -34106
rect 11074 -34509 11102 -34158
rect 11040 -34534 11102 -34509
rect 7298 -34687 7360 -34662
rect 7332 -35038 7360 -34687
rect 7298 -35090 7360 -35038
rect 7332 -35438 7360 -35090
rect 7298 -35462 7360 -35438
rect 8246 -34687 8308 -34662
rect 8280 -35038 8308 -34687
rect 8246 -35090 8308 -35038
rect 8280 -35438 8308 -35090
rect 8246 -35462 8308 -35438
rect 9182 -34687 9244 -34662
rect 9216 -35038 9244 -34687
rect 9182 -35090 9244 -35038
rect 9216 -35438 9244 -35090
rect 9182 -35462 9244 -35438
rect 10113 -34686 10175 -34661
rect 10147 -35037 10175 -34686
rect 10113 -35089 10175 -35037
rect 10147 -35437 10175 -35089
rect 10113 -35461 10175 -35437
rect 11040 -34687 11102 -34662
rect 11074 -35038 11102 -34687
rect 11040 -35090 11102 -35038
rect 11074 -35438 11102 -35090
rect 11040 -35462 11102 -35438
rect 12157 -34975 12407 -34958
rect 12157 -35036 12183 -34975
rect 12382 -35036 12407 -34975
rect 12923 -34971 13123 -34969
rect 12923 -35005 12954 -34971
rect 13086 -35005 13123 -34971
rect 12923 -35012 13123 -35005
rect 12157 -35054 12407 -35036
rect 12777 -35746 12820 -35715
rect 12777 -35878 12784 -35746
rect 12818 -35878 12820 -35746
rect 12777 -35915 12820 -35878
rect 12777 -36125 12820 -36094
rect 12777 -36257 12784 -36125
rect 12818 -36257 12820 -36125
rect 12777 -36294 12820 -36257
<< nsubdiff >>
rect 1795 6241 3005 6269
rect 1795 6169 1841 6241
rect 2963 6169 3005 6241
rect 1795 6143 3005 6169
rect 3401 6241 4611 6269
rect 3401 6169 3447 6241
rect 4569 6169 4611 6241
rect 3401 6143 4611 6169
rect 5105 6239 6315 6267
rect 5105 6167 5151 6239
rect 6273 6167 6315 6239
rect 5105 6141 6315 6167
rect 6943 5554 7560 5561
rect 6943 5507 6967 5554
rect 7536 5507 7560 5554
rect 6943 5495 7560 5507
rect 7809 5531 8023 5537
rect 7809 5497 7872 5531
rect 7963 5497 8023 5531
rect 7809 5471 8023 5497
rect -24042 4517 -22832 4545
rect -24042 4445 -24000 4517
rect -22878 4445 -22832 4517
rect -24042 4419 -22832 4445
rect -20751 4517 -19541 4545
rect -20751 4445 -20709 4517
rect -19587 4445 -19541 4517
rect -20751 4419 -19541 4445
rect -17460 4517 -16250 4545
rect -17460 4445 -17418 4517
rect -16296 4445 -16250 4517
rect -17460 4419 -16250 4445
rect -14169 4517 -12959 4545
rect -14169 4445 -14127 4517
rect -13005 4445 -12959 4517
rect -14169 4419 -12959 4445
rect -10878 4517 -9668 4545
rect -10878 4445 -10836 4517
rect -9714 4445 -9668 4517
rect -10878 4419 -9668 4445
rect -7588 4517 -6378 4545
rect -7588 4445 -7546 4517
rect -6424 4445 -6378 4517
rect -7588 4419 -6378 4445
rect -4297 4517 -3087 4545
rect -4297 4445 -4255 4517
rect -3133 4445 -3087 4517
rect -4297 4419 -3087 4445
rect -1006 4517 204 4545
rect -1006 4445 -964 4517
rect 158 4445 204 4517
rect -1006 4419 204 4445
rect 5658 3983 5872 3989
rect 5658 3949 5721 3983
rect 5812 3949 5872 3983
rect 5658 3923 5872 3949
rect 6098 3983 6312 3989
rect 6098 3949 6161 3983
rect 6252 3949 6312 3983
rect 6098 3923 6312 3949
rect 6538 3983 6752 3989
rect 6538 3949 6601 3983
rect 6692 3949 6752 3983
rect 6538 3923 6752 3949
rect 7138 3311 7964 3327
rect 7138 3276 7389 3311
rect 7677 3290 7964 3311
rect 8086 3311 8912 3327
rect 7677 3276 7963 3290
rect 7138 3273 7963 3276
rect 8086 3276 8337 3311
rect 8625 3290 8912 3311
rect 9022 3311 9848 3327
rect 8625 3276 8911 3290
rect 8086 3273 8911 3276
rect 9022 3276 9273 3311
rect 9561 3290 9848 3311
rect 9953 3311 10779 3327
rect 9561 3276 9847 3290
rect 9022 3273 9847 3276
rect 9953 3276 10204 3311
rect 10492 3290 10779 3311
rect 10880 3311 11706 3327
rect 10492 3276 10778 3290
rect 9953 3273 10778 3276
rect 10880 3276 11131 3311
rect 11419 3290 11706 3311
rect 11419 3276 11705 3290
rect 10880 3273 11705 3276
rect -24716 2733 -23506 2761
rect -24716 2661 -24670 2733
rect -23548 2661 -23506 2733
rect -24716 2635 -23506 2661
rect -23157 2733 -21947 2761
rect -23157 2661 -23111 2733
rect -21989 2661 -21947 2733
rect -23157 2635 -21947 2661
rect -21425 2733 -20215 2761
rect -21425 2661 -21379 2733
rect -20257 2661 -20215 2733
rect -21425 2635 -20215 2661
rect -19866 2733 -18656 2761
rect -19866 2661 -19820 2733
rect -18698 2661 -18656 2733
rect -19866 2635 -18656 2661
rect -18134 2733 -16924 2761
rect -18134 2661 -18088 2733
rect -16966 2661 -16924 2733
rect -18134 2635 -16924 2661
rect -16575 2733 -15365 2761
rect -16575 2661 -16529 2733
rect -15407 2661 -15365 2733
rect -16575 2635 -15365 2661
rect -14843 2733 -13633 2761
rect -14843 2661 -14797 2733
rect -13675 2661 -13633 2733
rect -14843 2635 -13633 2661
rect -13284 2733 -12074 2761
rect -13284 2661 -13238 2733
rect -12116 2661 -12074 2733
rect -13284 2635 -12074 2661
rect -11552 2733 -10342 2761
rect -11552 2661 -11506 2733
rect -10384 2661 -10342 2733
rect -11552 2635 -10342 2661
rect -9993 2733 -8783 2761
rect -9993 2661 -9947 2733
rect -8825 2661 -8783 2733
rect -9993 2635 -8783 2661
rect -8262 2733 -7052 2761
rect -8262 2661 -8216 2733
rect -7094 2661 -7052 2733
rect -8262 2635 -7052 2661
rect -6703 2733 -5493 2761
rect -6703 2661 -6657 2733
rect -5535 2661 -5493 2733
rect -6703 2635 -5493 2661
rect -4971 2733 -3761 2761
rect -4971 2661 -4925 2733
rect -3803 2661 -3761 2733
rect -4971 2635 -3761 2661
rect -3412 2733 -2202 2761
rect -3412 2661 -3366 2733
rect -2244 2661 -2202 2733
rect -3412 2635 -2202 2661
rect -1680 2733 -470 2761
rect -1680 2661 -1634 2733
rect -512 2661 -470 2733
rect -1680 2635 -470 2661
rect -121 2733 1089 2761
rect -121 2661 -75 2733
rect 1047 2661 1089 2733
rect -121 2635 1089 2661
rect 11783 2152 12203 2194
rect 11783 2101 11811 2152
rect 12168 2101 12203 2152
rect 11783 2063 12203 2101
rect 12923 1965 13137 1971
rect 12923 1931 12986 1965
rect 13077 1931 13137 1965
rect 12923 1905 13137 1931
rect -24593 988 -23976 995
rect -24593 941 -24569 988
rect -24000 941 -23976 988
rect -24593 929 -23976 941
rect -23484 988 -22867 995
rect -23484 941 -23460 988
rect -22891 941 -22867 988
rect -23484 929 -22867 941
rect -22602 988 -21985 995
rect -22602 941 -22578 988
rect -22009 941 -21985 988
rect -22602 929 -21985 941
rect -21302 988 -20685 995
rect -21302 941 -21278 988
rect -20709 941 -20685 988
rect -21302 929 -20685 941
rect -20193 988 -19576 995
rect -20193 941 -20169 988
rect -19600 941 -19576 988
rect -20193 929 -19576 941
rect -19311 988 -18694 995
rect -19311 941 -19287 988
rect -18718 941 -18694 988
rect -19311 929 -18694 941
rect -18011 988 -17394 995
rect -18011 941 -17987 988
rect -17418 941 -17394 988
rect -18011 929 -17394 941
rect -16902 988 -16285 995
rect -16902 941 -16878 988
rect -16309 941 -16285 988
rect -16902 929 -16285 941
rect -16020 988 -15403 995
rect -16020 941 -15996 988
rect -15427 941 -15403 988
rect -16020 929 -15403 941
rect -14720 988 -14103 995
rect -14720 941 -14696 988
rect -14127 941 -14103 988
rect -14720 929 -14103 941
rect -13611 988 -12994 995
rect -13611 941 -13587 988
rect -13018 941 -12994 988
rect -13611 929 -12994 941
rect -12729 988 -12112 995
rect -12729 941 -12705 988
rect -12136 941 -12112 988
rect -12729 929 -12112 941
rect -11429 988 -10812 995
rect -11429 941 -11405 988
rect -10836 941 -10812 988
rect -11429 929 -10812 941
rect -10320 988 -9703 995
rect -10320 941 -10296 988
rect -9727 941 -9703 988
rect -10320 929 -9703 941
rect -9438 988 -8821 995
rect -9438 941 -9414 988
rect -8845 941 -8821 988
rect -9438 929 -8821 941
rect -8139 988 -7522 995
rect -8139 941 -8115 988
rect -7546 941 -7522 988
rect -8139 929 -7522 941
rect -7030 988 -6413 995
rect -7030 941 -7006 988
rect -6437 941 -6413 988
rect -7030 929 -6413 941
rect -6148 988 -5531 995
rect -6148 941 -6124 988
rect -5555 941 -5531 988
rect -6148 929 -5531 941
rect -4848 988 -4231 995
rect -4848 941 -4824 988
rect -4255 941 -4231 988
rect -4848 929 -4231 941
rect -3739 988 -3122 995
rect -3739 941 -3715 988
rect -3146 941 -3122 988
rect -3739 929 -3122 941
rect -2857 988 -2240 995
rect -2857 941 -2833 988
rect -2264 941 -2240 988
rect -2857 929 -2240 941
rect -1557 988 -940 995
rect -1557 941 -1533 988
rect -964 941 -940 988
rect -1557 929 -940 941
rect -448 988 169 995
rect -448 941 -424 988
rect 145 941 169 988
rect -448 929 169 941
rect 434 988 1051 995
rect 434 941 458 988
rect 1027 941 1051 988
rect 434 929 1051 941
rect 7138 -24 7963 -21
rect 7138 -59 7389 -24
rect 7677 -38 7963 -24
rect 8086 -24 8911 -21
rect 7677 -59 7964 -38
rect 7138 -75 7964 -59
rect 8086 -59 8337 -24
rect 8625 -38 8911 -24
rect 9022 -24 9847 -21
rect 8625 -59 8912 -38
rect 8086 -75 8912 -59
rect 9022 -59 9273 -24
rect 9561 -38 9847 -24
rect 9953 -23 10778 -20
rect 9561 -59 9848 -38
rect 9022 -75 9848 -59
rect 9953 -58 10204 -23
rect 10492 -37 10778 -23
rect 10880 -24 11705 -21
rect 10492 -58 10779 -37
rect 9953 -74 10779 -58
rect 10880 -59 11131 -24
rect 11419 -38 11705 -24
rect 11419 -59 11706 -38
rect 10880 -75 11706 -59
rect 5658 -545 5872 -539
rect 5658 -579 5721 -545
rect 5812 -579 5872 -545
rect 5658 -605 5872 -579
rect 6098 -545 6312 -539
rect 6098 -579 6161 -545
rect 6252 -579 6312 -545
rect 6098 -605 6312 -579
rect 6538 -545 6752 -539
rect 6538 -579 6601 -545
rect 6692 -579 6752 -545
rect 6538 -605 6752 -579
rect 7138 -1217 7964 -1201
rect 7138 -1252 7389 -1217
rect 7677 -1238 7964 -1217
rect 8086 -1217 8912 -1201
rect 7677 -1252 7963 -1238
rect 7138 -1255 7963 -1252
rect 8086 -1252 8337 -1217
rect 8625 -1238 8912 -1217
rect 9022 -1217 9848 -1201
rect 8625 -1252 8911 -1238
rect 8086 -1255 8911 -1252
rect 9022 -1252 9273 -1217
rect 9561 -1238 9848 -1217
rect 9953 -1217 10779 -1201
rect 9561 -1252 9847 -1238
rect 9022 -1255 9847 -1252
rect 9953 -1252 10204 -1217
rect 10492 -1238 10779 -1217
rect 10880 -1217 11706 -1201
rect 10492 -1252 10778 -1238
rect 9953 -1255 10778 -1252
rect 10880 -1252 11131 -1217
rect 11419 -1238 11706 -1217
rect 11419 -1252 11705 -1238
rect 10880 -1255 11705 -1252
rect -23628 -2247 -23414 -2241
rect -23628 -2281 -23565 -2247
rect -23474 -2281 -23414 -2247
rect -24443 -2300 -23826 -2293
rect -24443 -2347 -24419 -2300
rect -23850 -2347 -23826 -2300
rect -24443 -2359 -23826 -2347
rect -23628 -2307 -23414 -2281
rect -21608 -2247 -21394 -2241
rect -21608 -2281 -21545 -2247
rect -21454 -2281 -21394 -2247
rect -22406 -2300 -21789 -2293
rect -22406 -2347 -22382 -2300
rect -21813 -2347 -21789 -2300
rect -22406 -2359 -21789 -2347
rect -21608 -2307 -21394 -2281
rect -19867 -2247 -19653 -2241
rect -19867 -2281 -19804 -2247
rect -19713 -2281 -19653 -2247
rect -20676 -2300 -20059 -2293
rect -20676 -2347 -20652 -2300
rect -20083 -2347 -20059 -2300
rect -20676 -2359 -20059 -2347
rect -19867 -2307 -19653 -2281
rect -18088 -2247 -17874 -2241
rect -18088 -2281 -18025 -2247
rect -17934 -2281 -17874 -2247
rect -18916 -2300 -18299 -2293
rect -18916 -2347 -18892 -2300
rect -18323 -2347 -18299 -2300
rect -18916 -2359 -18299 -2347
rect -18088 -2307 -17874 -2281
rect 11783 -2376 12203 -2334
rect 11783 -2427 11811 -2376
rect 12168 -2427 12203 -2376
rect 11783 -2465 12203 -2427
rect 12923 -2563 13137 -2557
rect 12923 -2597 12986 -2563
rect 13077 -2597 13137 -2563
rect 12923 -2623 13137 -2597
rect -20649 -3827 -19439 -3799
rect -20649 -3899 -20603 -3827
rect -19481 -3899 -19439 -3827
rect -20649 -3925 -19439 -3899
rect -19090 -3827 -17880 -3799
rect -19090 -3899 -19044 -3827
rect -17922 -3899 -17880 -3827
rect -19090 -3925 -17880 -3899
rect -17358 -3827 -16148 -3799
rect -17358 -3899 -17312 -3827
rect -16190 -3899 -16148 -3827
rect -17358 -3925 -16148 -3899
rect -15799 -3827 -14589 -3799
rect -15799 -3899 -15753 -3827
rect -14631 -3899 -14589 -3827
rect -15799 -3925 -14589 -3899
rect -14067 -3827 -12857 -3799
rect -14067 -3899 -14021 -3827
rect -12899 -3899 -12857 -3827
rect -14067 -3925 -12857 -3899
rect -12508 -3827 -11298 -3799
rect -12508 -3899 -12462 -3827
rect -11340 -3899 -11298 -3827
rect -12508 -3925 -11298 -3899
rect -10776 -3827 -9566 -3799
rect -10776 -3899 -10730 -3827
rect -9608 -3899 -9566 -3827
rect -10776 -3925 -9566 -3899
rect -9217 -3827 -8007 -3799
rect -9217 -3899 -9171 -3827
rect -8049 -3899 -8007 -3827
rect -9217 -3925 -8007 -3899
rect -23584 -4059 -23370 -4053
rect -23584 -4093 -23521 -4059
rect -23430 -4093 -23370 -4059
rect -24392 -4112 -23775 -4105
rect -24392 -4159 -24368 -4112
rect -23799 -4159 -23775 -4112
rect -24392 -4171 -23775 -4159
rect -23584 -4119 -23370 -4093
rect -21846 -4059 -21632 -4053
rect -21846 -4093 -21783 -4059
rect -21692 -4093 -21632 -4059
rect -22656 -4112 -22039 -4105
rect -22656 -4159 -22632 -4112
rect -22063 -4159 -22039 -4112
rect -22656 -4171 -22039 -4159
rect -21846 -4119 -21632 -4093
rect 7138 -4552 7963 -4549
rect 7138 -4587 7389 -4552
rect 7677 -4566 7963 -4552
rect 8086 -4552 8911 -4549
rect 7677 -4587 7964 -4566
rect 7138 -4603 7964 -4587
rect 8086 -4587 8337 -4552
rect 8625 -4566 8911 -4552
rect 9022 -4552 9847 -4549
rect 8625 -4587 8912 -4566
rect 8086 -4603 8912 -4587
rect 9022 -4587 9273 -4552
rect 9561 -4566 9847 -4552
rect 9953 -4551 10778 -4548
rect 9561 -4587 9848 -4566
rect 9022 -4603 9848 -4587
rect 9953 -4586 10204 -4551
rect 10492 -4565 10778 -4551
rect 10880 -4552 11705 -4549
rect 10492 -4586 10779 -4565
rect 9953 -4602 10779 -4586
rect 10880 -4587 11131 -4552
rect 11419 -4566 11705 -4552
rect 11419 -4587 11706 -4566
rect 10880 -4603 11706 -4587
rect 5658 -4973 5872 -4967
rect 5658 -5007 5721 -4973
rect 5812 -5007 5872 -4973
rect 5658 -5033 5872 -5007
rect 6098 -4973 6312 -4967
rect 6098 -5007 6161 -4973
rect 6252 -5007 6312 -4973
rect 6098 -5033 6312 -5007
rect -23586 -5351 -23372 -5345
rect -23586 -5385 -23523 -5351
rect -23432 -5385 -23372 -5351
rect -24392 -5404 -23775 -5397
rect -24392 -5451 -24368 -5404
rect -23799 -5451 -23775 -5404
rect -24392 -5463 -23775 -5451
rect -23586 -5411 -23372 -5385
rect -21852 -5351 -21638 -5345
rect -21852 -5385 -21789 -5351
rect -21698 -5385 -21638 -5351
rect 6538 -4973 6752 -4967
rect 6538 -5007 6601 -4973
rect 6692 -5007 6752 -4973
rect 6538 -5033 6752 -5007
rect -22656 -5404 -22039 -5397
rect -22656 -5451 -22632 -5404
rect -22063 -5451 -22039 -5404
rect -22656 -5463 -22039 -5451
rect -21852 -5411 -21638 -5385
rect -20526 -5572 -19909 -5565
rect -20526 -5619 -20502 -5572
rect -19933 -5619 -19909 -5572
rect -20526 -5631 -19909 -5619
rect -19417 -5572 -18800 -5565
rect -19417 -5619 -19393 -5572
rect -18824 -5619 -18800 -5572
rect -19417 -5631 -18800 -5619
rect -18535 -5572 -17918 -5565
rect -18535 -5619 -18511 -5572
rect -17942 -5619 -17918 -5572
rect -18535 -5631 -17918 -5619
rect -17235 -5572 -16618 -5565
rect -17235 -5619 -17211 -5572
rect -16642 -5619 -16618 -5572
rect -17235 -5631 -16618 -5619
rect -16126 -5572 -15509 -5565
rect -16126 -5619 -16102 -5572
rect -15533 -5619 -15509 -5572
rect -16126 -5631 -15509 -5619
rect -15244 -5572 -14627 -5565
rect -15244 -5619 -15220 -5572
rect -14651 -5619 -14627 -5572
rect -15244 -5631 -14627 -5619
rect -13944 -5572 -13327 -5565
rect -13944 -5619 -13920 -5572
rect -13351 -5619 -13327 -5572
rect -13944 -5631 -13327 -5619
rect -12835 -5572 -12218 -5565
rect -12835 -5619 -12811 -5572
rect -12242 -5619 -12218 -5572
rect -12835 -5631 -12218 -5619
rect -11953 -5572 -11336 -5565
rect -11953 -5619 -11929 -5572
rect -11360 -5619 -11336 -5572
rect -11953 -5631 -11336 -5619
rect -10653 -5572 -10036 -5565
rect -10653 -5619 -10629 -5572
rect -10060 -5619 -10036 -5572
rect -10653 -5631 -10036 -5619
rect -9544 -5572 -8927 -5565
rect -9544 -5619 -9520 -5572
rect -8951 -5619 -8927 -5572
rect -9544 -5631 -8927 -5619
rect -8662 -5572 -8045 -5565
rect -8662 -5619 -8638 -5572
rect -8069 -5619 -8045 -5572
rect -8662 -5631 -8045 -5619
rect 7138 -5645 7964 -5629
rect 7138 -5680 7389 -5645
rect 7677 -5666 7964 -5645
rect 8086 -5645 8912 -5629
rect 7677 -5680 7963 -5666
rect 7138 -5683 7963 -5680
rect 8086 -5680 8337 -5645
rect 8625 -5666 8912 -5645
rect 9022 -5645 9848 -5629
rect 8625 -5680 8911 -5666
rect 8086 -5683 8911 -5680
rect 9022 -5680 9273 -5645
rect 9561 -5666 9848 -5645
rect 9953 -5645 10779 -5629
rect 9561 -5680 9847 -5666
rect 9022 -5683 9847 -5680
rect 9953 -5680 10204 -5645
rect 10492 -5666 10779 -5645
rect 10880 -5645 11706 -5629
rect 10492 -5680 10778 -5666
rect 9953 -5683 10778 -5680
rect 10880 -5680 11131 -5645
rect 11419 -5666 11706 -5645
rect 11419 -5680 11705 -5666
rect 10880 -5683 11705 -5680
rect -20649 -7092 -19439 -7064
rect -20649 -7164 -20603 -7092
rect -19481 -7164 -19439 -7092
rect -20649 -7190 -19439 -7164
rect -19090 -7092 -17880 -7064
rect -19090 -7164 -19044 -7092
rect -17922 -7164 -17880 -7092
rect -19090 -7190 -17880 -7164
rect -17358 -7092 -16148 -7064
rect -17358 -7164 -17312 -7092
rect -16190 -7164 -16148 -7092
rect -17358 -7190 -16148 -7164
rect -15799 -7092 -14589 -7064
rect -15799 -7164 -15753 -7092
rect -14631 -7164 -14589 -7092
rect -15799 -7190 -14589 -7164
rect -14067 -7092 -12857 -7064
rect -14067 -7164 -14021 -7092
rect -12899 -7164 -12857 -7092
rect -14067 -7190 -12857 -7164
rect -12508 -7092 -11298 -7064
rect -12508 -7164 -12462 -7092
rect -11340 -7164 -11298 -7092
rect -12508 -7190 -11298 -7164
rect -10776 -7092 -9566 -7064
rect -10776 -7164 -10730 -7092
rect -9608 -7164 -9566 -7092
rect -10776 -7190 -9566 -7164
rect -9217 -7092 -8007 -7064
rect -9217 -7164 -9171 -7092
rect -8049 -7164 -8007 -7092
rect -9217 -7190 -8007 -7164
rect -23584 -7324 -23370 -7318
rect -23584 -7358 -23521 -7324
rect -23430 -7358 -23370 -7324
rect -24392 -7377 -23775 -7370
rect -24392 -7424 -24368 -7377
rect -23799 -7424 -23775 -7377
rect -24392 -7436 -23775 -7424
rect -23584 -7384 -23370 -7358
rect -21850 -7324 -21636 -7318
rect -21850 -7358 -21787 -7324
rect -21696 -7358 -21636 -7324
rect -22655 -7377 -22038 -7370
rect -22655 -7424 -22631 -7377
rect -22062 -7424 -22038 -7377
rect -22655 -7436 -22038 -7424
rect -21850 -7384 -21636 -7358
rect 11783 -6804 12203 -6762
rect 11783 -6855 11811 -6804
rect 12168 -6855 12203 -6804
rect 11783 -6893 12203 -6855
rect 12923 -6991 13137 -6985
rect 12923 -7025 12986 -6991
rect 13077 -7025 13137 -6991
rect 12923 -7051 13137 -7025
rect -23583 -8616 -23369 -8610
rect -23583 -8650 -23520 -8616
rect -23429 -8650 -23369 -8616
rect -24392 -8669 -23775 -8662
rect -24392 -8716 -24368 -8669
rect -23799 -8716 -23775 -8669
rect -24392 -8728 -23775 -8716
rect -23583 -8676 -23369 -8650
rect -21846 -8616 -21632 -8610
rect -21846 -8650 -21783 -8616
rect -21692 -8650 -21632 -8616
rect -22656 -8669 -22039 -8662
rect -22656 -8716 -22632 -8669
rect -22063 -8716 -22039 -8669
rect -22656 -8728 -22039 -8716
rect -21846 -8676 -21632 -8650
rect -20526 -8837 -19909 -8830
rect -20526 -8884 -20502 -8837
rect -19933 -8884 -19909 -8837
rect -20526 -8896 -19909 -8884
rect -19417 -8837 -18800 -8830
rect -19417 -8884 -19393 -8837
rect -18824 -8884 -18800 -8837
rect -19417 -8896 -18800 -8884
rect -18535 -8837 -17918 -8830
rect -18535 -8884 -18511 -8837
rect -17942 -8884 -17918 -8837
rect -18535 -8896 -17918 -8884
rect -17235 -8837 -16618 -8830
rect -17235 -8884 -17211 -8837
rect -16642 -8884 -16618 -8837
rect -17235 -8896 -16618 -8884
rect -16126 -8837 -15509 -8830
rect -16126 -8884 -16102 -8837
rect -15533 -8884 -15509 -8837
rect -16126 -8896 -15509 -8884
rect -15244 -8837 -14627 -8830
rect -15244 -8884 -15220 -8837
rect -14651 -8884 -14627 -8837
rect -15244 -8896 -14627 -8884
rect -13944 -8837 -13327 -8830
rect -13944 -8884 -13920 -8837
rect -13351 -8884 -13327 -8837
rect -13944 -8896 -13327 -8884
rect -12835 -8837 -12218 -8830
rect -12835 -8884 -12811 -8837
rect -12242 -8884 -12218 -8837
rect -12835 -8896 -12218 -8884
rect -11953 -8837 -11336 -8830
rect -11953 -8884 -11929 -8837
rect -11360 -8884 -11336 -8837
rect -11953 -8896 -11336 -8884
rect -10653 -8837 -10036 -8830
rect -10653 -8884 -10629 -8837
rect -10060 -8884 -10036 -8837
rect -10653 -8896 -10036 -8884
rect -9544 -8837 -8927 -8830
rect -9544 -8884 -9520 -8837
rect -8951 -8884 -8927 -8837
rect -9544 -8896 -8927 -8884
rect -8662 -8837 -8045 -8830
rect -8662 -8884 -8638 -8837
rect -8069 -8884 -8045 -8837
rect -8662 -8896 -8045 -8884
rect 7138 -8980 7963 -8977
rect 7138 -9015 7389 -8980
rect 7677 -8994 7963 -8980
rect 8086 -8980 8911 -8977
rect 7677 -9015 7964 -8994
rect 7138 -9031 7964 -9015
rect 8086 -9015 8337 -8980
rect 8625 -8994 8911 -8980
rect 9022 -8980 9847 -8977
rect 8625 -9015 8912 -8994
rect 8086 -9031 8912 -9015
rect 9022 -9015 9273 -8980
rect 9561 -8994 9847 -8980
rect 9953 -8979 10778 -8976
rect 9561 -9015 9848 -8994
rect 9022 -9031 9848 -9015
rect 9953 -9014 10204 -8979
rect 10492 -8993 10778 -8979
rect 10880 -8980 11705 -8977
rect 10492 -9014 10779 -8993
rect 9953 -9030 10779 -9014
rect 10880 -9015 11131 -8980
rect 11419 -8994 11705 -8980
rect 11419 -9015 11706 -8994
rect 10880 -9031 11706 -9015
rect 5658 -9601 5872 -9595
rect 5658 -9635 5721 -9601
rect 5812 -9635 5872 -9601
rect 5658 -9661 5872 -9635
rect 6098 -9601 6312 -9595
rect 6098 -9635 6161 -9601
rect 6252 -9635 6312 -9601
rect 6098 -9661 6312 -9635
rect 6538 -9601 6752 -9595
rect 6538 -9635 6601 -9601
rect 6692 -9635 6752 -9601
rect 6538 -9661 6752 -9635
rect 7138 -10273 7964 -10257
rect 7138 -10308 7389 -10273
rect 7677 -10294 7964 -10273
rect 8086 -10273 8912 -10257
rect 7677 -10308 7963 -10294
rect 7138 -10311 7963 -10308
rect 8086 -10308 8337 -10273
rect 8625 -10294 8912 -10273
rect 9022 -10273 9848 -10257
rect 8625 -10308 8911 -10294
rect 8086 -10311 8911 -10308
rect 9022 -10308 9273 -10273
rect 9561 -10294 9848 -10273
rect 9953 -10273 10779 -10257
rect 9561 -10308 9847 -10294
rect 9022 -10311 9847 -10308
rect 9953 -10308 10204 -10273
rect 10492 -10294 10779 -10273
rect 10880 -10273 11706 -10257
rect 10492 -10308 10778 -10294
rect 9953 -10311 10778 -10308
rect 10880 -10308 11131 -10273
rect 11419 -10294 11706 -10273
rect 11419 -10308 11705 -10294
rect 10880 -10311 11705 -10308
rect -20649 -10356 -19439 -10328
rect -20649 -10428 -20603 -10356
rect -19481 -10428 -19439 -10356
rect -20649 -10454 -19439 -10428
rect -19090 -10356 -17880 -10328
rect -19090 -10428 -19044 -10356
rect -17922 -10428 -17880 -10356
rect -19090 -10454 -17880 -10428
rect -17358 -10356 -16148 -10328
rect -17358 -10428 -17312 -10356
rect -16190 -10428 -16148 -10356
rect -17358 -10454 -16148 -10428
rect -15799 -10356 -14589 -10328
rect -15799 -10428 -15753 -10356
rect -14631 -10428 -14589 -10356
rect -15799 -10454 -14589 -10428
rect -14067 -10356 -12857 -10328
rect -14067 -10428 -14021 -10356
rect -12899 -10428 -12857 -10356
rect -14067 -10454 -12857 -10428
rect -12508 -10356 -11298 -10328
rect -12508 -10428 -12462 -10356
rect -11340 -10428 -11298 -10356
rect -12508 -10454 -11298 -10428
rect -10776 -10356 -9566 -10328
rect -10776 -10428 -10730 -10356
rect -9608 -10428 -9566 -10356
rect -10776 -10454 -9566 -10428
rect -9217 -10356 -8007 -10328
rect -9217 -10428 -9171 -10356
rect -8049 -10428 -8007 -10356
rect -9217 -10454 -8007 -10428
rect -23583 -10588 -23369 -10582
rect -23583 -10622 -23520 -10588
rect -23429 -10622 -23369 -10588
rect -24392 -10641 -23775 -10634
rect -24392 -10688 -24368 -10641
rect -23799 -10688 -23775 -10641
rect -24392 -10700 -23775 -10688
rect -23583 -10648 -23369 -10622
rect -21850 -10588 -21636 -10582
rect -21850 -10622 -21787 -10588
rect -21696 -10622 -21636 -10588
rect -22655 -10641 -22038 -10634
rect -22655 -10688 -22631 -10641
rect -22062 -10688 -22038 -10641
rect -22655 -10700 -22038 -10688
rect -21850 -10648 -21636 -10622
rect -23583 -11880 -23369 -11874
rect -23583 -11914 -23520 -11880
rect -23429 -11914 -23369 -11880
rect -24392 -11933 -23775 -11926
rect -24392 -11980 -24368 -11933
rect -23799 -11980 -23775 -11933
rect -24392 -11992 -23775 -11980
rect -23583 -11940 -23369 -11914
rect -21854 -11880 -21640 -11874
rect -21854 -11914 -21791 -11880
rect -21700 -11914 -21640 -11880
rect 11783 -11432 12203 -11390
rect 11783 -11483 11811 -11432
rect 12168 -11483 12203 -11432
rect 11783 -11521 12203 -11483
rect 12923 -11619 13137 -11613
rect 12923 -11653 12986 -11619
rect 13077 -11653 13137 -11619
rect 12923 -11679 13137 -11653
rect -22655 -11933 -22038 -11926
rect -22655 -11980 -22631 -11933
rect -22062 -11980 -22038 -11933
rect -22655 -11992 -22038 -11980
rect -21854 -11940 -21640 -11914
rect -20526 -12101 -19909 -12094
rect -20526 -12148 -20502 -12101
rect -19933 -12148 -19909 -12101
rect -20526 -12160 -19909 -12148
rect -19417 -12101 -18800 -12094
rect -19417 -12148 -19393 -12101
rect -18824 -12148 -18800 -12101
rect -19417 -12160 -18800 -12148
rect -18535 -12101 -17918 -12094
rect -18535 -12148 -18511 -12101
rect -17942 -12148 -17918 -12101
rect -18535 -12160 -17918 -12148
rect -17235 -12101 -16618 -12094
rect -17235 -12148 -17211 -12101
rect -16642 -12148 -16618 -12101
rect -17235 -12160 -16618 -12148
rect -16126 -12101 -15509 -12094
rect -16126 -12148 -16102 -12101
rect -15533 -12148 -15509 -12101
rect -16126 -12160 -15509 -12148
rect -15244 -12101 -14627 -12094
rect -15244 -12148 -15220 -12101
rect -14651 -12148 -14627 -12101
rect -15244 -12160 -14627 -12148
rect -13944 -12101 -13327 -12094
rect -13944 -12148 -13920 -12101
rect -13351 -12148 -13327 -12101
rect -13944 -12160 -13327 -12148
rect -12835 -12101 -12218 -12094
rect -12835 -12148 -12811 -12101
rect -12242 -12148 -12218 -12101
rect -12835 -12160 -12218 -12148
rect -11953 -12101 -11336 -12094
rect -11953 -12148 -11929 -12101
rect -11360 -12148 -11336 -12101
rect -11953 -12160 -11336 -12148
rect -10653 -12101 -10036 -12094
rect -10653 -12148 -10629 -12101
rect -10060 -12148 -10036 -12101
rect -10653 -12160 -10036 -12148
rect -9544 -12101 -8927 -12094
rect -9544 -12148 -9520 -12101
rect -8951 -12148 -8927 -12101
rect -9544 -12160 -8927 -12148
rect -8662 -12101 -8045 -12094
rect -8662 -12148 -8638 -12101
rect -8069 -12148 -8045 -12101
rect -8662 -12160 -8045 -12148
rect 7138 -13608 7963 -13605
rect 7138 -13643 7389 -13608
rect 7677 -13622 7963 -13608
rect 8086 -13608 8911 -13605
rect 7677 -13643 7964 -13622
rect 7138 -13659 7964 -13643
rect 8086 -13643 8337 -13608
rect 8625 -13622 8911 -13608
rect 9022 -13608 9847 -13605
rect 8625 -13643 8912 -13622
rect 8086 -13659 8912 -13643
rect 9022 -13643 9273 -13608
rect 9561 -13622 9847 -13608
rect 9953 -13607 10778 -13604
rect 9561 -13643 9848 -13622
rect 9022 -13659 9848 -13643
rect 9953 -13642 10204 -13607
rect 10492 -13621 10778 -13607
rect 10880 -13608 11705 -13605
rect 10492 -13642 10779 -13621
rect 9953 -13658 10779 -13642
rect 10880 -13643 11131 -13608
rect 11419 -13622 11705 -13608
rect 11419 -13643 11706 -13622
rect 10880 -13659 11706 -13643
rect -2178 -13878 -2112 -13818
rect -2178 -13969 -2172 -13878
rect -2138 -13969 -2112 -13878
rect -2178 -14032 -2112 -13969
rect 5658 -14129 5872 -14123
rect -12501 -14223 -12375 -14181
rect -24569 -14953 -24503 -14929
rect -24569 -15522 -24562 -14953
rect -24515 -15522 -24503 -14953
rect -17862 -15122 -17731 -15087
rect -24569 -15546 -24503 -15522
rect -17862 -15479 -17820 -15122
rect -17769 -15479 -17731 -15122
rect -12501 -15345 -12473 -14223
rect -12401 -15345 -12375 -14223
rect 5658 -14163 5721 -14129
rect 5812 -14163 5872 -14129
rect -12501 -15391 -12375 -15345
rect -4894 -14266 -4828 -14203
rect -4894 -14357 -4888 -14266
rect -4854 -14357 -4828 -14266
rect -4894 -14417 -4828 -14357
rect -2178 -14257 -2112 -14197
rect -2178 -14348 -2172 -14257
rect -2138 -14348 -2112 -14257
rect -2178 -14411 -2112 -14348
rect 5658 -14189 5872 -14163
rect 6098 -14129 6312 -14123
rect 6098 -14163 6161 -14129
rect 6252 -14163 6312 -14129
rect 6098 -14189 6312 -14163
rect 6538 -14129 6752 -14123
rect 6538 -14163 6601 -14129
rect 6692 -14163 6752 -14129
rect 6538 -14189 6752 -14163
rect -4894 -14706 -4828 -14643
rect -4894 -14797 -4888 -14706
rect -4854 -14797 -4828 -14706
rect -4894 -14857 -4828 -14797
rect -2178 -14697 -2112 -14637
rect -2178 -14788 -2172 -14697
rect -2138 -14788 -2112 -14697
rect -2178 -14851 -2112 -14788
rect 7138 -14801 7964 -14785
rect 7138 -14836 7389 -14801
rect 7677 -14822 7964 -14801
rect 8086 -14801 8912 -14785
rect 7677 -14836 7963 -14822
rect 7138 -14839 7963 -14836
rect 8086 -14836 8337 -14801
rect 8625 -14822 8912 -14801
rect 9022 -14801 9848 -14785
rect 8625 -14836 8911 -14822
rect 8086 -14839 8911 -14836
rect 9022 -14836 9273 -14801
rect 9561 -14822 9848 -14801
rect 9953 -14801 10779 -14785
rect 9561 -14836 9847 -14822
rect 9022 -14839 9847 -14836
rect 9953 -14836 10204 -14801
rect 10492 -14822 10779 -14801
rect 10880 -14801 11706 -14785
rect 10492 -14836 10778 -14822
rect 9953 -14839 10778 -14836
rect 10880 -14836 11131 -14801
rect 11419 -14822 11706 -14801
rect 11419 -14836 11705 -14822
rect 10880 -14839 11705 -14836
rect -4894 -15085 -4828 -15022
rect -4894 -15176 -4888 -15085
rect -4854 -15176 -4828 -15085
rect -4894 -15236 -4828 -15176
rect -2178 -15076 -2112 -15016
rect -2178 -15167 -2172 -15076
rect -2138 -15167 -2112 -15076
rect -2178 -15230 -2112 -15167
rect -8245 -15406 -8179 -15346
rect -17862 -15507 -17731 -15479
rect -8245 -15497 -8239 -15406
rect -8205 -15497 -8179 -15406
rect -8245 -15560 -8179 -15497
rect -4894 -15525 -4828 -15462
rect -4894 -15616 -4888 -15525
rect -4854 -15616 -4828 -15525
rect -4894 -15676 -4828 -15616
rect -2178 -15516 -2112 -15456
rect -2178 -15607 -2172 -15516
rect -2138 -15607 -2112 -15516
rect -2178 -15670 -2112 -15607
rect -8244 -15906 -8178 -15846
rect -8244 -15997 -8238 -15906
rect -8204 -15997 -8178 -15906
rect -8244 -16060 -8178 -15997
rect -4894 -15904 -4828 -15841
rect -4894 -15995 -4888 -15904
rect -4854 -15995 -4828 -15904
rect -4894 -16055 -4828 -15995
rect -2178 -15895 -2112 -15835
rect -2178 -15986 -2172 -15895
rect -2138 -15986 -2112 -15895
rect -24568 -16138 -24502 -16114
rect -24568 -16707 -24561 -16138
rect -24514 -16707 -24502 -16138
rect -2178 -16049 -2112 -15986
rect -17862 -16522 -17731 -16487
rect -24568 -16731 -24502 -16707
rect -17862 -16879 -17820 -16522
rect -17769 -16879 -17731 -16522
rect -8245 -16386 -8179 -16326
rect -8245 -16477 -8239 -16386
rect -8205 -16477 -8179 -16386
rect -8245 -16540 -8179 -16477
rect -4894 -16344 -4828 -16281
rect -4894 -16435 -4888 -16344
rect -4854 -16435 -4828 -16344
rect -4894 -16495 -4828 -16435
rect -2178 -16335 -2112 -16275
rect -2178 -16426 -2172 -16335
rect -2138 -16426 -2112 -16335
rect -2178 -16489 -2112 -16426
rect 11783 -15960 12203 -15918
rect 11783 -16011 11811 -15960
rect 12168 -16011 12203 -15960
rect 11783 -16049 12203 -16011
rect 12923 -16147 13137 -16141
rect 12923 -16181 12986 -16147
rect 13077 -16181 13137 -16147
rect 12923 -16207 13137 -16181
rect -4894 -16723 -4828 -16660
rect -4894 -16814 -4888 -16723
rect -4854 -16814 -4828 -16723
rect -17862 -16907 -17731 -16879
rect -8245 -16886 -8179 -16826
rect -8245 -16977 -8239 -16886
rect -8205 -16977 -8179 -16886
rect -12499 -17039 -12373 -16997
rect -24563 -17351 -24497 -17327
rect -24563 -17920 -24556 -17351
rect -24509 -17920 -24497 -17351
rect -24563 -17944 -24497 -17920
rect -17862 -17922 -17731 -17887
rect -21684 -18094 -21618 -18034
rect -21684 -18185 -21678 -18094
rect -21644 -18185 -21618 -18094
rect -21684 -18248 -21618 -18185
rect -17862 -18279 -17820 -17922
rect -17769 -18279 -17731 -17922
rect -16093 -17965 -16027 -17905
rect -16093 -18056 -16087 -17965
rect -16053 -18056 -16027 -17965
rect -16093 -18119 -16027 -18056
rect -12499 -18161 -12471 -17039
rect -12399 -18161 -12373 -17039
rect -12499 -18207 -12373 -18161
rect -8245 -17040 -8179 -16977
rect -4894 -16874 -4828 -16814
rect -2178 -16714 -2112 -16654
rect -2178 -16805 -2172 -16714
rect -2138 -16805 -2112 -16714
rect -2178 -16868 -2112 -16805
rect -4894 -17163 -4828 -17100
rect -4894 -17254 -4888 -17163
rect -4854 -17254 -4828 -17163
rect -8245 -17366 -8179 -17306
rect -8245 -17457 -8239 -17366
rect -8205 -17457 -8179 -17366
rect -8245 -17520 -8179 -17457
rect -4894 -17314 -4828 -17254
rect -2178 -17154 -2112 -17094
rect -2178 -17245 -2172 -17154
rect -2138 -17245 -2112 -17154
rect -2178 -17308 -2112 -17245
rect -4894 -17542 -4828 -17479
rect -4894 -17633 -4888 -17542
rect -4854 -17633 -4828 -17542
rect -4894 -17693 -4828 -17633
rect -2178 -17533 -2112 -17473
rect -2178 -17624 -2172 -17533
rect -2138 -17624 -2112 -17533
rect -2178 -17687 -2112 -17624
rect -8245 -17826 -8179 -17766
rect -8245 -17917 -8239 -17826
rect -8205 -17917 -8179 -17826
rect -8245 -17980 -8179 -17917
rect -4894 -17982 -4828 -17919
rect -4894 -18073 -4888 -17982
rect -4854 -18073 -4828 -17982
rect -4894 -18133 -4828 -18073
rect -2178 -17973 -2112 -17913
rect -2178 -18064 -2172 -17973
rect -2138 -18064 -2112 -17973
rect -2178 -18127 -2112 -18064
rect 15653 -17679 15763 -17667
rect 15653 -18033 15703 -17679
rect 15737 -18033 15763 -17679
rect 7138 -18136 7963 -18133
rect -17862 -18307 -17731 -18279
rect -8259 -18286 -8193 -18226
rect -24548 -18470 -24482 -18446
rect -24548 -19039 -24541 -18470
rect -24494 -19039 -24482 -18470
rect -16092 -18465 -16026 -18405
rect -21683 -18594 -21617 -18534
rect -21683 -18685 -21677 -18594
rect -21643 -18685 -21617 -18594
rect -21683 -18748 -21617 -18685
rect -16092 -18556 -16086 -18465
rect -16052 -18556 -16026 -18465
rect -16092 -18619 -16026 -18556
rect -8259 -18377 -8253 -18286
rect -8219 -18377 -8193 -18286
rect -8259 -18440 -8193 -18377
rect 7138 -18171 7389 -18136
rect 7677 -18150 7963 -18136
rect 8086 -18136 8911 -18133
rect 7677 -18171 7964 -18150
rect 7138 -18187 7964 -18171
rect 8086 -18171 8337 -18136
rect 8625 -18150 8911 -18136
rect 9022 -18136 9847 -18133
rect 8625 -18171 8912 -18150
rect 8086 -18187 8912 -18171
rect 9022 -18171 9273 -18136
rect 9561 -18150 9847 -18136
rect 9953 -18135 10778 -18132
rect 9561 -18171 9848 -18150
rect 9022 -18187 9848 -18171
rect 9953 -18170 10204 -18135
rect 10492 -18149 10778 -18135
rect 10880 -18136 11705 -18133
rect 10492 -18170 10779 -18149
rect 9953 -18186 10779 -18170
rect 10880 -18171 11131 -18136
rect 11419 -18150 11705 -18136
rect 11419 -18171 11706 -18150
rect 10880 -18187 11706 -18171
rect -4894 -18361 -4828 -18298
rect -4894 -18452 -4888 -18361
rect -4854 -18452 -4828 -18361
rect -4894 -18512 -4828 -18452
rect -2178 -18352 -2112 -18292
rect -2178 -18443 -2172 -18352
rect -2138 -18443 -2112 -18352
rect -2178 -18506 -2112 -18443
rect 15653 -18523 15763 -18033
rect 17298 -18162 17915 -18155
rect 17298 -18209 17322 -18162
rect 17891 -18209 17915 -18162
rect 17298 -18221 17915 -18209
rect 18096 -18187 18310 -18181
rect 18096 -18221 18159 -18187
rect 18250 -18221 18310 -18187
rect 18096 -18247 18310 -18221
rect -8257 -18766 -8191 -18706
rect -8257 -18857 -8251 -18766
rect -8217 -18857 -8191 -18766
rect -24548 -19063 -24482 -19039
rect -21684 -19074 -21618 -19014
rect -21684 -19165 -21678 -19074
rect -21644 -19165 -21618 -19074
rect -21684 -19228 -21618 -19165
rect -16093 -18945 -16027 -18885
rect -16093 -19036 -16087 -18945
rect -16053 -19036 -16027 -18945
rect -16093 -19099 -16027 -19036
rect -8257 -18920 -8191 -18857
rect 15653 -18649 15738 -18523
rect 5658 -18657 5872 -18651
rect 5658 -18691 5721 -18657
rect 5812 -18691 5872 -18657
rect 5658 -18717 5872 -18691
rect -4894 -18801 -4828 -18738
rect -4894 -18892 -4888 -18801
rect -4854 -18892 -4828 -18801
rect -4894 -18952 -4828 -18892
rect -2178 -18792 -2112 -18732
rect -2178 -18883 -2172 -18792
rect -2138 -18883 -2112 -18792
rect -2178 -18946 -2112 -18883
rect 6098 -18657 6312 -18651
rect 6098 -18691 6161 -18657
rect 6252 -18691 6312 -18657
rect 6098 -18717 6312 -18691
rect 6538 -18657 6752 -18651
rect 6538 -18691 6601 -18657
rect 6692 -18691 6752 -18657
rect 6538 -18717 6752 -18691
rect -17862 -19322 -17731 -19287
rect -21684 -19574 -21618 -19514
rect -24546 -19664 -24480 -19640
rect -24546 -20233 -24539 -19664
rect -24492 -20233 -24480 -19664
rect -21684 -19665 -21678 -19574
rect -21644 -19665 -21618 -19574
rect -21684 -19728 -21618 -19665
rect -17862 -19679 -17820 -19322
rect -17769 -19679 -17731 -19322
rect -4894 -19180 -4828 -19117
rect -4894 -19271 -4888 -19180
rect -4854 -19271 -4828 -19180
rect -4894 -19331 -4828 -19271
rect -2178 -19171 -2112 -19111
rect -2178 -19262 -2172 -19171
rect -2138 -19262 -2112 -19171
rect -2178 -19325 -2112 -19262
rect 15653 -19139 15763 -18649
rect 7138 -19329 7964 -19313
rect -16093 -19445 -16027 -19385
rect -16093 -19536 -16087 -19445
rect -16053 -19536 -16027 -19445
rect -16093 -19599 -16027 -19536
rect 7138 -19364 7389 -19329
rect 7677 -19350 7964 -19329
rect 8086 -19329 8912 -19313
rect 7677 -19364 7963 -19350
rect 7138 -19367 7963 -19364
rect 8086 -19364 8337 -19329
rect 8625 -19350 8912 -19329
rect 9022 -19329 9848 -19313
rect 8625 -19364 8911 -19350
rect 8086 -19367 8911 -19364
rect 9022 -19364 9273 -19329
rect 9561 -19350 9848 -19329
rect 9953 -19329 10779 -19313
rect 9561 -19364 9847 -19350
rect 9022 -19367 9847 -19364
rect 9953 -19364 10204 -19329
rect 10492 -19350 10779 -19329
rect 10880 -19329 11706 -19313
rect 10492 -19364 10778 -19350
rect 9953 -19367 10778 -19364
rect 10880 -19364 11131 -19329
rect 11419 -19350 11706 -19329
rect 11419 -19364 11705 -19350
rect 10880 -19367 11705 -19364
rect -4894 -19620 -4828 -19557
rect -17862 -19707 -17731 -19679
rect -4894 -19711 -4888 -19620
rect -4854 -19711 -4828 -19620
rect -4894 -19771 -4828 -19711
rect -2178 -19611 -2112 -19551
rect -2178 -19702 -2172 -19611
rect -2138 -19702 -2112 -19611
rect -2178 -19765 -2112 -19702
rect 15653 -19493 15703 -19139
rect 15737 -19493 15763 -19139
rect 15653 -19505 15763 -19493
rect -16093 -19925 -16027 -19865
rect -24546 -20257 -24480 -20233
rect -21684 -20054 -21618 -19994
rect -21684 -20145 -21678 -20054
rect -21644 -20145 -21618 -20054
rect -21684 -20208 -21618 -20145
rect -16093 -20016 -16087 -19925
rect -16053 -20016 -16027 -19925
rect -16093 -20079 -16027 -20016
rect -12499 -19996 -12373 -19954
rect -21684 -20514 -21618 -20454
rect -21684 -20605 -21678 -20514
rect -21644 -20605 -21618 -20514
rect -21684 -20668 -21618 -20605
rect -16093 -20385 -16027 -20325
rect -16093 -20476 -16087 -20385
rect -16053 -20476 -16027 -20385
rect -17862 -20722 -17731 -20687
rect -24515 -20864 -24449 -20840
rect -24515 -21433 -24508 -20864
rect -24461 -21433 -24449 -20864
rect -21698 -20974 -21632 -20914
rect -21698 -21065 -21692 -20974
rect -21658 -21065 -21632 -20974
rect -21698 -21128 -21632 -21065
rect -17862 -21079 -17820 -20722
rect -17769 -21079 -17731 -20722
rect -16093 -20539 -16027 -20476
rect -16107 -20845 -16041 -20785
rect -16107 -20936 -16101 -20845
rect -16067 -20936 -16041 -20845
rect -16107 -20999 -16041 -20936
rect -17862 -21107 -17731 -21079
rect -12499 -21118 -12471 -19996
rect -12399 -21118 -12373 -19996
rect -12499 -21164 -12373 -21118
rect -4894 -19999 -4828 -19936
rect -4894 -20090 -4888 -19999
rect -4854 -20090 -4828 -19999
rect -4894 -20150 -4828 -20090
rect -2178 -19990 -2112 -19930
rect -2178 -20081 -2172 -19990
rect -2138 -20081 -2112 -19990
rect -2178 -20144 -2112 -20081
rect -4894 -20439 -4828 -20376
rect -4894 -20530 -4888 -20439
rect -4854 -20530 -4828 -20439
rect -4894 -20590 -4828 -20530
rect -2178 -20430 -2112 -20370
rect -2178 -20521 -2172 -20430
rect -2138 -20521 -2112 -20430
rect -2178 -20584 -2112 -20521
rect -4894 -20818 -4828 -20755
rect -4894 -20909 -4888 -20818
rect -4854 -20909 -4828 -20818
rect -4894 -20969 -4828 -20909
rect 11783 -20488 12203 -20446
rect 11783 -20539 11811 -20488
rect 12168 -20539 12203 -20488
rect 11783 -20577 12203 -20539
rect 12923 -20675 13137 -20669
rect 12923 -20709 12986 -20675
rect 13077 -20709 13137 -20675
rect 12923 -20735 13137 -20709
rect -16105 -21325 -16039 -21265
rect -24515 -21457 -24449 -21433
rect -21696 -21454 -21630 -21394
rect -21696 -21545 -21690 -21454
rect -21656 -21545 -21630 -21454
rect -21696 -21608 -21630 -21545
rect -16105 -21416 -16099 -21325
rect -16065 -21416 -16039 -21325
rect -16105 -21479 -16039 -21416
rect -17862 -22122 -17731 -22087
rect -24516 -22167 -24450 -22143
rect -24516 -22736 -24509 -22167
rect -24462 -22736 -24450 -22167
rect -17862 -22479 -17820 -22122
rect -17769 -22479 -17731 -22122
rect -17862 -22507 -17731 -22479
rect -24516 -22760 -24450 -22736
rect -12499 -22575 -12373 -22533
rect -24516 -23476 -24450 -23452
rect -24516 -24045 -24509 -23476
rect -24462 -24045 -24450 -23476
rect -17862 -23522 -17731 -23487
rect -17862 -23879 -17820 -23522
rect -17769 -23879 -17731 -23522
rect -12499 -23697 -12471 -22575
rect -12399 -23697 -12373 -22575
rect -12499 -23743 -12373 -23697
rect 7138 -22664 7963 -22661
rect 7138 -22699 7389 -22664
rect 7677 -22678 7963 -22664
rect 8086 -22664 8911 -22661
rect 7677 -22699 7964 -22678
rect 7138 -22715 7964 -22699
rect 8086 -22699 8337 -22664
rect 8625 -22678 8911 -22664
rect 9022 -22664 9847 -22661
rect 8625 -22699 8912 -22678
rect 8086 -22715 8912 -22699
rect 9022 -22699 9273 -22664
rect 9561 -22678 9847 -22664
rect 9953 -22663 10778 -22660
rect 9561 -22699 9848 -22678
rect 9022 -22715 9848 -22699
rect 9953 -22698 10204 -22663
rect 10492 -22677 10778 -22663
rect 10880 -22664 11705 -22661
rect 10492 -22698 10779 -22677
rect 9953 -22714 10779 -22698
rect 10880 -22699 11131 -22664
rect 11419 -22678 11705 -22664
rect 11419 -22699 11706 -22678
rect 10880 -22715 11706 -22699
rect 5658 -23185 5872 -23179
rect 5658 -23219 5721 -23185
rect 5812 -23219 5872 -23185
rect 5658 -23245 5872 -23219
rect 6098 -23185 6312 -23179
rect 6098 -23219 6161 -23185
rect 6252 -23219 6312 -23185
rect 6098 -23245 6312 -23219
rect 6538 -23185 6752 -23179
rect 6538 -23219 6601 -23185
rect 6692 -23219 6752 -23185
rect 6538 -23245 6752 -23219
rect -17862 -23907 -17731 -23879
rect 7138 -23857 7964 -23841
rect -24516 -24069 -24450 -24045
rect 7138 -23892 7389 -23857
rect 7677 -23878 7964 -23857
rect 8086 -23857 8912 -23841
rect 7677 -23892 7963 -23878
rect 7138 -23895 7963 -23892
rect 8086 -23892 8337 -23857
rect 8625 -23878 8912 -23857
rect 9022 -23857 9848 -23841
rect 8625 -23892 8911 -23878
rect 8086 -23895 8911 -23892
rect 9022 -23892 9273 -23857
rect 9561 -23878 9848 -23857
rect 9953 -23857 10779 -23841
rect 9561 -23892 9847 -23878
rect 9022 -23895 9847 -23892
rect 9953 -23892 10204 -23857
rect 10492 -23878 10779 -23857
rect 10880 -23857 11706 -23841
rect 10492 -23892 10778 -23878
rect 9953 -23895 10778 -23892
rect 10880 -23892 11131 -23857
rect 11419 -23878 11706 -23857
rect 11419 -23892 11705 -23878
rect 10880 -23895 11705 -23892
rect -17862 -24922 -17731 -24887
rect -17862 -25279 -17820 -24922
rect -17769 -25279 -17731 -24922
rect -17862 -25307 -17731 -25279
rect -12499 -25343 -12373 -25301
rect -12499 -26465 -12471 -25343
rect -12399 -26465 -12373 -25343
rect -12499 -26511 -12373 -26465
rect 11783 -25016 12203 -24974
rect 11783 -25067 11811 -25016
rect 12168 -25067 12203 -25016
rect 11783 -25105 12203 -25067
rect 12923 -25203 13137 -25197
rect 12923 -25237 12986 -25203
rect 13077 -25237 13137 -25203
rect 12923 -25263 13137 -25237
rect 7138 -27192 7963 -27189
rect 7138 -27227 7389 -27192
rect 7677 -27206 7963 -27192
rect 8086 -27192 8911 -27189
rect 7677 -27227 7964 -27206
rect 7138 -27243 7964 -27227
rect 8086 -27227 8337 -27192
rect 8625 -27206 8911 -27192
rect 9022 -27192 9847 -27189
rect 8625 -27227 8912 -27206
rect 8086 -27243 8912 -27227
rect 9022 -27227 9273 -27192
rect 9561 -27206 9847 -27192
rect 9953 -27191 10778 -27188
rect 9561 -27227 9848 -27206
rect 9022 -27243 9848 -27227
rect 9953 -27226 10204 -27191
rect 10492 -27205 10778 -27191
rect 10880 -27192 11705 -27189
rect 10492 -27226 10779 -27205
rect 9953 -27242 10779 -27226
rect 10880 -27227 11131 -27192
rect 11419 -27206 11705 -27192
rect 11419 -27227 11706 -27206
rect 10880 -27243 11706 -27227
rect 5658 -27713 5872 -27707
rect 5658 -27747 5721 -27713
rect 5812 -27747 5872 -27713
rect 5658 -27773 5872 -27747
rect -12499 -27976 -12373 -27934
rect -12499 -29098 -12471 -27976
rect -12399 -29098 -12373 -27976
rect -12499 -29144 -12373 -29098
rect 6098 -27713 6312 -27707
rect 6098 -27747 6161 -27713
rect 6252 -27747 6312 -27713
rect 6098 -27773 6312 -27747
rect 6538 -27713 6752 -27707
rect 6538 -27747 6601 -27713
rect 6692 -27747 6752 -27713
rect 6538 -27773 6752 -27747
rect 7138 -28385 7964 -28369
rect 7138 -28420 7389 -28385
rect 7677 -28406 7964 -28385
rect 8086 -28385 8912 -28369
rect 7677 -28420 7963 -28406
rect 7138 -28423 7963 -28420
rect 8086 -28420 8337 -28385
rect 8625 -28406 8912 -28385
rect 9022 -28385 9848 -28369
rect 8625 -28420 8911 -28406
rect 8086 -28423 8911 -28420
rect 9022 -28420 9273 -28385
rect 9561 -28406 9848 -28385
rect 9953 -28385 10779 -28369
rect 9561 -28420 9847 -28406
rect 9022 -28423 9847 -28420
rect 9953 -28420 10204 -28385
rect 10492 -28406 10779 -28385
rect 10880 -28385 11706 -28369
rect 10492 -28420 10778 -28406
rect 9953 -28423 10778 -28420
rect 10880 -28420 11131 -28385
rect 11419 -28406 11706 -28385
rect 11419 -28420 11705 -28406
rect 10880 -28423 11705 -28420
rect 11783 -29544 12203 -29502
rect 11783 -29595 11811 -29544
rect 12168 -29595 12203 -29544
rect 11783 -29633 12203 -29595
rect 12923 -29731 13137 -29725
rect 12923 -29765 12986 -29731
rect 13077 -29765 13137 -29731
rect 12923 -29791 13137 -29765
rect -12499 -30585 -12373 -30543
rect -12499 -31707 -12471 -30585
rect -12399 -31707 -12373 -30585
rect -12499 -31753 -12373 -31707
rect 7138 -31720 7963 -31717
rect 7138 -31755 7389 -31720
rect 7677 -31734 7963 -31720
rect 8086 -31720 8911 -31717
rect 7677 -31755 7964 -31734
rect 7138 -31771 7964 -31755
rect 8086 -31755 8337 -31720
rect 8625 -31734 8911 -31720
rect 9022 -31720 9847 -31717
rect 8625 -31755 8912 -31734
rect 8086 -31771 8912 -31755
rect 9022 -31755 9273 -31720
rect 9561 -31734 9847 -31720
rect 9953 -31719 10778 -31716
rect 9561 -31755 9848 -31734
rect 9022 -31771 9848 -31755
rect 9953 -31754 10204 -31719
rect 10492 -31733 10778 -31719
rect 10880 -31720 11705 -31717
rect 10492 -31754 10779 -31733
rect 9953 -31770 10779 -31754
rect 10880 -31755 11131 -31720
rect 11419 -31734 11705 -31720
rect 11419 -31755 11706 -31734
rect 10880 -31771 11706 -31755
rect 5658 -32241 5872 -32235
rect 5658 -32275 5721 -32241
rect 5812 -32275 5872 -32241
rect 5658 -32301 5872 -32275
rect 6098 -32241 6312 -32235
rect 6098 -32275 6161 -32241
rect 6252 -32275 6312 -32241
rect 6098 -32301 6312 -32275
rect 6538 -32241 6752 -32235
rect 6538 -32275 6601 -32241
rect 6692 -32275 6752 -32241
rect 6538 -32301 6752 -32275
rect 7138 -32913 7964 -32897
rect 7138 -32948 7389 -32913
rect 7677 -32934 7964 -32913
rect 8086 -32913 8912 -32897
rect 7677 -32948 7963 -32934
rect 7138 -32951 7963 -32948
rect 8086 -32948 8337 -32913
rect 8625 -32934 8912 -32913
rect 9022 -32913 9848 -32897
rect 8625 -32948 8911 -32934
rect 8086 -32951 8911 -32948
rect 9022 -32948 9273 -32913
rect 9561 -32934 9848 -32913
rect 9953 -32913 10779 -32897
rect 9561 -32948 9847 -32934
rect 9022 -32951 9847 -32948
rect 9953 -32948 10204 -32913
rect 10492 -32934 10779 -32913
rect 10880 -32913 11706 -32897
rect 10492 -32948 10778 -32934
rect 9953 -32951 10778 -32948
rect 10880 -32948 11131 -32913
rect 11419 -32934 11706 -32913
rect 11419 -32948 11705 -32934
rect 10880 -32951 11705 -32948
rect -12501 -33205 -12375 -33163
rect -12501 -34327 -12473 -33205
rect -12401 -34327 -12375 -33205
rect -12501 -34373 -12375 -34327
rect 11783 -34072 12203 -34030
rect 11783 -34123 11811 -34072
rect 12168 -34123 12203 -34072
rect 11783 -34161 12203 -34123
rect 12923 -34259 13137 -34253
rect 12923 -34293 12986 -34259
rect 13077 -34293 13137 -34259
rect 12923 -34319 13137 -34293
rect 13470 -35778 13536 -35715
rect 13470 -35869 13496 -35778
rect 13530 -35869 13536 -35778
rect 13470 -35929 13536 -35869
rect 7138 -36248 7963 -36245
rect 7138 -36283 7389 -36248
rect 7677 -36262 7963 -36248
rect 8086 -36248 8911 -36245
rect 7677 -36283 7964 -36262
rect 7138 -36299 7964 -36283
rect 8086 -36283 8337 -36248
rect 8625 -36262 8911 -36248
rect 9022 -36248 9847 -36245
rect 8625 -36283 8912 -36262
rect 8086 -36299 8912 -36283
rect 9022 -36283 9273 -36248
rect 9561 -36262 9847 -36248
rect 9953 -36247 10778 -36244
rect 9561 -36283 9848 -36262
rect 9022 -36299 9848 -36283
rect 9953 -36282 10204 -36247
rect 10492 -36261 10778 -36247
rect 10880 -36248 11705 -36245
rect 10492 -36282 10779 -36261
rect 9953 -36298 10779 -36282
rect 10880 -36283 11131 -36248
rect 11419 -36262 11705 -36248
rect 11419 -36283 11706 -36262
rect 10880 -36299 11706 -36283
rect 13470 -36157 13536 -36094
rect 13470 -36248 13496 -36157
rect 13530 -36248 13536 -36157
rect 13470 -36308 13536 -36248
<< psubdiffcont >>
rect 1841 4792 2964 4838
rect 3447 4792 4570 4838
rect 5151 4790 6274 4836
rect 7200 4787 7535 4821
rect 7840 4785 7972 4819
rect 5689 3237 5821 3271
rect 6129 3237 6261 3271
rect 6569 3237 6701 3271
rect -24001 3068 -22878 3114
rect -20710 3068 -19587 3114
rect -17419 3068 -16296 3114
rect -14128 3068 -13005 3114
rect -10837 3068 -9714 3114
rect -7547 3068 -6424 3114
rect -4256 3068 -3133 3114
rect -965 3068 158 3114
rect 7298 2118 7332 2466
rect 7298 1715 7332 2066
rect 8246 2118 8280 2466
rect 8246 1715 8280 2066
rect 9182 2118 9216 2466
rect 9182 1715 9216 2066
rect 10113 2118 10147 2466
rect 10113 1715 10147 2066
rect 11040 2118 11074 2466
rect 11040 1715 11074 2066
rect -24670 1284 -23547 1330
rect -23111 1284 -21988 1330
rect -21379 1284 -20256 1330
rect -19820 1284 -18697 1330
rect -18088 1284 -16965 1330
rect -16529 1284 -15406 1330
rect -14797 1284 -13674 1330
rect -13238 1284 -12115 1330
rect -11506 1284 -10383 1330
rect -9947 1284 -8824 1330
rect -8216 1284 -7093 1330
rect -6657 1284 -5534 1330
rect -4925 1284 -3802 1330
rect -3366 1284 -2243 1330
rect -1634 1284 -511 1330
rect -75 1284 1048 1330
rect 7298 1186 7332 1537
rect 7298 786 7332 1134
rect 8246 1186 8280 1537
rect 8246 786 8280 1134
rect 9182 1186 9216 1537
rect 9182 786 9216 1134
rect 10113 1187 10147 1538
rect 10113 787 10147 1135
rect 11040 1186 11074 1537
rect 11040 786 11074 1134
rect 12183 1188 12382 1249
rect 12954 1219 13086 1253
rect -24336 221 -24001 255
rect -23227 221 -22892 255
rect -22345 221 -22010 255
rect -21045 221 -20710 255
rect -19936 221 -19601 255
rect -19054 221 -18719 255
rect -17754 221 -17419 255
rect -16645 221 -16310 255
rect -15763 221 -15428 255
rect -14463 221 -14128 255
rect -13354 221 -13019 255
rect -12472 221 -12137 255
rect -11172 221 -10837 255
rect -10063 221 -9728 255
rect -9181 221 -8846 255
rect -7882 221 -7547 255
rect -6773 221 -6438 255
rect -5891 221 -5556 255
rect -4591 221 -4256 255
rect -3482 221 -3147 255
rect -2600 221 -2265 255
rect -1300 221 -965 255
rect -191 221 144 255
rect 691 221 1026 255
rect 5689 -1291 5821 -1257
rect 6129 -1291 6261 -1257
rect 6569 -1291 6701 -1257
rect 7298 -2410 7332 -2062
rect 7298 -2813 7332 -2462
rect 8246 -2410 8280 -2062
rect 8246 -2813 8280 -2462
rect 9182 -2410 9216 -2062
rect 9182 -2813 9216 -2462
rect 10113 -2410 10147 -2062
rect 10113 -2813 10147 -2462
rect 11040 -2410 11074 -2062
rect 11040 -2813 11074 -2462
rect -23597 -2993 -23465 -2959
rect -24186 -3067 -23851 -3033
rect -21577 -2993 -21445 -2959
rect -22149 -3067 -21814 -3033
rect -19836 -2993 -19704 -2959
rect -20419 -3067 -20084 -3033
rect -18057 -2993 -17925 -2959
rect -18659 -3067 -18324 -3033
rect 7298 -3342 7332 -2991
rect 7298 -3742 7332 -3394
rect 8246 -3342 8280 -2991
rect 8246 -3742 8280 -3394
rect 9182 -3342 9216 -2991
rect 9182 -3742 9216 -3394
rect 10113 -3341 10147 -2990
rect 10113 -3741 10147 -3393
rect 11040 -3342 11074 -2991
rect 11040 -3742 11074 -3394
rect 12183 -3340 12382 -3279
rect 12954 -3309 13086 -3275
rect -23553 -4805 -23421 -4771
rect -24135 -4879 -23800 -4845
rect -21815 -4805 -21683 -4771
rect -22399 -4879 -22064 -4845
rect -20603 -5276 -19480 -5230
rect -19044 -5276 -17921 -5230
rect -17312 -5276 -16189 -5230
rect -15753 -5276 -14630 -5230
rect -14021 -5276 -12898 -5230
rect -12462 -5276 -11339 -5230
rect -10730 -5276 -9607 -5230
rect -9171 -5276 -8048 -5230
rect 5689 -5719 5821 -5685
rect 6129 -5719 6261 -5685
rect 6569 -5719 6701 -5685
rect -23555 -6097 -23423 -6063
rect -24135 -6171 -23800 -6137
rect -21821 -6097 -21689 -6063
rect -22399 -6171 -22064 -6137
rect -20269 -6339 -19934 -6305
rect -19160 -6339 -18825 -6305
rect -18278 -6339 -17943 -6305
rect -16978 -6339 -16643 -6305
rect -15869 -6339 -15534 -6305
rect -14987 -6339 -14652 -6305
rect -13687 -6339 -13352 -6305
rect -12578 -6339 -12243 -6305
rect -11696 -6339 -11361 -6305
rect -10396 -6339 -10061 -6305
rect -9287 -6339 -8952 -6305
rect -8405 -6339 -8070 -6305
rect 7298 -6838 7332 -6490
rect 7298 -7241 7332 -6890
rect 8246 -6838 8280 -6490
rect 8246 -7241 8280 -6890
rect 9182 -6838 9216 -6490
rect 9182 -7241 9216 -6890
rect 10113 -6838 10147 -6490
rect 10113 -7241 10147 -6890
rect 11040 -6838 11074 -6490
rect 11040 -7241 11074 -6890
rect 7298 -7770 7332 -7419
rect -23553 -8070 -23421 -8036
rect -24135 -8144 -23800 -8110
rect -21819 -8070 -21687 -8036
rect -22398 -8144 -22063 -8110
rect 7298 -8170 7332 -7822
rect 8246 -7770 8280 -7419
rect 8246 -8170 8280 -7822
rect 9182 -7770 9216 -7419
rect 9182 -8170 9216 -7822
rect 10113 -7769 10147 -7418
rect 10113 -8169 10147 -7821
rect 11040 -7770 11074 -7419
rect 11040 -8170 11074 -7822
rect -20603 -8541 -19480 -8495
rect -19044 -8541 -17921 -8495
rect -17312 -8541 -16189 -8495
rect -15753 -8541 -14630 -8495
rect -14021 -8541 -12898 -8495
rect -12462 -8541 -11339 -8495
rect -10730 -8541 -9607 -8495
rect -9171 -8541 -8048 -8495
rect 12183 -7768 12382 -7707
rect 12954 -7737 13086 -7703
rect -23552 -9362 -23420 -9328
rect -24135 -9436 -23800 -9402
rect -21815 -9362 -21683 -9328
rect -22399 -9436 -22064 -9402
rect -20269 -9604 -19934 -9570
rect -19160 -9604 -18825 -9570
rect -18278 -9604 -17943 -9570
rect -16978 -9604 -16643 -9570
rect -15869 -9604 -15534 -9570
rect -14987 -9604 -14652 -9570
rect -13687 -9604 -13352 -9570
rect -12578 -9604 -12243 -9570
rect -11696 -9604 -11361 -9570
rect -10396 -9604 -10061 -9570
rect -9287 -9604 -8952 -9570
rect -8405 -9604 -8070 -9570
rect 5689 -10347 5821 -10313
rect 6129 -10347 6261 -10313
rect 6569 -10347 6701 -10313
rect -23552 -11334 -23420 -11300
rect -24135 -11408 -23800 -11374
rect -21819 -11334 -21687 -11300
rect -22398 -11408 -22063 -11374
rect 7298 -11466 7332 -11118
rect -20603 -11805 -19480 -11759
rect -19044 -11805 -17921 -11759
rect -17312 -11805 -16189 -11759
rect -15753 -11805 -14630 -11759
rect -14021 -11805 -12898 -11759
rect -12462 -11805 -11339 -11759
rect -10730 -11805 -9607 -11759
rect -9171 -11805 -8048 -11759
rect 7298 -11869 7332 -11518
rect 8246 -11466 8280 -11118
rect 8246 -11869 8280 -11518
rect 9182 -11466 9216 -11118
rect 9182 -11869 9216 -11518
rect 10113 -11466 10147 -11118
rect 10113 -11869 10147 -11518
rect 11040 -11466 11074 -11118
rect 11040 -11869 11074 -11518
rect 7298 -12398 7332 -12047
rect -23552 -12626 -23420 -12592
rect -24135 -12700 -23800 -12666
rect -21823 -12626 -21691 -12592
rect -22398 -12700 -22063 -12666
rect -20269 -12868 -19934 -12834
rect -19160 -12868 -18825 -12834
rect -18278 -12868 -17943 -12834
rect -16978 -12868 -16643 -12834
rect -15869 -12868 -15534 -12834
rect -14987 -12868 -14652 -12834
rect -13687 -12868 -13352 -12834
rect -12578 -12868 -12243 -12834
rect -11696 -12868 -11361 -12834
rect -10396 -12868 -10061 -12834
rect -9287 -12868 -8952 -12834
rect 7298 -12798 7332 -12450
rect 8246 -12398 8280 -12047
rect 8246 -12798 8280 -12450
rect 9182 -12398 9216 -12047
rect 9182 -12798 9216 -12450
rect 10113 -12397 10147 -12046
rect 10113 -12797 10147 -12449
rect 11040 -12398 11074 -12047
rect 11040 -12798 11074 -12450
rect -8405 -12868 -8070 -12834
rect 12183 -12396 12382 -12335
rect 12954 -12365 13086 -12331
rect -1460 -14001 -1426 -13869
rect -23829 -15289 -23795 -14954
rect -16917 -15107 -16856 -14908
rect -11070 -15345 -11024 -14222
rect -4176 -14366 -4142 -14234
rect -1460 -14380 -1426 -14248
rect -4176 -14806 -4142 -14674
rect -1460 -14820 -1426 -14688
rect 5689 -14875 5821 -14841
rect 6129 -14875 6261 -14841
rect 6569 -14875 6701 -14841
rect -4176 -15185 -4142 -15053
rect -1460 -15199 -1426 -15067
rect -7527 -15529 -7493 -15397
rect -4176 -15625 -4142 -15493
rect -1460 -15639 -1426 -15507
rect -7526 -16029 -7492 -15897
rect -4176 -16004 -4142 -15872
rect -23828 -16474 -23794 -16139
rect -1460 -16018 -1426 -15886
rect 7298 -15994 7332 -15646
rect -16917 -16507 -16856 -16308
rect -7527 -16509 -7493 -16377
rect -4176 -16444 -4142 -16312
rect -1460 -16458 -1426 -16326
rect 7298 -16397 7332 -16046
rect 8246 -15994 8280 -15646
rect 8246 -16397 8280 -16046
rect 9182 -15994 9216 -15646
rect 9182 -16397 9216 -16046
rect 10113 -15994 10147 -15646
rect 10113 -16397 10147 -16046
rect 11040 -15994 11074 -15646
rect 11040 -16397 11074 -16046
rect -23823 -17687 -23789 -17352
rect -20966 -18217 -20932 -18085
rect -16917 -17907 -16856 -17708
rect -15375 -18088 -15341 -17956
rect -11068 -18161 -11022 -17038
rect -4176 -16823 -4142 -16691
rect -7527 -17009 -7493 -16877
rect -1460 -16837 -1426 -16705
rect 7298 -16926 7332 -16575
rect -4176 -17263 -4142 -17131
rect -1460 -17277 -1426 -17145
rect 7298 -17326 7332 -16978
rect -7527 -17489 -7493 -17357
rect 8246 -16926 8280 -16575
rect 8246 -17326 8280 -16978
rect 9182 -16926 9216 -16575
rect 9182 -17326 9216 -16978
rect 10113 -16925 10147 -16574
rect 10113 -17325 10147 -16977
rect 11040 -16926 11074 -16575
rect 11040 -17326 11074 -16978
rect -4176 -17642 -4142 -17510
rect -1460 -17656 -1426 -17524
rect 12183 -16924 12382 -16863
rect 12954 -16893 13086 -16859
rect 16211 -16927 16541 -16814
rect -7527 -17949 -7493 -17817
rect -4176 -18082 -4142 -17950
rect -1460 -18096 -1426 -17964
rect -23808 -18806 -23774 -18471
rect -20965 -18717 -20931 -18585
rect -15374 -18588 -15340 -18456
rect -7541 -18409 -7507 -18277
rect -4176 -18461 -4142 -18329
rect -1460 -18475 -1426 -18343
rect -20966 -19197 -20932 -19065
rect -7539 -18889 -7505 -18757
rect -15375 -19068 -15341 -18936
rect -4176 -18901 -4142 -18769
rect -1460 -18915 -1426 -18783
rect -23806 -20000 -23772 -19665
rect -20966 -19697 -20932 -19565
rect -16917 -19307 -16856 -19108
rect -4176 -19280 -4142 -19148
rect -1460 -19294 -1426 -19162
rect 5689 -19403 5821 -19369
rect 6129 -19403 6261 -19369
rect 6569 -19403 6701 -19369
rect -15375 -19568 -15341 -19436
rect -4176 -19720 -4142 -19588
rect -1460 -19734 -1426 -19602
rect 17555 -18929 17890 -18895
rect 18127 -18933 18259 -18899
rect -20966 -20177 -20932 -20045
rect -15375 -20048 -15341 -19916
rect -20966 -20637 -20932 -20505
rect -23775 -21200 -23741 -20865
rect -20980 -21097 -20946 -20965
rect -16917 -20707 -16856 -20508
rect -15375 -20508 -15341 -20376
rect -15389 -20968 -15355 -20836
rect -11068 -21118 -11022 -19995
rect -4176 -20099 -4142 -19967
rect -1460 -20113 -1426 -19981
rect -4176 -20539 -4142 -20407
rect -1460 -20553 -1426 -20421
rect 7298 -20522 7332 -20174
rect -4176 -20918 -4142 -20786
rect 7298 -20925 7332 -20574
rect 8246 -20522 8280 -20174
rect 8246 -20925 8280 -20574
rect 9182 -20522 9216 -20174
rect 9182 -20925 9216 -20574
rect 10113 -20522 10147 -20174
rect 10113 -20925 10147 -20574
rect 11040 -20522 11074 -20174
rect 11040 -20925 11074 -20574
rect 16211 -20358 16541 -20245
rect -20978 -21577 -20944 -21445
rect -15387 -21448 -15353 -21316
rect 7298 -21454 7332 -21103
rect 7298 -21854 7332 -21506
rect 8246 -21454 8280 -21103
rect 8246 -21854 8280 -21506
rect 9182 -21454 9216 -21103
rect 9182 -21854 9216 -21506
rect 10113 -21453 10147 -21102
rect 10113 -21853 10147 -21505
rect 11040 -21454 11074 -21103
rect 11040 -21854 11074 -21506
rect -23776 -22503 -23742 -22168
rect -16917 -22107 -16856 -21908
rect 12183 -21452 12382 -21391
rect 12954 -21421 13086 -21387
rect -23776 -23812 -23742 -23477
rect -16917 -23507 -16856 -23308
rect -11068 -23697 -11022 -22574
rect 5689 -23931 5821 -23897
rect 6129 -23931 6261 -23897
rect 6569 -23931 6701 -23897
rect -16917 -24907 -16856 -24708
rect 7298 -25050 7332 -24702
rect -11068 -26465 -11022 -25342
rect 7298 -25453 7332 -25102
rect 8246 -25050 8280 -24702
rect 8246 -25453 8280 -25102
rect 9182 -25050 9216 -24702
rect 9182 -25453 9216 -25102
rect 10113 -25050 10147 -24702
rect 10113 -25453 10147 -25102
rect 11040 -25050 11074 -24702
rect 11040 -25453 11074 -25102
rect 7298 -25982 7332 -25631
rect 7298 -26382 7332 -26034
rect 8246 -25982 8280 -25631
rect 8246 -26382 8280 -26034
rect 9182 -25982 9216 -25631
rect 9182 -26382 9216 -26034
rect 10113 -25981 10147 -25630
rect 10113 -26381 10147 -26033
rect 11040 -25982 11074 -25631
rect 11040 -26382 11074 -26034
rect 12183 -25980 12382 -25919
rect 12954 -25949 13086 -25915
rect -11068 -29098 -11022 -27975
rect 5689 -28459 5821 -28425
rect 6129 -28459 6261 -28425
rect 6569 -28459 6701 -28425
rect 7298 -29578 7332 -29230
rect 7298 -29981 7332 -29630
rect 8246 -29578 8280 -29230
rect 8246 -29981 8280 -29630
rect 9182 -29578 9216 -29230
rect 9182 -29981 9216 -29630
rect 10113 -29578 10147 -29230
rect 10113 -29981 10147 -29630
rect 11040 -29578 11074 -29230
rect 11040 -29981 11074 -29630
rect 7298 -30510 7332 -30159
rect -11068 -31707 -11022 -30584
rect 7298 -30910 7332 -30562
rect 8246 -30510 8280 -30159
rect 8246 -30910 8280 -30562
rect 9182 -30510 9216 -30159
rect 9182 -30910 9216 -30562
rect 10113 -30509 10147 -30158
rect 10113 -30909 10147 -30561
rect 11040 -30510 11074 -30159
rect 11040 -30910 11074 -30562
rect 12183 -30508 12382 -30447
rect 12954 -30477 13086 -30443
rect 5689 -32987 5821 -32953
rect 6129 -32987 6261 -32953
rect 6569 -32987 6701 -32953
rect -11070 -34327 -11024 -33204
rect 7298 -34106 7332 -33758
rect 7298 -34509 7332 -34158
rect 8246 -34106 8280 -33758
rect 8246 -34509 8280 -34158
rect 9182 -34106 9216 -33758
rect 9182 -34509 9216 -34158
rect 10113 -34106 10147 -33758
rect 10113 -34509 10147 -34158
rect 11040 -34106 11074 -33758
rect 11040 -34509 11074 -34158
rect 7298 -35038 7332 -34687
rect 7298 -35438 7332 -35090
rect 8246 -35038 8280 -34687
rect 8246 -35438 8280 -35090
rect 9182 -35038 9216 -34687
rect 9182 -35438 9216 -35090
rect 10113 -35037 10147 -34686
rect 10113 -35437 10147 -35089
rect 11040 -35038 11074 -34687
rect 11040 -35438 11074 -35090
rect 12183 -35036 12382 -34975
rect 12954 -35005 13086 -34971
rect 12784 -35878 12818 -35746
rect 12784 -36257 12818 -36125
<< nsubdiffcont >>
rect 1841 6169 2963 6241
rect 3447 6169 4569 6241
rect 5151 6167 6273 6239
rect 6967 5507 7536 5554
rect 7872 5497 7963 5531
rect -24000 4445 -22878 4517
rect -20709 4445 -19587 4517
rect -17418 4445 -16296 4517
rect -14127 4445 -13005 4517
rect -10836 4445 -9714 4517
rect -7546 4445 -6424 4517
rect -4255 4445 -3133 4517
rect -964 4445 158 4517
rect 5721 3949 5812 3983
rect 6161 3949 6252 3983
rect 6601 3949 6692 3983
rect 7389 3276 7677 3311
rect 8337 3276 8625 3311
rect 9273 3276 9561 3311
rect 10204 3276 10492 3311
rect 11131 3276 11419 3311
rect -24670 2661 -23548 2733
rect -23111 2661 -21989 2733
rect -21379 2661 -20257 2733
rect -19820 2661 -18698 2733
rect -18088 2661 -16966 2733
rect -16529 2661 -15407 2733
rect -14797 2661 -13675 2733
rect -13238 2661 -12116 2733
rect -11506 2661 -10384 2733
rect -9947 2661 -8825 2733
rect -8216 2661 -7094 2733
rect -6657 2661 -5535 2733
rect -4925 2661 -3803 2733
rect -3366 2661 -2244 2733
rect -1634 2661 -512 2733
rect -75 2661 1047 2733
rect 11811 2101 12168 2152
rect 12986 1931 13077 1965
rect -24569 941 -24000 988
rect -23460 941 -22891 988
rect -22578 941 -22009 988
rect -21278 941 -20709 988
rect -20169 941 -19600 988
rect -19287 941 -18718 988
rect -17987 941 -17418 988
rect -16878 941 -16309 988
rect -15996 941 -15427 988
rect -14696 941 -14127 988
rect -13587 941 -13018 988
rect -12705 941 -12136 988
rect -11405 941 -10836 988
rect -10296 941 -9727 988
rect -9414 941 -8845 988
rect -8115 941 -7546 988
rect -7006 941 -6437 988
rect -6124 941 -5555 988
rect -4824 941 -4255 988
rect -3715 941 -3146 988
rect -2833 941 -2264 988
rect -1533 941 -964 988
rect -424 941 145 988
rect 458 941 1027 988
rect 7389 -59 7677 -24
rect 8337 -59 8625 -24
rect 9273 -59 9561 -24
rect 10204 -58 10492 -23
rect 11131 -59 11419 -24
rect 5721 -579 5812 -545
rect 6161 -579 6252 -545
rect 6601 -579 6692 -545
rect 7389 -1252 7677 -1217
rect 8337 -1252 8625 -1217
rect 9273 -1252 9561 -1217
rect 10204 -1252 10492 -1217
rect 11131 -1252 11419 -1217
rect -23565 -2281 -23474 -2247
rect -24419 -2347 -23850 -2300
rect -21545 -2281 -21454 -2247
rect -22382 -2347 -21813 -2300
rect -19804 -2281 -19713 -2247
rect -20652 -2347 -20083 -2300
rect -18025 -2281 -17934 -2247
rect -18892 -2347 -18323 -2300
rect 11811 -2427 12168 -2376
rect 12986 -2597 13077 -2563
rect -20603 -3899 -19481 -3827
rect -19044 -3899 -17922 -3827
rect -17312 -3899 -16190 -3827
rect -15753 -3899 -14631 -3827
rect -14021 -3899 -12899 -3827
rect -12462 -3899 -11340 -3827
rect -10730 -3899 -9608 -3827
rect -9171 -3899 -8049 -3827
rect -23521 -4093 -23430 -4059
rect -24368 -4159 -23799 -4112
rect -21783 -4093 -21692 -4059
rect -22632 -4159 -22063 -4112
rect 7389 -4587 7677 -4552
rect 8337 -4587 8625 -4552
rect 9273 -4587 9561 -4552
rect 10204 -4586 10492 -4551
rect 11131 -4587 11419 -4552
rect 5721 -5007 5812 -4973
rect 6161 -5007 6252 -4973
rect -23523 -5385 -23432 -5351
rect -24368 -5451 -23799 -5404
rect -21789 -5385 -21698 -5351
rect 6601 -5007 6692 -4973
rect -22632 -5451 -22063 -5404
rect -20502 -5619 -19933 -5572
rect -19393 -5619 -18824 -5572
rect -18511 -5619 -17942 -5572
rect -17211 -5619 -16642 -5572
rect -16102 -5619 -15533 -5572
rect -15220 -5619 -14651 -5572
rect -13920 -5619 -13351 -5572
rect -12811 -5619 -12242 -5572
rect -11929 -5619 -11360 -5572
rect -10629 -5619 -10060 -5572
rect -9520 -5619 -8951 -5572
rect -8638 -5619 -8069 -5572
rect 7389 -5680 7677 -5645
rect 8337 -5680 8625 -5645
rect 9273 -5680 9561 -5645
rect 10204 -5680 10492 -5645
rect 11131 -5680 11419 -5645
rect -20603 -7164 -19481 -7092
rect -19044 -7164 -17922 -7092
rect -17312 -7164 -16190 -7092
rect -15753 -7164 -14631 -7092
rect -14021 -7164 -12899 -7092
rect -12462 -7164 -11340 -7092
rect -10730 -7164 -9608 -7092
rect -9171 -7164 -8049 -7092
rect -23521 -7358 -23430 -7324
rect -24368 -7424 -23799 -7377
rect -21787 -7358 -21696 -7324
rect -22631 -7424 -22062 -7377
rect 11811 -6855 12168 -6804
rect 12986 -7025 13077 -6991
rect -23520 -8650 -23429 -8616
rect -24368 -8716 -23799 -8669
rect -21783 -8650 -21692 -8616
rect -22632 -8716 -22063 -8669
rect -20502 -8884 -19933 -8837
rect -19393 -8884 -18824 -8837
rect -18511 -8884 -17942 -8837
rect -17211 -8884 -16642 -8837
rect -16102 -8884 -15533 -8837
rect -15220 -8884 -14651 -8837
rect -13920 -8884 -13351 -8837
rect -12811 -8884 -12242 -8837
rect -11929 -8884 -11360 -8837
rect -10629 -8884 -10060 -8837
rect -9520 -8884 -8951 -8837
rect -8638 -8884 -8069 -8837
rect 7389 -9015 7677 -8980
rect 8337 -9015 8625 -8980
rect 9273 -9015 9561 -8980
rect 10204 -9014 10492 -8979
rect 11131 -9015 11419 -8980
rect 5721 -9635 5812 -9601
rect 6161 -9635 6252 -9601
rect 6601 -9635 6692 -9601
rect 7389 -10308 7677 -10273
rect 8337 -10308 8625 -10273
rect 9273 -10308 9561 -10273
rect 10204 -10308 10492 -10273
rect 11131 -10308 11419 -10273
rect -20603 -10428 -19481 -10356
rect -19044 -10428 -17922 -10356
rect -17312 -10428 -16190 -10356
rect -15753 -10428 -14631 -10356
rect -14021 -10428 -12899 -10356
rect -12462 -10428 -11340 -10356
rect -10730 -10428 -9608 -10356
rect -9171 -10428 -8049 -10356
rect -23520 -10622 -23429 -10588
rect -24368 -10688 -23799 -10641
rect -21787 -10622 -21696 -10588
rect -22631 -10688 -22062 -10641
rect -23520 -11914 -23429 -11880
rect -24368 -11980 -23799 -11933
rect -21791 -11914 -21700 -11880
rect 11811 -11483 12168 -11432
rect 12986 -11653 13077 -11619
rect -22631 -11980 -22062 -11933
rect -20502 -12148 -19933 -12101
rect -19393 -12148 -18824 -12101
rect -18511 -12148 -17942 -12101
rect -17211 -12148 -16642 -12101
rect -16102 -12148 -15533 -12101
rect -15220 -12148 -14651 -12101
rect -13920 -12148 -13351 -12101
rect -12811 -12148 -12242 -12101
rect -11929 -12148 -11360 -12101
rect -10629 -12148 -10060 -12101
rect -9520 -12148 -8951 -12101
rect -8638 -12148 -8069 -12101
rect 7389 -13643 7677 -13608
rect 8337 -13643 8625 -13608
rect 9273 -13643 9561 -13608
rect 10204 -13642 10492 -13607
rect 11131 -13643 11419 -13608
rect -2172 -13969 -2138 -13878
rect -24562 -15522 -24515 -14953
rect -17820 -15479 -17769 -15122
rect -12473 -15345 -12401 -14223
rect 5721 -14163 5812 -14129
rect -4888 -14357 -4854 -14266
rect -2172 -14348 -2138 -14257
rect 6161 -14163 6252 -14129
rect 6601 -14163 6692 -14129
rect -4888 -14797 -4854 -14706
rect -2172 -14788 -2138 -14697
rect 7389 -14836 7677 -14801
rect 8337 -14836 8625 -14801
rect 9273 -14836 9561 -14801
rect 10204 -14836 10492 -14801
rect 11131 -14836 11419 -14801
rect -4888 -15176 -4854 -15085
rect -2172 -15167 -2138 -15076
rect -8239 -15497 -8205 -15406
rect -4888 -15616 -4854 -15525
rect -2172 -15607 -2138 -15516
rect -8238 -15997 -8204 -15906
rect -4888 -15995 -4854 -15904
rect -2172 -15986 -2138 -15895
rect -24561 -16707 -24514 -16138
rect -17820 -16879 -17769 -16522
rect -8239 -16477 -8205 -16386
rect -4888 -16435 -4854 -16344
rect -2172 -16426 -2138 -16335
rect 11811 -16011 12168 -15960
rect 12986 -16181 13077 -16147
rect -4888 -16814 -4854 -16723
rect -8239 -16977 -8205 -16886
rect -24556 -17920 -24509 -17351
rect -21678 -18185 -21644 -18094
rect -17820 -18279 -17769 -17922
rect -16087 -18056 -16053 -17965
rect -12471 -18161 -12399 -17039
rect -2172 -16805 -2138 -16714
rect -4888 -17254 -4854 -17163
rect -8239 -17457 -8205 -17366
rect -2172 -17245 -2138 -17154
rect -4888 -17633 -4854 -17542
rect -2172 -17624 -2138 -17533
rect -8239 -17917 -8205 -17826
rect -4888 -18073 -4854 -17982
rect -2172 -18064 -2138 -17973
rect 15703 -18033 15737 -17679
rect -24541 -19039 -24494 -18470
rect -21677 -18685 -21643 -18594
rect -16086 -18556 -16052 -18465
rect -8253 -18377 -8219 -18286
rect 7389 -18171 7677 -18136
rect 8337 -18171 8625 -18136
rect 9273 -18171 9561 -18136
rect 10204 -18170 10492 -18135
rect 11131 -18171 11419 -18136
rect -4888 -18452 -4854 -18361
rect -2172 -18443 -2138 -18352
rect 17322 -18209 17891 -18162
rect 18159 -18221 18250 -18187
rect -8251 -18857 -8217 -18766
rect -21678 -19165 -21644 -19074
rect -16087 -19036 -16053 -18945
rect 5721 -18691 5812 -18657
rect -4888 -18892 -4854 -18801
rect -2172 -18883 -2138 -18792
rect 6161 -18691 6252 -18657
rect 6601 -18691 6692 -18657
rect -24539 -20233 -24492 -19664
rect -21678 -19665 -21644 -19574
rect -17820 -19679 -17769 -19322
rect -4888 -19271 -4854 -19180
rect -2172 -19262 -2138 -19171
rect -16087 -19536 -16053 -19445
rect 7389 -19364 7677 -19329
rect 8337 -19364 8625 -19329
rect 9273 -19364 9561 -19329
rect 10204 -19364 10492 -19329
rect 11131 -19364 11419 -19329
rect -4888 -19711 -4854 -19620
rect -2172 -19702 -2138 -19611
rect 15703 -19493 15737 -19139
rect -21678 -20145 -21644 -20054
rect -16087 -20016 -16053 -19925
rect -21678 -20605 -21644 -20514
rect -16087 -20476 -16053 -20385
rect -24508 -21433 -24461 -20864
rect -21692 -21065 -21658 -20974
rect -17820 -21079 -17769 -20722
rect -16101 -20936 -16067 -20845
rect -12471 -21118 -12399 -19996
rect -4888 -20090 -4854 -19999
rect -2172 -20081 -2138 -19990
rect -4888 -20530 -4854 -20439
rect -2172 -20521 -2138 -20430
rect -4888 -20909 -4854 -20818
rect 11811 -20539 12168 -20488
rect 12986 -20709 13077 -20675
rect -21690 -21545 -21656 -21454
rect -16099 -21416 -16065 -21325
rect -24509 -22736 -24462 -22167
rect -17820 -22479 -17769 -22122
rect -24509 -24045 -24462 -23476
rect -17820 -23879 -17769 -23522
rect -12471 -23697 -12399 -22575
rect 7389 -22699 7677 -22664
rect 8337 -22699 8625 -22664
rect 9273 -22699 9561 -22664
rect 10204 -22698 10492 -22663
rect 11131 -22699 11419 -22664
rect 5721 -23219 5812 -23185
rect 6161 -23219 6252 -23185
rect 6601 -23219 6692 -23185
rect 7389 -23892 7677 -23857
rect 8337 -23892 8625 -23857
rect 9273 -23892 9561 -23857
rect 10204 -23892 10492 -23857
rect 11131 -23892 11419 -23857
rect -17820 -25279 -17769 -24922
rect -12471 -26465 -12399 -25343
rect 11811 -25067 12168 -25016
rect 12986 -25237 13077 -25203
rect 7389 -27227 7677 -27192
rect 8337 -27227 8625 -27192
rect 9273 -27227 9561 -27192
rect 10204 -27226 10492 -27191
rect 11131 -27227 11419 -27192
rect 5721 -27747 5812 -27713
rect -12471 -29098 -12399 -27976
rect 6161 -27747 6252 -27713
rect 6601 -27747 6692 -27713
rect 7389 -28420 7677 -28385
rect 8337 -28420 8625 -28385
rect 9273 -28420 9561 -28385
rect 10204 -28420 10492 -28385
rect 11131 -28420 11419 -28385
rect 11811 -29595 12168 -29544
rect 12986 -29765 13077 -29731
rect -12471 -31707 -12399 -30585
rect 7389 -31755 7677 -31720
rect 8337 -31755 8625 -31720
rect 9273 -31755 9561 -31720
rect 10204 -31754 10492 -31719
rect 11131 -31755 11419 -31720
rect 5721 -32275 5812 -32241
rect 6161 -32275 6252 -32241
rect 6601 -32275 6692 -32241
rect 7389 -32948 7677 -32913
rect 8337 -32948 8625 -32913
rect 9273 -32948 9561 -32913
rect 10204 -32948 10492 -32913
rect 11131 -32948 11419 -32913
rect -12473 -34327 -12401 -33205
rect 11811 -34123 12168 -34072
rect 12986 -34293 13077 -34259
rect 13496 -35869 13530 -35778
rect 7389 -36283 7677 -36248
rect 8337 -36283 8625 -36248
rect 9273 -36283 9561 -36248
rect 10204 -36282 10492 -36247
rect 11131 -36283 11419 -36248
rect 13496 -36248 13530 -36157
<< poly >>
rect 1765 6084 1795 6110
rect 1857 6084 1887 6115
rect 1953 6084 1983 6115
rect 2049 6084 2079 6115
rect 2145 6084 2175 6115
rect 2241 6084 2271 6115
rect 2337 6084 2367 6115
rect 2433 6084 2463 6115
rect 2529 6084 2559 6115
rect 2625 6084 2655 6115
rect 2721 6084 2751 6115
rect 2817 6084 2847 6115
rect 2913 6084 2943 6115
rect 3005 6084 3035 6110
rect 3371 6084 3401 6110
rect 3463 6084 3493 6115
rect 3559 6084 3589 6115
rect 3655 6084 3685 6115
rect 3751 6084 3781 6115
rect 3847 6084 3877 6115
rect 3943 6084 3973 6115
rect 4039 6084 4069 6115
rect 4135 6084 4165 6115
rect 4231 6084 4261 6115
rect 4327 6084 4357 6115
rect 4423 6084 4453 6115
rect 4519 6084 4549 6115
rect 4611 6084 4641 6110
rect 5075 6082 5105 6108
rect 5167 6082 5197 6113
rect 5263 6082 5293 6113
rect 5359 6082 5389 6113
rect 5455 6082 5485 6113
rect 5551 6082 5581 6113
rect 5647 6082 5677 6113
rect 5743 6082 5773 6113
rect 5839 6082 5869 6113
rect 5935 6082 5965 6113
rect 6031 6082 6061 6113
rect 6127 6082 6157 6113
rect 6223 6082 6253 6113
rect 6315 6082 6345 6108
rect 1765 5503 1795 5534
rect 1857 5503 1887 5534
rect 1953 5503 1983 5534
rect 2049 5503 2079 5534
rect 2145 5504 2175 5534
rect 2241 5504 2271 5534
rect 2337 5504 2367 5534
rect 1732 5353 2081 5503
rect 2145 5475 2367 5504
rect 2145 5430 2175 5475
rect 2305 5430 2367 5475
rect 2145 5411 2367 5430
rect 2433 5503 2463 5534
rect 2529 5503 2559 5534
rect 2625 5503 2655 5534
rect 2433 5470 2655 5503
rect 2433 5425 2506 5470
rect 2636 5425 2655 5470
rect 2433 5410 2655 5425
rect 2721 5503 2751 5534
rect 2817 5503 2847 5534
rect 2913 5503 2943 5534
rect 3005 5503 3035 5534
rect 3371 5503 3401 5534
rect 3463 5503 3493 5534
rect 3559 5503 3589 5534
rect 3655 5503 3685 5534
rect 3751 5504 3781 5534
rect 3847 5504 3877 5534
rect 3943 5504 3973 5534
rect 1557 5343 2655 5353
rect 1557 5254 1573 5343
rect 1662 5254 2655 5343
rect 1557 5244 2655 5254
rect 1732 5069 1808 5244
rect 1857 5154 2079 5179
rect 1857 5109 1900 5154
rect 2030 5109 2079 5154
rect 1765 5044 1795 5069
rect 1857 5066 2079 5109
rect 1857 5044 1887 5066
rect 1953 5044 1983 5066
rect 2049 5044 2079 5066
rect 2145 5146 2367 5174
rect 2145 5101 2183 5146
rect 2313 5101 2367 5146
rect 2145 5066 2367 5101
rect 2145 5044 2175 5066
rect 2241 5044 2271 5066
rect 2337 5044 2367 5066
rect 2433 5066 2655 5244
rect 2433 5044 2463 5066
rect 2529 5044 2559 5066
rect 2625 5044 2655 5066
rect 2721 5346 3035 5503
rect 3338 5353 3687 5503
rect 3751 5475 3973 5504
rect 3751 5430 3781 5475
rect 3911 5430 3973 5475
rect 3751 5411 3973 5430
rect 4039 5503 4069 5534
rect 4135 5503 4165 5534
rect 4231 5503 4261 5534
rect 4039 5470 4261 5503
rect 4039 5425 4112 5470
rect 4242 5425 4261 5470
rect 4039 5410 4261 5425
rect 4327 5503 4357 5534
rect 4423 5503 4453 5534
rect 4519 5503 4549 5534
rect 4611 5503 4641 5534
rect 2721 5291 2753 5346
rect 2818 5291 3035 5346
rect 2721 5066 3035 5291
rect 3171 5343 4261 5353
rect 3171 5254 3187 5343
rect 3276 5254 4261 5343
rect 3171 5244 4261 5254
rect 3338 5069 3414 5244
rect 3463 5154 3685 5179
rect 3463 5109 3506 5154
rect 3636 5109 3685 5154
rect 2721 5044 2751 5066
rect 2817 5044 2847 5066
rect 2913 5044 2943 5066
rect 3005 5044 3035 5066
rect 3371 5044 3401 5069
rect 3463 5066 3685 5109
rect 3463 5044 3493 5066
rect 3559 5044 3589 5066
rect 3655 5044 3685 5066
rect 3751 5146 3973 5174
rect 3751 5101 3789 5146
rect 3919 5101 3973 5146
rect 3751 5066 3973 5101
rect 3751 5044 3781 5066
rect 3847 5044 3877 5066
rect 3943 5044 3973 5066
rect 4039 5066 4261 5244
rect 4039 5044 4069 5066
rect 4135 5044 4165 5066
rect 4231 5044 4261 5066
rect 4327 5346 4641 5503
rect 5075 5501 5105 5532
rect 5167 5501 5197 5532
rect 5263 5501 5293 5532
rect 5359 5501 5389 5532
rect 5455 5502 5485 5532
rect 5551 5502 5581 5532
rect 5647 5502 5677 5532
rect 5042 5351 5391 5501
rect 5455 5473 5677 5502
rect 5455 5428 5485 5473
rect 5615 5428 5677 5473
rect 5455 5409 5677 5428
rect 5743 5501 5773 5532
rect 5839 5501 5869 5532
rect 5935 5501 5965 5532
rect 5743 5468 5965 5501
rect 5743 5423 5816 5468
rect 5946 5423 5965 5468
rect 5743 5408 5965 5423
rect 6031 5501 6061 5532
rect 6127 5501 6157 5532
rect 6223 5501 6253 5532
rect 6315 5501 6345 5532
rect 4327 5291 4359 5346
rect 4424 5291 4641 5346
rect 4327 5066 4641 5291
rect 4855 5341 5965 5351
rect 4855 5252 4871 5341
rect 4960 5252 5965 5341
rect 4855 5242 5965 5252
rect 5042 5067 5118 5242
rect 5167 5152 5389 5177
rect 5167 5107 5210 5152
rect 5340 5107 5389 5152
rect 4327 5044 4357 5066
rect 4423 5044 4453 5066
rect 4519 5044 4549 5066
rect 4611 5044 4641 5066
rect 5075 5042 5105 5067
rect 5167 5064 5389 5107
rect 5167 5042 5197 5064
rect 5263 5042 5293 5064
rect 5359 5042 5389 5064
rect 5455 5144 5677 5172
rect 5455 5099 5493 5144
rect 5623 5099 5677 5144
rect 5455 5064 5677 5099
rect 5455 5042 5485 5064
rect 5551 5042 5581 5064
rect 5647 5042 5677 5064
rect 5743 5064 5965 5242
rect 5743 5042 5773 5064
rect 5839 5042 5869 5064
rect 5935 5042 5965 5064
rect 6031 5344 6345 5501
rect 7001 5441 7031 5472
rect 7097 5441 7127 5472
rect 7193 5441 7223 5472
rect 7289 5441 7319 5472
rect 7385 5441 7415 5472
rect 7481 5441 7511 5472
rect 6031 5289 6063 5344
rect 6128 5289 6345 5344
rect 6031 5064 6345 5289
rect 7712 5411 7778 5427
rect 7001 5201 7031 5227
rect 7097 5201 7127 5227
rect 7193 5201 7223 5227
rect 6031 5042 6061 5064
rect 6127 5042 6157 5064
rect 6223 5042 6253 5064
rect 6315 5042 6345 5064
rect 7000 5180 7223 5201
rect 7000 5145 7017 5180
rect 7051 5171 7223 5180
rect 7289 5201 7319 5227
rect 7385 5201 7415 5227
rect 7481 5201 7511 5227
rect 7289 5180 7511 5201
rect 7051 5145 7067 5171
rect 7000 5134 7067 5145
rect 7289 5145 7306 5180
rect 7340 5171 7511 5180
rect 7712 5185 7728 5411
rect 7762 5409 7778 5411
rect 7762 5379 7809 5409
rect 8023 5379 8049 5409
rect 7762 5313 7778 5379
rect 7762 5283 7809 5313
rect 8023 5283 8049 5313
rect 7762 5217 7778 5283
rect 7762 5187 7809 5217
rect 8023 5187 8049 5217
rect 7762 5185 7778 5187
rect 7340 5145 7356 5171
rect 7712 5169 7778 5185
rect 7289 5134 7356 5145
rect 1765 4888 1795 4914
rect 1857 4888 1887 4914
rect 1953 4888 1983 4914
rect 2049 4888 2079 4914
rect 2145 4888 2175 4914
rect 2241 4888 2271 4914
rect 2337 4888 2367 4914
rect 2433 4888 2463 4914
rect 2529 4888 2559 4914
rect 2625 4888 2655 4914
rect 2721 4888 2751 4914
rect 2817 4888 2847 4914
rect 2913 4888 2943 4914
rect 3005 4888 3035 4914
rect 3371 4888 3401 4914
rect 3463 4888 3493 4914
rect 3559 4888 3589 4914
rect 3655 4888 3685 4914
rect 3751 4888 3781 4914
rect 3847 4888 3877 4914
rect 3943 4888 3973 4914
rect 4039 4888 4069 4914
rect 4135 4888 4165 4914
rect 4231 4888 4261 4914
rect 4327 4888 4357 4914
rect 4423 4888 4453 4914
rect 4519 4888 4549 4914
rect 4611 4888 4641 4914
rect 7000 4939 7043 5134
rect 7085 5056 7151 5072
rect 7085 5021 7101 5056
rect 7135 5035 7151 5056
rect 7135 5021 7173 5035
rect 7085 5005 7173 5021
rect 7573 5005 7599 5035
rect 7712 4965 7779 4981
rect 7000 4923 7173 4939
rect 5075 4886 5105 4912
rect 5167 4886 5197 4912
rect 5263 4886 5293 4912
rect 5359 4886 5389 4912
rect 5455 4886 5485 4912
rect 5551 4886 5581 4912
rect 5647 4886 5677 4912
rect 5743 4886 5773 4912
rect 5839 4886 5869 4912
rect 5935 4886 5965 4912
rect 6031 4886 6061 4912
rect 6127 4886 6157 4912
rect 6223 4886 6253 4912
rect 6315 4886 6345 4912
rect 7000 4888 7101 4923
rect 7135 4909 7173 4923
rect 7573 4909 7599 4939
rect 7712 4931 7728 4965
rect 7762 4963 7779 4965
rect 7762 4933 7809 4963
rect 8009 4933 8035 4963
rect 7762 4931 7779 4933
rect 7712 4915 7779 4931
rect 7135 4888 7151 4909
rect 7000 4872 7151 4888
rect -24072 4360 -24042 4386
rect -23980 4360 -23950 4391
rect -23884 4360 -23854 4391
rect -23788 4360 -23758 4391
rect -23692 4360 -23662 4391
rect -23596 4360 -23566 4391
rect -23500 4360 -23470 4391
rect -23404 4360 -23374 4391
rect -23308 4360 -23278 4391
rect -23212 4360 -23182 4391
rect -23116 4360 -23086 4391
rect -23020 4360 -22990 4391
rect -22924 4360 -22894 4391
rect -22832 4360 -22802 4386
rect -20781 4360 -20751 4386
rect -20689 4360 -20659 4391
rect -20593 4360 -20563 4391
rect -20497 4360 -20467 4391
rect -20401 4360 -20371 4391
rect -20305 4360 -20275 4391
rect -20209 4360 -20179 4391
rect -20113 4360 -20083 4391
rect -20017 4360 -19987 4391
rect -19921 4360 -19891 4391
rect -19825 4360 -19795 4391
rect -19729 4360 -19699 4391
rect -19633 4360 -19603 4391
rect -19541 4360 -19511 4386
rect -17490 4360 -17460 4386
rect -17398 4360 -17368 4391
rect -17302 4360 -17272 4391
rect -17206 4360 -17176 4391
rect -17110 4360 -17080 4391
rect -17014 4360 -16984 4391
rect -16918 4360 -16888 4391
rect -16822 4360 -16792 4391
rect -16726 4360 -16696 4391
rect -16630 4360 -16600 4391
rect -16534 4360 -16504 4391
rect -16438 4360 -16408 4391
rect -16342 4360 -16312 4391
rect -16250 4360 -16220 4386
rect -14199 4360 -14169 4386
rect -14107 4360 -14077 4391
rect -14011 4360 -13981 4391
rect -13915 4360 -13885 4391
rect -13819 4360 -13789 4391
rect -13723 4360 -13693 4391
rect -13627 4360 -13597 4391
rect -13531 4360 -13501 4391
rect -13435 4360 -13405 4391
rect -13339 4360 -13309 4391
rect -13243 4360 -13213 4391
rect -13147 4360 -13117 4391
rect -13051 4360 -13021 4391
rect -12959 4360 -12929 4386
rect -10908 4360 -10878 4386
rect -10816 4360 -10786 4391
rect -10720 4360 -10690 4391
rect -10624 4360 -10594 4391
rect -10528 4360 -10498 4391
rect -10432 4360 -10402 4391
rect -10336 4360 -10306 4391
rect -10240 4360 -10210 4391
rect -10144 4360 -10114 4391
rect -10048 4360 -10018 4391
rect -9952 4360 -9922 4391
rect -9856 4360 -9826 4391
rect -9760 4360 -9730 4391
rect -9668 4360 -9638 4386
rect -7618 4360 -7588 4386
rect -7526 4360 -7496 4391
rect -7430 4360 -7400 4391
rect -7334 4360 -7304 4391
rect -7238 4360 -7208 4391
rect -7142 4360 -7112 4391
rect -7046 4360 -7016 4391
rect -6950 4360 -6920 4391
rect -6854 4360 -6824 4391
rect -6758 4360 -6728 4391
rect -6662 4360 -6632 4391
rect -6566 4360 -6536 4391
rect -6470 4360 -6440 4391
rect -6378 4360 -6348 4386
rect -4327 4360 -4297 4386
rect -4235 4360 -4205 4391
rect -4139 4360 -4109 4391
rect -4043 4360 -4013 4391
rect -3947 4360 -3917 4391
rect -3851 4360 -3821 4391
rect -3755 4360 -3725 4391
rect -3659 4360 -3629 4391
rect -3563 4360 -3533 4391
rect -3467 4360 -3437 4391
rect -3371 4360 -3341 4391
rect -3275 4360 -3245 4391
rect -3179 4360 -3149 4391
rect -3087 4360 -3057 4386
rect -1036 4360 -1006 4386
rect -944 4360 -914 4391
rect -848 4360 -818 4391
rect -752 4360 -722 4391
rect -656 4360 -626 4391
rect -560 4360 -530 4391
rect -464 4360 -434 4391
rect -368 4360 -338 4391
rect -272 4360 -242 4391
rect -176 4360 -146 4391
rect -80 4360 -50 4391
rect 16 4360 46 4391
rect 112 4360 142 4391
rect 204 4360 234 4386
rect 5561 3863 5627 3879
rect -24072 3779 -24042 3810
rect -23980 3779 -23950 3810
rect -23884 3779 -23854 3810
rect -23788 3779 -23758 3810
rect -24072 3622 -23758 3779
rect -23692 3779 -23662 3810
rect -23596 3779 -23566 3810
rect -23500 3779 -23470 3810
rect -23692 3746 -23470 3779
rect -23692 3701 -23673 3746
rect -23543 3701 -23470 3746
rect -23692 3686 -23470 3701
rect -23404 3780 -23374 3810
rect -23308 3780 -23278 3810
rect -23212 3780 -23182 3810
rect -23404 3751 -23182 3780
rect -23116 3779 -23086 3810
rect -23020 3779 -22990 3810
rect -22924 3779 -22894 3810
rect -22832 3779 -22802 3810
rect -22712 3779 -22461 3784
rect -23404 3706 -23342 3751
rect -23212 3706 -23182 3751
rect -23404 3687 -23182 3706
rect -23118 3767 -22461 3779
rect -23118 3629 -22680 3767
rect -24072 3567 -23855 3622
rect -23790 3567 -23758 3622
rect -24072 3342 -23758 3567
rect -24072 3320 -24042 3342
rect -23980 3320 -23950 3342
rect -23884 3320 -23854 3342
rect -23788 3320 -23758 3342
rect -23692 3547 -22680 3629
rect -22488 3547 -22461 3767
rect -23692 3521 -22461 3547
rect -20781 3779 -20751 3810
rect -20689 3779 -20659 3810
rect -20593 3779 -20563 3810
rect -20497 3779 -20467 3810
rect -20781 3622 -20467 3779
rect -20401 3779 -20371 3810
rect -20305 3779 -20275 3810
rect -20209 3779 -20179 3810
rect -20401 3746 -20179 3779
rect -20401 3701 -20382 3746
rect -20252 3701 -20179 3746
rect -20401 3686 -20179 3701
rect -20113 3780 -20083 3810
rect -20017 3780 -19987 3810
rect -19921 3780 -19891 3810
rect -20113 3751 -19891 3780
rect -19825 3779 -19795 3810
rect -19729 3779 -19699 3810
rect -19633 3779 -19603 3810
rect -19541 3779 -19511 3810
rect -19421 3779 -19170 3784
rect -20113 3706 -20051 3751
rect -19921 3706 -19891 3751
rect -20113 3687 -19891 3706
rect -19827 3767 -19170 3779
rect -19827 3629 -19389 3767
rect -20781 3567 -20564 3622
rect -20499 3567 -20467 3622
rect -23692 3520 -22471 3521
rect -23692 3342 -23470 3520
rect -23692 3320 -23662 3342
rect -23596 3320 -23566 3342
rect -23500 3320 -23470 3342
rect -23404 3422 -23182 3450
rect -23404 3377 -23350 3422
rect -23220 3377 -23182 3422
rect -23404 3342 -23182 3377
rect -23404 3320 -23374 3342
rect -23308 3320 -23278 3342
rect -23212 3320 -23182 3342
rect -23116 3430 -22894 3455
rect -23116 3385 -23067 3430
rect -22937 3385 -22894 3430
rect -23116 3342 -22894 3385
rect -22845 3345 -22769 3520
rect -23116 3320 -23086 3342
rect -23020 3320 -22990 3342
rect -22924 3320 -22894 3342
rect -22832 3320 -22802 3345
rect -20781 3342 -20467 3567
rect -20781 3320 -20751 3342
rect -20689 3320 -20659 3342
rect -20593 3320 -20563 3342
rect -20497 3320 -20467 3342
rect -20401 3547 -19389 3629
rect -19197 3547 -19170 3767
rect -20401 3521 -19170 3547
rect -17490 3779 -17460 3810
rect -17398 3779 -17368 3810
rect -17302 3779 -17272 3810
rect -17206 3779 -17176 3810
rect -17490 3622 -17176 3779
rect -17110 3779 -17080 3810
rect -17014 3779 -16984 3810
rect -16918 3779 -16888 3810
rect -17110 3746 -16888 3779
rect -17110 3701 -17091 3746
rect -16961 3701 -16888 3746
rect -17110 3686 -16888 3701
rect -16822 3780 -16792 3810
rect -16726 3780 -16696 3810
rect -16630 3780 -16600 3810
rect -16822 3751 -16600 3780
rect -16534 3779 -16504 3810
rect -16438 3779 -16408 3810
rect -16342 3779 -16312 3810
rect -16250 3779 -16220 3810
rect -16130 3779 -15879 3784
rect -16822 3706 -16760 3751
rect -16630 3706 -16600 3751
rect -16822 3687 -16600 3706
rect -16536 3767 -15879 3779
rect -16536 3629 -16098 3767
rect -17490 3567 -17273 3622
rect -17208 3567 -17176 3622
rect -20401 3520 -19180 3521
rect -20401 3342 -20179 3520
rect -20401 3320 -20371 3342
rect -20305 3320 -20275 3342
rect -20209 3320 -20179 3342
rect -20113 3422 -19891 3450
rect -20113 3377 -20059 3422
rect -19929 3377 -19891 3422
rect -20113 3342 -19891 3377
rect -20113 3320 -20083 3342
rect -20017 3320 -19987 3342
rect -19921 3320 -19891 3342
rect -19825 3430 -19603 3455
rect -19825 3385 -19776 3430
rect -19646 3385 -19603 3430
rect -19825 3342 -19603 3385
rect -19554 3345 -19478 3520
rect -19825 3320 -19795 3342
rect -19729 3320 -19699 3342
rect -19633 3320 -19603 3342
rect -19541 3320 -19511 3345
rect -17490 3342 -17176 3567
rect -17490 3320 -17460 3342
rect -17398 3320 -17368 3342
rect -17302 3320 -17272 3342
rect -17206 3320 -17176 3342
rect -17110 3547 -16098 3629
rect -15906 3547 -15879 3767
rect -17110 3521 -15879 3547
rect -14199 3779 -14169 3810
rect -14107 3779 -14077 3810
rect -14011 3779 -13981 3810
rect -13915 3779 -13885 3810
rect -14199 3622 -13885 3779
rect -13819 3779 -13789 3810
rect -13723 3779 -13693 3810
rect -13627 3779 -13597 3810
rect -13819 3746 -13597 3779
rect -13819 3701 -13800 3746
rect -13670 3701 -13597 3746
rect -13819 3686 -13597 3701
rect -13531 3780 -13501 3810
rect -13435 3780 -13405 3810
rect -13339 3780 -13309 3810
rect -13531 3751 -13309 3780
rect -13243 3779 -13213 3810
rect -13147 3779 -13117 3810
rect -13051 3779 -13021 3810
rect -12959 3779 -12929 3810
rect -12839 3779 -12588 3784
rect -13531 3706 -13469 3751
rect -13339 3706 -13309 3751
rect -13531 3687 -13309 3706
rect -13245 3767 -12588 3779
rect -13245 3629 -12807 3767
rect -14199 3567 -13982 3622
rect -13917 3567 -13885 3622
rect -17110 3520 -15889 3521
rect -17110 3342 -16888 3520
rect -17110 3320 -17080 3342
rect -17014 3320 -16984 3342
rect -16918 3320 -16888 3342
rect -16822 3422 -16600 3450
rect -16822 3377 -16768 3422
rect -16638 3377 -16600 3422
rect -16822 3342 -16600 3377
rect -16822 3320 -16792 3342
rect -16726 3320 -16696 3342
rect -16630 3320 -16600 3342
rect -16534 3430 -16312 3455
rect -16534 3385 -16485 3430
rect -16355 3385 -16312 3430
rect -16534 3342 -16312 3385
rect -16263 3345 -16187 3520
rect -16534 3320 -16504 3342
rect -16438 3320 -16408 3342
rect -16342 3320 -16312 3342
rect -16250 3320 -16220 3345
rect -14199 3342 -13885 3567
rect -14199 3320 -14169 3342
rect -14107 3320 -14077 3342
rect -14011 3320 -13981 3342
rect -13915 3320 -13885 3342
rect -13819 3547 -12807 3629
rect -12615 3547 -12588 3767
rect -13819 3521 -12588 3547
rect -10908 3779 -10878 3810
rect -10816 3779 -10786 3810
rect -10720 3779 -10690 3810
rect -10624 3779 -10594 3810
rect -10908 3622 -10594 3779
rect -10528 3779 -10498 3810
rect -10432 3779 -10402 3810
rect -10336 3779 -10306 3810
rect -10528 3746 -10306 3779
rect -10528 3701 -10509 3746
rect -10379 3701 -10306 3746
rect -10528 3686 -10306 3701
rect -10240 3780 -10210 3810
rect -10144 3780 -10114 3810
rect -10048 3780 -10018 3810
rect -10240 3751 -10018 3780
rect -9952 3779 -9922 3810
rect -9856 3779 -9826 3810
rect -9760 3779 -9730 3810
rect -9668 3779 -9638 3810
rect -9548 3779 -9297 3784
rect -10240 3706 -10178 3751
rect -10048 3706 -10018 3751
rect -10240 3687 -10018 3706
rect -9954 3767 -9297 3779
rect -9954 3629 -9516 3767
rect -10908 3567 -10691 3622
rect -10626 3567 -10594 3622
rect -13819 3520 -12598 3521
rect -13819 3342 -13597 3520
rect -13819 3320 -13789 3342
rect -13723 3320 -13693 3342
rect -13627 3320 -13597 3342
rect -13531 3422 -13309 3450
rect -13531 3377 -13477 3422
rect -13347 3377 -13309 3422
rect -13531 3342 -13309 3377
rect -13531 3320 -13501 3342
rect -13435 3320 -13405 3342
rect -13339 3320 -13309 3342
rect -13243 3430 -13021 3455
rect -13243 3385 -13194 3430
rect -13064 3385 -13021 3430
rect -13243 3342 -13021 3385
rect -12972 3345 -12896 3520
rect -13243 3320 -13213 3342
rect -13147 3320 -13117 3342
rect -13051 3320 -13021 3342
rect -12959 3320 -12929 3345
rect -10908 3342 -10594 3567
rect -10908 3320 -10878 3342
rect -10816 3320 -10786 3342
rect -10720 3320 -10690 3342
rect -10624 3320 -10594 3342
rect -10528 3547 -9516 3629
rect -9324 3547 -9297 3767
rect -10528 3521 -9297 3547
rect -7618 3779 -7588 3810
rect -7526 3779 -7496 3810
rect -7430 3779 -7400 3810
rect -7334 3779 -7304 3810
rect -7618 3622 -7304 3779
rect -7238 3779 -7208 3810
rect -7142 3779 -7112 3810
rect -7046 3779 -7016 3810
rect -7238 3746 -7016 3779
rect -7238 3701 -7219 3746
rect -7089 3701 -7016 3746
rect -7238 3686 -7016 3701
rect -6950 3780 -6920 3810
rect -6854 3780 -6824 3810
rect -6758 3780 -6728 3810
rect -6950 3751 -6728 3780
rect -6662 3779 -6632 3810
rect -6566 3779 -6536 3810
rect -6470 3779 -6440 3810
rect -6378 3779 -6348 3810
rect -6258 3779 -6007 3784
rect -6950 3706 -6888 3751
rect -6758 3706 -6728 3751
rect -6950 3687 -6728 3706
rect -6664 3767 -6007 3779
rect -6664 3629 -6226 3767
rect -7618 3567 -7401 3622
rect -7336 3567 -7304 3622
rect -10528 3520 -9307 3521
rect -10528 3342 -10306 3520
rect -10528 3320 -10498 3342
rect -10432 3320 -10402 3342
rect -10336 3320 -10306 3342
rect -10240 3422 -10018 3450
rect -10240 3377 -10186 3422
rect -10056 3377 -10018 3422
rect -10240 3342 -10018 3377
rect -10240 3320 -10210 3342
rect -10144 3320 -10114 3342
rect -10048 3320 -10018 3342
rect -9952 3430 -9730 3455
rect -9952 3385 -9903 3430
rect -9773 3385 -9730 3430
rect -9952 3342 -9730 3385
rect -9681 3345 -9605 3520
rect -9952 3320 -9922 3342
rect -9856 3320 -9826 3342
rect -9760 3320 -9730 3342
rect -9668 3320 -9638 3345
rect -7618 3342 -7304 3567
rect -7618 3320 -7588 3342
rect -7526 3320 -7496 3342
rect -7430 3320 -7400 3342
rect -7334 3320 -7304 3342
rect -7238 3547 -6226 3629
rect -6034 3547 -6007 3767
rect -7238 3521 -6007 3547
rect -4327 3779 -4297 3810
rect -4235 3779 -4205 3810
rect -4139 3779 -4109 3810
rect -4043 3779 -4013 3810
rect -4327 3622 -4013 3779
rect -3947 3779 -3917 3810
rect -3851 3779 -3821 3810
rect -3755 3779 -3725 3810
rect -3947 3746 -3725 3779
rect -3947 3701 -3928 3746
rect -3798 3701 -3725 3746
rect -3947 3686 -3725 3701
rect -3659 3780 -3629 3810
rect -3563 3780 -3533 3810
rect -3467 3780 -3437 3810
rect -3659 3751 -3437 3780
rect -3371 3779 -3341 3810
rect -3275 3779 -3245 3810
rect -3179 3779 -3149 3810
rect -3087 3779 -3057 3810
rect -2967 3779 -2716 3784
rect -3659 3706 -3597 3751
rect -3467 3706 -3437 3751
rect -3659 3687 -3437 3706
rect -3373 3767 -2716 3779
rect -3373 3629 -2935 3767
rect -4327 3567 -4110 3622
rect -4045 3567 -4013 3622
rect -7238 3520 -6017 3521
rect -7238 3342 -7016 3520
rect -7238 3320 -7208 3342
rect -7142 3320 -7112 3342
rect -7046 3320 -7016 3342
rect -6950 3422 -6728 3450
rect -6950 3377 -6896 3422
rect -6766 3377 -6728 3422
rect -6950 3342 -6728 3377
rect -6950 3320 -6920 3342
rect -6854 3320 -6824 3342
rect -6758 3320 -6728 3342
rect -6662 3430 -6440 3455
rect -6662 3385 -6613 3430
rect -6483 3385 -6440 3430
rect -6662 3342 -6440 3385
rect -6391 3345 -6315 3520
rect -6662 3320 -6632 3342
rect -6566 3320 -6536 3342
rect -6470 3320 -6440 3342
rect -6378 3320 -6348 3345
rect -4327 3342 -4013 3567
rect -4327 3320 -4297 3342
rect -4235 3320 -4205 3342
rect -4139 3320 -4109 3342
rect -4043 3320 -4013 3342
rect -3947 3547 -2935 3629
rect -2743 3547 -2716 3767
rect -3947 3521 -2716 3547
rect -1036 3779 -1006 3810
rect -944 3779 -914 3810
rect -848 3779 -818 3810
rect -752 3779 -722 3810
rect -1036 3622 -722 3779
rect -656 3779 -626 3810
rect -560 3779 -530 3810
rect -464 3779 -434 3810
rect -656 3746 -434 3779
rect -656 3701 -637 3746
rect -507 3701 -434 3746
rect -656 3686 -434 3701
rect -368 3780 -338 3810
rect -272 3780 -242 3810
rect -176 3780 -146 3810
rect -368 3751 -146 3780
rect -80 3779 -50 3810
rect 16 3779 46 3810
rect 112 3779 142 3810
rect 204 3779 234 3810
rect 324 3779 575 3784
rect -368 3706 -306 3751
rect -176 3706 -146 3751
rect -368 3687 -146 3706
rect -82 3767 575 3779
rect -82 3629 356 3767
rect -1036 3567 -819 3622
rect -754 3567 -722 3622
rect -3947 3520 -2726 3521
rect -3947 3342 -3725 3520
rect -3947 3320 -3917 3342
rect -3851 3320 -3821 3342
rect -3755 3320 -3725 3342
rect -3659 3422 -3437 3450
rect -3659 3377 -3605 3422
rect -3475 3377 -3437 3422
rect -3659 3342 -3437 3377
rect -3659 3320 -3629 3342
rect -3563 3320 -3533 3342
rect -3467 3320 -3437 3342
rect -3371 3430 -3149 3455
rect -3371 3385 -3322 3430
rect -3192 3385 -3149 3430
rect -3371 3342 -3149 3385
rect -3100 3345 -3024 3520
rect -3371 3320 -3341 3342
rect -3275 3320 -3245 3342
rect -3179 3320 -3149 3342
rect -3087 3320 -3057 3345
rect -1036 3342 -722 3567
rect -1036 3320 -1006 3342
rect -944 3320 -914 3342
rect -848 3320 -818 3342
rect -752 3320 -722 3342
rect -656 3547 356 3629
rect 548 3547 575 3767
rect 5561 3637 5577 3863
rect 5611 3861 5627 3863
rect 6001 3863 6067 3879
rect 5611 3831 5658 3861
rect 5872 3831 5898 3861
rect 5611 3765 5627 3831
rect 5611 3735 5658 3765
rect 5872 3735 5898 3765
rect 5611 3669 5627 3735
rect 5611 3639 5658 3669
rect 5872 3639 5898 3669
rect 5611 3637 5627 3639
rect 5561 3621 5627 3637
rect 6001 3637 6017 3863
rect 6051 3861 6067 3863
rect 6441 3863 6507 3879
rect 6051 3831 6098 3861
rect 6312 3831 6338 3861
rect 6051 3765 6067 3831
rect 6051 3735 6098 3765
rect 6312 3735 6338 3765
rect 6051 3669 6067 3735
rect 6051 3639 6098 3669
rect 6312 3639 6338 3669
rect 6051 3637 6067 3639
rect 6001 3621 6067 3637
rect 6441 3637 6457 3863
rect 6491 3861 6507 3863
rect 6491 3831 6538 3861
rect 6752 3831 6778 3861
rect 6491 3765 6507 3831
rect 6491 3735 6538 3765
rect 6752 3735 6778 3765
rect 6491 3669 6507 3735
rect 6491 3639 6538 3669
rect 6752 3639 6778 3669
rect 6491 3637 6507 3639
rect 6441 3621 6507 3637
rect -656 3521 575 3547
rect -656 3520 565 3521
rect -656 3342 -434 3520
rect -656 3320 -626 3342
rect -560 3320 -530 3342
rect -464 3320 -434 3342
rect -368 3422 -146 3450
rect -368 3377 -314 3422
rect -184 3377 -146 3422
rect -368 3342 -146 3377
rect -368 3320 -338 3342
rect -272 3320 -242 3342
rect -176 3320 -146 3342
rect -80 3430 142 3455
rect -80 3385 -31 3430
rect 99 3385 142 3430
rect -80 3342 142 3385
rect 191 3345 267 3520
rect 5561 3417 5628 3433
rect 5561 3383 5577 3417
rect 5611 3415 5628 3417
rect 6001 3417 6068 3433
rect 5611 3385 5658 3415
rect 5858 3385 5884 3415
rect 5611 3383 5628 3385
rect 5561 3367 5628 3383
rect -80 3320 -50 3342
rect 16 3320 46 3342
rect 112 3320 142 3342
rect 204 3320 234 3345
rect 6001 3383 6017 3417
rect 6051 3415 6068 3417
rect 6441 3417 6508 3433
rect 6051 3385 6098 3415
rect 6298 3385 6324 3415
rect 6051 3383 6068 3385
rect 6001 3367 6068 3383
rect 6441 3383 6457 3417
rect 6491 3415 6508 3417
rect 6491 3385 6538 3415
rect 6738 3385 6764 3415
rect 6491 3383 6508 3385
rect 6441 3367 6508 3383
rect 7200 3219 7230 3245
rect 7296 3219 7326 3245
rect 7392 3219 7422 3245
rect 7488 3219 7518 3245
rect 7584 3219 7614 3245
rect 7680 3219 7710 3245
rect 7776 3219 7806 3245
rect 7872 3219 7902 3245
rect 8148 3219 8178 3245
rect 8244 3219 8274 3245
rect 8340 3219 8370 3245
rect 8436 3219 8466 3245
rect 8532 3219 8562 3245
rect 8628 3219 8658 3245
rect 8724 3219 8754 3245
rect 8820 3219 8850 3245
rect 9084 3219 9114 3245
rect 9180 3219 9210 3245
rect 9276 3219 9306 3245
rect 9372 3219 9402 3245
rect 9468 3219 9498 3245
rect 9564 3219 9594 3245
rect 9660 3219 9690 3245
rect 9756 3219 9786 3245
rect 10015 3219 10045 3245
rect 10111 3219 10141 3245
rect 10207 3219 10237 3245
rect 10303 3219 10333 3245
rect 10399 3219 10429 3245
rect 10495 3219 10525 3245
rect 10591 3219 10621 3245
rect 10687 3219 10717 3245
rect 10942 3219 10972 3245
rect 11038 3219 11068 3245
rect 11134 3219 11164 3245
rect 11230 3219 11260 3245
rect 11326 3219 11356 3245
rect 11422 3219 11452 3245
rect 11518 3219 11548 3245
rect 11614 3219 11644 3245
rect -24072 3164 -24042 3190
rect -23980 3164 -23950 3190
rect -23884 3164 -23854 3190
rect -23788 3164 -23758 3190
rect -23692 3164 -23662 3190
rect -23596 3164 -23566 3190
rect -23500 3164 -23470 3190
rect -23404 3164 -23374 3190
rect -23308 3164 -23278 3190
rect -23212 3164 -23182 3190
rect -23116 3164 -23086 3190
rect -23020 3164 -22990 3190
rect -22924 3164 -22894 3190
rect -22832 3164 -22802 3190
rect -20781 3164 -20751 3190
rect -20689 3164 -20659 3190
rect -20593 3164 -20563 3190
rect -20497 3164 -20467 3190
rect -20401 3164 -20371 3190
rect -20305 3164 -20275 3190
rect -20209 3164 -20179 3190
rect -20113 3164 -20083 3190
rect -20017 3164 -19987 3190
rect -19921 3164 -19891 3190
rect -19825 3164 -19795 3190
rect -19729 3164 -19699 3190
rect -19633 3164 -19603 3190
rect -19541 3164 -19511 3190
rect -17490 3164 -17460 3190
rect -17398 3164 -17368 3190
rect -17302 3164 -17272 3190
rect -17206 3164 -17176 3190
rect -17110 3164 -17080 3190
rect -17014 3164 -16984 3190
rect -16918 3164 -16888 3190
rect -16822 3164 -16792 3190
rect -16726 3164 -16696 3190
rect -16630 3164 -16600 3190
rect -16534 3164 -16504 3190
rect -16438 3164 -16408 3190
rect -16342 3164 -16312 3190
rect -16250 3164 -16220 3190
rect -14199 3164 -14169 3190
rect -14107 3164 -14077 3190
rect -14011 3164 -13981 3190
rect -13915 3164 -13885 3190
rect -13819 3164 -13789 3190
rect -13723 3164 -13693 3190
rect -13627 3164 -13597 3190
rect -13531 3164 -13501 3190
rect -13435 3164 -13405 3190
rect -13339 3164 -13309 3190
rect -13243 3164 -13213 3190
rect -13147 3164 -13117 3190
rect -13051 3164 -13021 3190
rect -12959 3164 -12929 3190
rect -10908 3164 -10878 3190
rect -10816 3164 -10786 3190
rect -10720 3164 -10690 3190
rect -10624 3164 -10594 3190
rect -10528 3164 -10498 3190
rect -10432 3164 -10402 3190
rect -10336 3164 -10306 3190
rect -10240 3164 -10210 3190
rect -10144 3164 -10114 3190
rect -10048 3164 -10018 3190
rect -9952 3164 -9922 3190
rect -9856 3164 -9826 3190
rect -9760 3164 -9730 3190
rect -9668 3164 -9638 3190
rect -7618 3164 -7588 3190
rect -7526 3164 -7496 3190
rect -7430 3164 -7400 3190
rect -7334 3164 -7304 3190
rect -7238 3164 -7208 3190
rect -7142 3164 -7112 3190
rect -7046 3164 -7016 3190
rect -6950 3164 -6920 3190
rect -6854 3164 -6824 3190
rect -6758 3164 -6728 3190
rect -6662 3164 -6632 3190
rect -6566 3164 -6536 3190
rect -6470 3164 -6440 3190
rect -6378 3164 -6348 3190
rect -4327 3164 -4297 3190
rect -4235 3164 -4205 3190
rect -4139 3164 -4109 3190
rect -4043 3164 -4013 3190
rect -3947 3164 -3917 3190
rect -3851 3164 -3821 3190
rect -3755 3164 -3725 3190
rect -3659 3164 -3629 3190
rect -3563 3164 -3533 3190
rect -3467 3164 -3437 3190
rect -3371 3164 -3341 3190
rect -3275 3164 -3245 3190
rect -3179 3164 -3149 3190
rect -3087 3164 -3057 3190
rect -1036 3164 -1006 3190
rect -944 3164 -914 3190
rect -848 3164 -818 3190
rect -752 3164 -722 3190
rect -656 3164 -626 3190
rect -560 3164 -530 3190
rect -464 3164 -434 3190
rect -368 3164 -338 3190
rect -272 3164 -242 3190
rect -176 3164 -146 3190
rect -80 3164 -50 3190
rect 16 3164 46 3190
rect 112 3164 142 3190
rect 204 3164 234 3190
rect 7200 2866 7230 2897
rect 7296 2866 7326 2897
rect 7392 2866 7422 2897
rect 7488 2866 7518 2897
rect 7584 2866 7614 2897
rect 7680 2866 7710 2897
rect 7776 2866 7806 2897
rect 7872 2866 7902 2897
rect 8148 2866 8178 2897
rect 8244 2866 8274 2897
rect 8340 2866 8370 2897
rect 8436 2866 8466 2897
rect 8532 2866 8562 2897
rect 8628 2866 8658 2897
rect 8724 2866 8754 2897
rect 8820 2866 8850 2897
rect 9084 2866 9114 2897
rect 9180 2866 9210 2897
rect 9276 2866 9306 2897
rect 9372 2866 9402 2897
rect 9468 2866 9498 2897
rect 9564 2866 9594 2897
rect 9660 2866 9690 2897
rect 9756 2866 9786 2897
rect 10015 2866 10045 2897
rect 10111 2866 10141 2897
rect 10207 2866 10237 2897
rect 10303 2866 10333 2897
rect 10399 2866 10429 2897
rect 10495 2866 10525 2897
rect 10591 2866 10621 2897
rect 10687 2866 10717 2897
rect 10942 2866 10972 2897
rect 11038 2866 11068 2897
rect 11134 2866 11164 2897
rect 11230 2866 11260 2897
rect 11326 2866 11356 2897
rect 11422 2866 11452 2897
rect 11518 2866 11548 2897
rect 11614 2866 11644 2897
rect 7182 2850 7326 2866
rect 7182 2816 7198 2850
rect 7232 2816 7326 2850
rect 7182 2800 7326 2816
rect 7374 2850 7518 2866
rect 7374 2816 7390 2850
rect 7424 2816 7518 2850
rect -24746 2576 -24716 2602
rect -24654 2576 -24624 2607
rect -24558 2576 -24528 2607
rect -24462 2576 -24432 2607
rect -24366 2576 -24336 2607
rect -24270 2576 -24240 2607
rect -24174 2576 -24144 2607
rect -24078 2576 -24048 2607
rect -23982 2576 -23952 2607
rect -23886 2576 -23856 2607
rect -23790 2576 -23760 2607
rect -23694 2576 -23664 2607
rect -23598 2576 -23568 2607
rect -23506 2576 -23476 2602
rect -23187 2576 -23157 2602
rect -23095 2576 -23065 2607
rect -22999 2576 -22969 2607
rect -22903 2576 -22873 2607
rect -22807 2576 -22777 2607
rect -22711 2576 -22681 2607
rect -22615 2576 -22585 2607
rect -22519 2576 -22489 2607
rect -22423 2576 -22393 2607
rect -22327 2576 -22297 2607
rect -22231 2576 -22201 2607
rect -22135 2576 -22105 2607
rect -22039 2576 -22009 2607
rect -21947 2576 -21917 2602
rect -21455 2576 -21425 2602
rect -21363 2576 -21333 2607
rect -21267 2576 -21237 2607
rect -21171 2576 -21141 2607
rect -21075 2576 -21045 2607
rect -20979 2576 -20949 2607
rect -20883 2576 -20853 2607
rect -20787 2576 -20757 2607
rect -20691 2576 -20661 2607
rect -20595 2576 -20565 2607
rect -20499 2576 -20469 2607
rect -20403 2576 -20373 2607
rect -20307 2576 -20277 2607
rect -20215 2576 -20185 2602
rect -19896 2576 -19866 2602
rect -19804 2576 -19774 2607
rect -19708 2576 -19678 2607
rect -19612 2576 -19582 2607
rect -19516 2576 -19486 2607
rect -19420 2576 -19390 2607
rect -19324 2576 -19294 2607
rect -19228 2576 -19198 2607
rect -19132 2576 -19102 2607
rect -19036 2576 -19006 2607
rect -18940 2576 -18910 2607
rect -18844 2576 -18814 2607
rect -18748 2576 -18718 2607
rect -18656 2576 -18626 2602
rect -18164 2576 -18134 2602
rect -18072 2576 -18042 2607
rect -17976 2576 -17946 2607
rect -17880 2576 -17850 2607
rect -17784 2576 -17754 2607
rect -17688 2576 -17658 2607
rect -17592 2576 -17562 2607
rect -17496 2576 -17466 2607
rect -17400 2576 -17370 2607
rect -17304 2576 -17274 2607
rect -17208 2576 -17178 2607
rect -17112 2576 -17082 2607
rect -17016 2576 -16986 2607
rect -16924 2576 -16894 2602
rect -16605 2576 -16575 2602
rect -16513 2576 -16483 2607
rect -16417 2576 -16387 2607
rect -16321 2576 -16291 2607
rect -16225 2576 -16195 2607
rect -16129 2576 -16099 2607
rect -16033 2576 -16003 2607
rect -15937 2576 -15907 2607
rect -15841 2576 -15811 2607
rect -15745 2576 -15715 2607
rect -15649 2576 -15619 2607
rect -15553 2576 -15523 2607
rect -15457 2576 -15427 2607
rect -15365 2576 -15335 2602
rect -14873 2576 -14843 2602
rect -14781 2576 -14751 2607
rect -14685 2576 -14655 2607
rect -14589 2576 -14559 2607
rect -14493 2576 -14463 2607
rect -14397 2576 -14367 2607
rect -14301 2576 -14271 2607
rect -14205 2576 -14175 2607
rect -14109 2576 -14079 2607
rect -14013 2576 -13983 2607
rect -13917 2576 -13887 2607
rect -13821 2576 -13791 2607
rect -13725 2576 -13695 2607
rect -13633 2576 -13603 2602
rect -13314 2576 -13284 2602
rect -13222 2576 -13192 2607
rect -13126 2576 -13096 2607
rect -13030 2576 -13000 2607
rect -12934 2576 -12904 2607
rect -12838 2576 -12808 2607
rect -12742 2576 -12712 2607
rect -12646 2576 -12616 2607
rect -12550 2576 -12520 2607
rect -12454 2576 -12424 2607
rect -12358 2576 -12328 2607
rect -12262 2576 -12232 2607
rect -12166 2576 -12136 2607
rect -12074 2576 -12044 2602
rect -11582 2576 -11552 2602
rect -11490 2576 -11460 2607
rect -11394 2576 -11364 2607
rect -11298 2576 -11268 2607
rect -11202 2576 -11172 2607
rect -11106 2576 -11076 2607
rect -11010 2576 -10980 2607
rect -10914 2576 -10884 2607
rect -10818 2576 -10788 2607
rect -10722 2576 -10692 2607
rect -10626 2576 -10596 2607
rect -10530 2576 -10500 2607
rect -10434 2576 -10404 2607
rect -10342 2576 -10312 2602
rect -10023 2576 -9993 2602
rect -9931 2576 -9901 2607
rect -9835 2576 -9805 2607
rect -9739 2576 -9709 2607
rect -9643 2576 -9613 2607
rect -9547 2576 -9517 2607
rect -9451 2576 -9421 2607
rect -9355 2576 -9325 2607
rect -9259 2576 -9229 2607
rect -9163 2576 -9133 2607
rect -9067 2576 -9037 2607
rect -8971 2576 -8941 2607
rect -8875 2576 -8845 2607
rect -8783 2576 -8753 2602
rect -8292 2576 -8262 2602
rect -8200 2576 -8170 2607
rect -8104 2576 -8074 2607
rect -8008 2576 -7978 2607
rect -7912 2576 -7882 2607
rect -7816 2576 -7786 2607
rect -7720 2576 -7690 2607
rect -7624 2576 -7594 2607
rect -7528 2576 -7498 2607
rect -7432 2576 -7402 2607
rect -7336 2576 -7306 2607
rect -7240 2576 -7210 2607
rect -7144 2576 -7114 2607
rect -7052 2576 -7022 2602
rect -6733 2576 -6703 2602
rect -6641 2576 -6611 2607
rect -6545 2576 -6515 2607
rect -6449 2576 -6419 2607
rect -6353 2576 -6323 2607
rect -6257 2576 -6227 2607
rect -6161 2576 -6131 2607
rect -6065 2576 -6035 2607
rect -5969 2576 -5939 2607
rect -5873 2576 -5843 2607
rect -5777 2576 -5747 2607
rect -5681 2576 -5651 2607
rect -5585 2576 -5555 2607
rect -5493 2576 -5463 2602
rect -5001 2576 -4971 2602
rect -4909 2576 -4879 2607
rect -4813 2576 -4783 2607
rect -4717 2576 -4687 2607
rect -4621 2576 -4591 2607
rect -4525 2576 -4495 2607
rect -4429 2576 -4399 2607
rect -4333 2576 -4303 2607
rect -4237 2576 -4207 2607
rect -4141 2576 -4111 2607
rect -4045 2576 -4015 2607
rect -3949 2576 -3919 2607
rect -3853 2576 -3823 2607
rect -3761 2576 -3731 2602
rect -3442 2576 -3412 2602
rect -3350 2576 -3320 2607
rect -3254 2576 -3224 2607
rect -3158 2576 -3128 2607
rect -3062 2576 -3032 2607
rect -2966 2576 -2936 2607
rect -2870 2576 -2840 2607
rect -2774 2576 -2744 2607
rect -2678 2576 -2648 2607
rect -2582 2576 -2552 2607
rect -2486 2576 -2456 2607
rect -2390 2576 -2360 2607
rect -2294 2576 -2264 2607
rect -2202 2576 -2172 2602
rect -1710 2576 -1680 2602
rect -1618 2576 -1588 2607
rect -1522 2576 -1492 2607
rect -1426 2576 -1396 2607
rect -1330 2576 -1300 2607
rect -1234 2576 -1204 2607
rect -1138 2576 -1108 2607
rect -1042 2576 -1012 2607
rect -946 2576 -916 2607
rect -850 2576 -820 2607
rect -754 2576 -724 2607
rect -658 2576 -628 2607
rect -562 2576 -532 2607
rect -470 2576 -440 2602
rect -151 2576 -121 2602
rect -59 2576 -29 2607
rect 37 2576 67 2607
rect 133 2576 163 2607
rect 229 2576 259 2607
rect 325 2576 355 2607
rect 421 2576 451 2607
rect 517 2576 547 2607
rect 613 2576 643 2607
rect 709 2576 739 2607
rect 805 2576 835 2607
rect 901 2576 931 2607
rect 997 2576 1027 2607
rect 1089 2576 1119 2602
rect 7238 2553 7268 2800
rect 7374 2733 7518 2816
rect 7566 2850 7710 2866
rect 7566 2816 7582 2850
rect 7616 2816 7710 2850
rect 7566 2800 7710 2816
rect 7758 2850 7902 2866
rect 7758 2816 7774 2850
rect 7808 2816 7902 2850
rect 7758 2800 7902 2816
rect 8130 2850 8274 2866
rect 8130 2816 8146 2850
rect 8180 2816 8274 2850
rect 8130 2800 8274 2816
rect 8322 2850 8466 2866
rect 8322 2816 8338 2850
rect 8372 2816 8466 2850
rect 7584 2775 7644 2800
rect 7374 2595 7548 2733
rect 7238 2523 7452 2553
rect 7422 2490 7452 2523
rect 7518 2490 7548 2595
rect 7590 2513 7644 2775
rect 7758 2670 7848 2800
rect 7614 2490 7644 2513
rect 7710 2640 7848 2670
rect 7710 2490 7740 2640
rect 8186 2553 8216 2800
rect 8322 2733 8466 2816
rect 8514 2850 8658 2866
rect 8514 2816 8530 2850
rect 8564 2816 8658 2850
rect 8514 2800 8658 2816
rect 8706 2850 8850 2866
rect 8706 2816 8722 2850
rect 8756 2816 8850 2850
rect 8706 2800 8850 2816
rect 9066 2850 9210 2866
rect 9066 2816 9082 2850
rect 9116 2816 9210 2850
rect 9066 2800 9210 2816
rect 9258 2850 9402 2866
rect 9258 2816 9274 2850
rect 9308 2816 9402 2850
rect 8532 2775 8592 2800
rect 8322 2595 8496 2733
rect 8186 2523 8400 2553
rect 8370 2490 8400 2523
rect 8466 2490 8496 2595
rect 8538 2513 8592 2775
rect 8706 2670 8796 2800
rect 8562 2490 8592 2513
rect 8658 2640 8796 2670
rect 8658 2490 8688 2640
rect 9122 2553 9152 2800
rect 9258 2733 9402 2816
rect 9450 2850 9594 2866
rect 9450 2816 9466 2850
rect 9500 2816 9594 2850
rect 9450 2800 9594 2816
rect 9642 2850 9786 2866
rect 9642 2816 9658 2850
rect 9692 2816 9786 2850
rect 9642 2800 9786 2816
rect 9997 2850 10141 2866
rect 9997 2816 10013 2850
rect 10047 2816 10141 2850
rect 9997 2800 10141 2816
rect 10189 2850 10333 2866
rect 10189 2816 10205 2850
rect 10239 2816 10333 2850
rect 9468 2775 9528 2800
rect 9258 2595 9432 2733
rect 9122 2523 9336 2553
rect 9306 2490 9336 2523
rect 9402 2490 9432 2595
rect 9474 2513 9528 2775
rect 9642 2670 9732 2800
rect 9498 2490 9528 2513
rect 9594 2640 9732 2670
rect 9594 2490 9624 2640
rect 10053 2553 10083 2800
rect 10189 2733 10333 2816
rect 10381 2850 10525 2866
rect 10381 2816 10397 2850
rect 10431 2816 10525 2850
rect 10381 2800 10525 2816
rect 10573 2850 10717 2866
rect 10573 2816 10589 2850
rect 10623 2816 10717 2850
rect 10573 2800 10717 2816
rect 10924 2850 11068 2866
rect 10924 2816 10940 2850
rect 10974 2816 11068 2850
rect 10924 2800 11068 2816
rect 11116 2850 11260 2866
rect 11116 2816 11132 2850
rect 11166 2816 11260 2850
rect 10399 2775 10459 2800
rect 10189 2595 10363 2733
rect 10053 2523 10267 2553
rect 10237 2490 10267 2523
rect 10333 2490 10363 2595
rect 10405 2513 10459 2775
rect 10573 2670 10663 2800
rect 10429 2490 10459 2513
rect 10525 2640 10663 2670
rect 10525 2490 10555 2640
rect 10980 2553 11010 2800
rect 11116 2733 11260 2816
rect 11308 2850 11452 2866
rect 11308 2816 11324 2850
rect 11358 2816 11452 2850
rect 11308 2800 11452 2816
rect 11500 2850 11644 2866
rect 11500 2816 11516 2850
rect 11550 2816 11644 2850
rect 11500 2800 11644 2816
rect 11326 2775 11386 2800
rect 11116 2595 11290 2733
rect 10980 2523 11194 2553
rect 11164 2490 11194 2523
rect 11260 2490 11290 2595
rect 11332 2513 11386 2775
rect 11500 2670 11590 2800
rect 11356 2490 11386 2513
rect 11452 2640 11590 2670
rect 11452 2490 11482 2640
rect -24746 1995 -24716 2026
rect -24654 1995 -24624 2026
rect -24558 1995 -24528 2026
rect -24462 1995 -24432 2026
rect -24366 1996 -24336 2026
rect -24270 1996 -24240 2026
rect -24174 1996 -24144 2026
rect -24940 1938 -24430 1995
rect -24940 1828 -24921 1938
rect -24874 1845 -24430 1938
rect -24366 1967 -24144 1996
rect -24366 1922 -24336 1967
rect -24206 1922 -24144 1967
rect -24366 1903 -24144 1922
rect -24078 1995 -24048 2026
rect -23982 1995 -23952 2026
rect -23886 1995 -23856 2026
rect -24078 1962 -23856 1995
rect -24078 1917 -24005 1962
rect -23875 1917 -23856 1962
rect -24078 1902 -23856 1917
rect -23790 1995 -23760 2026
rect -23694 1995 -23664 2026
rect -23598 1995 -23568 2026
rect -23506 1995 -23476 2026
rect -23187 1995 -23157 2026
rect -23095 1995 -23065 2026
rect -22999 1995 -22969 2026
rect -22903 1995 -22873 2026
rect -22807 1996 -22777 2026
rect -22711 1996 -22681 2026
rect -22615 1996 -22585 2026
rect -24874 1828 -23856 1845
rect -24940 1736 -23856 1828
rect -24779 1561 -24703 1736
rect -24654 1646 -24432 1671
rect -24654 1601 -24611 1646
rect -24481 1601 -24432 1646
rect -24746 1536 -24716 1561
rect -24654 1558 -24432 1601
rect -24654 1536 -24624 1558
rect -24558 1536 -24528 1558
rect -24462 1536 -24432 1558
rect -24366 1638 -24144 1666
rect -24366 1593 -24328 1638
rect -24198 1593 -24144 1638
rect -24366 1558 -24144 1593
rect -24366 1536 -24336 1558
rect -24270 1536 -24240 1558
rect -24174 1536 -24144 1558
rect -24078 1558 -23856 1736
rect -24078 1536 -24048 1558
rect -23982 1536 -23952 1558
rect -23886 1536 -23856 1558
rect -23790 1838 -23476 1995
rect -23220 1908 -22871 1995
rect -23790 1783 -23758 1838
rect -23693 1783 -23476 1838
rect -23790 1558 -23476 1783
rect -23409 1893 -22871 1908
rect -22807 1967 -22585 1996
rect -22807 1922 -22777 1967
rect -22647 1922 -22585 1967
rect -22807 1903 -22585 1922
rect -22519 1995 -22489 2026
rect -22423 1995 -22393 2026
rect -22327 1995 -22297 2026
rect -22519 1962 -22297 1995
rect -22519 1917 -22446 1962
rect -22316 1917 -22297 1962
rect -22519 1902 -22297 1917
rect -22231 1995 -22201 2026
rect -22135 1995 -22105 2026
rect -22039 1995 -22009 2026
rect -21947 1995 -21917 2026
rect -21455 1995 -21425 2026
rect -21363 1995 -21333 2026
rect -21267 1995 -21237 2026
rect -21171 1995 -21141 2026
rect -21075 1996 -21045 2026
rect -20979 1996 -20949 2026
rect -20883 1996 -20853 2026
rect -23409 1753 -23364 1893
rect -23291 1845 -22871 1893
rect -23291 1753 -22297 1845
rect -23409 1736 -22297 1753
rect -23220 1561 -23144 1736
rect -23095 1646 -22873 1671
rect -23095 1601 -23052 1646
rect -22922 1601 -22873 1646
rect -23790 1536 -23760 1558
rect -23694 1536 -23664 1558
rect -23598 1536 -23568 1558
rect -23506 1536 -23476 1558
rect -23187 1536 -23157 1561
rect -23095 1558 -22873 1601
rect -23095 1536 -23065 1558
rect -22999 1536 -22969 1558
rect -22903 1536 -22873 1558
rect -22807 1638 -22585 1666
rect -22807 1593 -22769 1638
rect -22639 1593 -22585 1638
rect -22807 1558 -22585 1593
rect -22807 1536 -22777 1558
rect -22711 1536 -22681 1558
rect -22615 1536 -22585 1558
rect -22519 1558 -22297 1736
rect -22519 1536 -22489 1558
rect -22423 1536 -22393 1558
rect -22327 1536 -22297 1558
rect -22231 1838 -21917 1995
rect -22231 1783 -22199 1838
rect -22134 1783 -21917 1838
rect -22231 1558 -21917 1783
rect -21649 1938 -21139 1995
rect -21649 1828 -21630 1938
rect -21583 1845 -21139 1938
rect -21075 1967 -20853 1996
rect -21075 1922 -21045 1967
rect -20915 1922 -20853 1967
rect -21075 1903 -20853 1922
rect -20787 1995 -20757 2026
rect -20691 1995 -20661 2026
rect -20595 1995 -20565 2026
rect -20787 1962 -20565 1995
rect -20787 1917 -20714 1962
rect -20584 1917 -20565 1962
rect -20787 1902 -20565 1917
rect -20499 1995 -20469 2026
rect -20403 1995 -20373 2026
rect -20307 1995 -20277 2026
rect -20215 1995 -20185 2026
rect -19896 1995 -19866 2026
rect -19804 1995 -19774 2026
rect -19708 1995 -19678 2026
rect -19612 1995 -19582 2026
rect -19516 1996 -19486 2026
rect -19420 1996 -19390 2026
rect -19324 1996 -19294 2026
rect -21583 1828 -20565 1845
rect -21649 1736 -20565 1828
rect -21488 1561 -21412 1736
rect -21363 1646 -21141 1671
rect -21363 1601 -21320 1646
rect -21190 1601 -21141 1646
rect -22231 1536 -22201 1558
rect -22135 1536 -22105 1558
rect -22039 1536 -22009 1558
rect -21947 1536 -21917 1558
rect -21455 1536 -21425 1561
rect -21363 1558 -21141 1601
rect -21363 1536 -21333 1558
rect -21267 1536 -21237 1558
rect -21171 1536 -21141 1558
rect -21075 1638 -20853 1666
rect -21075 1593 -21037 1638
rect -20907 1593 -20853 1638
rect -21075 1558 -20853 1593
rect -21075 1536 -21045 1558
rect -20979 1536 -20949 1558
rect -20883 1536 -20853 1558
rect -20787 1558 -20565 1736
rect -20787 1536 -20757 1558
rect -20691 1536 -20661 1558
rect -20595 1536 -20565 1558
rect -20499 1838 -20185 1995
rect -19929 1908 -19580 1995
rect -20499 1783 -20467 1838
rect -20402 1783 -20185 1838
rect -20499 1558 -20185 1783
rect -20118 1893 -19580 1908
rect -19516 1967 -19294 1996
rect -19516 1922 -19486 1967
rect -19356 1922 -19294 1967
rect -19516 1903 -19294 1922
rect -19228 1995 -19198 2026
rect -19132 1995 -19102 2026
rect -19036 1995 -19006 2026
rect -19228 1962 -19006 1995
rect -19228 1917 -19155 1962
rect -19025 1917 -19006 1962
rect -19228 1902 -19006 1917
rect -18940 1995 -18910 2026
rect -18844 1995 -18814 2026
rect -18748 1995 -18718 2026
rect -18656 1995 -18626 2026
rect -18164 1995 -18134 2026
rect -18072 1995 -18042 2026
rect -17976 1995 -17946 2026
rect -17880 1995 -17850 2026
rect -17784 1996 -17754 2026
rect -17688 1996 -17658 2026
rect -17592 1996 -17562 2026
rect -20118 1753 -20073 1893
rect -20000 1845 -19580 1893
rect -20000 1753 -19006 1845
rect -20118 1736 -19006 1753
rect -19929 1561 -19853 1736
rect -19804 1646 -19582 1671
rect -19804 1601 -19761 1646
rect -19631 1601 -19582 1646
rect -20499 1536 -20469 1558
rect -20403 1536 -20373 1558
rect -20307 1536 -20277 1558
rect -20215 1536 -20185 1558
rect -19896 1536 -19866 1561
rect -19804 1558 -19582 1601
rect -19804 1536 -19774 1558
rect -19708 1536 -19678 1558
rect -19612 1536 -19582 1558
rect -19516 1638 -19294 1666
rect -19516 1593 -19478 1638
rect -19348 1593 -19294 1638
rect -19516 1558 -19294 1593
rect -19516 1536 -19486 1558
rect -19420 1536 -19390 1558
rect -19324 1536 -19294 1558
rect -19228 1558 -19006 1736
rect -19228 1536 -19198 1558
rect -19132 1536 -19102 1558
rect -19036 1536 -19006 1558
rect -18940 1838 -18626 1995
rect -18940 1783 -18908 1838
rect -18843 1783 -18626 1838
rect -18940 1558 -18626 1783
rect -18358 1938 -17848 1995
rect -18358 1828 -18339 1938
rect -18292 1845 -17848 1938
rect -17784 1967 -17562 1996
rect -17784 1922 -17754 1967
rect -17624 1922 -17562 1967
rect -17784 1903 -17562 1922
rect -17496 1995 -17466 2026
rect -17400 1995 -17370 2026
rect -17304 1995 -17274 2026
rect -17496 1962 -17274 1995
rect -17496 1917 -17423 1962
rect -17293 1917 -17274 1962
rect -17496 1902 -17274 1917
rect -17208 1995 -17178 2026
rect -17112 1995 -17082 2026
rect -17016 1995 -16986 2026
rect -16924 1995 -16894 2026
rect -16605 1995 -16575 2026
rect -16513 1995 -16483 2026
rect -16417 1995 -16387 2026
rect -16321 1995 -16291 2026
rect -16225 1996 -16195 2026
rect -16129 1996 -16099 2026
rect -16033 1996 -16003 2026
rect -18292 1828 -17274 1845
rect -18358 1736 -17274 1828
rect -18197 1561 -18121 1736
rect -18072 1646 -17850 1671
rect -18072 1601 -18029 1646
rect -17899 1601 -17850 1646
rect -18940 1536 -18910 1558
rect -18844 1536 -18814 1558
rect -18748 1536 -18718 1558
rect -18656 1536 -18626 1558
rect -18164 1536 -18134 1561
rect -18072 1558 -17850 1601
rect -18072 1536 -18042 1558
rect -17976 1536 -17946 1558
rect -17880 1536 -17850 1558
rect -17784 1638 -17562 1666
rect -17784 1593 -17746 1638
rect -17616 1593 -17562 1638
rect -17784 1558 -17562 1593
rect -17784 1536 -17754 1558
rect -17688 1536 -17658 1558
rect -17592 1536 -17562 1558
rect -17496 1558 -17274 1736
rect -17496 1536 -17466 1558
rect -17400 1536 -17370 1558
rect -17304 1536 -17274 1558
rect -17208 1838 -16894 1995
rect -16638 1908 -16289 1995
rect -17208 1783 -17176 1838
rect -17111 1783 -16894 1838
rect -17208 1558 -16894 1783
rect -16827 1893 -16289 1908
rect -16225 1967 -16003 1996
rect -16225 1922 -16195 1967
rect -16065 1922 -16003 1967
rect -16225 1903 -16003 1922
rect -15937 1995 -15907 2026
rect -15841 1995 -15811 2026
rect -15745 1995 -15715 2026
rect -15937 1962 -15715 1995
rect -15937 1917 -15864 1962
rect -15734 1917 -15715 1962
rect -15937 1902 -15715 1917
rect -15649 1995 -15619 2026
rect -15553 1995 -15523 2026
rect -15457 1995 -15427 2026
rect -15365 1995 -15335 2026
rect -14873 1995 -14843 2026
rect -14781 1995 -14751 2026
rect -14685 1995 -14655 2026
rect -14589 1995 -14559 2026
rect -14493 1996 -14463 2026
rect -14397 1996 -14367 2026
rect -14301 1996 -14271 2026
rect -16827 1753 -16782 1893
rect -16709 1845 -16289 1893
rect -16709 1753 -15715 1845
rect -16827 1736 -15715 1753
rect -16638 1561 -16562 1736
rect -16513 1646 -16291 1671
rect -16513 1601 -16470 1646
rect -16340 1601 -16291 1646
rect -17208 1536 -17178 1558
rect -17112 1536 -17082 1558
rect -17016 1536 -16986 1558
rect -16924 1536 -16894 1558
rect -16605 1536 -16575 1561
rect -16513 1558 -16291 1601
rect -16513 1536 -16483 1558
rect -16417 1536 -16387 1558
rect -16321 1536 -16291 1558
rect -16225 1638 -16003 1666
rect -16225 1593 -16187 1638
rect -16057 1593 -16003 1638
rect -16225 1558 -16003 1593
rect -16225 1536 -16195 1558
rect -16129 1536 -16099 1558
rect -16033 1536 -16003 1558
rect -15937 1558 -15715 1736
rect -15937 1536 -15907 1558
rect -15841 1536 -15811 1558
rect -15745 1536 -15715 1558
rect -15649 1838 -15335 1995
rect -15649 1783 -15617 1838
rect -15552 1783 -15335 1838
rect -15649 1558 -15335 1783
rect -15067 1938 -14557 1995
rect -15067 1828 -15048 1938
rect -15001 1845 -14557 1938
rect -14493 1967 -14271 1996
rect -14493 1922 -14463 1967
rect -14333 1922 -14271 1967
rect -14493 1903 -14271 1922
rect -14205 1995 -14175 2026
rect -14109 1995 -14079 2026
rect -14013 1995 -13983 2026
rect -14205 1962 -13983 1995
rect -14205 1917 -14132 1962
rect -14002 1917 -13983 1962
rect -14205 1902 -13983 1917
rect -13917 1995 -13887 2026
rect -13821 1995 -13791 2026
rect -13725 1995 -13695 2026
rect -13633 1995 -13603 2026
rect -13314 1995 -13284 2026
rect -13222 1995 -13192 2026
rect -13126 1995 -13096 2026
rect -13030 1995 -13000 2026
rect -12934 1996 -12904 2026
rect -12838 1996 -12808 2026
rect -12742 1996 -12712 2026
rect -15001 1828 -13983 1845
rect -15067 1736 -13983 1828
rect -14906 1561 -14830 1736
rect -14781 1646 -14559 1671
rect -14781 1601 -14738 1646
rect -14608 1601 -14559 1646
rect -15649 1536 -15619 1558
rect -15553 1536 -15523 1558
rect -15457 1536 -15427 1558
rect -15365 1536 -15335 1558
rect -14873 1536 -14843 1561
rect -14781 1558 -14559 1601
rect -14781 1536 -14751 1558
rect -14685 1536 -14655 1558
rect -14589 1536 -14559 1558
rect -14493 1638 -14271 1666
rect -14493 1593 -14455 1638
rect -14325 1593 -14271 1638
rect -14493 1558 -14271 1593
rect -14493 1536 -14463 1558
rect -14397 1536 -14367 1558
rect -14301 1536 -14271 1558
rect -14205 1558 -13983 1736
rect -14205 1536 -14175 1558
rect -14109 1536 -14079 1558
rect -14013 1536 -13983 1558
rect -13917 1838 -13603 1995
rect -13347 1908 -12998 1995
rect -13917 1783 -13885 1838
rect -13820 1783 -13603 1838
rect -13917 1558 -13603 1783
rect -13536 1893 -12998 1908
rect -12934 1967 -12712 1996
rect -12934 1922 -12904 1967
rect -12774 1922 -12712 1967
rect -12934 1903 -12712 1922
rect -12646 1995 -12616 2026
rect -12550 1995 -12520 2026
rect -12454 1995 -12424 2026
rect -12646 1962 -12424 1995
rect -12646 1917 -12573 1962
rect -12443 1917 -12424 1962
rect -12646 1902 -12424 1917
rect -12358 1995 -12328 2026
rect -12262 1995 -12232 2026
rect -12166 1995 -12136 2026
rect -12074 1995 -12044 2026
rect -11582 1995 -11552 2026
rect -11490 1995 -11460 2026
rect -11394 1995 -11364 2026
rect -11298 1995 -11268 2026
rect -11202 1996 -11172 2026
rect -11106 1996 -11076 2026
rect -11010 1996 -10980 2026
rect -13536 1753 -13491 1893
rect -13418 1845 -12998 1893
rect -13418 1753 -12424 1845
rect -13536 1736 -12424 1753
rect -13347 1561 -13271 1736
rect -13222 1646 -13000 1671
rect -13222 1601 -13179 1646
rect -13049 1601 -13000 1646
rect -13917 1536 -13887 1558
rect -13821 1536 -13791 1558
rect -13725 1536 -13695 1558
rect -13633 1536 -13603 1558
rect -13314 1536 -13284 1561
rect -13222 1558 -13000 1601
rect -13222 1536 -13192 1558
rect -13126 1536 -13096 1558
rect -13030 1536 -13000 1558
rect -12934 1638 -12712 1666
rect -12934 1593 -12896 1638
rect -12766 1593 -12712 1638
rect -12934 1558 -12712 1593
rect -12934 1536 -12904 1558
rect -12838 1536 -12808 1558
rect -12742 1536 -12712 1558
rect -12646 1558 -12424 1736
rect -12646 1536 -12616 1558
rect -12550 1536 -12520 1558
rect -12454 1536 -12424 1558
rect -12358 1838 -12044 1995
rect -12358 1783 -12326 1838
rect -12261 1783 -12044 1838
rect -12358 1558 -12044 1783
rect -11776 1938 -11266 1995
rect -11776 1828 -11757 1938
rect -11710 1845 -11266 1938
rect -11202 1967 -10980 1996
rect -11202 1922 -11172 1967
rect -11042 1922 -10980 1967
rect -11202 1903 -10980 1922
rect -10914 1995 -10884 2026
rect -10818 1995 -10788 2026
rect -10722 1995 -10692 2026
rect -10914 1962 -10692 1995
rect -10914 1917 -10841 1962
rect -10711 1917 -10692 1962
rect -10914 1902 -10692 1917
rect -10626 1995 -10596 2026
rect -10530 1995 -10500 2026
rect -10434 1995 -10404 2026
rect -10342 1995 -10312 2026
rect -10023 1995 -9993 2026
rect -9931 1995 -9901 2026
rect -9835 1995 -9805 2026
rect -9739 1995 -9709 2026
rect -9643 1996 -9613 2026
rect -9547 1996 -9517 2026
rect -9451 1996 -9421 2026
rect -11710 1828 -10692 1845
rect -11776 1736 -10692 1828
rect -11615 1561 -11539 1736
rect -11490 1646 -11268 1671
rect -11490 1601 -11447 1646
rect -11317 1601 -11268 1646
rect -12358 1536 -12328 1558
rect -12262 1536 -12232 1558
rect -12166 1536 -12136 1558
rect -12074 1536 -12044 1558
rect -11582 1536 -11552 1561
rect -11490 1558 -11268 1601
rect -11490 1536 -11460 1558
rect -11394 1536 -11364 1558
rect -11298 1536 -11268 1558
rect -11202 1638 -10980 1666
rect -11202 1593 -11164 1638
rect -11034 1593 -10980 1638
rect -11202 1558 -10980 1593
rect -11202 1536 -11172 1558
rect -11106 1536 -11076 1558
rect -11010 1536 -10980 1558
rect -10914 1558 -10692 1736
rect -10914 1536 -10884 1558
rect -10818 1536 -10788 1558
rect -10722 1536 -10692 1558
rect -10626 1838 -10312 1995
rect -10056 1908 -9707 1995
rect -10626 1783 -10594 1838
rect -10529 1783 -10312 1838
rect -10626 1558 -10312 1783
rect -10245 1893 -9707 1908
rect -9643 1967 -9421 1996
rect -9643 1922 -9613 1967
rect -9483 1922 -9421 1967
rect -9643 1903 -9421 1922
rect -9355 1995 -9325 2026
rect -9259 1995 -9229 2026
rect -9163 1995 -9133 2026
rect -9355 1962 -9133 1995
rect -9355 1917 -9282 1962
rect -9152 1917 -9133 1962
rect -9355 1902 -9133 1917
rect -9067 1995 -9037 2026
rect -8971 1995 -8941 2026
rect -8875 1995 -8845 2026
rect -8783 1995 -8753 2026
rect -8292 1995 -8262 2026
rect -8200 1995 -8170 2026
rect -8104 1995 -8074 2026
rect -8008 1995 -7978 2026
rect -7912 1996 -7882 2026
rect -7816 1996 -7786 2026
rect -7720 1996 -7690 2026
rect -10245 1753 -10200 1893
rect -10127 1845 -9707 1893
rect -10127 1753 -9133 1845
rect -10245 1736 -9133 1753
rect -10056 1561 -9980 1736
rect -9931 1646 -9709 1671
rect -9931 1601 -9888 1646
rect -9758 1601 -9709 1646
rect -10626 1536 -10596 1558
rect -10530 1536 -10500 1558
rect -10434 1536 -10404 1558
rect -10342 1536 -10312 1558
rect -10023 1536 -9993 1561
rect -9931 1558 -9709 1601
rect -9931 1536 -9901 1558
rect -9835 1536 -9805 1558
rect -9739 1536 -9709 1558
rect -9643 1638 -9421 1666
rect -9643 1593 -9605 1638
rect -9475 1593 -9421 1638
rect -9643 1558 -9421 1593
rect -9643 1536 -9613 1558
rect -9547 1536 -9517 1558
rect -9451 1536 -9421 1558
rect -9355 1558 -9133 1736
rect -9355 1536 -9325 1558
rect -9259 1536 -9229 1558
rect -9163 1536 -9133 1558
rect -9067 1838 -8753 1995
rect -9067 1783 -9035 1838
rect -8970 1783 -8753 1838
rect -9067 1558 -8753 1783
rect -8486 1938 -7976 1995
rect -8486 1828 -8467 1938
rect -8420 1845 -7976 1938
rect -7912 1967 -7690 1996
rect -7912 1922 -7882 1967
rect -7752 1922 -7690 1967
rect -7912 1903 -7690 1922
rect -7624 1995 -7594 2026
rect -7528 1995 -7498 2026
rect -7432 1995 -7402 2026
rect -7624 1962 -7402 1995
rect -7624 1917 -7551 1962
rect -7421 1917 -7402 1962
rect -7624 1902 -7402 1917
rect -7336 1995 -7306 2026
rect -7240 1995 -7210 2026
rect -7144 1995 -7114 2026
rect -7052 1995 -7022 2026
rect -6733 1995 -6703 2026
rect -6641 1995 -6611 2026
rect -6545 1995 -6515 2026
rect -6449 1995 -6419 2026
rect -6353 1996 -6323 2026
rect -6257 1996 -6227 2026
rect -6161 1996 -6131 2026
rect -8420 1828 -7402 1845
rect -8486 1736 -7402 1828
rect -8325 1561 -8249 1736
rect -8200 1646 -7978 1671
rect -8200 1601 -8157 1646
rect -8027 1601 -7978 1646
rect -9067 1536 -9037 1558
rect -8971 1536 -8941 1558
rect -8875 1536 -8845 1558
rect -8783 1536 -8753 1558
rect -8292 1536 -8262 1561
rect -8200 1558 -7978 1601
rect -8200 1536 -8170 1558
rect -8104 1536 -8074 1558
rect -8008 1536 -7978 1558
rect -7912 1638 -7690 1666
rect -7912 1593 -7874 1638
rect -7744 1593 -7690 1638
rect -7912 1558 -7690 1593
rect -7912 1536 -7882 1558
rect -7816 1536 -7786 1558
rect -7720 1536 -7690 1558
rect -7624 1558 -7402 1736
rect -7624 1536 -7594 1558
rect -7528 1536 -7498 1558
rect -7432 1536 -7402 1558
rect -7336 1838 -7022 1995
rect -6766 1908 -6417 1995
rect -7336 1783 -7304 1838
rect -7239 1783 -7022 1838
rect -7336 1558 -7022 1783
rect -6955 1893 -6417 1908
rect -6353 1967 -6131 1996
rect -6353 1922 -6323 1967
rect -6193 1922 -6131 1967
rect -6353 1903 -6131 1922
rect -6065 1995 -6035 2026
rect -5969 1995 -5939 2026
rect -5873 1995 -5843 2026
rect -6065 1962 -5843 1995
rect -6065 1917 -5992 1962
rect -5862 1917 -5843 1962
rect -6065 1902 -5843 1917
rect -5777 1995 -5747 2026
rect -5681 1995 -5651 2026
rect -5585 1995 -5555 2026
rect -5493 1995 -5463 2026
rect -5001 1995 -4971 2026
rect -4909 1995 -4879 2026
rect -4813 1995 -4783 2026
rect -4717 1995 -4687 2026
rect -4621 1996 -4591 2026
rect -4525 1996 -4495 2026
rect -4429 1996 -4399 2026
rect -6955 1753 -6910 1893
rect -6837 1845 -6417 1893
rect -6837 1753 -5843 1845
rect -6955 1736 -5843 1753
rect -6766 1561 -6690 1736
rect -6641 1646 -6419 1671
rect -6641 1601 -6598 1646
rect -6468 1601 -6419 1646
rect -7336 1536 -7306 1558
rect -7240 1536 -7210 1558
rect -7144 1536 -7114 1558
rect -7052 1536 -7022 1558
rect -6733 1536 -6703 1561
rect -6641 1558 -6419 1601
rect -6641 1536 -6611 1558
rect -6545 1536 -6515 1558
rect -6449 1536 -6419 1558
rect -6353 1638 -6131 1666
rect -6353 1593 -6315 1638
rect -6185 1593 -6131 1638
rect -6353 1558 -6131 1593
rect -6353 1536 -6323 1558
rect -6257 1536 -6227 1558
rect -6161 1536 -6131 1558
rect -6065 1558 -5843 1736
rect -6065 1536 -6035 1558
rect -5969 1536 -5939 1558
rect -5873 1536 -5843 1558
rect -5777 1838 -5463 1995
rect -5777 1783 -5745 1838
rect -5680 1783 -5463 1838
rect -5777 1558 -5463 1783
rect -5195 1938 -4685 1995
rect -5195 1828 -5176 1938
rect -5129 1845 -4685 1938
rect -4621 1967 -4399 1996
rect -4621 1922 -4591 1967
rect -4461 1922 -4399 1967
rect -4621 1903 -4399 1922
rect -4333 1995 -4303 2026
rect -4237 1995 -4207 2026
rect -4141 1995 -4111 2026
rect -4333 1962 -4111 1995
rect -4333 1917 -4260 1962
rect -4130 1917 -4111 1962
rect -4333 1902 -4111 1917
rect -4045 1995 -4015 2026
rect -3949 1995 -3919 2026
rect -3853 1995 -3823 2026
rect -3761 1995 -3731 2026
rect -3442 1995 -3412 2026
rect -3350 1995 -3320 2026
rect -3254 1995 -3224 2026
rect -3158 1995 -3128 2026
rect -3062 1996 -3032 2026
rect -2966 1996 -2936 2026
rect -2870 1996 -2840 2026
rect -5129 1828 -4111 1845
rect -5195 1736 -4111 1828
rect -5034 1561 -4958 1736
rect -4909 1646 -4687 1671
rect -4909 1601 -4866 1646
rect -4736 1601 -4687 1646
rect -5777 1536 -5747 1558
rect -5681 1536 -5651 1558
rect -5585 1536 -5555 1558
rect -5493 1536 -5463 1558
rect -5001 1536 -4971 1561
rect -4909 1558 -4687 1601
rect -4909 1536 -4879 1558
rect -4813 1536 -4783 1558
rect -4717 1536 -4687 1558
rect -4621 1638 -4399 1666
rect -4621 1593 -4583 1638
rect -4453 1593 -4399 1638
rect -4621 1558 -4399 1593
rect -4621 1536 -4591 1558
rect -4525 1536 -4495 1558
rect -4429 1536 -4399 1558
rect -4333 1558 -4111 1736
rect -4333 1536 -4303 1558
rect -4237 1536 -4207 1558
rect -4141 1536 -4111 1558
rect -4045 1838 -3731 1995
rect -3475 1908 -3126 1995
rect -4045 1783 -4013 1838
rect -3948 1783 -3731 1838
rect -4045 1558 -3731 1783
rect -3664 1893 -3126 1908
rect -3062 1967 -2840 1996
rect -3062 1922 -3032 1967
rect -2902 1922 -2840 1967
rect -3062 1903 -2840 1922
rect -2774 1995 -2744 2026
rect -2678 1995 -2648 2026
rect -2582 1995 -2552 2026
rect -2774 1962 -2552 1995
rect -2774 1917 -2701 1962
rect -2571 1917 -2552 1962
rect -2774 1902 -2552 1917
rect -2486 1995 -2456 2026
rect -2390 1995 -2360 2026
rect -2294 1995 -2264 2026
rect -2202 1995 -2172 2026
rect -1710 1995 -1680 2026
rect -1618 1995 -1588 2026
rect -1522 1995 -1492 2026
rect -1426 1995 -1396 2026
rect -1330 1996 -1300 2026
rect -1234 1996 -1204 2026
rect -1138 1996 -1108 2026
rect -3664 1753 -3619 1893
rect -3546 1845 -3126 1893
rect -3546 1753 -2552 1845
rect -3664 1736 -2552 1753
rect -3475 1561 -3399 1736
rect -3350 1646 -3128 1671
rect -3350 1601 -3307 1646
rect -3177 1601 -3128 1646
rect -4045 1536 -4015 1558
rect -3949 1536 -3919 1558
rect -3853 1536 -3823 1558
rect -3761 1536 -3731 1558
rect -3442 1536 -3412 1561
rect -3350 1558 -3128 1601
rect -3350 1536 -3320 1558
rect -3254 1536 -3224 1558
rect -3158 1536 -3128 1558
rect -3062 1638 -2840 1666
rect -3062 1593 -3024 1638
rect -2894 1593 -2840 1638
rect -3062 1558 -2840 1593
rect -3062 1536 -3032 1558
rect -2966 1536 -2936 1558
rect -2870 1536 -2840 1558
rect -2774 1558 -2552 1736
rect -2774 1536 -2744 1558
rect -2678 1536 -2648 1558
rect -2582 1536 -2552 1558
rect -2486 1838 -2172 1995
rect -2486 1783 -2454 1838
rect -2389 1783 -2172 1838
rect -2486 1558 -2172 1783
rect -1904 1938 -1394 1995
rect -1904 1828 -1885 1938
rect -1838 1845 -1394 1938
rect -1330 1967 -1108 1996
rect -1330 1922 -1300 1967
rect -1170 1922 -1108 1967
rect -1330 1903 -1108 1922
rect -1042 1995 -1012 2026
rect -946 1995 -916 2026
rect -850 1995 -820 2026
rect -1042 1962 -820 1995
rect -1042 1917 -969 1962
rect -839 1917 -820 1962
rect -1042 1902 -820 1917
rect -754 1995 -724 2026
rect -658 1995 -628 2026
rect -562 1995 -532 2026
rect -470 1995 -440 2026
rect -151 1995 -121 2026
rect -59 1995 -29 2026
rect 37 1995 67 2026
rect 133 1995 163 2026
rect 229 1996 259 2026
rect 325 1996 355 2026
rect 421 1996 451 2026
rect -1838 1828 -820 1845
rect -1904 1736 -820 1828
rect -1743 1561 -1667 1736
rect -1618 1646 -1396 1671
rect -1618 1601 -1575 1646
rect -1445 1601 -1396 1646
rect -2486 1536 -2456 1558
rect -2390 1536 -2360 1558
rect -2294 1536 -2264 1558
rect -2202 1536 -2172 1558
rect -1710 1536 -1680 1561
rect -1618 1558 -1396 1601
rect -1618 1536 -1588 1558
rect -1522 1536 -1492 1558
rect -1426 1536 -1396 1558
rect -1330 1638 -1108 1666
rect -1330 1593 -1292 1638
rect -1162 1593 -1108 1638
rect -1330 1558 -1108 1593
rect -1330 1536 -1300 1558
rect -1234 1536 -1204 1558
rect -1138 1536 -1108 1558
rect -1042 1558 -820 1736
rect -1042 1536 -1012 1558
rect -946 1536 -916 1558
rect -850 1536 -820 1558
rect -754 1838 -440 1995
rect -184 1908 165 1995
rect -754 1783 -722 1838
rect -657 1783 -440 1838
rect -754 1558 -440 1783
rect -373 1893 165 1908
rect 229 1967 451 1996
rect 229 1922 259 1967
rect 389 1922 451 1967
rect 229 1903 451 1922
rect 517 1995 547 2026
rect 613 1995 643 2026
rect 709 1995 739 2026
rect 517 1962 739 1995
rect 517 1917 590 1962
rect 720 1917 739 1962
rect 517 1902 739 1917
rect 805 1995 835 2026
rect 901 1995 931 2026
rect 997 1995 1027 2026
rect 1089 1995 1119 2026
rect -373 1753 -328 1893
rect -255 1845 165 1893
rect -255 1753 739 1845
rect -373 1736 739 1753
rect -184 1561 -108 1736
rect -59 1646 163 1671
rect -59 1601 -16 1646
rect 114 1601 163 1646
rect -754 1536 -724 1558
rect -658 1536 -628 1558
rect -562 1536 -532 1558
rect -470 1536 -440 1558
rect -151 1536 -121 1561
rect -59 1558 163 1601
rect -59 1536 -29 1558
rect 37 1536 67 1558
rect 133 1536 163 1558
rect 229 1638 451 1666
rect 229 1593 267 1638
rect 397 1593 451 1638
rect 229 1558 451 1593
rect 229 1536 259 1558
rect 325 1536 355 1558
rect 421 1536 451 1558
rect 517 1558 739 1736
rect 517 1536 547 1558
rect 613 1536 643 1558
rect 709 1536 739 1558
rect 805 1838 1119 1995
rect 805 1783 837 1838
rect 902 1783 1119 1838
rect 805 1558 1119 1783
rect 11835 2009 11865 2035
rect 11931 2009 11961 2035
rect 12027 2009 12057 2035
rect 12123 2009 12153 2035
rect 12219 2009 12249 2035
rect 12315 2009 12345 2035
rect 12411 2009 12441 2035
rect 12507 2009 12537 2035
rect 12603 2009 12633 2035
rect 12699 2009 12729 2035
rect 12826 1845 12892 1861
rect 11835 1727 11865 1753
rect 11931 1727 11961 1753
rect 12027 1727 12057 1753
rect 12123 1727 12153 1753
rect 12219 1727 12249 1753
rect 11835 1703 12249 1727
rect 7422 1664 7452 1690
rect 7518 1664 7548 1690
rect 7614 1664 7644 1690
rect 7710 1664 7740 1690
rect 8370 1664 8400 1690
rect 8466 1664 8496 1690
rect 8562 1664 8592 1690
rect 8658 1664 8688 1690
rect 9306 1664 9336 1690
rect 9402 1664 9432 1690
rect 9498 1664 9528 1690
rect 9594 1664 9624 1690
rect 10237 1664 10267 1690
rect 10333 1664 10363 1690
rect 10429 1664 10459 1690
rect 10525 1664 10555 1690
rect 11164 1664 11194 1690
rect 11260 1664 11290 1690
rect 11356 1664 11386 1690
rect 11452 1664 11482 1690
rect 11835 1669 12170 1703
rect 12204 1669 12249 1703
rect 11835 1656 12249 1669
rect 7422 1562 7452 1588
rect 7518 1562 7548 1588
rect 7614 1562 7644 1588
rect 7710 1562 7740 1588
rect 8370 1562 8400 1588
rect 8466 1562 8496 1588
rect 8562 1562 8592 1588
rect 8658 1562 8688 1588
rect 9306 1562 9336 1588
rect 9402 1562 9432 1588
rect 9498 1562 9528 1588
rect 9594 1562 9624 1588
rect 10237 1563 10267 1589
rect 10333 1563 10363 1589
rect 10429 1563 10459 1589
rect 10525 1563 10555 1589
rect 805 1536 835 1558
rect 901 1536 931 1558
rect 997 1536 1027 1558
rect 1089 1536 1119 1558
rect -24746 1380 -24716 1406
rect -24654 1380 -24624 1406
rect -24558 1380 -24528 1406
rect -24462 1380 -24432 1406
rect -24366 1380 -24336 1406
rect -24270 1380 -24240 1406
rect -24174 1380 -24144 1406
rect -24078 1380 -24048 1406
rect -23982 1380 -23952 1406
rect -23886 1380 -23856 1406
rect -23790 1380 -23760 1406
rect -23694 1380 -23664 1406
rect -23598 1380 -23568 1406
rect -23506 1380 -23476 1406
rect -23187 1380 -23157 1406
rect -23095 1380 -23065 1406
rect -22999 1380 -22969 1406
rect -22903 1380 -22873 1406
rect -22807 1380 -22777 1406
rect -22711 1380 -22681 1406
rect -22615 1380 -22585 1406
rect -22519 1380 -22489 1406
rect -22423 1380 -22393 1406
rect -22327 1380 -22297 1406
rect -22231 1380 -22201 1406
rect -22135 1380 -22105 1406
rect -22039 1380 -22009 1406
rect -21947 1380 -21917 1406
rect -21455 1380 -21425 1406
rect -21363 1380 -21333 1406
rect -21267 1380 -21237 1406
rect -21171 1380 -21141 1406
rect -21075 1380 -21045 1406
rect -20979 1380 -20949 1406
rect -20883 1380 -20853 1406
rect -20787 1380 -20757 1406
rect -20691 1380 -20661 1406
rect -20595 1380 -20565 1406
rect -20499 1380 -20469 1406
rect -20403 1380 -20373 1406
rect -20307 1380 -20277 1406
rect -20215 1380 -20185 1406
rect -19896 1380 -19866 1406
rect -19804 1380 -19774 1406
rect -19708 1380 -19678 1406
rect -19612 1380 -19582 1406
rect -19516 1380 -19486 1406
rect -19420 1380 -19390 1406
rect -19324 1380 -19294 1406
rect -19228 1380 -19198 1406
rect -19132 1380 -19102 1406
rect -19036 1380 -19006 1406
rect -18940 1380 -18910 1406
rect -18844 1380 -18814 1406
rect -18748 1380 -18718 1406
rect -18656 1380 -18626 1406
rect -18164 1380 -18134 1406
rect -18072 1380 -18042 1406
rect -17976 1380 -17946 1406
rect -17880 1380 -17850 1406
rect -17784 1380 -17754 1406
rect -17688 1380 -17658 1406
rect -17592 1380 -17562 1406
rect -17496 1380 -17466 1406
rect -17400 1380 -17370 1406
rect -17304 1380 -17274 1406
rect -17208 1380 -17178 1406
rect -17112 1380 -17082 1406
rect -17016 1380 -16986 1406
rect -16924 1380 -16894 1406
rect -16605 1380 -16575 1406
rect -16513 1380 -16483 1406
rect -16417 1380 -16387 1406
rect -16321 1380 -16291 1406
rect -16225 1380 -16195 1406
rect -16129 1380 -16099 1406
rect -16033 1380 -16003 1406
rect -15937 1380 -15907 1406
rect -15841 1380 -15811 1406
rect -15745 1380 -15715 1406
rect -15649 1380 -15619 1406
rect -15553 1380 -15523 1406
rect -15457 1380 -15427 1406
rect -15365 1380 -15335 1406
rect -14873 1380 -14843 1406
rect -14781 1380 -14751 1406
rect -14685 1380 -14655 1406
rect -14589 1380 -14559 1406
rect -14493 1380 -14463 1406
rect -14397 1380 -14367 1406
rect -14301 1380 -14271 1406
rect -14205 1380 -14175 1406
rect -14109 1380 -14079 1406
rect -14013 1380 -13983 1406
rect -13917 1380 -13887 1406
rect -13821 1380 -13791 1406
rect -13725 1380 -13695 1406
rect -13633 1380 -13603 1406
rect -13314 1380 -13284 1406
rect -13222 1380 -13192 1406
rect -13126 1380 -13096 1406
rect -13030 1380 -13000 1406
rect -12934 1380 -12904 1406
rect -12838 1380 -12808 1406
rect -12742 1380 -12712 1406
rect -12646 1380 -12616 1406
rect -12550 1380 -12520 1406
rect -12454 1380 -12424 1406
rect -12358 1380 -12328 1406
rect -12262 1380 -12232 1406
rect -12166 1380 -12136 1406
rect -12074 1380 -12044 1406
rect -11582 1380 -11552 1406
rect -11490 1380 -11460 1406
rect -11394 1380 -11364 1406
rect -11298 1380 -11268 1406
rect -11202 1380 -11172 1406
rect -11106 1380 -11076 1406
rect -11010 1380 -10980 1406
rect -10914 1380 -10884 1406
rect -10818 1380 -10788 1406
rect -10722 1380 -10692 1406
rect -10626 1380 -10596 1406
rect -10530 1380 -10500 1406
rect -10434 1380 -10404 1406
rect -10342 1380 -10312 1406
rect -10023 1380 -9993 1406
rect -9931 1380 -9901 1406
rect -9835 1380 -9805 1406
rect -9739 1380 -9709 1406
rect -9643 1380 -9613 1406
rect -9547 1380 -9517 1406
rect -9451 1380 -9421 1406
rect -9355 1380 -9325 1406
rect -9259 1380 -9229 1406
rect -9163 1380 -9133 1406
rect -9067 1380 -9037 1406
rect -8971 1380 -8941 1406
rect -8875 1380 -8845 1406
rect -8783 1380 -8753 1406
rect -8292 1380 -8262 1406
rect -8200 1380 -8170 1406
rect -8104 1380 -8074 1406
rect -8008 1380 -7978 1406
rect -7912 1380 -7882 1406
rect -7816 1380 -7786 1406
rect -7720 1380 -7690 1406
rect -7624 1380 -7594 1406
rect -7528 1380 -7498 1406
rect -7432 1380 -7402 1406
rect -7336 1380 -7306 1406
rect -7240 1380 -7210 1406
rect -7144 1380 -7114 1406
rect -7052 1380 -7022 1406
rect -6733 1380 -6703 1406
rect -6641 1380 -6611 1406
rect -6545 1380 -6515 1406
rect -6449 1380 -6419 1406
rect -6353 1380 -6323 1406
rect -6257 1380 -6227 1406
rect -6161 1380 -6131 1406
rect -6065 1380 -6035 1406
rect -5969 1380 -5939 1406
rect -5873 1380 -5843 1406
rect -5777 1380 -5747 1406
rect -5681 1380 -5651 1406
rect -5585 1380 -5555 1406
rect -5493 1380 -5463 1406
rect -5001 1380 -4971 1406
rect -4909 1380 -4879 1406
rect -4813 1380 -4783 1406
rect -4717 1380 -4687 1406
rect -4621 1380 -4591 1406
rect -4525 1380 -4495 1406
rect -4429 1380 -4399 1406
rect -4333 1380 -4303 1406
rect -4237 1380 -4207 1406
rect -4141 1380 -4111 1406
rect -4045 1380 -4015 1406
rect -3949 1380 -3919 1406
rect -3853 1380 -3823 1406
rect -3761 1380 -3731 1406
rect -3442 1380 -3412 1406
rect -3350 1380 -3320 1406
rect -3254 1380 -3224 1406
rect -3158 1380 -3128 1406
rect -3062 1380 -3032 1406
rect -2966 1380 -2936 1406
rect -2870 1380 -2840 1406
rect -2774 1380 -2744 1406
rect -2678 1380 -2648 1406
rect -2582 1380 -2552 1406
rect -2486 1380 -2456 1406
rect -2390 1380 -2360 1406
rect -2294 1380 -2264 1406
rect -2202 1380 -2172 1406
rect -1710 1380 -1680 1406
rect -1618 1380 -1588 1406
rect -1522 1380 -1492 1406
rect -1426 1380 -1396 1406
rect -1330 1380 -1300 1406
rect -1234 1380 -1204 1406
rect -1138 1380 -1108 1406
rect -1042 1380 -1012 1406
rect -946 1380 -916 1406
rect -850 1380 -820 1406
rect -754 1380 -724 1406
rect -658 1380 -628 1406
rect -562 1380 -532 1406
rect -470 1380 -440 1406
rect -151 1380 -121 1406
rect -59 1380 -29 1406
rect 37 1380 67 1406
rect 133 1380 163 1406
rect 229 1380 259 1406
rect 325 1380 355 1406
rect 421 1380 451 1406
rect 517 1380 547 1406
rect 613 1380 643 1406
rect 709 1380 739 1406
rect 805 1380 835 1406
rect 901 1380 931 1406
rect 997 1380 1027 1406
rect 1089 1380 1119 1406
rect -24535 875 -24505 906
rect -24439 875 -24409 906
rect -24343 875 -24313 906
rect -24247 875 -24217 906
rect -24151 875 -24121 906
rect -24055 875 -24025 906
rect -23426 875 -23396 906
rect -23330 875 -23300 906
rect -23234 875 -23204 906
rect -23138 875 -23108 906
rect -23042 875 -23012 906
rect -22946 875 -22916 906
rect -22544 875 -22514 906
rect -22448 875 -22418 906
rect -22352 875 -22322 906
rect -22256 875 -22226 906
rect -22160 875 -22130 906
rect -22064 875 -22034 906
rect -21244 875 -21214 906
rect -21148 875 -21118 906
rect -21052 875 -21022 906
rect -20956 875 -20926 906
rect -20860 875 -20830 906
rect -20764 875 -20734 906
rect -20135 875 -20105 906
rect -20039 875 -20009 906
rect -19943 875 -19913 906
rect -19847 875 -19817 906
rect -19751 875 -19721 906
rect -19655 875 -19625 906
rect -19253 875 -19223 906
rect -19157 875 -19127 906
rect -19061 875 -19031 906
rect -18965 875 -18935 906
rect -18869 875 -18839 906
rect -18773 875 -18743 906
rect -17953 875 -17923 906
rect -17857 875 -17827 906
rect -17761 875 -17731 906
rect -17665 875 -17635 906
rect -17569 875 -17539 906
rect -17473 875 -17443 906
rect -16844 875 -16814 906
rect -16748 875 -16718 906
rect -16652 875 -16622 906
rect -16556 875 -16526 906
rect -16460 875 -16430 906
rect -16364 875 -16334 906
rect -15962 875 -15932 906
rect -15866 875 -15836 906
rect -15770 875 -15740 906
rect -15674 875 -15644 906
rect -15578 875 -15548 906
rect -15482 875 -15452 906
rect -14662 875 -14632 906
rect -14566 875 -14536 906
rect -14470 875 -14440 906
rect -14374 875 -14344 906
rect -14278 875 -14248 906
rect -14182 875 -14152 906
rect -13553 875 -13523 906
rect -13457 875 -13427 906
rect -13361 875 -13331 906
rect -13265 875 -13235 906
rect -13169 875 -13139 906
rect -13073 875 -13043 906
rect -12671 875 -12641 906
rect -12575 875 -12545 906
rect -12479 875 -12449 906
rect -12383 875 -12353 906
rect -12287 875 -12257 906
rect -12191 875 -12161 906
rect -11371 875 -11341 906
rect -11275 875 -11245 906
rect -11179 875 -11149 906
rect -11083 875 -11053 906
rect -10987 875 -10957 906
rect -10891 875 -10861 906
rect -10262 875 -10232 906
rect -10166 875 -10136 906
rect -10070 875 -10040 906
rect -9974 875 -9944 906
rect -9878 875 -9848 906
rect -9782 875 -9752 906
rect -9380 875 -9350 906
rect -9284 875 -9254 906
rect -9188 875 -9158 906
rect -9092 875 -9062 906
rect -8996 875 -8966 906
rect -8900 875 -8870 906
rect -8081 875 -8051 906
rect -7985 875 -7955 906
rect -7889 875 -7859 906
rect -7793 875 -7763 906
rect -7697 875 -7667 906
rect -7601 875 -7571 906
rect -6972 875 -6942 906
rect -6876 875 -6846 906
rect -6780 875 -6750 906
rect -6684 875 -6654 906
rect -6588 875 -6558 906
rect -6492 875 -6462 906
rect -6090 875 -6060 906
rect -5994 875 -5964 906
rect -5898 875 -5868 906
rect -5802 875 -5772 906
rect -5706 875 -5676 906
rect -5610 875 -5580 906
rect -4790 875 -4760 906
rect -4694 875 -4664 906
rect -4598 875 -4568 906
rect -4502 875 -4472 906
rect -4406 875 -4376 906
rect -4310 875 -4280 906
rect -3681 875 -3651 906
rect -3585 875 -3555 906
rect -3489 875 -3459 906
rect -3393 875 -3363 906
rect -3297 875 -3267 906
rect -3201 875 -3171 906
rect -2799 875 -2769 906
rect -2703 875 -2673 906
rect -2607 875 -2577 906
rect -2511 875 -2481 906
rect -2415 875 -2385 906
rect -2319 875 -2289 906
rect -1499 875 -1469 906
rect -1403 875 -1373 906
rect -1307 875 -1277 906
rect -1211 875 -1181 906
rect -1115 875 -1085 906
rect -1019 875 -989 906
rect -390 875 -360 906
rect -294 875 -264 906
rect -198 875 -168 906
rect -102 875 -72 906
rect -6 875 24 906
rect 90 875 120 906
rect 492 875 522 906
rect 588 875 618 906
rect 684 875 714 906
rect 780 875 810 906
rect 876 875 906 906
rect 972 875 1002 906
rect 11164 1562 11194 1588
rect 11260 1562 11290 1588
rect 11356 1562 11386 1588
rect 11452 1562 11482 1588
rect 7422 729 7452 762
rect 7238 699 7452 729
rect -24535 635 -24505 661
rect -24439 635 -24409 661
rect -24343 635 -24313 661
rect -24536 614 -24313 635
rect -24536 579 -24519 614
rect -24485 605 -24313 614
rect -24247 635 -24217 661
rect -24151 635 -24121 661
rect -24055 635 -24025 661
rect -23426 635 -23396 661
rect -23330 635 -23300 661
rect -23234 635 -23204 661
rect -24247 614 -24025 635
rect -24485 579 -24469 605
rect -24536 568 -24469 579
rect -24247 579 -24230 614
rect -24196 605 -24025 614
rect -23427 614 -23204 635
rect -24196 579 -24180 605
rect -24247 568 -24180 579
rect -23427 579 -23410 614
rect -23376 605 -23204 614
rect -23138 635 -23108 661
rect -23042 635 -23012 661
rect -22946 635 -22916 661
rect -22544 635 -22514 661
rect -22448 635 -22418 661
rect -22352 635 -22322 661
rect -23138 614 -22916 635
rect -23376 579 -23360 605
rect -23427 568 -23360 579
rect -23138 579 -23121 614
rect -23087 605 -22916 614
rect -22545 614 -22322 635
rect -23087 579 -23071 605
rect -23138 568 -23071 579
rect -22545 579 -22528 614
rect -22494 605 -22322 614
rect -22256 635 -22226 661
rect -22160 635 -22130 661
rect -22064 635 -22034 661
rect -21244 635 -21214 661
rect -21148 635 -21118 661
rect -21052 635 -21022 661
rect -22256 614 -22034 635
rect -22494 579 -22478 605
rect -22545 568 -22478 579
rect -22256 579 -22239 614
rect -22205 605 -22034 614
rect -21245 614 -21022 635
rect -22205 579 -22189 605
rect -22256 568 -22189 579
rect -21245 579 -21228 614
rect -21194 605 -21022 614
rect -20956 635 -20926 661
rect -20860 635 -20830 661
rect -20764 635 -20734 661
rect -20135 635 -20105 661
rect -20039 635 -20009 661
rect -19943 635 -19913 661
rect -20956 614 -20734 635
rect -21194 579 -21178 605
rect -21245 568 -21178 579
rect -20956 579 -20939 614
rect -20905 605 -20734 614
rect -20136 614 -19913 635
rect -20905 579 -20889 605
rect -20956 568 -20889 579
rect -20136 579 -20119 614
rect -20085 605 -19913 614
rect -19847 635 -19817 661
rect -19751 635 -19721 661
rect -19655 635 -19625 661
rect -19253 635 -19223 661
rect -19157 635 -19127 661
rect -19061 635 -19031 661
rect -19847 614 -19625 635
rect -20085 579 -20069 605
rect -20136 568 -20069 579
rect -19847 579 -19830 614
rect -19796 605 -19625 614
rect -19254 614 -19031 635
rect -19796 579 -19780 605
rect -19847 568 -19780 579
rect -19254 579 -19237 614
rect -19203 605 -19031 614
rect -18965 635 -18935 661
rect -18869 635 -18839 661
rect -18773 635 -18743 661
rect -17953 635 -17923 661
rect -17857 635 -17827 661
rect -17761 635 -17731 661
rect -18965 614 -18743 635
rect -19203 579 -19187 605
rect -19254 568 -19187 579
rect -18965 579 -18948 614
rect -18914 605 -18743 614
rect -17954 614 -17731 635
rect -18914 579 -18898 605
rect -18965 568 -18898 579
rect -17954 579 -17937 614
rect -17903 605 -17731 614
rect -17665 635 -17635 661
rect -17569 635 -17539 661
rect -17473 635 -17443 661
rect -16844 635 -16814 661
rect -16748 635 -16718 661
rect -16652 635 -16622 661
rect -17665 614 -17443 635
rect -17903 579 -17887 605
rect -17954 568 -17887 579
rect -17665 579 -17648 614
rect -17614 605 -17443 614
rect -16845 614 -16622 635
rect -17614 579 -17598 605
rect -17665 568 -17598 579
rect -16845 579 -16828 614
rect -16794 605 -16622 614
rect -16556 635 -16526 661
rect -16460 635 -16430 661
rect -16364 635 -16334 661
rect -15962 635 -15932 661
rect -15866 635 -15836 661
rect -15770 635 -15740 661
rect -16556 614 -16334 635
rect -16794 579 -16778 605
rect -16845 568 -16778 579
rect -16556 579 -16539 614
rect -16505 605 -16334 614
rect -15963 614 -15740 635
rect -16505 579 -16489 605
rect -16556 568 -16489 579
rect -15963 579 -15946 614
rect -15912 605 -15740 614
rect -15674 635 -15644 661
rect -15578 635 -15548 661
rect -15482 635 -15452 661
rect -14662 635 -14632 661
rect -14566 635 -14536 661
rect -14470 635 -14440 661
rect -15674 614 -15452 635
rect -15912 579 -15896 605
rect -15963 568 -15896 579
rect -15674 579 -15657 614
rect -15623 605 -15452 614
rect -14663 614 -14440 635
rect -15623 579 -15607 605
rect -15674 568 -15607 579
rect -14663 579 -14646 614
rect -14612 605 -14440 614
rect -14374 635 -14344 661
rect -14278 635 -14248 661
rect -14182 635 -14152 661
rect -13553 635 -13523 661
rect -13457 635 -13427 661
rect -13361 635 -13331 661
rect -14374 614 -14152 635
rect -14612 579 -14596 605
rect -14663 568 -14596 579
rect -14374 579 -14357 614
rect -14323 605 -14152 614
rect -13554 614 -13331 635
rect -14323 579 -14307 605
rect -14374 568 -14307 579
rect -13554 579 -13537 614
rect -13503 605 -13331 614
rect -13265 635 -13235 661
rect -13169 635 -13139 661
rect -13073 635 -13043 661
rect -12671 635 -12641 661
rect -12575 635 -12545 661
rect -12479 635 -12449 661
rect -13265 614 -13043 635
rect -13503 579 -13487 605
rect -13554 568 -13487 579
rect -13265 579 -13248 614
rect -13214 605 -13043 614
rect -12672 614 -12449 635
rect -13214 579 -13198 605
rect -13265 568 -13198 579
rect -12672 579 -12655 614
rect -12621 605 -12449 614
rect -12383 635 -12353 661
rect -12287 635 -12257 661
rect -12191 635 -12161 661
rect -11371 635 -11341 661
rect -11275 635 -11245 661
rect -11179 635 -11149 661
rect -12383 614 -12161 635
rect -12621 579 -12605 605
rect -12672 568 -12605 579
rect -12383 579 -12366 614
rect -12332 605 -12161 614
rect -11372 614 -11149 635
rect -12332 579 -12316 605
rect -12383 568 -12316 579
rect -11372 579 -11355 614
rect -11321 605 -11149 614
rect -11083 635 -11053 661
rect -10987 635 -10957 661
rect -10891 635 -10861 661
rect -10262 635 -10232 661
rect -10166 635 -10136 661
rect -10070 635 -10040 661
rect -11083 614 -10861 635
rect -11321 579 -11305 605
rect -11372 568 -11305 579
rect -11083 579 -11066 614
rect -11032 605 -10861 614
rect -10263 614 -10040 635
rect -11032 579 -11016 605
rect -11083 568 -11016 579
rect -10263 579 -10246 614
rect -10212 605 -10040 614
rect -9974 635 -9944 661
rect -9878 635 -9848 661
rect -9782 635 -9752 661
rect -9380 635 -9350 661
rect -9284 635 -9254 661
rect -9188 635 -9158 661
rect -9974 614 -9752 635
rect -10212 579 -10196 605
rect -10263 568 -10196 579
rect -9974 579 -9957 614
rect -9923 605 -9752 614
rect -9381 614 -9158 635
rect -9923 579 -9907 605
rect -9974 568 -9907 579
rect -9381 579 -9364 614
rect -9330 605 -9158 614
rect -9092 635 -9062 661
rect -8996 635 -8966 661
rect -8900 635 -8870 661
rect -8081 635 -8051 661
rect -7985 635 -7955 661
rect -7889 635 -7859 661
rect -9092 614 -8870 635
rect -9330 579 -9314 605
rect -9381 568 -9314 579
rect -9092 579 -9075 614
rect -9041 605 -8870 614
rect -8082 614 -7859 635
rect -9041 579 -9025 605
rect -9092 568 -9025 579
rect -8082 579 -8065 614
rect -8031 605 -7859 614
rect -7793 635 -7763 661
rect -7697 635 -7667 661
rect -7601 635 -7571 661
rect -6972 635 -6942 661
rect -6876 635 -6846 661
rect -6780 635 -6750 661
rect -7793 614 -7571 635
rect -8031 579 -8015 605
rect -8082 568 -8015 579
rect -7793 579 -7776 614
rect -7742 605 -7571 614
rect -6973 614 -6750 635
rect -7742 579 -7726 605
rect -7793 568 -7726 579
rect -6973 579 -6956 614
rect -6922 605 -6750 614
rect -6684 635 -6654 661
rect -6588 635 -6558 661
rect -6492 635 -6462 661
rect -6090 635 -6060 661
rect -5994 635 -5964 661
rect -5898 635 -5868 661
rect -6684 614 -6462 635
rect -6922 579 -6906 605
rect -6973 568 -6906 579
rect -6684 579 -6667 614
rect -6633 605 -6462 614
rect -6091 614 -5868 635
rect -6633 579 -6617 605
rect -6684 568 -6617 579
rect -6091 579 -6074 614
rect -6040 605 -5868 614
rect -5802 635 -5772 661
rect -5706 635 -5676 661
rect -5610 635 -5580 661
rect -4790 635 -4760 661
rect -4694 635 -4664 661
rect -4598 635 -4568 661
rect -5802 614 -5580 635
rect -6040 579 -6024 605
rect -6091 568 -6024 579
rect -5802 579 -5785 614
rect -5751 605 -5580 614
rect -4791 614 -4568 635
rect -5751 579 -5735 605
rect -5802 568 -5735 579
rect -4791 579 -4774 614
rect -4740 605 -4568 614
rect -4502 635 -4472 661
rect -4406 635 -4376 661
rect -4310 635 -4280 661
rect -3681 635 -3651 661
rect -3585 635 -3555 661
rect -3489 635 -3459 661
rect -4502 614 -4280 635
rect -4740 579 -4724 605
rect -4791 568 -4724 579
rect -4502 579 -4485 614
rect -4451 605 -4280 614
rect -3682 614 -3459 635
rect -4451 579 -4435 605
rect -4502 568 -4435 579
rect -3682 579 -3665 614
rect -3631 605 -3459 614
rect -3393 635 -3363 661
rect -3297 635 -3267 661
rect -3201 635 -3171 661
rect -2799 635 -2769 661
rect -2703 635 -2673 661
rect -2607 635 -2577 661
rect -3393 614 -3171 635
rect -3631 579 -3615 605
rect -3682 568 -3615 579
rect -3393 579 -3376 614
rect -3342 605 -3171 614
rect -2800 614 -2577 635
rect -3342 579 -3326 605
rect -3393 568 -3326 579
rect -2800 579 -2783 614
rect -2749 605 -2577 614
rect -2511 635 -2481 661
rect -2415 635 -2385 661
rect -2319 635 -2289 661
rect -1499 635 -1469 661
rect -1403 635 -1373 661
rect -1307 635 -1277 661
rect -2511 614 -2289 635
rect -2749 579 -2733 605
rect -2800 568 -2733 579
rect -2511 579 -2494 614
rect -2460 605 -2289 614
rect -1500 614 -1277 635
rect -2460 579 -2444 605
rect -2511 568 -2444 579
rect -1500 579 -1483 614
rect -1449 605 -1277 614
rect -1211 635 -1181 661
rect -1115 635 -1085 661
rect -1019 635 -989 661
rect -390 635 -360 661
rect -294 635 -264 661
rect -198 635 -168 661
rect -1211 614 -989 635
rect -1449 579 -1433 605
rect -1500 568 -1433 579
rect -1211 579 -1194 614
rect -1160 605 -989 614
rect -391 614 -168 635
rect -1160 579 -1144 605
rect -1211 568 -1144 579
rect -391 579 -374 614
rect -340 605 -168 614
rect -102 635 -72 661
rect -6 635 24 661
rect 90 635 120 661
rect 492 635 522 661
rect 588 635 618 661
rect 684 635 714 661
rect -102 614 120 635
rect -340 579 -324 605
rect -391 568 -324 579
rect -102 579 -85 614
rect -51 605 120 614
rect 491 614 714 635
rect -51 579 -35 605
rect -102 568 -35 579
rect 491 579 508 614
rect 542 605 714 614
rect 780 635 810 661
rect 876 635 906 661
rect 972 635 1002 661
rect 780 614 1002 635
rect 542 579 558 605
rect 491 568 558 579
rect 780 579 797 614
rect 831 605 1002 614
rect 831 579 847 605
rect 780 568 847 579
rect -24536 373 -24493 568
rect -24451 490 -24385 506
rect -24451 455 -24435 490
rect -24401 469 -24385 490
rect -24401 455 -24363 469
rect -24451 439 -24363 455
rect -23963 439 -23937 469
rect -23427 373 -23384 568
rect -23342 490 -23276 506
rect -23342 455 -23326 490
rect -23292 469 -23276 490
rect -23292 455 -23254 469
rect -23342 439 -23254 455
rect -22854 439 -22828 469
rect -22545 373 -22502 568
rect -22460 490 -22394 506
rect -22460 455 -22444 490
rect -22410 469 -22394 490
rect -22410 455 -22372 469
rect -22460 439 -22372 455
rect -21972 439 -21946 469
rect -21245 373 -21202 568
rect -21160 490 -21094 506
rect -21160 455 -21144 490
rect -21110 469 -21094 490
rect -21110 455 -21072 469
rect -21160 439 -21072 455
rect -20672 439 -20646 469
rect -20136 373 -20093 568
rect -20051 490 -19985 506
rect -20051 455 -20035 490
rect -20001 469 -19985 490
rect -20001 455 -19963 469
rect -20051 439 -19963 455
rect -19563 439 -19537 469
rect -19254 373 -19211 568
rect -19169 490 -19103 506
rect -19169 455 -19153 490
rect -19119 469 -19103 490
rect -19119 455 -19081 469
rect -19169 439 -19081 455
rect -18681 439 -18655 469
rect -17954 373 -17911 568
rect -17869 490 -17803 506
rect -17869 455 -17853 490
rect -17819 469 -17803 490
rect -17819 455 -17781 469
rect -17869 439 -17781 455
rect -17381 439 -17355 469
rect -16845 373 -16802 568
rect -16760 490 -16694 506
rect -16760 455 -16744 490
rect -16710 469 -16694 490
rect -16710 455 -16672 469
rect -16760 439 -16672 455
rect -16272 439 -16246 469
rect -15963 373 -15920 568
rect -15878 490 -15812 506
rect -15878 455 -15862 490
rect -15828 469 -15812 490
rect -15828 455 -15790 469
rect -15878 439 -15790 455
rect -15390 439 -15364 469
rect -14663 373 -14620 568
rect -14578 490 -14512 506
rect -14578 455 -14562 490
rect -14528 469 -14512 490
rect -14528 455 -14490 469
rect -14578 439 -14490 455
rect -14090 439 -14064 469
rect -13554 373 -13511 568
rect -13469 490 -13403 506
rect -13469 455 -13453 490
rect -13419 469 -13403 490
rect -13419 455 -13381 469
rect -13469 439 -13381 455
rect -12981 439 -12955 469
rect -12672 373 -12629 568
rect -12587 490 -12521 506
rect -12587 455 -12571 490
rect -12537 469 -12521 490
rect -12537 455 -12499 469
rect -12587 439 -12499 455
rect -12099 439 -12073 469
rect -11372 373 -11329 568
rect -11287 490 -11221 506
rect -11287 455 -11271 490
rect -11237 469 -11221 490
rect -11237 455 -11199 469
rect -11287 439 -11199 455
rect -10799 439 -10773 469
rect -10263 373 -10220 568
rect -10178 490 -10112 506
rect -10178 455 -10162 490
rect -10128 469 -10112 490
rect -10128 455 -10090 469
rect -10178 439 -10090 455
rect -9690 439 -9664 469
rect -9381 373 -9338 568
rect -9296 490 -9230 506
rect -9296 455 -9280 490
rect -9246 469 -9230 490
rect -9246 455 -9208 469
rect -9296 439 -9208 455
rect -8808 439 -8782 469
rect -8082 373 -8039 568
rect -7997 490 -7931 506
rect -7997 455 -7981 490
rect -7947 469 -7931 490
rect -7947 455 -7909 469
rect -7997 439 -7909 455
rect -7509 439 -7483 469
rect -6973 373 -6930 568
rect -6888 490 -6822 506
rect -6888 455 -6872 490
rect -6838 469 -6822 490
rect -6838 455 -6800 469
rect -6888 439 -6800 455
rect -6400 439 -6374 469
rect -6091 373 -6048 568
rect -6006 490 -5940 506
rect -6006 455 -5990 490
rect -5956 469 -5940 490
rect -5956 455 -5918 469
rect -6006 439 -5918 455
rect -5518 439 -5492 469
rect -4791 373 -4748 568
rect -4706 490 -4640 506
rect -4706 455 -4690 490
rect -4656 469 -4640 490
rect -4656 455 -4618 469
rect -4706 439 -4618 455
rect -4218 439 -4192 469
rect -3682 373 -3639 568
rect -3597 490 -3531 506
rect -3597 455 -3581 490
rect -3547 469 -3531 490
rect -3547 455 -3509 469
rect -3597 439 -3509 455
rect -3109 439 -3083 469
rect -2800 373 -2757 568
rect -2715 490 -2649 506
rect -2715 455 -2699 490
rect -2665 469 -2649 490
rect -2665 455 -2627 469
rect -2715 439 -2627 455
rect -2227 439 -2201 469
rect -1500 373 -1457 568
rect -1415 490 -1349 506
rect -1415 455 -1399 490
rect -1365 469 -1349 490
rect -1365 455 -1327 469
rect -1415 439 -1327 455
rect -927 439 -901 469
rect -391 373 -348 568
rect -306 490 -240 506
rect -306 455 -290 490
rect -256 469 -240 490
rect -256 455 -218 469
rect -306 439 -218 455
rect 182 439 208 469
rect 491 373 534 568
rect 576 490 642 506
rect 576 455 592 490
rect 626 469 642 490
rect 626 455 664 469
rect 576 439 664 455
rect 1064 439 1090 469
rect 7238 452 7268 699
rect 7518 657 7548 762
rect 7614 739 7644 762
rect 7374 519 7548 657
rect 7182 436 7326 452
rect 7182 402 7198 436
rect 7232 402 7326 436
rect 7182 386 7326 402
rect 7374 436 7518 519
rect 7590 477 7644 739
rect 7710 612 7740 762
rect 8370 729 8400 762
rect 8186 699 8400 729
rect 7710 582 7848 612
rect 7584 452 7644 477
rect 7758 452 7848 582
rect 8186 452 8216 699
rect 8466 657 8496 762
rect 8562 739 8592 762
rect 8322 519 8496 657
rect 7374 402 7390 436
rect 7424 402 7518 436
rect 7374 386 7518 402
rect 7566 436 7710 452
rect 7566 402 7582 436
rect 7616 402 7710 436
rect 7566 386 7710 402
rect 7758 436 7902 452
rect 7758 402 7774 436
rect 7808 402 7902 436
rect 7758 386 7902 402
rect 8130 436 8274 452
rect 8130 402 8146 436
rect 8180 402 8274 436
rect 8130 386 8274 402
rect 8322 436 8466 519
rect 8538 477 8592 739
rect 8658 612 8688 762
rect 9306 729 9336 762
rect 9122 699 9336 729
rect 8658 582 8796 612
rect 8532 452 8592 477
rect 8706 452 8796 582
rect 9122 452 9152 699
rect 9402 657 9432 762
rect 9498 739 9528 762
rect 9258 519 9432 657
rect 8322 402 8338 436
rect 8372 402 8466 436
rect 8322 386 8466 402
rect 8514 436 8658 452
rect 8514 402 8530 436
rect 8564 402 8658 436
rect 8514 386 8658 402
rect 8706 436 8850 452
rect 8706 402 8722 436
rect 8756 402 8850 436
rect 8706 386 8850 402
rect 9066 436 9210 452
rect 9066 402 9082 436
rect 9116 402 9210 436
rect 9066 386 9210 402
rect 9258 436 9402 519
rect 9474 477 9528 739
rect 9594 612 9624 762
rect 10237 730 10267 763
rect 10053 700 10267 730
rect 9594 582 9732 612
rect 9468 452 9528 477
rect 9642 452 9732 582
rect 10053 453 10083 700
rect 10333 658 10363 763
rect 10429 740 10459 763
rect 10189 520 10363 658
rect 9258 402 9274 436
rect 9308 402 9402 436
rect 9258 386 9402 402
rect 9450 436 9594 452
rect 9450 402 9466 436
rect 9500 402 9594 436
rect 9450 386 9594 402
rect 9642 436 9786 452
rect 9642 402 9658 436
rect 9692 402 9786 436
rect 9642 386 9786 402
rect 9997 437 10141 453
rect 9997 403 10013 437
rect 10047 403 10141 437
rect 9997 387 10141 403
rect 10189 437 10333 520
rect 10405 478 10459 740
rect 10525 613 10555 763
rect 12219 1520 12249 1656
rect 12315 1727 12345 1753
rect 12411 1727 12441 1753
rect 12507 1727 12537 1753
rect 12603 1727 12633 1753
rect 12699 1727 12729 1753
rect 12315 1656 12729 1727
rect 12315 1614 12345 1656
rect 12826 1619 12842 1845
rect 12876 1843 12892 1845
rect 12876 1813 12923 1843
rect 13137 1813 13163 1843
rect 12876 1747 12892 1813
rect 12876 1717 12923 1747
rect 13137 1717 13163 1747
rect 12876 1651 12892 1717
rect 12876 1621 12923 1651
rect 13137 1621 13163 1651
rect 12876 1619 12892 1621
rect 12297 1598 12363 1614
rect 12826 1603 12892 1619
rect 12297 1564 12313 1598
rect 12347 1564 12363 1598
rect 12297 1548 12363 1564
rect 12315 1520 12345 1548
rect 12826 1399 12893 1415
rect 12826 1365 12842 1399
rect 12876 1397 12893 1399
rect 12876 1367 12923 1397
rect 13123 1367 13149 1397
rect 12876 1365 12893 1367
rect 12826 1349 12893 1365
rect 12219 1294 12249 1320
rect 12315 1294 12345 1320
rect 11164 729 11194 762
rect 10980 699 11194 729
rect 10525 583 10663 613
rect 10399 453 10459 478
rect 10573 453 10663 583
rect 10189 403 10205 437
rect 10239 403 10333 437
rect 10189 387 10333 403
rect 10381 437 10525 453
rect 10381 403 10397 437
rect 10431 403 10525 437
rect 10381 387 10525 403
rect 10573 437 10717 453
rect 10980 452 11010 699
rect 11260 657 11290 762
rect 11356 739 11386 762
rect 11116 519 11290 657
rect 10573 403 10589 437
rect 10623 403 10717 437
rect 10573 387 10717 403
rect -24536 357 -24363 373
rect -24536 322 -24435 357
rect -24401 343 -24363 357
rect -23963 343 -23937 373
rect -23427 357 -23254 373
rect -24401 322 -24385 343
rect -24536 306 -24385 322
rect -23427 322 -23326 357
rect -23292 343 -23254 357
rect -22854 343 -22828 373
rect -22545 357 -22372 373
rect -23292 322 -23276 343
rect -23427 306 -23276 322
rect -22545 322 -22444 357
rect -22410 343 -22372 357
rect -21972 343 -21946 373
rect -21245 357 -21072 373
rect -22410 322 -22394 343
rect -22545 306 -22394 322
rect -21245 322 -21144 357
rect -21110 343 -21072 357
rect -20672 343 -20646 373
rect -20136 357 -19963 373
rect -21110 322 -21094 343
rect -21245 306 -21094 322
rect -20136 322 -20035 357
rect -20001 343 -19963 357
rect -19563 343 -19537 373
rect -19254 357 -19081 373
rect -20001 322 -19985 343
rect -20136 306 -19985 322
rect -19254 322 -19153 357
rect -19119 343 -19081 357
rect -18681 343 -18655 373
rect -17954 357 -17781 373
rect -19119 322 -19103 343
rect -19254 306 -19103 322
rect -17954 322 -17853 357
rect -17819 343 -17781 357
rect -17381 343 -17355 373
rect -16845 357 -16672 373
rect -17819 322 -17803 343
rect -17954 306 -17803 322
rect -16845 322 -16744 357
rect -16710 343 -16672 357
rect -16272 343 -16246 373
rect -15963 357 -15790 373
rect -16710 322 -16694 343
rect -16845 306 -16694 322
rect -15963 322 -15862 357
rect -15828 343 -15790 357
rect -15390 343 -15364 373
rect -14663 357 -14490 373
rect -15828 322 -15812 343
rect -15963 306 -15812 322
rect -14663 322 -14562 357
rect -14528 343 -14490 357
rect -14090 343 -14064 373
rect -13554 357 -13381 373
rect -14528 322 -14512 343
rect -14663 306 -14512 322
rect -13554 322 -13453 357
rect -13419 343 -13381 357
rect -12981 343 -12955 373
rect -12672 357 -12499 373
rect -13419 322 -13403 343
rect -13554 306 -13403 322
rect -12672 322 -12571 357
rect -12537 343 -12499 357
rect -12099 343 -12073 373
rect -11372 357 -11199 373
rect -12537 322 -12521 343
rect -12672 306 -12521 322
rect -11372 322 -11271 357
rect -11237 343 -11199 357
rect -10799 343 -10773 373
rect -10263 357 -10090 373
rect -11237 322 -11221 343
rect -11372 306 -11221 322
rect -10263 322 -10162 357
rect -10128 343 -10090 357
rect -9690 343 -9664 373
rect -9381 357 -9208 373
rect -10128 322 -10112 343
rect -10263 306 -10112 322
rect -9381 322 -9280 357
rect -9246 343 -9208 357
rect -8808 343 -8782 373
rect -8082 357 -7909 373
rect -9246 322 -9230 343
rect -9381 306 -9230 322
rect -8082 322 -7981 357
rect -7947 343 -7909 357
rect -7509 343 -7483 373
rect -6973 357 -6800 373
rect -7947 322 -7931 343
rect -8082 306 -7931 322
rect -6973 322 -6872 357
rect -6838 343 -6800 357
rect -6400 343 -6374 373
rect -6091 357 -5918 373
rect -6838 322 -6822 343
rect -6973 306 -6822 322
rect -6091 322 -5990 357
rect -5956 343 -5918 357
rect -5518 343 -5492 373
rect -4791 357 -4618 373
rect -5956 322 -5940 343
rect -6091 306 -5940 322
rect -4791 322 -4690 357
rect -4656 343 -4618 357
rect -4218 343 -4192 373
rect -3682 357 -3509 373
rect -4656 322 -4640 343
rect -4791 306 -4640 322
rect -3682 322 -3581 357
rect -3547 343 -3509 357
rect -3109 343 -3083 373
rect -2800 357 -2627 373
rect -3547 322 -3531 343
rect -3682 306 -3531 322
rect -2800 322 -2699 357
rect -2665 343 -2627 357
rect -2227 343 -2201 373
rect -1500 357 -1327 373
rect -2665 322 -2649 343
rect -2800 306 -2649 322
rect -1500 322 -1399 357
rect -1365 343 -1327 357
rect -927 343 -901 373
rect -391 357 -218 373
rect -1365 322 -1349 343
rect -1500 306 -1349 322
rect -391 322 -290 357
rect -256 343 -218 357
rect 182 343 208 373
rect 491 357 664 373
rect -256 322 -240 343
rect -391 306 -240 322
rect 491 322 592 357
rect 626 343 664 357
rect 1064 343 1090 373
rect 7200 355 7230 386
rect 7296 355 7326 386
rect 7392 355 7422 386
rect 7488 355 7518 386
rect 7584 355 7614 386
rect 7680 355 7710 386
rect 7776 355 7806 386
rect 7872 355 7902 386
rect 8148 355 8178 386
rect 8244 355 8274 386
rect 8340 355 8370 386
rect 8436 355 8466 386
rect 8532 355 8562 386
rect 8628 355 8658 386
rect 8724 355 8754 386
rect 8820 355 8850 386
rect 9084 355 9114 386
rect 9180 355 9210 386
rect 9276 355 9306 386
rect 9372 355 9402 386
rect 9468 355 9498 386
rect 9564 355 9594 386
rect 9660 355 9690 386
rect 9756 355 9786 386
rect 10015 356 10045 387
rect 10111 356 10141 387
rect 10207 356 10237 387
rect 10303 356 10333 387
rect 10399 356 10429 387
rect 10495 356 10525 387
rect 10591 356 10621 387
rect 10687 356 10717 387
rect 10924 436 11068 452
rect 10924 402 10940 436
rect 10974 402 11068 436
rect 10924 386 11068 402
rect 11116 436 11260 519
rect 11332 477 11386 739
rect 11452 612 11482 762
rect 11452 582 11590 612
rect 11326 452 11386 477
rect 11500 452 11590 582
rect 11116 402 11132 436
rect 11166 402 11260 436
rect 11116 386 11260 402
rect 11308 436 11452 452
rect 11308 402 11324 436
rect 11358 402 11452 436
rect 11308 386 11452 402
rect 11500 436 11644 452
rect 11500 402 11516 436
rect 11550 402 11644 436
rect 11500 386 11644 402
rect 626 322 642 343
rect 491 306 642 322
rect 10942 355 10972 386
rect 11038 355 11068 386
rect 11134 355 11164 386
rect 11230 355 11260 386
rect 11326 355 11356 386
rect 11422 355 11452 386
rect 11518 355 11548 386
rect 11614 355 11644 386
rect 7200 7 7230 33
rect 7296 7 7326 33
rect 7392 7 7422 33
rect 7488 7 7518 33
rect 7584 7 7614 33
rect 7680 7 7710 33
rect 7776 7 7806 33
rect 7872 7 7902 33
rect 8148 7 8178 33
rect 8244 7 8274 33
rect 8340 7 8370 33
rect 8436 7 8466 33
rect 8532 7 8562 33
rect 8628 7 8658 33
rect 8724 7 8754 33
rect 8820 7 8850 33
rect 9084 7 9114 33
rect 9180 7 9210 33
rect 9276 7 9306 33
rect 9372 7 9402 33
rect 9468 7 9498 33
rect 9564 7 9594 33
rect 9660 7 9690 33
rect 9756 7 9786 33
rect 10015 8 10045 34
rect 10111 8 10141 34
rect 10207 8 10237 34
rect 10303 8 10333 34
rect 10399 8 10429 34
rect 10495 8 10525 34
rect 10591 8 10621 34
rect 10687 8 10717 34
rect 10942 7 10972 33
rect 11038 7 11068 33
rect 11134 7 11164 33
rect 11230 7 11260 33
rect 11326 7 11356 33
rect 11422 7 11452 33
rect 11518 7 11548 33
rect 11614 7 11644 33
rect 5561 -665 5627 -649
rect 5561 -891 5577 -665
rect 5611 -667 5627 -665
rect 6001 -665 6067 -649
rect 5611 -697 5658 -667
rect 5872 -697 5898 -667
rect 5611 -763 5627 -697
rect 5611 -793 5658 -763
rect 5872 -793 5898 -763
rect 5611 -859 5627 -793
rect 5611 -889 5658 -859
rect 5872 -889 5898 -859
rect 5611 -891 5627 -889
rect 5561 -907 5627 -891
rect 6001 -891 6017 -665
rect 6051 -667 6067 -665
rect 6441 -665 6507 -649
rect 6051 -697 6098 -667
rect 6312 -697 6338 -667
rect 6051 -763 6067 -697
rect 6051 -793 6098 -763
rect 6312 -793 6338 -763
rect 6051 -859 6067 -793
rect 6051 -889 6098 -859
rect 6312 -889 6338 -859
rect 6051 -891 6067 -889
rect 6001 -907 6067 -891
rect 6441 -891 6457 -665
rect 6491 -667 6507 -665
rect 6491 -697 6538 -667
rect 6752 -697 6778 -667
rect 6491 -763 6507 -697
rect 6491 -793 6538 -763
rect 6752 -793 6778 -763
rect 6491 -859 6507 -793
rect 6491 -889 6538 -859
rect 6752 -889 6778 -859
rect 6491 -891 6507 -889
rect 6441 -907 6507 -891
rect 5561 -1111 5628 -1095
rect 5561 -1145 5577 -1111
rect 5611 -1113 5628 -1111
rect 6001 -1111 6068 -1095
rect 5611 -1143 5658 -1113
rect 5858 -1143 5884 -1113
rect 5611 -1145 5628 -1143
rect 5561 -1161 5628 -1145
rect 6001 -1145 6017 -1111
rect 6051 -1113 6068 -1111
rect 6441 -1111 6508 -1095
rect 6051 -1143 6098 -1113
rect 6298 -1143 6324 -1113
rect 6051 -1145 6068 -1143
rect 6001 -1161 6068 -1145
rect 6441 -1145 6457 -1111
rect 6491 -1113 6508 -1111
rect 6491 -1143 6538 -1113
rect 6738 -1143 6764 -1113
rect 6491 -1145 6508 -1143
rect 6441 -1161 6508 -1145
rect 7200 -1309 7230 -1283
rect 7296 -1309 7326 -1283
rect 7392 -1309 7422 -1283
rect 7488 -1309 7518 -1283
rect 7584 -1309 7614 -1283
rect 7680 -1309 7710 -1283
rect 7776 -1309 7806 -1283
rect 7872 -1309 7902 -1283
rect 8148 -1309 8178 -1283
rect 8244 -1309 8274 -1283
rect 8340 -1309 8370 -1283
rect 8436 -1309 8466 -1283
rect 8532 -1309 8562 -1283
rect 8628 -1309 8658 -1283
rect 8724 -1309 8754 -1283
rect 8820 -1309 8850 -1283
rect 9084 -1309 9114 -1283
rect 9180 -1309 9210 -1283
rect 9276 -1309 9306 -1283
rect 9372 -1309 9402 -1283
rect 9468 -1309 9498 -1283
rect 9564 -1309 9594 -1283
rect 9660 -1309 9690 -1283
rect 9756 -1309 9786 -1283
rect 10015 -1309 10045 -1283
rect 10111 -1309 10141 -1283
rect 10207 -1309 10237 -1283
rect 10303 -1309 10333 -1283
rect 10399 -1309 10429 -1283
rect 10495 -1309 10525 -1283
rect 10591 -1309 10621 -1283
rect 10687 -1309 10717 -1283
rect 10942 -1309 10972 -1283
rect 11038 -1309 11068 -1283
rect 11134 -1309 11164 -1283
rect 11230 -1309 11260 -1283
rect 11326 -1309 11356 -1283
rect 11422 -1309 11452 -1283
rect 11518 -1309 11548 -1283
rect 11614 -1309 11644 -1283
rect 7200 -1662 7230 -1631
rect 7296 -1662 7326 -1631
rect 7392 -1662 7422 -1631
rect 7488 -1662 7518 -1631
rect 7584 -1662 7614 -1631
rect 7680 -1662 7710 -1631
rect 7776 -1662 7806 -1631
rect 7872 -1662 7902 -1631
rect 8148 -1662 8178 -1631
rect 8244 -1662 8274 -1631
rect 8340 -1662 8370 -1631
rect 8436 -1662 8466 -1631
rect 8532 -1662 8562 -1631
rect 8628 -1662 8658 -1631
rect 8724 -1662 8754 -1631
rect 8820 -1662 8850 -1631
rect 9084 -1662 9114 -1631
rect 9180 -1662 9210 -1631
rect 9276 -1662 9306 -1631
rect 9372 -1662 9402 -1631
rect 9468 -1662 9498 -1631
rect 9564 -1662 9594 -1631
rect 9660 -1662 9690 -1631
rect 9756 -1662 9786 -1631
rect 10015 -1662 10045 -1631
rect 10111 -1662 10141 -1631
rect 10207 -1662 10237 -1631
rect 10303 -1662 10333 -1631
rect 10399 -1662 10429 -1631
rect 10495 -1662 10525 -1631
rect 10591 -1662 10621 -1631
rect 10687 -1662 10717 -1631
rect 10942 -1662 10972 -1631
rect 11038 -1662 11068 -1631
rect 11134 -1662 11164 -1631
rect 11230 -1662 11260 -1631
rect 11326 -1662 11356 -1631
rect 11422 -1662 11452 -1631
rect 11518 -1662 11548 -1631
rect 11614 -1662 11644 -1631
rect 7182 -1678 7326 -1662
rect 7182 -1712 7198 -1678
rect 7232 -1712 7326 -1678
rect 7182 -1728 7326 -1712
rect 7374 -1678 7518 -1662
rect 7374 -1712 7390 -1678
rect 7424 -1712 7518 -1678
rect 7238 -1975 7268 -1728
rect 7374 -1795 7518 -1712
rect 7566 -1678 7710 -1662
rect 7566 -1712 7582 -1678
rect 7616 -1712 7710 -1678
rect 7566 -1728 7710 -1712
rect 7758 -1678 7902 -1662
rect 7758 -1712 7774 -1678
rect 7808 -1712 7902 -1678
rect 7758 -1728 7902 -1712
rect 8130 -1678 8274 -1662
rect 8130 -1712 8146 -1678
rect 8180 -1712 8274 -1678
rect 8130 -1728 8274 -1712
rect 8322 -1678 8466 -1662
rect 8322 -1712 8338 -1678
rect 8372 -1712 8466 -1678
rect 7584 -1753 7644 -1728
rect 7374 -1933 7548 -1795
rect 7238 -2005 7452 -1975
rect 7422 -2038 7452 -2005
rect 7518 -2038 7548 -1933
rect 7590 -2015 7644 -1753
rect 7758 -1858 7848 -1728
rect 7614 -2038 7644 -2015
rect 7710 -1888 7848 -1858
rect 7710 -2038 7740 -1888
rect 8186 -1975 8216 -1728
rect 8322 -1795 8466 -1712
rect 8514 -1678 8658 -1662
rect 8514 -1712 8530 -1678
rect 8564 -1712 8658 -1678
rect 8514 -1728 8658 -1712
rect 8706 -1678 8850 -1662
rect 8706 -1712 8722 -1678
rect 8756 -1712 8850 -1678
rect 8706 -1728 8850 -1712
rect 9066 -1678 9210 -1662
rect 9066 -1712 9082 -1678
rect 9116 -1712 9210 -1678
rect 9066 -1728 9210 -1712
rect 9258 -1678 9402 -1662
rect 9258 -1712 9274 -1678
rect 9308 -1712 9402 -1678
rect 8532 -1753 8592 -1728
rect 8322 -1933 8496 -1795
rect 8186 -2005 8400 -1975
rect 8370 -2038 8400 -2005
rect 8466 -2038 8496 -1933
rect 8538 -2015 8592 -1753
rect 8706 -1858 8796 -1728
rect 8562 -2038 8592 -2015
rect 8658 -1888 8796 -1858
rect 8658 -2038 8688 -1888
rect 9122 -1975 9152 -1728
rect 9258 -1795 9402 -1712
rect 9450 -1678 9594 -1662
rect 9450 -1712 9466 -1678
rect 9500 -1712 9594 -1678
rect 9450 -1728 9594 -1712
rect 9642 -1678 9786 -1662
rect 9642 -1712 9658 -1678
rect 9692 -1712 9786 -1678
rect 9642 -1728 9786 -1712
rect 9997 -1678 10141 -1662
rect 9997 -1712 10013 -1678
rect 10047 -1712 10141 -1678
rect 9997 -1728 10141 -1712
rect 10189 -1678 10333 -1662
rect 10189 -1712 10205 -1678
rect 10239 -1712 10333 -1678
rect 9468 -1753 9528 -1728
rect 9258 -1933 9432 -1795
rect 9122 -2005 9336 -1975
rect 9306 -2038 9336 -2005
rect 9402 -2038 9432 -1933
rect 9474 -2015 9528 -1753
rect 9642 -1858 9732 -1728
rect 9498 -2038 9528 -2015
rect 9594 -1888 9732 -1858
rect 9594 -2038 9624 -1888
rect 10053 -1975 10083 -1728
rect 10189 -1795 10333 -1712
rect 10381 -1678 10525 -1662
rect 10381 -1712 10397 -1678
rect 10431 -1712 10525 -1678
rect 10381 -1728 10525 -1712
rect 10573 -1678 10717 -1662
rect 10573 -1712 10589 -1678
rect 10623 -1712 10717 -1678
rect 10573 -1728 10717 -1712
rect 10924 -1678 11068 -1662
rect 10924 -1712 10940 -1678
rect 10974 -1712 11068 -1678
rect 10924 -1728 11068 -1712
rect 11116 -1678 11260 -1662
rect 11116 -1712 11132 -1678
rect 11166 -1712 11260 -1678
rect 10399 -1753 10459 -1728
rect 10189 -1933 10363 -1795
rect 10053 -2005 10267 -1975
rect 10237 -2038 10267 -2005
rect 10333 -2038 10363 -1933
rect 10405 -2015 10459 -1753
rect 10573 -1858 10663 -1728
rect 10429 -2038 10459 -2015
rect 10525 -1888 10663 -1858
rect 10525 -2038 10555 -1888
rect 10980 -1975 11010 -1728
rect 11116 -1795 11260 -1712
rect 11308 -1678 11452 -1662
rect 11308 -1712 11324 -1678
rect 11358 -1712 11452 -1678
rect 11308 -1728 11452 -1712
rect 11500 -1678 11644 -1662
rect 11500 -1712 11516 -1678
rect 11550 -1712 11644 -1678
rect 11500 -1728 11644 -1712
rect 11326 -1753 11386 -1728
rect 11116 -1933 11290 -1795
rect 10980 -2005 11194 -1975
rect 11164 -2038 11194 -2005
rect 11260 -2038 11290 -1933
rect 11332 -2015 11386 -1753
rect 11500 -1858 11590 -1728
rect 11356 -2038 11386 -2015
rect 11452 -1888 11590 -1858
rect 11452 -2038 11482 -1888
rect -23725 -2367 -23659 -2351
rect -24385 -2413 -24355 -2382
rect -24289 -2413 -24259 -2382
rect -24193 -2413 -24163 -2382
rect -24097 -2413 -24067 -2382
rect -24001 -2413 -23971 -2382
rect -23905 -2413 -23875 -2382
rect -23725 -2593 -23709 -2367
rect -23675 -2369 -23659 -2367
rect -21705 -2367 -21639 -2351
rect -23675 -2399 -23628 -2369
rect -23414 -2399 -23388 -2369
rect -23675 -2465 -23659 -2399
rect -22348 -2413 -22318 -2382
rect -22252 -2413 -22222 -2382
rect -22156 -2413 -22126 -2382
rect -22060 -2413 -22030 -2382
rect -21964 -2413 -21934 -2382
rect -21868 -2413 -21838 -2382
rect -23675 -2495 -23628 -2465
rect -23414 -2495 -23388 -2465
rect -23675 -2561 -23659 -2495
rect -23675 -2591 -23628 -2561
rect -23414 -2591 -23388 -2561
rect -23675 -2593 -23659 -2591
rect -23725 -2609 -23659 -2593
rect -24385 -2653 -24355 -2627
rect -24289 -2653 -24259 -2627
rect -24193 -2653 -24163 -2627
rect -24386 -2674 -24163 -2653
rect -24386 -2709 -24369 -2674
rect -24335 -2683 -24163 -2674
rect -24097 -2653 -24067 -2627
rect -24001 -2653 -23971 -2627
rect -23905 -2653 -23875 -2627
rect -21705 -2593 -21689 -2367
rect -21655 -2369 -21639 -2367
rect -19964 -2367 -19898 -2351
rect -21655 -2399 -21608 -2369
rect -21394 -2399 -21368 -2369
rect -21655 -2465 -21639 -2399
rect -20618 -2413 -20588 -2382
rect -20522 -2413 -20492 -2382
rect -20426 -2413 -20396 -2382
rect -20330 -2413 -20300 -2382
rect -20234 -2413 -20204 -2382
rect -20138 -2413 -20108 -2382
rect -21655 -2495 -21608 -2465
rect -21394 -2495 -21368 -2465
rect -21655 -2561 -21639 -2495
rect -21655 -2591 -21608 -2561
rect -21394 -2591 -21368 -2561
rect -21655 -2593 -21639 -2591
rect -21705 -2609 -21639 -2593
rect -22348 -2653 -22318 -2627
rect -22252 -2653 -22222 -2627
rect -22156 -2653 -22126 -2627
rect -24097 -2674 -23875 -2653
rect -24335 -2709 -24319 -2683
rect -24386 -2720 -24319 -2709
rect -24097 -2709 -24080 -2674
rect -24046 -2683 -23875 -2674
rect -22349 -2674 -22126 -2653
rect -24046 -2709 -24030 -2683
rect -24097 -2720 -24030 -2709
rect -22349 -2709 -22332 -2674
rect -22298 -2683 -22126 -2674
rect -22060 -2653 -22030 -2627
rect -21964 -2653 -21934 -2627
rect -21868 -2653 -21838 -2627
rect -19964 -2593 -19948 -2367
rect -19914 -2369 -19898 -2367
rect -18185 -2367 -18119 -2351
rect -19914 -2399 -19867 -2369
rect -19653 -2399 -19627 -2369
rect -19914 -2465 -19898 -2399
rect -18858 -2413 -18828 -2382
rect -18762 -2413 -18732 -2382
rect -18666 -2413 -18636 -2382
rect -18570 -2413 -18540 -2382
rect -18474 -2413 -18444 -2382
rect -18378 -2413 -18348 -2382
rect -19914 -2495 -19867 -2465
rect -19653 -2495 -19627 -2465
rect -19914 -2561 -19898 -2495
rect -19914 -2591 -19867 -2561
rect -19653 -2591 -19627 -2561
rect -19914 -2593 -19898 -2591
rect -19964 -2609 -19898 -2593
rect -20618 -2653 -20588 -2627
rect -20522 -2653 -20492 -2627
rect -20426 -2653 -20396 -2627
rect -22060 -2674 -21838 -2653
rect -22298 -2709 -22282 -2683
rect -22349 -2720 -22282 -2709
rect -22060 -2709 -22043 -2674
rect -22009 -2683 -21838 -2674
rect -20619 -2674 -20396 -2653
rect -22009 -2709 -21993 -2683
rect -22060 -2720 -21993 -2709
rect -20619 -2709 -20602 -2674
rect -20568 -2683 -20396 -2674
rect -20330 -2653 -20300 -2627
rect -20234 -2653 -20204 -2627
rect -20138 -2653 -20108 -2627
rect -18185 -2593 -18169 -2367
rect -18135 -2369 -18119 -2367
rect -18135 -2399 -18088 -2369
rect -17874 -2399 -17848 -2369
rect -18135 -2465 -18119 -2399
rect -18135 -2495 -18088 -2465
rect -17874 -2495 -17848 -2465
rect -18135 -2561 -18119 -2495
rect -18135 -2591 -18088 -2561
rect -17874 -2591 -17848 -2561
rect -18135 -2593 -18119 -2591
rect -18185 -2609 -18119 -2593
rect -18858 -2653 -18828 -2627
rect -18762 -2653 -18732 -2627
rect -18666 -2653 -18636 -2627
rect -20330 -2674 -20108 -2653
rect -20568 -2709 -20552 -2683
rect -20619 -2720 -20552 -2709
rect -20330 -2709 -20313 -2674
rect -20279 -2683 -20108 -2674
rect -18859 -2674 -18636 -2653
rect -20279 -2709 -20263 -2683
rect -20330 -2720 -20263 -2709
rect -18859 -2709 -18842 -2674
rect -18808 -2683 -18636 -2674
rect -18570 -2653 -18540 -2627
rect -18474 -2653 -18444 -2627
rect -18378 -2653 -18348 -2627
rect -18570 -2674 -18348 -2653
rect -18808 -2709 -18792 -2683
rect -18859 -2720 -18792 -2709
rect -18570 -2709 -18553 -2674
rect -18519 -2683 -18348 -2674
rect -18519 -2709 -18503 -2683
rect -18570 -2720 -18503 -2709
rect -24386 -2915 -24343 -2720
rect -24301 -2798 -24235 -2782
rect -24301 -2833 -24285 -2798
rect -24251 -2819 -24235 -2798
rect -23725 -2813 -23658 -2797
rect -24251 -2833 -24213 -2819
rect -24301 -2849 -24213 -2833
rect -23813 -2849 -23787 -2819
rect -23725 -2847 -23709 -2813
rect -23675 -2815 -23658 -2813
rect -23675 -2845 -23628 -2815
rect -23428 -2845 -23402 -2815
rect -23675 -2847 -23658 -2845
rect -23725 -2863 -23658 -2847
rect -22349 -2915 -22306 -2720
rect -22264 -2798 -22198 -2782
rect -22264 -2833 -22248 -2798
rect -22214 -2819 -22198 -2798
rect -21705 -2813 -21638 -2797
rect -22214 -2833 -22176 -2819
rect -22264 -2849 -22176 -2833
rect -21776 -2849 -21750 -2819
rect -21705 -2847 -21689 -2813
rect -21655 -2815 -21638 -2813
rect -21655 -2845 -21608 -2815
rect -21408 -2845 -21382 -2815
rect -21655 -2847 -21638 -2845
rect -21705 -2863 -21638 -2847
rect -20619 -2915 -20576 -2720
rect -20534 -2798 -20468 -2782
rect -20534 -2833 -20518 -2798
rect -20484 -2819 -20468 -2798
rect -19964 -2813 -19897 -2797
rect -20484 -2833 -20446 -2819
rect -20534 -2849 -20446 -2833
rect -20046 -2849 -20020 -2819
rect -19964 -2847 -19948 -2813
rect -19914 -2815 -19897 -2813
rect -19914 -2845 -19867 -2815
rect -19667 -2845 -19641 -2815
rect -19914 -2847 -19897 -2845
rect -19964 -2863 -19897 -2847
rect -18859 -2915 -18816 -2720
rect -18774 -2798 -18708 -2782
rect -18774 -2833 -18758 -2798
rect -18724 -2819 -18708 -2798
rect -18185 -2813 -18118 -2797
rect -18724 -2833 -18686 -2819
rect -18774 -2849 -18686 -2833
rect -18286 -2849 -18260 -2819
rect -18185 -2847 -18169 -2813
rect -18135 -2815 -18118 -2813
rect -18135 -2845 -18088 -2815
rect -17888 -2845 -17862 -2815
rect 11835 -2519 11865 -2493
rect 11931 -2519 11961 -2493
rect 12027 -2519 12057 -2493
rect 12123 -2519 12153 -2493
rect 12219 -2519 12249 -2493
rect 12315 -2519 12345 -2493
rect 12411 -2519 12441 -2493
rect 12507 -2519 12537 -2493
rect 12603 -2519 12633 -2493
rect 12699 -2519 12729 -2493
rect 12826 -2683 12892 -2667
rect 11835 -2801 11865 -2775
rect 11931 -2801 11961 -2775
rect 12027 -2801 12057 -2775
rect 12123 -2801 12153 -2775
rect 12219 -2801 12249 -2775
rect 11835 -2825 12249 -2801
rect -18135 -2847 -18118 -2845
rect -18185 -2863 -18118 -2847
rect 7422 -2864 7452 -2838
rect 7518 -2864 7548 -2838
rect 7614 -2864 7644 -2838
rect 7710 -2864 7740 -2838
rect 8370 -2864 8400 -2838
rect 8466 -2864 8496 -2838
rect 8562 -2864 8592 -2838
rect 8658 -2864 8688 -2838
rect 9306 -2864 9336 -2838
rect 9402 -2864 9432 -2838
rect 9498 -2864 9528 -2838
rect 9594 -2864 9624 -2838
rect 10237 -2864 10267 -2838
rect 10333 -2864 10363 -2838
rect 10429 -2864 10459 -2838
rect 10525 -2864 10555 -2838
rect 11164 -2864 11194 -2838
rect 11260 -2864 11290 -2838
rect 11356 -2864 11386 -2838
rect 11452 -2864 11482 -2838
rect 11835 -2859 12170 -2825
rect 12204 -2859 12249 -2825
rect 11835 -2872 12249 -2859
rect -24386 -2931 -24213 -2915
rect -24386 -2966 -24285 -2931
rect -24251 -2945 -24213 -2931
rect -23813 -2945 -23787 -2915
rect -22349 -2931 -22176 -2915
rect -24251 -2966 -24235 -2945
rect -24386 -2982 -24235 -2966
rect -22349 -2966 -22248 -2931
rect -22214 -2945 -22176 -2931
rect -21776 -2945 -21750 -2915
rect -20619 -2931 -20446 -2915
rect -22214 -2966 -22198 -2945
rect -22349 -2982 -22198 -2966
rect -20619 -2966 -20518 -2931
rect -20484 -2945 -20446 -2931
rect -20046 -2945 -20020 -2915
rect -18859 -2931 -18686 -2915
rect -20484 -2966 -20468 -2945
rect -20619 -2982 -20468 -2966
rect -18859 -2966 -18758 -2931
rect -18724 -2945 -18686 -2931
rect -18286 -2945 -18260 -2915
rect -18724 -2966 -18708 -2945
rect -18859 -2982 -18708 -2966
rect 7422 -2966 7452 -2940
rect 7518 -2966 7548 -2940
rect 7614 -2966 7644 -2940
rect 7710 -2966 7740 -2940
rect 8370 -2966 8400 -2940
rect 8466 -2966 8496 -2940
rect 8562 -2966 8592 -2940
rect 8658 -2966 8688 -2940
rect 9306 -2966 9336 -2940
rect 9402 -2966 9432 -2940
rect 9498 -2966 9528 -2940
rect 9594 -2966 9624 -2940
rect 10237 -2965 10267 -2939
rect 10333 -2965 10363 -2939
rect 10429 -2965 10459 -2939
rect 10525 -2965 10555 -2939
rect 11164 -2966 11194 -2940
rect 11260 -2966 11290 -2940
rect 11356 -2966 11386 -2940
rect 11452 -2966 11482 -2940
rect 7422 -3799 7452 -3766
rect 7238 -3829 7452 -3799
rect -20679 -3984 -20649 -3958
rect -20587 -3984 -20557 -3953
rect -20491 -3984 -20461 -3953
rect -20395 -3984 -20365 -3953
rect -20299 -3984 -20269 -3953
rect -20203 -3984 -20173 -3953
rect -20107 -3984 -20077 -3953
rect -20011 -3984 -19981 -3953
rect -19915 -3984 -19885 -3953
rect -19819 -3984 -19789 -3953
rect -19723 -3984 -19693 -3953
rect -19627 -3984 -19597 -3953
rect -19531 -3984 -19501 -3953
rect -19439 -3984 -19409 -3958
rect -19120 -3984 -19090 -3958
rect -19028 -3984 -18998 -3953
rect -18932 -3984 -18902 -3953
rect -18836 -3984 -18806 -3953
rect -18740 -3984 -18710 -3953
rect -18644 -3984 -18614 -3953
rect -18548 -3984 -18518 -3953
rect -18452 -3984 -18422 -3953
rect -18356 -3984 -18326 -3953
rect -18260 -3984 -18230 -3953
rect -18164 -3984 -18134 -3953
rect -18068 -3984 -18038 -3953
rect -17972 -3984 -17942 -3953
rect -17880 -3984 -17850 -3958
rect -17388 -3984 -17358 -3958
rect -17296 -3984 -17266 -3953
rect -17200 -3984 -17170 -3953
rect -17104 -3984 -17074 -3953
rect -17008 -3984 -16978 -3953
rect -16912 -3984 -16882 -3953
rect -16816 -3984 -16786 -3953
rect -16720 -3984 -16690 -3953
rect -16624 -3984 -16594 -3953
rect -16528 -3984 -16498 -3953
rect -16432 -3984 -16402 -3953
rect -16336 -3984 -16306 -3953
rect -16240 -3984 -16210 -3953
rect -16148 -3984 -16118 -3958
rect -15829 -3984 -15799 -3958
rect -15737 -3984 -15707 -3953
rect -15641 -3984 -15611 -3953
rect -15545 -3984 -15515 -3953
rect -15449 -3984 -15419 -3953
rect -15353 -3984 -15323 -3953
rect -15257 -3984 -15227 -3953
rect -15161 -3984 -15131 -3953
rect -15065 -3984 -15035 -3953
rect -14969 -3984 -14939 -3953
rect -14873 -3984 -14843 -3953
rect -14777 -3984 -14747 -3953
rect -14681 -3984 -14651 -3953
rect -14589 -3984 -14559 -3958
rect -14097 -3984 -14067 -3958
rect -14005 -3984 -13975 -3953
rect -13909 -3984 -13879 -3953
rect -13813 -3984 -13783 -3953
rect -13717 -3984 -13687 -3953
rect -13621 -3984 -13591 -3953
rect -13525 -3984 -13495 -3953
rect -13429 -3984 -13399 -3953
rect -13333 -3984 -13303 -3953
rect -13237 -3984 -13207 -3953
rect -13141 -3984 -13111 -3953
rect -13045 -3984 -13015 -3953
rect -12949 -3984 -12919 -3953
rect -12857 -3984 -12827 -3958
rect -12538 -3984 -12508 -3958
rect -12446 -3984 -12416 -3953
rect -12350 -3984 -12320 -3953
rect -12254 -3984 -12224 -3953
rect -12158 -3984 -12128 -3953
rect -12062 -3984 -12032 -3953
rect -11966 -3984 -11936 -3953
rect -11870 -3984 -11840 -3953
rect -11774 -3984 -11744 -3953
rect -11678 -3984 -11648 -3953
rect -11582 -3984 -11552 -3953
rect -11486 -3984 -11456 -3953
rect -11390 -3984 -11360 -3953
rect -11298 -3984 -11268 -3958
rect -10806 -3984 -10776 -3958
rect -10714 -3984 -10684 -3953
rect -10618 -3984 -10588 -3953
rect -10522 -3984 -10492 -3953
rect -10426 -3984 -10396 -3953
rect -10330 -3984 -10300 -3953
rect -10234 -3984 -10204 -3953
rect -10138 -3984 -10108 -3953
rect -10042 -3984 -10012 -3953
rect -9946 -3984 -9916 -3953
rect -9850 -3984 -9820 -3953
rect -9754 -3984 -9724 -3953
rect -9658 -3984 -9628 -3953
rect -9566 -3984 -9536 -3958
rect -9247 -3984 -9217 -3958
rect -9155 -3984 -9125 -3953
rect -9059 -3984 -9029 -3953
rect -8963 -3984 -8933 -3953
rect -8867 -3984 -8837 -3953
rect -8771 -3984 -8741 -3953
rect -8675 -3984 -8645 -3953
rect -8579 -3984 -8549 -3953
rect -8483 -3984 -8453 -3953
rect -8387 -3984 -8357 -3953
rect -8291 -3984 -8261 -3953
rect -8195 -3984 -8165 -3953
rect -8099 -3984 -8069 -3953
rect -8007 -3984 -7977 -3958
rect -23681 -4179 -23615 -4163
rect -24334 -4225 -24304 -4194
rect -24238 -4225 -24208 -4194
rect -24142 -4225 -24112 -4194
rect -24046 -4225 -24016 -4194
rect -23950 -4225 -23920 -4194
rect -23854 -4225 -23824 -4194
rect -23681 -4405 -23665 -4179
rect -23631 -4181 -23615 -4179
rect -21943 -4179 -21877 -4163
rect -23631 -4211 -23584 -4181
rect -23370 -4211 -23344 -4181
rect -23631 -4277 -23615 -4211
rect -22598 -4225 -22568 -4194
rect -22502 -4225 -22472 -4194
rect -22406 -4225 -22376 -4194
rect -22310 -4225 -22280 -4194
rect -22214 -4225 -22184 -4194
rect -22118 -4225 -22088 -4194
rect -23631 -4307 -23584 -4277
rect -23370 -4307 -23344 -4277
rect -23631 -4373 -23615 -4307
rect -23631 -4403 -23584 -4373
rect -23370 -4403 -23344 -4373
rect -23631 -4405 -23615 -4403
rect -23681 -4421 -23615 -4405
rect -24334 -4465 -24304 -4439
rect -24238 -4465 -24208 -4439
rect -24142 -4465 -24112 -4439
rect -24335 -4486 -24112 -4465
rect -24335 -4521 -24318 -4486
rect -24284 -4495 -24112 -4486
rect -24046 -4465 -24016 -4439
rect -23950 -4465 -23920 -4439
rect -23854 -4465 -23824 -4439
rect -21943 -4405 -21927 -4179
rect -21893 -4181 -21877 -4179
rect -21893 -4211 -21846 -4181
rect -21632 -4211 -21606 -4181
rect -21893 -4277 -21877 -4211
rect -21893 -4307 -21846 -4277
rect -21632 -4307 -21606 -4277
rect -21893 -4373 -21877 -4307
rect -21893 -4403 -21846 -4373
rect -21632 -4403 -21606 -4373
rect -21893 -4405 -21877 -4403
rect -21943 -4421 -21877 -4405
rect -22598 -4465 -22568 -4439
rect -22502 -4465 -22472 -4439
rect -22406 -4465 -22376 -4439
rect -24046 -4486 -23824 -4465
rect -24284 -4521 -24268 -4495
rect -24335 -4532 -24268 -4521
rect -24046 -4521 -24029 -4486
rect -23995 -4495 -23824 -4486
rect -22599 -4486 -22376 -4465
rect -23995 -4521 -23979 -4495
rect -24046 -4532 -23979 -4521
rect -22599 -4521 -22582 -4486
rect -22548 -4495 -22376 -4486
rect -22310 -4465 -22280 -4439
rect -22214 -4465 -22184 -4439
rect -22118 -4465 -22088 -4439
rect -22310 -4486 -22088 -4465
rect -22548 -4521 -22532 -4495
rect -22599 -4532 -22532 -4521
rect -22310 -4521 -22293 -4486
rect -22259 -4495 -22088 -4486
rect -22259 -4521 -22243 -4495
rect -22310 -4532 -22243 -4521
rect -24335 -4727 -24292 -4532
rect -24250 -4610 -24184 -4594
rect -24250 -4645 -24234 -4610
rect -24200 -4631 -24184 -4610
rect -23681 -4625 -23614 -4609
rect -24200 -4645 -24162 -4631
rect -24250 -4661 -24162 -4645
rect -23762 -4661 -23736 -4631
rect -23681 -4659 -23665 -4625
rect -23631 -4627 -23614 -4625
rect -23631 -4657 -23584 -4627
rect -23384 -4657 -23358 -4627
rect -23631 -4659 -23614 -4657
rect -23681 -4675 -23614 -4659
rect -22599 -4727 -22556 -4532
rect 7238 -4076 7268 -3829
rect 7518 -3871 7548 -3766
rect 7614 -3789 7644 -3766
rect 7374 -4009 7548 -3871
rect 7182 -4092 7326 -4076
rect 7182 -4126 7198 -4092
rect 7232 -4126 7326 -4092
rect 7182 -4142 7326 -4126
rect 7374 -4092 7518 -4009
rect 7590 -4051 7644 -3789
rect 7710 -3916 7740 -3766
rect 8370 -3799 8400 -3766
rect 8186 -3829 8400 -3799
rect 7710 -3946 7848 -3916
rect 7584 -4076 7644 -4051
rect 7758 -4076 7848 -3946
rect 8186 -4076 8216 -3829
rect 8466 -3871 8496 -3766
rect 8562 -3789 8592 -3766
rect 8322 -4009 8496 -3871
rect 7374 -4126 7390 -4092
rect 7424 -4126 7518 -4092
rect 7374 -4142 7518 -4126
rect 7566 -4092 7710 -4076
rect 7566 -4126 7582 -4092
rect 7616 -4126 7710 -4092
rect 7566 -4142 7710 -4126
rect 7758 -4092 7902 -4076
rect 7758 -4126 7774 -4092
rect 7808 -4126 7902 -4092
rect 7758 -4142 7902 -4126
rect 8130 -4092 8274 -4076
rect 8130 -4126 8146 -4092
rect 8180 -4126 8274 -4092
rect 8130 -4142 8274 -4126
rect 8322 -4092 8466 -4009
rect 8538 -4051 8592 -3789
rect 8658 -3916 8688 -3766
rect 9306 -3799 9336 -3766
rect 9122 -3829 9336 -3799
rect 8658 -3946 8796 -3916
rect 8532 -4076 8592 -4051
rect 8706 -4076 8796 -3946
rect 9122 -4076 9152 -3829
rect 9402 -3871 9432 -3766
rect 9498 -3789 9528 -3766
rect 9258 -4009 9432 -3871
rect 8322 -4126 8338 -4092
rect 8372 -4126 8466 -4092
rect 8322 -4142 8466 -4126
rect 8514 -4092 8658 -4076
rect 8514 -4126 8530 -4092
rect 8564 -4126 8658 -4092
rect 8514 -4142 8658 -4126
rect 8706 -4092 8850 -4076
rect 8706 -4126 8722 -4092
rect 8756 -4126 8850 -4092
rect 8706 -4142 8850 -4126
rect 9066 -4092 9210 -4076
rect 9066 -4126 9082 -4092
rect 9116 -4126 9210 -4092
rect 9066 -4142 9210 -4126
rect 9258 -4092 9402 -4009
rect 9474 -4051 9528 -3789
rect 9594 -3916 9624 -3766
rect 10237 -3798 10267 -3765
rect 10053 -3828 10267 -3798
rect 9594 -3946 9732 -3916
rect 9468 -4076 9528 -4051
rect 9642 -4076 9732 -3946
rect 10053 -4075 10083 -3828
rect 10333 -3870 10363 -3765
rect 10429 -3788 10459 -3765
rect 10189 -4008 10363 -3870
rect 9258 -4126 9274 -4092
rect 9308 -4126 9402 -4092
rect 9258 -4142 9402 -4126
rect 9450 -4092 9594 -4076
rect 9450 -4126 9466 -4092
rect 9500 -4126 9594 -4092
rect 9450 -4142 9594 -4126
rect 9642 -4092 9786 -4076
rect 9642 -4126 9658 -4092
rect 9692 -4126 9786 -4092
rect 9642 -4142 9786 -4126
rect 9997 -4091 10141 -4075
rect 9997 -4125 10013 -4091
rect 10047 -4125 10141 -4091
rect 9997 -4141 10141 -4125
rect 10189 -4091 10333 -4008
rect 10405 -4050 10459 -3788
rect 10525 -3915 10555 -3765
rect 12219 -3008 12249 -2872
rect 12315 -2801 12345 -2775
rect 12411 -2801 12441 -2775
rect 12507 -2801 12537 -2775
rect 12603 -2801 12633 -2775
rect 12699 -2801 12729 -2775
rect 12315 -2872 12729 -2801
rect 12315 -2914 12345 -2872
rect 12826 -2909 12842 -2683
rect 12876 -2685 12892 -2683
rect 12876 -2715 12923 -2685
rect 13137 -2715 13163 -2685
rect 12876 -2781 12892 -2715
rect 12876 -2811 12923 -2781
rect 13137 -2811 13163 -2781
rect 12876 -2877 12892 -2811
rect 12876 -2907 12923 -2877
rect 13137 -2907 13163 -2877
rect 12876 -2909 12892 -2907
rect 12297 -2930 12363 -2914
rect 12826 -2925 12892 -2909
rect 12297 -2964 12313 -2930
rect 12347 -2964 12363 -2930
rect 12297 -2980 12363 -2964
rect 12315 -3008 12345 -2980
rect 12826 -3129 12893 -3113
rect 12826 -3163 12842 -3129
rect 12876 -3131 12893 -3129
rect 12876 -3161 12923 -3131
rect 13123 -3161 13149 -3131
rect 12876 -3163 12893 -3161
rect 12826 -3179 12893 -3163
rect 12219 -3234 12249 -3208
rect 12315 -3234 12345 -3208
rect 11164 -3799 11194 -3766
rect 10980 -3829 11194 -3799
rect 10525 -3945 10663 -3915
rect 10399 -4075 10459 -4050
rect 10573 -4075 10663 -3945
rect 10189 -4125 10205 -4091
rect 10239 -4125 10333 -4091
rect 10189 -4141 10333 -4125
rect 10381 -4091 10525 -4075
rect 10381 -4125 10397 -4091
rect 10431 -4125 10525 -4091
rect 10381 -4141 10525 -4125
rect 10573 -4091 10717 -4075
rect 10980 -4076 11010 -3829
rect 11260 -3871 11290 -3766
rect 11356 -3789 11386 -3766
rect 11116 -4009 11290 -3871
rect 10573 -4125 10589 -4091
rect 10623 -4125 10717 -4091
rect 10573 -4141 10717 -4125
rect 7200 -4173 7230 -4142
rect 7296 -4173 7326 -4142
rect 7392 -4173 7422 -4142
rect 7488 -4173 7518 -4142
rect 7584 -4173 7614 -4142
rect 7680 -4173 7710 -4142
rect 7776 -4173 7806 -4142
rect 7872 -4173 7902 -4142
rect 8148 -4173 8178 -4142
rect 8244 -4173 8274 -4142
rect 8340 -4173 8370 -4142
rect 8436 -4173 8466 -4142
rect 8532 -4173 8562 -4142
rect 8628 -4173 8658 -4142
rect 8724 -4173 8754 -4142
rect 8820 -4173 8850 -4142
rect 9084 -4173 9114 -4142
rect 9180 -4173 9210 -4142
rect 9276 -4173 9306 -4142
rect 9372 -4173 9402 -4142
rect 9468 -4173 9498 -4142
rect 9564 -4173 9594 -4142
rect 9660 -4173 9690 -4142
rect 9756 -4173 9786 -4142
rect 10015 -4172 10045 -4141
rect 10111 -4172 10141 -4141
rect 10207 -4172 10237 -4141
rect 10303 -4172 10333 -4141
rect 10399 -4172 10429 -4141
rect 10495 -4172 10525 -4141
rect 10591 -4172 10621 -4141
rect 10687 -4172 10717 -4141
rect 10924 -4092 11068 -4076
rect 10924 -4126 10940 -4092
rect 10974 -4126 11068 -4092
rect 10924 -4142 11068 -4126
rect 11116 -4092 11260 -4009
rect 11332 -4051 11386 -3789
rect 11452 -3916 11482 -3766
rect 11452 -3946 11590 -3916
rect 11326 -4076 11386 -4051
rect 11500 -4076 11590 -3946
rect 11116 -4126 11132 -4092
rect 11166 -4126 11260 -4092
rect 11116 -4142 11260 -4126
rect 11308 -4092 11452 -4076
rect 11308 -4126 11324 -4092
rect 11358 -4126 11452 -4092
rect 11308 -4142 11452 -4126
rect 11500 -4092 11644 -4076
rect 11500 -4126 11516 -4092
rect 11550 -4126 11644 -4092
rect 11500 -4142 11644 -4126
rect 10942 -4173 10972 -4142
rect 11038 -4173 11068 -4142
rect 11134 -4173 11164 -4142
rect 11230 -4173 11260 -4142
rect 11326 -4173 11356 -4142
rect 11422 -4173 11452 -4142
rect 11518 -4173 11548 -4142
rect 11614 -4173 11644 -4142
rect 7200 -4521 7230 -4495
rect 7296 -4521 7326 -4495
rect 7392 -4521 7422 -4495
rect 7488 -4521 7518 -4495
rect 7584 -4521 7614 -4495
rect 7680 -4521 7710 -4495
rect 7776 -4521 7806 -4495
rect 7872 -4521 7902 -4495
rect 8148 -4521 8178 -4495
rect 8244 -4521 8274 -4495
rect 8340 -4521 8370 -4495
rect 8436 -4521 8466 -4495
rect 8532 -4521 8562 -4495
rect 8628 -4521 8658 -4495
rect 8724 -4521 8754 -4495
rect 8820 -4521 8850 -4495
rect 9084 -4521 9114 -4495
rect 9180 -4521 9210 -4495
rect 9276 -4521 9306 -4495
rect 9372 -4521 9402 -4495
rect 9468 -4521 9498 -4495
rect 9564 -4521 9594 -4495
rect 9660 -4521 9690 -4495
rect 9756 -4521 9786 -4495
rect 10015 -4520 10045 -4494
rect 10111 -4520 10141 -4494
rect 10207 -4520 10237 -4494
rect 10303 -4520 10333 -4494
rect 10399 -4520 10429 -4494
rect 10495 -4520 10525 -4494
rect 10591 -4520 10621 -4494
rect 10687 -4520 10717 -4494
rect 10942 -4521 10972 -4495
rect 11038 -4521 11068 -4495
rect 11134 -4521 11164 -4495
rect 11230 -4521 11260 -4495
rect 11326 -4521 11356 -4495
rect 11422 -4521 11452 -4495
rect 11518 -4521 11548 -4495
rect 11614 -4521 11644 -4495
rect -20679 -4565 -20649 -4534
rect -20587 -4565 -20557 -4534
rect -20491 -4565 -20461 -4534
rect -20395 -4565 -20365 -4534
rect -20299 -4564 -20269 -4534
rect -20203 -4564 -20173 -4534
rect -20107 -4564 -20077 -4534
rect -22514 -4610 -22448 -4594
rect -22514 -4645 -22498 -4610
rect -22464 -4631 -22448 -4610
rect -21943 -4625 -21876 -4609
rect -22464 -4645 -22426 -4631
rect -22514 -4661 -22426 -4645
rect -22026 -4661 -22000 -4631
rect -21943 -4659 -21927 -4625
rect -21893 -4627 -21876 -4625
rect -20873 -4622 -20363 -4565
rect -21893 -4657 -21846 -4627
rect -21646 -4657 -21620 -4627
rect -21893 -4659 -21876 -4657
rect -21943 -4675 -21876 -4659
rect -24335 -4743 -24162 -4727
rect -24335 -4778 -24234 -4743
rect -24200 -4757 -24162 -4743
rect -23762 -4757 -23736 -4727
rect -22599 -4743 -22426 -4727
rect -24200 -4778 -24184 -4757
rect -24335 -4794 -24184 -4778
rect -22599 -4778 -22498 -4743
rect -22464 -4757 -22426 -4743
rect -22026 -4757 -22000 -4727
rect -20873 -4732 -20854 -4622
rect -20807 -4715 -20363 -4622
rect -20299 -4593 -20077 -4564
rect -20299 -4638 -20269 -4593
rect -20139 -4638 -20077 -4593
rect -20299 -4657 -20077 -4638
rect -20011 -4565 -19981 -4534
rect -19915 -4565 -19885 -4534
rect -19819 -4565 -19789 -4534
rect -20011 -4598 -19789 -4565
rect -20011 -4643 -19938 -4598
rect -19808 -4643 -19789 -4598
rect -20011 -4658 -19789 -4643
rect -19723 -4565 -19693 -4534
rect -19627 -4565 -19597 -4534
rect -19531 -4565 -19501 -4534
rect -19439 -4565 -19409 -4534
rect -19120 -4565 -19090 -4534
rect -19028 -4565 -18998 -4534
rect -18932 -4565 -18902 -4534
rect -18836 -4565 -18806 -4534
rect -18740 -4564 -18710 -4534
rect -18644 -4564 -18614 -4534
rect -18548 -4564 -18518 -4534
rect -20807 -4732 -19789 -4715
rect -22464 -4778 -22448 -4757
rect -22599 -4794 -22448 -4778
rect -20873 -4824 -19789 -4732
rect -20712 -4999 -20636 -4824
rect -20587 -4914 -20365 -4889
rect -20587 -4959 -20544 -4914
rect -20414 -4959 -20365 -4914
rect -20679 -5024 -20649 -4999
rect -20587 -5002 -20365 -4959
rect -20587 -5024 -20557 -5002
rect -20491 -5024 -20461 -5002
rect -20395 -5024 -20365 -5002
rect -20299 -4922 -20077 -4894
rect -20299 -4967 -20261 -4922
rect -20131 -4967 -20077 -4922
rect -20299 -5002 -20077 -4967
rect -20299 -5024 -20269 -5002
rect -20203 -5024 -20173 -5002
rect -20107 -5024 -20077 -5002
rect -20011 -5002 -19789 -4824
rect -20011 -5024 -19981 -5002
rect -19915 -5024 -19885 -5002
rect -19819 -5024 -19789 -5002
rect -19723 -4722 -19409 -4565
rect -19153 -4652 -18804 -4565
rect -19723 -4777 -19691 -4722
rect -19626 -4777 -19409 -4722
rect -19723 -5002 -19409 -4777
rect -19342 -4667 -18804 -4652
rect -18740 -4593 -18518 -4564
rect -18740 -4638 -18710 -4593
rect -18580 -4638 -18518 -4593
rect -18740 -4657 -18518 -4638
rect -18452 -4565 -18422 -4534
rect -18356 -4565 -18326 -4534
rect -18260 -4565 -18230 -4534
rect -18452 -4598 -18230 -4565
rect -18452 -4643 -18379 -4598
rect -18249 -4643 -18230 -4598
rect -18452 -4658 -18230 -4643
rect -18164 -4565 -18134 -4534
rect -18068 -4565 -18038 -4534
rect -17972 -4565 -17942 -4534
rect -17880 -4565 -17850 -4534
rect -17388 -4565 -17358 -4534
rect -17296 -4565 -17266 -4534
rect -17200 -4565 -17170 -4534
rect -17104 -4565 -17074 -4534
rect -17008 -4564 -16978 -4534
rect -16912 -4564 -16882 -4534
rect -16816 -4564 -16786 -4534
rect -19342 -4807 -19297 -4667
rect -19224 -4715 -18804 -4667
rect -19224 -4807 -18230 -4715
rect -19342 -4824 -18230 -4807
rect -19153 -4999 -19077 -4824
rect -19028 -4914 -18806 -4889
rect -19028 -4959 -18985 -4914
rect -18855 -4959 -18806 -4914
rect -19723 -5024 -19693 -5002
rect -19627 -5024 -19597 -5002
rect -19531 -5024 -19501 -5002
rect -19439 -5024 -19409 -5002
rect -19120 -5024 -19090 -4999
rect -19028 -5002 -18806 -4959
rect -19028 -5024 -18998 -5002
rect -18932 -5024 -18902 -5002
rect -18836 -5024 -18806 -5002
rect -18740 -4922 -18518 -4894
rect -18740 -4967 -18702 -4922
rect -18572 -4967 -18518 -4922
rect -18740 -5002 -18518 -4967
rect -18740 -5024 -18710 -5002
rect -18644 -5024 -18614 -5002
rect -18548 -5024 -18518 -5002
rect -18452 -5002 -18230 -4824
rect -18452 -5024 -18422 -5002
rect -18356 -5024 -18326 -5002
rect -18260 -5024 -18230 -5002
rect -18164 -4722 -17850 -4565
rect -18164 -4777 -18132 -4722
rect -18067 -4777 -17850 -4722
rect -18164 -5002 -17850 -4777
rect -17582 -4622 -17072 -4565
rect -17582 -4732 -17563 -4622
rect -17516 -4715 -17072 -4622
rect -17008 -4593 -16786 -4564
rect -17008 -4638 -16978 -4593
rect -16848 -4638 -16786 -4593
rect -17008 -4657 -16786 -4638
rect -16720 -4565 -16690 -4534
rect -16624 -4565 -16594 -4534
rect -16528 -4565 -16498 -4534
rect -16720 -4598 -16498 -4565
rect -16720 -4643 -16647 -4598
rect -16517 -4643 -16498 -4598
rect -16720 -4658 -16498 -4643
rect -16432 -4565 -16402 -4534
rect -16336 -4565 -16306 -4534
rect -16240 -4565 -16210 -4534
rect -16148 -4565 -16118 -4534
rect -15829 -4565 -15799 -4534
rect -15737 -4565 -15707 -4534
rect -15641 -4565 -15611 -4534
rect -15545 -4565 -15515 -4534
rect -15449 -4564 -15419 -4534
rect -15353 -4564 -15323 -4534
rect -15257 -4564 -15227 -4534
rect -17516 -4732 -16498 -4715
rect -17582 -4824 -16498 -4732
rect -17421 -4999 -17345 -4824
rect -17296 -4914 -17074 -4889
rect -17296 -4959 -17253 -4914
rect -17123 -4959 -17074 -4914
rect -18164 -5024 -18134 -5002
rect -18068 -5024 -18038 -5002
rect -17972 -5024 -17942 -5002
rect -17880 -5024 -17850 -5002
rect -17388 -5024 -17358 -4999
rect -17296 -5002 -17074 -4959
rect -17296 -5024 -17266 -5002
rect -17200 -5024 -17170 -5002
rect -17104 -5024 -17074 -5002
rect -17008 -4922 -16786 -4894
rect -17008 -4967 -16970 -4922
rect -16840 -4967 -16786 -4922
rect -17008 -5002 -16786 -4967
rect -17008 -5024 -16978 -5002
rect -16912 -5024 -16882 -5002
rect -16816 -5024 -16786 -5002
rect -16720 -5002 -16498 -4824
rect -16720 -5024 -16690 -5002
rect -16624 -5024 -16594 -5002
rect -16528 -5024 -16498 -5002
rect -16432 -4722 -16118 -4565
rect -15862 -4652 -15513 -4565
rect -16432 -4777 -16400 -4722
rect -16335 -4777 -16118 -4722
rect -16432 -5002 -16118 -4777
rect -16051 -4667 -15513 -4652
rect -15449 -4593 -15227 -4564
rect -15449 -4638 -15419 -4593
rect -15289 -4638 -15227 -4593
rect -15449 -4657 -15227 -4638
rect -15161 -4565 -15131 -4534
rect -15065 -4565 -15035 -4534
rect -14969 -4565 -14939 -4534
rect -15161 -4598 -14939 -4565
rect -15161 -4643 -15088 -4598
rect -14958 -4643 -14939 -4598
rect -15161 -4658 -14939 -4643
rect -14873 -4565 -14843 -4534
rect -14777 -4565 -14747 -4534
rect -14681 -4565 -14651 -4534
rect -14589 -4565 -14559 -4534
rect -14097 -4565 -14067 -4534
rect -14005 -4565 -13975 -4534
rect -13909 -4565 -13879 -4534
rect -13813 -4565 -13783 -4534
rect -13717 -4564 -13687 -4534
rect -13621 -4564 -13591 -4534
rect -13525 -4564 -13495 -4534
rect -16051 -4807 -16006 -4667
rect -15933 -4715 -15513 -4667
rect -15933 -4807 -14939 -4715
rect -16051 -4824 -14939 -4807
rect -15862 -4999 -15786 -4824
rect -15737 -4914 -15515 -4889
rect -15737 -4959 -15694 -4914
rect -15564 -4959 -15515 -4914
rect -16432 -5024 -16402 -5002
rect -16336 -5024 -16306 -5002
rect -16240 -5024 -16210 -5002
rect -16148 -5024 -16118 -5002
rect -15829 -5024 -15799 -4999
rect -15737 -5002 -15515 -4959
rect -15737 -5024 -15707 -5002
rect -15641 -5024 -15611 -5002
rect -15545 -5024 -15515 -5002
rect -15449 -4922 -15227 -4894
rect -15449 -4967 -15411 -4922
rect -15281 -4967 -15227 -4922
rect -15449 -5002 -15227 -4967
rect -15449 -5024 -15419 -5002
rect -15353 -5024 -15323 -5002
rect -15257 -5024 -15227 -5002
rect -15161 -5002 -14939 -4824
rect -15161 -5024 -15131 -5002
rect -15065 -5024 -15035 -5002
rect -14969 -5024 -14939 -5002
rect -14873 -4722 -14559 -4565
rect -14873 -4777 -14841 -4722
rect -14776 -4777 -14559 -4722
rect -14873 -5002 -14559 -4777
rect -14291 -4622 -13781 -4565
rect -14291 -4732 -14272 -4622
rect -14225 -4715 -13781 -4622
rect -13717 -4593 -13495 -4564
rect -13717 -4638 -13687 -4593
rect -13557 -4638 -13495 -4593
rect -13717 -4657 -13495 -4638
rect -13429 -4565 -13399 -4534
rect -13333 -4565 -13303 -4534
rect -13237 -4565 -13207 -4534
rect -13429 -4598 -13207 -4565
rect -13429 -4643 -13356 -4598
rect -13226 -4643 -13207 -4598
rect -13429 -4658 -13207 -4643
rect -13141 -4565 -13111 -4534
rect -13045 -4565 -13015 -4534
rect -12949 -4565 -12919 -4534
rect -12857 -4565 -12827 -4534
rect -12538 -4565 -12508 -4534
rect -12446 -4565 -12416 -4534
rect -12350 -4565 -12320 -4534
rect -12254 -4565 -12224 -4534
rect -12158 -4564 -12128 -4534
rect -12062 -4564 -12032 -4534
rect -11966 -4564 -11936 -4534
rect -14225 -4732 -13207 -4715
rect -14291 -4824 -13207 -4732
rect -14130 -4999 -14054 -4824
rect -14005 -4914 -13783 -4889
rect -14005 -4959 -13962 -4914
rect -13832 -4959 -13783 -4914
rect -14873 -5024 -14843 -5002
rect -14777 -5024 -14747 -5002
rect -14681 -5024 -14651 -5002
rect -14589 -5024 -14559 -5002
rect -14097 -5024 -14067 -4999
rect -14005 -5002 -13783 -4959
rect -14005 -5024 -13975 -5002
rect -13909 -5024 -13879 -5002
rect -13813 -5024 -13783 -5002
rect -13717 -4922 -13495 -4894
rect -13717 -4967 -13679 -4922
rect -13549 -4967 -13495 -4922
rect -13717 -5002 -13495 -4967
rect -13717 -5024 -13687 -5002
rect -13621 -5024 -13591 -5002
rect -13525 -5024 -13495 -5002
rect -13429 -5002 -13207 -4824
rect -13429 -5024 -13399 -5002
rect -13333 -5024 -13303 -5002
rect -13237 -5024 -13207 -5002
rect -13141 -4722 -12827 -4565
rect -12571 -4652 -12222 -4565
rect -13141 -4777 -13109 -4722
rect -13044 -4777 -12827 -4722
rect -13141 -5002 -12827 -4777
rect -12760 -4667 -12222 -4652
rect -12158 -4593 -11936 -4564
rect -12158 -4638 -12128 -4593
rect -11998 -4638 -11936 -4593
rect -12158 -4657 -11936 -4638
rect -11870 -4565 -11840 -4534
rect -11774 -4565 -11744 -4534
rect -11678 -4565 -11648 -4534
rect -11870 -4598 -11648 -4565
rect -11870 -4643 -11797 -4598
rect -11667 -4643 -11648 -4598
rect -11870 -4658 -11648 -4643
rect -11582 -4565 -11552 -4534
rect -11486 -4565 -11456 -4534
rect -11390 -4565 -11360 -4534
rect -11298 -4565 -11268 -4534
rect -10806 -4565 -10776 -4534
rect -10714 -4565 -10684 -4534
rect -10618 -4565 -10588 -4534
rect -10522 -4565 -10492 -4534
rect -10426 -4564 -10396 -4534
rect -10330 -4564 -10300 -4534
rect -10234 -4564 -10204 -4534
rect -12760 -4807 -12715 -4667
rect -12642 -4715 -12222 -4667
rect -12642 -4807 -11648 -4715
rect -12760 -4824 -11648 -4807
rect -12571 -4999 -12495 -4824
rect -12446 -4914 -12224 -4889
rect -12446 -4959 -12403 -4914
rect -12273 -4959 -12224 -4914
rect -13141 -5024 -13111 -5002
rect -13045 -5024 -13015 -5002
rect -12949 -5024 -12919 -5002
rect -12857 -5024 -12827 -5002
rect -12538 -5024 -12508 -4999
rect -12446 -5002 -12224 -4959
rect -12446 -5024 -12416 -5002
rect -12350 -5024 -12320 -5002
rect -12254 -5024 -12224 -5002
rect -12158 -4922 -11936 -4894
rect -12158 -4967 -12120 -4922
rect -11990 -4967 -11936 -4922
rect -12158 -5002 -11936 -4967
rect -12158 -5024 -12128 -5002
rect -12062 -5024 -12032 -5002
rect -11966 -5024 -11936 -5002
rect -11870 -5002 -11648 -4824
rect -11870 -5024 -11840 -5002
rect -11774 -5024 -11744 -5002
rect -11678 -5024 -11648 -5002
rect -11582 -4722 -11268 -4565
rect -11582 -4777 -11550 -4722
rect -11485 -4777 -11268 -4722
rect -11582 -5002 -11268 -4777
rect -11000 -4622 -10490 -4565
rect -11000 -4732 -10981 -4622
rect -10934 -4715 -10490 -4622
rect -10426 -4593 -10204 -4564
rect -10426 -4638 -10396 -4593
rect -10266 -4638 -10204 -4593
rect -10426 -4657 -10204 -4638
rect -10138 -4565 -10108 -4534
rect -10042 -4565 -10012 -4534
rect -9946 -4565 -9916 -4534
rect -10138 -4598 -9916 -4565
rect -10138 -4643 -10065 -4598
rect -9935 -4643 -9916 -4598
rect -10138 -4658 -9916 -4643
rect -9850 -4565 -9820 -4534
rect -9754 -4565 -9724 -4534
rect -9658 -4565 -9628 -4534
rect -9566 -4565 -9536 -4534
rect -9247 -4565 -9217 -4534
rect -9155 -4565 -9125 -4534
rect -9059 -4565 -9029 -4534
rect -8963 -4565 -8933 -4534
rect -8867 -4564 -8837 -4534
rect -8771 -4564 -8741 -4534
rect -8675 -4564 -8645 -4534
rect -10934 -4732 -9916 -4715
rect -11000 -4824 -9916 -4732
rect -10839 -4999 -10763 -4824
rect -10714 -4914 -10492 -4889
rect -10714 -4959 -10671 -4914
rect -10541 -4959 -10492 -4914
rect -11582 -5024 -11552 -5002
rect -11486 -5024 -11456 -5002
rect -11390 -5024 -11360 -5002
rect -11298 -5024 -11268 -5002
rect -10806 -5024 -10776 -4999
rect -10714 -5002 -10492 -4959
rect -10714 -5024 -10684 -5002
rect -10618 -5024 -10588 -5002
rect -10522 -5024 -10492 -5002
rect -10426 -4922 -10204 -4894
rect -10426 -4967 -10388 -4922
rect -10258 -4967 -10204 -4922
rect -10426 -5002 -10204 -4967
rect -10426 -5024 -10396 -5002
rect -10330 -5024 -10300 -5002
rect -10234 -5024 -10204 -5002
rect -10138 -5002 -9916 -4824
rect -10138 -5024 -10108 -5002
rect -10042 -5024 -10012 -5002
rect -9946 -5024 -9916 -5002
rect -9850 -4722 -9536 -4565
rect -9280 -4652 -8931 -4565
rect -9850 -4777 -9818 -4722
rect -9753 -4777 -9536 -4722
rect -9850 -5002 -9536 -4777
rect -9469 -4667 -8931 -4652
rect -8867 -4593 -8645 -4564
rect -8867 -4638 -8837 -4593
rect -8707 -4638 -8645 -4593
rect -8867 -4657 -8645 -4638
rect -8579 -4565 -8549 -4534
rect -8483 -4565 -8453 -4534
rect -8387 -4565 -8357 -4534
rect -8579 -4598 -8357 -4565
rect -8579 -4643 -8506 -4598
rect -8376 -4643 -8357 -4598
rect -8579 -4658 -8357 -4643
rect -8291 -4565 -8261 -4534
rect -8195 -4565 -8165 -4534
rect -8099 -4565 -8069 -4534
rect -8007 -4565 -7977 -4534
rect -9469 -4807 -9424 -4667
rect -9351 -4715 -8931 -4667
rect -9351 -4807 -8357 -4715
rect -9469 -4824 -8357 -4807
rect -9280 -4999 -9204 -4824
rect -9155 -4914 -8933 -4889
rect -9155 -4959 -9112 -4914
rect -8982 -4959 -8933 -4914
rect -9850 -5024 -9820 -5002
rect -9754 -5024 -9724 -5002
rect -9658 -5024 -9628 -5002
rect -9566 -5024 -9536 -5002
rect -9247 -5024 -9217 -4999
rect -9155 -5002 -8933 -4959
rect -9155 -5024 -9125 -5002
rect -9059 -5024 -9029 -5002
rect -8963 -5024 -8933 -5002
rect -8867 -4922 -8645 -4894
rect -8867 -4967 -8829 -4922
rect -8699 -4967 -8645 -4922
rect -8867 -5002 -8645 -4967
rect -8867 -5024 -8837 -5002
rect -8771 -5024 -8741 -5002
rect -8675 -5024 -8645 -5002
rect -8579 -5002 -8357 -4824
rect -8579 -5024 -8549 -5002
rect -8483 -5024 -8453 -5002
rect -8387 -5024 -8357 -5002
rect -8291 -4722 -7977 -4565
rect -8291 -4777 -8259 -4722
rect -8194 -4777 -7977 -4722
rect -8291 -5002 -7977 -4777
rect -8291 -5024 -8261 -5002
rect -8195 -5024 -8165 -5002
rect -8099 -5024 -8069 -5002
rect -8007 -5024 -7977 -5002
rect 5561 -5093 5627 -5077
rect -20679 -5180 -20649 -5154
rect -20587 -5180 -20557 -5154
rect -20491 -5180 -20461 -5154
rect -20395 -5180 -20365 -5154
rect -20299 -5180 -20269 -5154
rect -20203 -5180 -20173 -5154
rect -20107 -5180 -20077 -5154
rect -20011 -5180 -19981 -5154
rect -19915 -5180 -19885 -5154
rect -19819 -5180 -19789 -5154
rect -19723 -5180 -19693 -5154
rect -19627 -5180 -19597 -5154
rect -19531 -5180 -19501 -5154
rect -19439 -5180 -19409 -5154
rect -19120 -5180 -19090 -5154
rect -19028 -5180 -18998 -5154
rect -18932 -5180 -18902 -5154
rect -18836 -5180 -18806 -5154
rect -18740 -5180 -18710 -5154
rect -18644 -5180 -18614 -5154
rect -18548 -5180 -18518 -5154
rect -18452 -5180 -18422 -5154
rect -18356 -5180 -18326 -5154
rect -18260 -5180 -18230 -5154
rect -18164 -5180 -18134 -5154
rect -18068 -5180 -18038 -5154
rect -17972 -5180 -17942 -5154
rect -17880 -5180 -17850 -5154
rect -17388 -5180 -17358 -5154
rect -17296 -5180 -17266 -5154
rect -17200 -5180 -17170 -5154
rect -17104 -5180 -17074 -5154
rect -17008 -5180 -16978 -5154
rect -16912 -5180 -16882 -5154
rect -16816 -5180 -16786 -5154
rect -16720 -5180 -16690 -5154
rect -16624 -5180 -16594 -5154
rect -16528 -5180 -16498 -5154
rect -16432 -5180 -16402 -5154
rect -16336 -5180 -16306 -5154
rect -16240 -5180 -16210 -5154
rect -16148 -5180 -16118 -5154
rect -15829 -5180 -15799 -5154
rect -15737 -5180 -15707 -5154
rect -15641 -5180 -15611 -5154
rect -15545 -5180 -15515 -5154
rect -15449 -5180 -15419 -5154
rect -15353 -5180 -15323 -5154
rect -15257 -5180 -15227 -5154
rect -15161 -5180 -15131 -5154
rect -15065 -5180 -15035 -5154
rect -14969 -5180 -14939 -5154
rect -14873 -5180 -14843 -5154
rect -14777 -5180 -14747 -5154
rect -14681 -5180 -14651 -5154
rect -14589 -5180 -14559 -5154
rect -14097 -5180 -14067 -5154
rect -14005 -5180 -13975 -5154
rect -13909 -5180 -13879 -5154
rect -13813 -5180 -13783 -5154
rect -13717 -5180 -13687 -5154
rect -13621 -5180 -13591 -5154
rect -13525 -5180 -13495 -5154
rect -13429 -5180 -13399 -5154
rect -13333 -5180 -13303 -5154
rect -13237 -5180 -13207 -5154
rect -13141 -5180 -13111 -5154
rect -13045 -5180 -13015 -5154
rect -12949 -5180 -12919 -5154
rect -12857 -5180 -12827 -5154
rect -12538 -5180 -12508 -5154
rect -12446 -5180 -12416 -5154
rect -12350 -5180 -12320 -5154
rect -12254 -5180 -12224 -5154
rect -12158 -5180 -12128 -5154
rect -12062 -5180 -12032 -5154
rect -11966 -5180 -11936 -5154
rect -11870 -5180 -11840 -5154
rect -11774 -5180 -11744 -5154
rect -11678 -5180 -11648 -5154
rect -11582 -5180 -11552 -5154
rect -11486 -5180 -11456 -5154
rect -11390 -5180 -11360 -5154
rect -11298 -5180 -11268 -5154
rect -10806 -5180 -10776 -5154
rect -10714 -5180 -10684 -5154
rect -10618 -5180 -10588 -5154
rect -10522 -5180 -10492 -5154
rect -10426 -5180 -10396 -5154
rect -10330 -5180 -10300 -5154
rect -10234 -5180 -10204 -5154
rect -10138 -5180 -10108 -5154
rect -10042 -5180 -10012 -5154
rect -9946 -5180 -9916 -5154
rect -9850 -5180 -9820 -5154
rect -9754 -5180 -9724 -5154
rect -9658 -5180 -9628 -5154
rect -9566 -5180 -9536 -5154
rect -9247 -5180 -9217 -5154
rect -9155 -5180 -9125 -5154
rect -9059 -5180 -9029 -5154
rect -8963 -5180 -8933 -5154
rect -8867 -5180 -8837 -5154
rect -8771 -5180 -8741 -5154
rect -8675 -5180 -8645 -5154
rect -8579 -5180 -8549 -5154
rect -8483 -5180 -8453 -5154
rect -8387 -5180 -8357 -5154
rect -8291 -5180 -8261 -5154
rect -8195 -5180 -8165 -5154
rect -8099 -5180 -8069 -5154
rect -8007 -5180 -7977 -5154
rect 5561 -5319 5577 -5093
rect 5611 -5095 5627 -5093
rect 6001 -5093 6067 -5077
rect 5611 -5125 5658 -5095
rect 5872 -5125 5898 -5095
rect 5611 -5191 5627 -5125
rect 5611 -5221 5658 -5191
rect 5872 -5221 5898 -5191
rect 5611 -5287 5627 -5221
rect 5611 -5317 5658 -5287
rect 5872 -5317 5898 -5287
rect 5611 -5319 5627 -5317
rect 5561 -5335 5627 -5319
rect 6001 -5319 6017 -5093
rect 6051 -5095 6067 -5093
rect 6441 -5093 6507 -5077
rect 6051 -5125 6098 -5095
rect 6312 -5125 6338 -5095
rect 6051 -5191 6067 -5125
rect 6051 -5221 6098 -5191
rect 6312 -5221 6338 -5191
rect 6051 -5287 6067 -5221
rect 6051 -5317 6098 -5287
rect 6312 -5317 6338 -5287
rect 6051 -5319 6067 -5317
rect 6001 -5335 6067 -5319
rect 6441 -5319 6457 -5093
rect 6491 -5095 6507 -5093
rect 6491 -5125 6538 -5095
rect 6752 -5125 6778 -5095
rect 6491 -5191 6507 -5125
rect 6491 -5221 6538 -5191
rect 6752 -5221 6778 -5191
rect 6491 -5287 6507 -5221
rect 6491 -5317 6538 -5287
rect 6752 -5317 6778 -5287
rect 6491 -5319 6507 -5317
rect 6441 -5335 6507 -5319
rect -23683 -5471 -23617 -5455
rect -24334 -5517 -24304 -5486
rect -24238 -5517 -24208 -5486
rect -24142 -5517 -24112 -5486
rect -24046 -5517 -24016 -5486
rect -23950 -5517 -23920 -5486
rect -23854 -5517 -23824 -5486
rect -23683 -5697 -23667 -5471
rect -23633 -5473 -23617 -5471
rect -21949 -5471 -21883 -5455
rect -23633 -5503 -23586 -5473
rect -23372 -5503 -23346 -5473
rect -23633 -5569 -23617 -5503
rect -22598 -5517 -22568 -5486
rect -22502 -5517 -22472 -5486
rect -22406 -5517 -22376 -5486
rect -22310 -5517 -22280 -5486
rect -22214 -5517 -22184 -5486
rect -22118 -5517 -22088 -5486
rect -23633 -5599 -23586 -5569
rect -23372 -5599 -23346 -5569
rect -23633 -5665 -23617 -5599
rect -23633 -5695 -23586 -5665
rect -23372 -5695 -23346 -5665
rect -23633 -5697 -23617 -5695
rect -23683 -5713 -23617 -5697
rect -24334 -5757 -24304 -5731
rect -24238 -5757 -24208 -5731
rect -24142 -5757 -24112 -5731
rect -24335 -5778 -24112 -5757
rect -24335 -5813 -24318 -5778
rect -24284 -5787 -24112 -5778
rect -24046 -5757 -24016 -5731
rect -23950 -5757 -23920 -5731
rect -23854 -5757 -23824 -5731
rect -21949 -5697 -21933 -5471
rect -21899 -5473 -21883 -5471
rect -21899 -5503 -21852 -5473
rect -21638 -5503 -21612 -5473
rect -21899 -5569 -21883 -5503
rect 5561 -5539 5628 -5523
rect -21899 -5599 -21852 -5569
rect -21638 -5599 -21612 -5569
rect -21899 -5665 -21883 -5599
rect 5561 -5573 5577 -5539
rect 5611 -5541 5628 -5539
rect 6001 -5539 6068 -5523
rect 5611 -5571 5658 -5541
rect 5858 -5571 5884 -5541
rect 5611 -5573 5628 -5571
rect 5561 -5589 5628 -5573
rect 6001 -5573 6017 -5539
rect 6051 -5541 6068 -5539
rect 6441 -5539 6508 -5523
rect 6051 -5571 6098 -5541
rect 6298 -5571 6324 -5541
rect 6051 -5573 6068 -5571
rect 6001 -5589 6068 -5573
rect 6441 -5573 6457 -5539
rect 6491 -5541 6508 -5539
rect 6491 -5571 6538 -5541
rect 6738 -5571 6764 -5541
rect 6491 -5573 6508 -5571
rect 6441 -5589 6508 -5573
rect -21899 -5695 -21852 -5665
rect -21638 -5695 -21612 -5665
rect -20468 -5685 -20438 -5654
rect -20372 -5685 -20342 -5654
rect -20276 -5685 -20246 -5654
rect -20180 -5685 -20150 -5654
rect -20084 -5685 -20054 -5654
rect -19988 -5685 -19958 -5654
rect -19359 -5685 -19329 -5654
rect -19263 -5685 -19233 -5654
rect -19167 -5685 -19137 -5654
rect -19071 -5685 -19041 -5654
rect -18975 -5685 -18945 -5654
rect -18879 -5685 -18849 -5654
rect -18477 -5685 -18447 -5654
rect -18381 -5685 -18351 -5654
rect -18285 -5685 -18255 -5654
rect -18189 -5685 -18159 -5654
rect -18093 -5685 -18063 -5654
rect -17997 -5685 -17967 -5654
rect -17177 -5685 -17147 -5654
rect -17081 -5685 -17051 -5654
rect -16985 -5685 -16955 -5654
rect -16889 -5685 -16859 -5654
rect -16793 -5685 -16763 -5654
rect -16697 -5685 -16667 -5654
rect -16068 -5685 -16038 -5654
rect -15972 -5685 -15942 -5654
rect -15876 -5685 -15846 -5654
rect -15780 -5685 -15750 -5654
rect -15684 -5685 -15654 -5654
rect -15588 -5685 -15558 -5654
rect -15186 -5685 -15156 -5654
rect -15090 -5685 -15060 -5654
rect -14994 -5685 -14964 -5654
rect -14898 -5685 -14868 -5654
rect -14802 -5685 -14772 -5654
rect -14706 -5685 -14676 -5654
rect -13886 -5685 -13856 -5654
rect -13790 -5685 -13760 -5654
rect -13694 -5685 -13664 -5654
rect -13598 -5685 -13568 -5654
rect -13502 -5685 -13472 -5654
rect -13406 -5685 -13376 -5654
rect -12777 -5685 -12747 -5654
rect -12681 -5685 -12651 -5654
rect -12585 -5685 -12555 -5654
rect -12489 -5685 -12459 -5654
rect -12393 -5685 -12363 -5654
rect -12297 -5685 -12267 -5654
rect -11895 -5685 -11865 -5654
rect -11799 -5685 -11769 -5654
rect -11703 -5685 -11673 -5654
rect -11607 -5685 -11577 -5654
rect -11511 -5685 -11481 -5654
rect -11415 -5685 -11385 -5654
rect -10595 -5685 -10565 -5654
rect -10499 -5685 -10469 -5654
rect -10403 -5685 -10373 -5654
rect -10307 -5685 -10277 -5654
rect -10211 -5685 -10181 -5654
rect -10115 -5685 -10085 -5654
rect -9486 -5685 -9456 -5654
rect -9390 -5685 -9360 -5654
rect -9294 -5685 -9264 -5654
rect -9198 -5685 -9168 -5654
rect -9102 -5685 -9072 -5654
rect -9006 -5685 -8976 -5654
rect -8604 -5685 -8574 -5654
rect -8508 -5685 -8478 -5654
rect -8412 -5685 -8382 -5654
rect -8316 -5685 -8286 -5654
rect -8220 -5685 -8190 -5654
rect -8124 -5685 -8094 -5654
rect -21899 -5697 -21883 -5695
rect -21949 -5713 -21883 -5697
rect -22598 -5757 -22568 -5731
rect -22502 -5757 -22472 -5731
rect -22406 -5757 -22376 -5731
rect -24046 -5778 -23824 -5757
rect -24284 -5813 -24268 -5787
rect -24335 -5824 -24268 -5813
rect -24046 -5813 -24029 -5778
rect -23995 -5787 -23824 -5778
rect -22599 -5778 -22376 -5757
rect -23995 -5813 -23979 -5787
rect -24046 -5824 -23979 -5813
rect -22599 -5813 -22582 -5778
rect -22548 -5787 -22376 -5778
rect -22310 -5757 -22280 -5731
rect -22214 -5757 -22184 -5731
rect -22118 -5757 -22088 -5731
rect -22310 -5778 -22088 -5757
rect -22548 -5813 -22532 -5787
rect -22599 -5824 -22532 -5813
rect -22310 -5813 -22293 -5778
rect -22259 -5787 -22088 -5778
rect -22259 -5813 -22243 -5787
rect -22310 -5824 -22243 -5813
rect -24335 -6019 -24292 -5824
rect -24250 -5902 -24184 -5886
rect -24250 -5937 -24234 -5902
rect -24200 -5923 -24184 -5902
rect -23683 -5917 -23616 -5901
rect -24200 -5937 -24162 -5923
rect -24250 -5953 -24162 -5937
rect -23762 -5953 -23736 -5923
rect -23683 -5951 -23667 -5917
rect -23633 -5919 -23616 -5917
rect -23633 -5949 -23586 -5919
rect -23386 -5949 -23360 -5919
rect -23633 -5951 -23616 -5949
rect -23683 -5967 -23616 -5951
rect -22599 -6019 -22556 -5824
rect -22514 -5902 -22448 -5886
rect -22514 -5937 -22498 -5902
rect -22464 -5923 -22448 -5902
rect -21949 -5917 -21882 -5901
rect -22464 -5937 -22426 -5923
rect -22514 -5953 -22426 -5937
rect -22026 -5953 -22000 -5923
rect -21949 -5951 -21933 -5917
rect -21899 -5919 -21882 -5917
rect 7200 -5737 7230 -5711
rect 7296 -5737 7326 -5711
rect 7392 -5737 7422 -5711
rect 7488 -5737 7518 -5711
rect 7584 -5737 7614 -5711
rect 7680 -5737 7710 -5711
rect 7776 -5737 7806 -5711
rect 7872 -5737 7902 -5711
rect 8148 -5737 8178 -5711
rect 8244 -5737 8274 -5711
rect 8340 -5737 8370 -5711
rect 8436 -5737 8466 -5711
rect 8532 -5737 8562 -5711
rect 8628 -5737 8658 -5711
rect 8724 -5737 8754 -5711
rect 8820 -5737 8850 -5711
rect 9084 -5737 9114 -5711
rect 9180 -5737 9210 -5711
rect 9276 -5737 9306 -5711
rect 9372 -5737 9402 -5711
rect 9468 -5737 9498 -5711
rect 9564 -5737 9594 -5711
rect 9660 -5737 9690 -5711
rect 9756 -5737 9786 -5711
rect 10015 -5737 10045 -5711
rect 10111 -5737 10141 -5711
rect 10207 -5737 10237 -5711
rect 10303 -5737 10333 -5711
rect 10399 -5737 10429 -5711
rect 10495 -5737 10525 -5711
rect 10591 -5737 10621 -5711
rect 10687 -5737 10717 -5711
rect 10942 -5737 10972 -5711
rect 11038 -5737 11068 -5711
rect 11134 -5737 11164 -5711
rect 11230 -5737 11260 -5711
rect 11326 -5737 11356 -5711
rect 11422 -5737 11452 -5711
rect 11518 -5737 11548 -5711
rect 11614 -5737 11644 -5711
rect -21899 -5949 -21852 -5919
rect -21652 -5949 -21626 -5919
rect -20468 -5925 -20438 -5899
rect -20372 -5925 -20342 -5899
rect -20276 -5925 -20246 -5899
rect -20469 -5946 -20246 -5925
rect -21899 -5951 -21882 -5949
rect -21949 -5967 -21882 -5951
rect -20469 -5981 -20452 -5946
rect -20418 -5955 -20246 -5946
rect -20180 -5925 -20150 -5899
rect -20084 -5925 -20054 -5899
rect -19988 -5925 -19958 -5899
rect -19359 -5925 -19329 -5899
rect -19263 -5925 -19233 -5899
rect -19167 -5925 -19137 -5899
rect -20180 -5946 -19958 -5925
rect -20418 -5981 -20402 -5955
rect -20469 -5992 -20402 -5981
rect -20180 -5981 -20163 -5946
rect -20129 -5955 -19958 -5946
rect -19360 -5946 -19137 -5925
rect -20129 -5981 -20113 -5955
rect -20180 -5992 -20113 -5981
rect -19360 -5981 -19343 -5946
rect -19309 -5955 -19137 -5946
rect -19071 -5925 -19041 -5899
rect -18975 -5925 -18945 -5899
rect -18879 -5925 -18849 -5899
rect -18477 -5925 -18447 -5899
rect -18381 -5925 -18351 -5899
rect -18285 -5925 -18255 -5899
rect -19071 -5946 -18849 -5925
rect -19309 -5981 -19293 -5955
rect -19360 -5992 -19293 -5981
rect -19071 -5981 -19054 -5946
rect -19020 -5955 -18849 -5946
rect -18478 -5946 -18255 -5925
rect -19020 -5981 -19004 -5955
rect -19071 -5992 -19004 -5981
rect -18478 -5981 -18461 -5946
rect -18427 -5955 -18255 -5946
rect -18189 -5925 -18159 -5899
rect -18093 -5925 -18063 -5899
rect -17997 -5925 -17967 -5899
rect -17177 -5925 -17147 -5899
rect -17081 -5925 -17051 -5899
rect -16985 -5925 -16955 -5899
rect -18189 -5946 -17967 -5925
rect -18427 -5981 -18411 -5955
rect -18478 -5992 -18411 -5981
rect -18189 -5981 -18172 -5946
rect -18138 -5955 -17967 -5946
rect -17178 -5946 -16955 -5925
rect -18138 -5981 -18122 -5955
rect -18189 -5992 -18122 -5981
rect -17178 -5981 -17161 -5946
rect -17127 -5955 -16955 -5946
rect -16889 -5925 -16859 -5899
rect -16793 -5925 -16763 -5899
rect -16697 -5925 -16667 -5899
rect -16068 -5925 -16038 -5899
rect -15972 -5925 -15942 -5899
rect -15876 -5925 -15846 -5899
rect -16889 -5946 -16667 -5925
rect -17127 -5981 -17111 -5955
rect -17178 -5992 -17111 -5981
rect -16889 -5981 -16872 -5946
rect -16838 -5955 -16667 -5946
rect -16069 -5946 -15846 -5925
rect -16838 -5981 -16822 -5955
rect -16889 -5992 -16822 -5981
rect -16069 -5981 -16052 -5946
rect -16018 -5955 -15846 -5946
rect -15780 -5925 -15750 -5899
rect -15684 -5925 -15654 -5899
rect -15588 -5925 -15558 -5899
rect -15186 -5925 -15156 -5899
rect -15090 -5925 -15060 -5899
rect -14994 -5925 -14964 -5899
rect -15780 -5946 -15558 -5925
rect -16018 -5981 -16002 -5955
rect -16069 -5992 -16002 -5981
rect -15780 -5981 -15763 -5946
rect -15729 -5955 -15558 -5946
rect -15187 -5946 -14964 -5925
rect -15729 -5981 -15713 -5955
rect -15780 -5992 -15713 -5981
rect -15187 -5981 -15170 -5946
rect -15136 -5955 -14964 -5946
rect -14898 -5925 -14868 -5899
rect -14802 -5925 -14772 -5899
rect -14706 -5925 -14676 -5899
rect -13886 -5925 -13856 -5899
rect -13790 -5925 -13760 -5899
rect -13694 -5925 -13664 -5899
rect -14898 -5946 -14676 -5925
rect -15136 -5981 -15120 -5955
rect -15187 -5992 -15120 -5981
rect -14898 -5981 -14881 -5946
rect -14847 -5955 -14676 -5946
rect -13887 -5946 -13664 -5925
rect -14847 -5981 -14831 -5955
rect -14898 -5992 -14831 -5981
rect -13887 -5981 -13870 -5946
rect -13836 -5955 -13664 -5946
rect -13598 -5925 -13568 -5899
rect -13502 -5925 -13472 -5899
rect -13406 -5925 -13376 -5899
rect -12777 -5925 -12747 -5899
rect -12681 -5925 -12651 -5899
rect -12585 -5925 -12555 -5899
rect -13598 -5946 -13376 -5925
rect -13836 -5981 -13820 -5955
rect -13887 -5992 -13820 -5981
rect -13598 -5981 -13581 -5946
rect -13547 -5955 -13376 -5946
rect -12778 -5946 -12555 -5925
rect -13547 -5981 -13531 -5955
rect -13598 -5992 -13531 -5981
rect -12778 -5981 -12761 -5946
rect -12727 -5955 -12555 -5946
rect -12489 -5925 -12459 -5899
rect -12393 -5925 -12363 -5899
rect -12297 -5925 -12267 -5899
rect -11895 -5925 -11865 -5899
rect -11799 -5925 -11769 -5899
rect -11703 -5925 -11673 -5899
rect -12489 -5946 -12267 -5925
rect -12727 -5981 -12711 -5955
rect -12778 -5992 -12711 -5981
rect -12489 -5981 -12472 -5946
rect -12438 -5955 -12267 -5946
rect -11896 -5946 -11673 -5925
rect -12438 -5981 -12422 -5955
rect -12489 -5992 -12422 -5981
rect -11896 -5981 -11879 -5946
rect -11845 -5955 -11673 -5946
rect -11607 -5925 -11577 -5899
rect -11511 -5925 -11481 -5899
rect -11415 -5925 -11385 -5899
rect -10595 -5925 -10565 -5899
rect -10499 -5925 -10469 -5899
rect -10403 -5925 -10373 -5899
rect -11607 -5946 -11385 -5925
rect -11845 -5981 -11829 -5955
rect -11896 -5992 -11829 -5981
rect -11607 -5981 -11590 -5946
rect -11556 -5955 -11385 -5946
rect -10596 -5946 -10373 -5925
rect -11556 -5981 -11540 -5955
rect -11607 -5992 -11540 -5981
rect -10596 -5981 -10579 -5946
rect -10545 -5955 -10373 -5946
rect -10307 -5925 -10277 -5899
rect -10211 -5925 -10181 -5899
rect -10115 -5925 -10085 -5899
rect -9486 -5925 -9456 -5899
rect -9390 -5925 -9360 -5899
rect -9294 -5925 -9264 -5899
rect -10307 -5946 -10085 -5925
rect -10545 -5981 -10529 -5955
rect -10596 -5992 -10529 -5981
rect -10307 -5981 -10290 -5946
rect -10256 -5955 -10085 -5946
rect -9487 -5946 -9264 -5925
rect -10256 -5981 -10240 -5955
rect -10307 -5992 -10240 -5981
rect -9487 -5981 -9470 -5946
rect -9436 -5955 -9264 -5946
rect -9198 -5925 -9168 -5899
rect -9102 -5925 -9072 -5899
rect -9006 -5925 -8976 -5899
rect -8604 -5925 -8574 -5899
rect -8508 -5925 -8478 -5899
rect -8412 -5925 -8382 -5899
rect -9198 -5946 -8976 -5925
rect -9436 -5981 -9420 -5955
rect -9487 -5992 -9420 -5981
rect -9198 -5981 -9181 -5946
rect -9147 -5955 -8976 -5946
rect -8605 -5946 -8382 -5925
rect -9147 -5981 -9131 -5955
rect -9198 -5992 -9131 -5981
rect -8605 -5981 -8588 -5946
rect -8554 -5955 -8382 -5946
rect -8316 -5925 -8286 -5899
rect -8220 -5925 -8190 -5899
rect -8124 -5925 -8094 -5899
rect -8316 -5946 -8094 -5925
rect -8554 -5981 -8538 -5955
rect -8605 -5992 -8538 -5981
rect -8316 -5981 -8299 -5946
rect -8265 -5955 -8094 -5946
rect -8265 -5981 -8249 -5955
rect -8316 -5992 -8249 -5981
rect -24335 -6035 -24162 -6019
rect -24335 -6070 -24234 -6035
rect -24200 -6049 -24162 -6035
rect -23762 -6049 -23736 -6019
rect -22599 -6035 -22426 -6019
rect -24200 -6070 -24184 -6049
rect -24335 -6086 -24184 -6070
rect -22599 -6070 -22498 -6035
rect -22464 -6049 -22426 -6035
rect -22026 -6049 -22000 -6019
rect -22464 -6070 -22448 -6049
rect -22599 -6086 -22448 -6070
rect -20469 -6187 -20426 -5992
rect -20384 -6070 -20318 -6054
rect -20384 -6105 -20368 -6070
rect -20334 -6091 -20318 -6070
rect -20334 -6105 -20296 -6091
rect -20384 -6121 -20296 -6105
rect -19896 -6121 -19870 -6091
rect -19360 -6187 -19317 -5992
rect -19275 -6070 -19209 -6054
rect -19275 -6105 -19259 -6070
rect -19225 -6091 -19209 -6070
rect -19225 -6105 -19187 -6091
rect -19275 -6121 -19187 -6105
rect -18787 -6121 -18761 -6091
rect -18478 -6187 -18435 -5992
rect -18393 -6070 -18327 -6054
rect -18393 -6105 -18377 -6070
rect -18343 -6091 -18327 -6070
rect -18343 -6105 -18305 -6091
rect -18393 -6121 -18305 -6105
rect -17905 -6121 -17879 -6091
rect -17178 -6187 -17135 -5992
rect -17093 -6070 -17027 -6054
rect -17093 -6105 -17077 -6070
rect -17043 -6091 -17027 -6070
rect -17043 -6105 -17005 -6091
rect -17093 -6121 -17005 -6105
rect -16605 -6121 -16579 -6091
rect -16069 -6187 -16026 -5992
rect -15984 -6070 -15918 -6054
rect -15984 -6105 -15968 -6070
rect -15934 -6091 -15918 -6070
rect -15934 -6105 -15896 -6091
rect -15984 -6121 -15896 -6105
rect -15496 -6121 -15470 -6091
rect -15187 -6187 -15144 -5992
rect -15102 -6070 -15036 -6054
rect -15102 -6105 -15086 -6070
rect -15052 -6091 -15036 -6070
rect -15052 -6105 -15014 -6091
rect -15102 -6121 -15014 -6105
rect -14614 -6121 -14588 -6091
rect -13887 -6187 -13844 -5992
rect -13802 -6070 -13736 -6054
rect -13802 -6105 -13786 -6070
rect -13752 -6091 -13736 -6070
rect -13752 -6105 -13714 -6091
rect -13802 -6121 -13714 -6105
rect -13314 -6121 -13288 -6091
rect -12778 -6187 -12735 -5992
rect -12693 -6070 -12627 -6054
rect -12693 -6105 -12677 -6070
rect -12643 -6091 -12627 -6070
rect -12643 -6105 -12605 -6091
rect -12693 -6121 -12605 -6105
rect -12205 -6121 -12179 -6091
rect -11896 -6187 -11853 -5992
rect -11811 -6070 -11745 -6054
rect -11811 -6105 -11795 -6070
rect -11761 -6091 -11745 -6070
rect -11761 -6105 -11723 -6091
rect -11811 -6121 -11723 -6105
rect -11323 -6121 -11297 -6091
rect -10596 -6187 -10553 -5992
rect -10511 -6070 -10445 -6054
rect -10511 -6105 -10495 -6070
rect -10461 -6091 -10445 -6070
rect -10461 -6105 -10423 -6091
rect -10511 -6121 -10423 -6105
rect -10023 -6121 -9997 -6091
rect -9487 -6187 -9444 -5992
rect -9402 -6070 -9336 -6054
rect -9402 -6105 -9386 -6070
rect -9352 -6091 -9336 -6070
rect -9352 -6105 -9314 -6091
rect -9402 -6121 -9314 -6105
rect -8914 -6121 -8888 -6091
rect -8605 -6187 -8562 -5992
rect -8520 -6070 -8454 -6054
rect -8520 -6105 -8504 -6070
rect -8470 -6091 -8454 -6070
rect 7200 -6090 7230 -6059
rect 7296 -6090 7326 -6059
rect 7392 -6090 7422 -6059
rect 7488 -6090 7518 -6059
rect 7584 -6090 7614 -6059
rect 7680 -6090 7710 -6059
rect 7776 -6090 7806 -6059
rect 7872 -6090 7902 -6059
rect 8148 -6090 8178 -6059
rect 8244 -6090 8274 -6059
rect 8340 -6090 8370 -6059
rect 8436 -6090 8466 -6059
rect 8532 -6090 8562 -6059
rect 8628 -6090 8658 -6059
rect 8724 -6090 8754 -6059
rect 8820 -6090 8850 -6059
rect 9084 -6090 9114 -6059
rect 9180 -6090 9210 -6059
rect 9276 -6090 9306 -6059
rect 9372 -6090 9402 -6059
rect 9468 -6090 9498 -6059
rect 9564 -6090 9594 -6059
rect 9660 -6090 9690 -6059
rect 9756 -6090 9786 -6059
rect 10015 -6090 10045 -6059
rect 10111 -6090 10141 -6059
rect 10207 -6090 10237 -6059
rect 10303 -6090 10333 -6059
rect 10399 -6090 10429 -6059
rect 10495 -6090 10525 -6059
rect 10591 -6090 10621 -6059
rect 10687 -6090 10717 -6059
rect 10942 -6090 10972 -6059
rect 11038 -6090 11068 -6059
rect 11134 -6090 11164 -6059
rect 11230 -6090 11260 -6059
rect 11326 -6090 11356 -6059
rect 11422 -6090 11452 -6059
rect 11518 -6090 11548 -6059
rect 11614 -6090 11644 -6059
rect -8470 -6105 -8432 -6091
rect -8520 -6121 -8432 -6105
rect -8032 -6121 -8006 -6091
rect 7182 -6106 7326 -6090
rect 7182 -6140 7198 -6106
rect 7232 -6140 7326 -6106
rect 7182 -6156 7326 -6140
rect 7374 -6106 7518 -6090
rect 7374 -6140 7390 -6106
rect 7424 -6140 7518 -6106
rect -20469 -6203 -20296 -6187
rect -20469 -6238 -20368 -6203
rect -20334 -6217 -20296 -6203
rect -19896 -6217 -19870 -6187
rect -19360 -6203 -19187 -6187
rect -20334 -6238 -20318 -6217
rect -20469 -6254 -20318 -6238
rect -19360 -6238 -19259 -6203
rect -19225 -6217 -19187 -6203
rect -18787 -6217 -18761 -6187
rect -18478 -6203 -18305 -6187
rect -19225 -6238 -19209 -6217
rect -19360 -6254 -19209 -6238
rect -18478 -6238 -18377 -6203
rect -18343 -6217 -18305 -6203
rect -17905 -6217 -17879 -6187
rect -17178 -6203 -17005 -6187
rect -18343 -6238 -18327 -6217
rect -18478 -6254 -18327 -6238
rect -17178 -6238 -17077 -6203
rect -17043 -6217 -17005 -6203
rect -16605 -6217 -16579 -6187
rect -16069 -6203 -15896 -6187
rect -17043 -6238 -17027 -6217
rect -17178 -6254 -17027 -6238
rect -16069 -6238 -15968 -6203
rect -15934 -6217 -15896 -6203
rect -15496 -6217 -15470 -6187
rect -15187 -6203 -15014 -6187
rect -15934 -6238 -15918 -6217
rect -16069 -6254 -15918 -6238
rect -15187 -6238 -15086 -6203
rect -15052 -6217 -15014 -6203
rect -14614 -6217 -14588 -6187
rect -13887 -6203 -13714 -6187
rect -15052 -6238 -15036 -6217
rect -15187 -6254 -15036 -6238
rect -13887 -6238 -13786 -6203
rect -13752 -6217 -13714 -6203
rect -13314 -6217 -13288 -6187
rect -12778 -6203 -12605 -6187
rect -13752 -6238 -13736 -6217
rect -13887 -6254 -13736 -6238
rect -12778 -6238 -12677 -6203
rect -12643 -6217 -12605 -6203
rect -12205 -6217 -12179 -6187
rect -11896 -6203 -11723 -6187
rect -12643 -6238 -12627 -6217
rect -12778 -6254 -12627 -6238
rect -11896 -6238 -11795 -6203
rect -11761 -6217 -11723 -6203
rect -11323 -6217 -11297 -6187
rect -10596 -6203 -10423 -6187
rect -11761 -6238 -11745 -6217
rect -11896 -6254 -11745 -6238
rect -10596 -6238 -10495 -6203
rect -10461 -6217 -10423 -6203
rect -10023 -6217 -9997 -6187
rect -9487 -6203 -9314 -6187
rect -10461 -6238 -10445 -6217
rect -10596 -6254 -10445 -6238
rect -9487 -6238 -9386 -6203
rect -9352 -6217 -9314 -6203
rect -8914 -6217 -8888 -6187
rect -8605 -6203 -8432 -6187
rect -9352 -6238 -9336 -6217
rect -9487 -6254 -9336 -6238
rect -8605 -6238 -8504 -6203
rect -8470 -6217 -8432 -6203
rect -8032 -6217 -8006 -6187
rect -8470 -6238 -8454 -6217
rect -8605 -6254 -8454 -6238
rect 7238 -6403 7268 -6156
rect 7374 -6223 7518 -6140
rect 7566 -6106 7710 -6090
rect 7566 -6140 7582 -6106
rect 7616 -6140 7710 -6106
rect 7566 -6156 7710 -6140
rect 7758 -6106 7902 -6090
rect 7758 -6140 7774 -6106
rect 7808 -6140 7902 -6106
rect 7758 -6156 7902 -6140
rect 8130 -6106 8274 -6090
rect 8130 -6140 8146 -6106
rect 8180 -6140 8274 -6106
rect 8130 -6156 8274 -6140
rect 8322 -6106 8466 -6090
rect 8322 -6140 8338 -6106
rect 8372 -6140 8466 -6106
rect 7584 -6181 7644 -6156
rect 7374 -6361 7548 -6223
rect 7238 -6433 7452 -6403
rect 7422 -6466 7452 -6433
rect 7518 -6466 7548 -6361
rect 7590 -6443 7644 -6181
rect 7758 -6286 7848 -6156
rect 7614 -6466 7644 -6443
rect 7710 -6316 7848 -6286
rect 7710 -6466 7740 -6316
rect 8186 -6403 8216 -6156
rect 8322 -6223 8466 -6140
rect 8514 -6106 8658 -6090
rect 8514 -6140 8530 -6106
rect 8564 -6140 8658 -6106
rect 8514 -6156 8658 -6140
rect 8706 -6106 8850 -6090
rect 8706 -6140 8722 -6106
rect 8756 -6140 8850 -6106
rect 8706 -6156 8850 -6140
rect 9066 -6106 9210 -6090
rect 9066 -6140 9082 -6106
rect 9116 -6140 9210 -6106
rect 9066 -6156 9210 -6140
rect 9258 -6106 9402 -6090
rect 9258 -6140 9274 -6106
rect 9308 -6140 9402 -6106
rect 8532 -6181 8592 -6156
rect 8322 -6361 8496 -6223
rect 8186 -6433 8400 -6403
rect 8370 -6466 8400 -6433
rect 8466 -6466 8496 -6361
rect 8538 -6443 8592 -6181
rect 8706 -6286 8796 -6156
rect 8562 -6466 8592 -6443
rect 8658 -6316 8796 -6286
rect 8658 -6466 8688 -6316
rect 9122 -6403 9152 -6156
rect 9258 -6223 9402 -6140
rect 9450 -6106 9594 -6090
rect 9450 -6140 9466 -6106
rect 9500 -6140 9594 -6106
rect 9450 -6156 9594 -6140
rect 9642 -6106 9786 -6090
rect 9642 -6140 9658 -6106
rect 9692 -6140 9786 -6106
rect 9642 -6156 9786 -6140
rect 9997 -6106 10141 -6090
rect 9997 -6140 10013 -6106
rect 10047 -6140 10141 -6106
rect 9997 -6156 10141 -6140
rect 10189 -6106 10333 -6090
rect 10189 -6140 10205 -6106
rect 10239 -6140 10333 -6106
rect 9468 -6181 9528 -6156
rect 9258 -6361 9432 -6223
rect 9122 -6433 9336 -6403
rect 9306 -6466 9336 -6433
rect 9402 -6466 9432 -6361
rect 9474 -6443 9528 -6181
rect 9642 -6286 9732 -6156
rect 9498 -6466 9528 -6443
rect 9594 -6316 9732 -6286
rect 9594 -6466 9624 -6316
rect 10053 -6403 10083 -6156
rect 10189 -6223 10333 -6140
rect 10381 -6106 10525 -6090
rect 10381 -6140 10397 -6106
rect 10431 -6140 10525 -6106
rect 10381 -6156 10525 -6140
rect 10573 -6106 10717 -6090
rect 10573 -6140 10589 -6106
rect 10623 -6140 10717 -6106
rect 10573 -6156 10717 -6140
rect 10924 -6106 11068 -6090
rect 10924 -6140 10940 -6106
rect 10974 -6140 11068 -6106
rect 10924 -6156 11068 -6140
rect 11116 -6106 11260 -6090
rect 11116 -6140 11132 -6106
rect 11166 -6140 11260 -6106
rect 10399 -6181 10459 -6156
rect 10189 -6361 10363 -6223
rect 10053 -6433 10267 -6403
rect 10237 -6466 10267 -6433
rect 10333 -6466 10363 -6361
rect 10405 -6443 10459 -6181
rect 10573 -6286 10663 -6156
rect 10429 -6466 10459 -6443
rect 10525 -6316 10663 -6286
rect 10525 -6466 10555 -6316
rect 10980 -6403 11010 -6156
rect 11116 -6223 11260 -6140
rect 11308 -6106 11452 -6090
rect 11308 -6140 11324 -6106
rect 11358 -6140 11452 -6106
rect 11308 -6156 11452 -6140
rect 11500 -6106 11644 -6090
rect 11500 -6140 11516 -6106
rect 11550 -6140 11644 -6106
rect 11500 -6156 11644 -6140
rect 11326 -6181 11386 -6156
rect 11116 -6361 11290 -6223
rect 10980 -6433 11194 -6403
rect 11164 -6466 11194 -6433
rect 11260 -6466 11290 -6361
rect 11332 -6443 11386 -6181
rect 11500 -6286 11590 -6156
rect 11356 -6466 11386 -6443
rect 11452 -6316 11590 -6286
rect 11452 -6466 11482 -6316
rect -20679 -7249 -20649 -7223
rect -20587 -7249 -20557 -7218
rect -20491 -7249 -20461 -7218
rect -20395 -7249 -20365 -7218
rect -20299 -7249 -20269 -7218
rect -20203 -7249 -20173 -7218
rect -20107 -7249 -20077 -7218
rect -20011 -7249 -19981 -7218
rect -19915 -7249 -19885 -7218
rect -19819 -7249 -19789 -7218
rect -19723 -7249 -19693 -7218
rect -19627 -7249 -19597 -7218
rect -19531 -7249 -19501 -7218
rect -19439 -7249 -19409 -7223
rect -19120 -7249 -19090 -7223
rect -19028 -7249 -18998 -7218
rect -18932 -7249 -18902 -7218
rect -18836 -7249 -18806 -7218
rect -18740 -7249 -18710 -7218
rect -18644 -7249 -18614 -7218
rect -18548 -7249 -18518 -7218
rect -18452 -7249 -18422 -7218
rect -18356 -7249 -18326 -7218
rect -18260 -7249 -18230 -7218
rect -18164 -7249 -18134 -7218
rect -18068 -7249 -18038 -7218
rect -17972 -7249 -17942 -7218
rect -17880 -7249 -17850 -7223
rect -17388 -7249 -17358 -7223
rect -17296 -7249 -17266 -7218
rect -17200 -7249 -17170 -7218
rect -17104 -7249 -17074 -7218
rect -17008 -7249 -16978 -7218
rect -16912 -7249 -16882 -7218
rect -16816 -7249 -16786 -7218
rect -16720 -7249 -16690 -7218
rect -16624 -7249 -16594 -7218
rect -16528 -7249 -16498 -7218
rect -16432 -7249 -16402 -7218
rect -16336 -7249 -16306 -7218
rect -16240 -7249 -16210 -7218
rect -16148 -7249 -16118 -7223
rect -15829 -7249 -15799 -7223
rect -15737 -7249 -15707 -7218
rect -15641 -7249 -15611 -7218
rect -15545 -7249 -15515 -7218
rect -15449 -7249 -15419 -7218
rect -15353 -7249 -15323 -7218
rect -15257 -7249 -15227 -7218
rect -15161 -7249 -15131 -7218
rect -15065 -7249 -15035 -7218
rect -14969 -7249 -14939 -7218
rect -14873 -7249 -14843 -7218
rect -14777 -7249 -14747 -7218
rect -14681 -7249 -14651 -7218
rect -14589 -7249 -14559 -7223
rect -14097 -7249 -14067 -7223
rect -14005 -7249 -13975 -7218
rect -13909 -7249 -13879 -7218
rect -13813 -7249 -13783 -7218
rect -13717 -7249 -13687 -7218
rect -13621 -7249 -13591 -7218
rect -13525 -7249 -13495 -7218
rect -13429 -7249 -13399 -7218
rect -13333 -7249 -13303 -7218
rect -13237 -7249 -13207 -7218
rect -13141 -7249 -13111 -7218
rect -13045 -7249 -13015 -7218
rect -12949 -7249 -12919 -7218
rect -12857 -7249 -12827 -7223
rect -12538 -7249 -12508 -7223
rect -12446 -7249 -12416 -7218
rect -12350 -7249 -12320 -7218
rect -12254 -7249 -12224 -7218
rect -12158 -7249 -12128 -7218
rect -12062 -7249 -12032 -7218
rect -11966 -7249 -11936 -7218
rect -11870 -7249 -11840 -7218
rect -11774 -7249 -11744 -7218
rect -11678 -7249 -11648 -7218
rect -11582 -7249 -11552 -7218
rect -11486 -7249 -11456 -7218
rect -11390 -7249 -11360 -7218
rect -11298 -7249 -11268 -7223
rect -10806 -7249 -10776 -7223
rect -10714 -7249 -10684 -7218
rect -10618 -7249 -10588 -7218
rect -10522 -7249 -10492 -7218
rect -10426 -7249 -10396 -7218
rect -10330 -7249 -10300 -7218
rect -10234 -7249 -10204 -7218
rect -10138 -7249 -10108 -7218
rect -10042 -7249 -10012 -7218
rect -9946 -7249 -9916 -7218
rect -9850 -7249 -9820 -7218
rect -9754 -7249 -9724 -7218
rect -9658 -7249 -9628 -7218
rect -9566 -7249 -9536 -7223
rect -9247 -7249 -9217 -7223
rect -9155 -7249 -9125 -7218
rect -9059 -7249 -9029 -7218
rect -8963 -7249 -8933 -7218
rect -8867 -7249 -8837 -7218
rect -8771 -7249 -8741 -7218
rect -8675 -7249 -8645 -7218
rect -8579 -7249 -8549 -7218
rect -8483 -7249 -8453 -7218
rect -8387 -7249 -8357 -7218
rect -8291 -7249 -8261 -7218
rect -8195 -7249 -8165 -7218
rect -8099 -7249 -8069 -7218
rect -8007 -7249 -7977 -7223
rect -23681 -7444 -23615 -7428
rect -24334 -7490 -24304 -7459
rect -24238 -7490 -24208 -7459
rect -24142 -7490 -24112 -7459
rect -24046 -7490 -24016 -7459
rect -23950 -7490 -23920 -7459
rect -23854 -7490 -23824 -7459
rect -23681 -7670 -23665 -7444
rect -23631 -7446 -23615 -7444
rect -21947 -7444 -21881 -7428
rect -23631 -7476 -23584 -7446
rect -23370 -7476 -23344 -7446
rect -23631 -7542 -23615 -7476
rect -22597 -7490 -22567 -7459
rect -22501 -7490 -22471 -7459
rect -22405 -7490 -22375 -7459
rect -22309 -7490 -22279 -7459
rect -22213 -7490 -22183 -7459
rect -22117 -7490 -22087 -7459
rect -23631 -7572 -23584 -7542
rect -23370 -7572 -23344 -7542
rect -23631 -7638 -23615 -7572
rect -23631 -7668 -23584 -7638
rect -23370 -7668 -23344 -7638
rect -23631 -7670 -23615 -7668
rect -23681 -7686 -23615 -7670
rect -24334 -7730 -24304 -7704
rect -24238 -7730 -24208 -7704
rect -24142 -7730 -24112 -7704
rect -24335 -7751 -24112 -7730
rect -24335 -7786 -24318 -7751
rect -24284 -7760 -24112 -7751
rect -24046 -7730 -24016 -7704
rect -23950 -7730 -23920 -7704
rect -23854 -7730 -23824 -7704
rect -21947 -7670 -21931 -7444
rect -21897 -7446 -21881 -7444
rect -21897 -7476 -21850 -7446
rect -21636 -7476 -21610 -7446
rect -21897 -7542 -21881 -7476
rect -21897 -7572 -21850 -7542
rect -21636 -7572 -21610 -7542
rect -21897 -7638 -21881 -7572
rect -21897 -7668 -21850 -7638
rect -21636 -7668 -21610 -7638
rect -21897 -7670 -21881 -7668
rect -21947 -7686 -21881 -7670
rect -22597 -7730 -22567 -7704
rect -22501 -7730 -22471 -7704
rect -22405 -7730 -22375 -7704
rect -24046 -7751 -23824 -7730
rect -24284 -7786 -24268 -7760
rect -24335 -7797 -24268 -7786
rect -24046 -7786 -24029 -7751
rect -23995 -7760 -23824 -7751
rect -22598 -7751 -22375 -7730
rect -23995 -7786 -23979 -7760
rect -24046 -7797 -23979 -7786
rect -22598 -7786 -22581 -7751
rect -22547 -7760 -22375 -7751
rect -22309 -7730 -22279 -7704
rect -22213 -7730 -22183 -7704
rect -22117 -7730 -22087 -7704
rect -22309 -7751 -22087 -7730
rect -22547 -7786 -22531 -7760
rect -22598 -7797 -22531 -7786
rect -22309 -7786 -22292 -7751
rect -22258 -7760 -22087 -7751
rect -22258 -7786 -22242 -7760
rect -22309 -7797 -22242 -7786
rect -24335 -7992 -24292 -7797
rect -24250 -7875 -24184 -7859
rect -24250 -7910 -24234 -7875
rect -24200 -7896 -24184 -7875
rect -23681 -7890 -23614 -7874
rect -24200 -7910 -24162 -7896
rect -24250 -7926 -24162 -7910
rect -23762 -7926 -23736 -7896
rect -23681 -7924 -23665 -7890
rect -23631 -7892 -23614 -7890
rect -23631 -7922 -23584 -7892
rect -23384 -7922 -23358 -7892
rect -23631 -7924 -23614 -7922
rect -23681 -7940 -23614 -7924
rect -22598 -7992 -22555 -7797
rect 11835 -6947 11865 -6921
rect 11931 -6947 11961 -6921
rect 12027 -6947 12057 -6921
rect 12123 -6947 12153 -6921
rect 12219 -6947 12249 -6921
rect 12315 -6947 12345 -6921
rect 12411 -6947 12441 -6921
rect 12507 -6947 12537 -6921
rect 12603 -6947 12633 -6921
rect 12699 -6947 12729 -6921
rect 12826 -7111 12892 -7095
rect 11835 -7229 11865 -7203
rect 11931 -7229 11961 -7203
rect 12027 -7229 12057 -7203
rect 12123 -7229 12153 -7203
rect 12219 -7229 12249 -7203
rect 11835 -7253 12249 -7229
rect 7422 -7292 7452 -7266
rect 7518 -7292 7548 -7266
rect 7614 -7292 7644 -7266
rect 7710 -7292 7740 -7266
rect 8370 -7292 8400 -7266
rect 8466 -7292 8496 -7266
rect 8562 -7292 8592 -7266
rect 8658 -7292 8688 -7266
rect 9306 -7292 9336 -7266
rect 9402 -7292 9432 -7266
rect 9498 -7292 9528 -7266
rect 9594 -7292 9624 -7266
rect 10237 -7292 10267 -7266
rect 10333 -7292 10363 -7266
rect 10429 -7292 10459 -7266
rect 10525 -7292 10555 -7266
rect 11164 -7292 11194 -7266
rect 11260 -7292 11290 -7266
rect 11356 -7292 11386 -7266
rect 11452 -7292 11482 -7266
rect 11835 -7287 12170 -7253
rect 12204 -7287 12249 -7253
rect 11835 -7300 12249 -7287
rect 7422 -7394 7452 -7368
rect 7518 -7394 7548 -7368
rect 7614 -7394 7644 -7368
rect 7710 -7394 7740 -7368
rect 8370 -7394 8400 -7368
rect 8466 -7394 8496 -7368
rect 8562 -7394 8592 -7368
rect 8658 -7394 8688 -7368
rect 9306 -7394 9336 -7368
rect 9402 -7394 9432 -7368
rect 9498 -7394 9528 -7368
rect 9594 -7394 9624 -7368
rect 10237 -7393 10267 -7367
rect 10333 -7393 10363 -7367
rect 10429 -7393 10459 -7367
rect 10525 -7393 10555 -7367
rect -20679 -7830 -20649 -7799
rect -20587 -7830 -20557 -7799
rect -20491 -7830 -20461 -7799
rect -20395 -7830 -20365 -7799
rect -20299 -7829 -20269 -7799
rect -20203 -7829 -20173 -7799
rect -20107 -7829 -20077 -7799
rect -22513 -7875 -22447 -7859
rect -22513 -7910 -22497 -7875
rect -22463 -7896 -22447 -7875
rect -21947 -7890 -21880 -7874
rect -22463 -7910 -22425 -7896
rect -22513 -7926 -22425 -7910
rect -22025 -7926 -21999 -7896
rect -21947 -7924 -21931 -7890
rect -21897 -7892 -21880 -7890
rect -20873 -7887 -20363 -7830
rect -21897 -7922 -21850 -7892
rect -21650 -7922 -21624 -7892
rect -21897 -7924 -21880 -7922
rect -21947 -7940 -21880 -7924
rect -24335 -8008 -24162 -7992
rect -24335 -8043 -24234 -8008
rect -24200 -8022 -24162 -8008
rect -23762 -8022 -23736 -7992
rect -22598 -8008 -22425 -7992
rect -24200 -8043 -24184 -8022
rect -24335 -8059 -24184 -8043
rect -22598 -8043 -22497 -8008
rect -22463 -8022 -22425 -8008
rect -22025 -8022 -21999 -7992
rect -20873 -7997 -20854 -7887
rect -20807 -7980 -20363 -7887
rect -20299 -7858 -20077 -7829
rect -20299 -7903 -20269 -7858
rect -20139 -7903 -20077 -7858
rect -20299 -7922 -20077 -7903
rect -20011 -7830 -19981 -7799
rect -19915 -7830 -19885 -7799
rect -19819 -7830 -19789 -7799
rect -20011 -7863 -19789 -7830
rect -20011 -7908 -19938 -7863
rect -19808 -7908 -19789 -7863
rect -20011 -7923 -19789 -7908
rect -19723 -7830 -19693 -7799
rect -19627 -7830 -19597 -7799
rect -19531 -7830 -19501 -7799
rect -19439 -7830 -19409 -7799
rect -19120 -7830 -19090 -7799
rect -19028 -7830 -18998 -7799
rect -18932 -7830 -18902 -7799
rect -18836 -7830 -18806 -7799
rect -18740 -7829 -18710 -7799
rect -18644 -7829 -18614 -7799
rect -18548 -7829 -18518 -7799
rect -20807 -7997 -19789 -7980
rect -22463 -8043 -22447 -8022
rect -22598 -8059 -22447 -8043
rect -20873 -8089 -19789 -7997
rect -20712 -8264 -20636 -8089
rect -20587 -8179 -20365 -8154
rect -20587 -8224 -20544 -8179
rect -20414 -8224 -20365 -8179
rect -20679 -8289 -20649 -8264
rect -20587 -8267 -20365 -8224
rect -20587 -8289 -20557 -8267
rect -20491 -8289 -20461 -8267
rect -20395 -8289 -20365 -8267
rect -20299 -8187 -20077 -8159
rect -20299 -8232 -20261 -8187
rect -20131 -8232 -20077 -8187
rect -20299 -8267 -20077 -8232
rect -20299 -8289 -20269 -8267
rect -20203 -8289 -20173 -8267
rect -20107 -8289 -20077 -8267
rect -20011 -8267 -19789 -8089
rect -20011 -8289 -19981 -8267
rect -19915 -8289 -19885 -8267
rect -19819 -8289 -19789 -8267
rect -19723 -7987 -19409 -7830
rect -19153 -7917 -18804 -7830
rect -19723 -8042 -19691 -7987
rect -19626 -8042 -19409 -7987
rect -19723 -8267 -19409 -8042
rect -19342 -7932 -18804 -7917
rect -18740 -7858 -18518 -7829
rect -18740 -7903 -18710 -7858
rect -18580 -7903 -18518 -7858
rect -18740 -7922 -18518 -7903
rect -18452 -7830 -18422 -7799
rect -18356 -7830 -18326 -7799
rect -18260 -7830 -18230 -7799
rect -18452 -7863 -18230 -7830
rect -18452 -7908 -18379 -7863
rect -18249 -7908 -18230 -7863
rect -18452 -7923 -18230 -7908
rect -18164 -7830 -18134 -7799
rect -18068 -7830 -18038 -7799
rect -17972 -7830 -17942 -7799
rect -17880 -7830 -17850 -7799
rect -17388 -7830 -17358 -7799
rect -17296 -7830 -17266 -7799
rect -17200 -7830 -17170 -7799
rect -17104 -7830 -17074 -7799
rect -17008 -7829 -16978 -7799
rect -16912 -7829 -16882 -7799
rect -16816 -7829 -16786 -7799
rect -19342 -8072 -19297 -7932
rect -19224 -7980 -18804 -7932
rect -19224 -8072 -18230 -7980
rect -19342 -8089 -18230 -8072
rect -19153 -8264 -19077 -8089
rect -19028 -8179 -18806 -8154
rect -19028 -8224 -18985 -8179
rect -18855 -8224 -18806 -8179
rect -19723 -8289 -19693 -8267
rect -19627 -8289 -19597 -8267
rect -19531 -8289 -19501 -8267
rect -19439 -8289 -19409 -8267
rect -19120 -8289 -19090 -8264
rect -19028 -8267 -18806 -8224
rect -19028 -8289 -18998 -8267
rect -18932 -8289 -18902 -8267
rect -18836 -8289 -18806 -8267
rect -18740 -8187 -18518 -8159
rect -18740 -8232 -18702 -8187
rect -18572 -8232 -18518 -8187
rect -18740 -8267 -18518 -8232
rect -18740 -8289 -18710 -8267
rect -18644 -8289 -18614 -8267
rect -18548 -8289 -18518 -8267
rect -18452 -8267 -18230 -8089
rect -18452 -8289 -18422 -8267
rect -18356 -8289 -18326 -8267
rect -18260 -8289 -18230 -8267
rect -18164 -7987 -17850 -7830
rect -18164 -8042 -18132 -7987
rect -18067 -8042 -17850 -7987
rect -18164 -8267 -17850 -8042
rect -17582 -7887 -17072 -7830
rect -17582 -7997 -17563 -7887
rect -17516 -7980 -17072 -7887
rect -17008 -7858 -16786 -7829
rect -17008 -7903 -16978 -7858
rect -16848 -7903 -16786 -7858
rect -17008 -7922 -16786 -7903
rect -16720 -7830 -16690 -7799
rect -16624 -7830 -16594 -7799
rect -16528 -7830 -16498 -7799
rect -16720 -7863 -16498 -7830
rect -16720 -7908 -16647 -7863
rect -16517 -7908 -16498 -7863
rect -16720 -7923 -16498 -7908
rect -16432 -7830 -16402 -7799
rect -16336 -7830 -16306 -7799
rect -16240 -7830 -16210 -7799
rect -16148 -7830 -16118 -7799
rect -15829 -7830 -15799 -7799
rect -15737 -7830 -15707 -7799
rect -15641 -7830 -15611 -7799
rect -15545 -7830 -15515 -7799
rect -15449 -7829 -15419 -7799
rect -15353 -7829 -15323 -7799
rect -15257 -7829 -15227 -7799
rect -17516 -7997 -16498 -7980
rect -17582 -8089 -16498 -7997
rect -17421 -8264 -17345 -8089
rect -17296 -8179 -17074 -8154
rect -17296 -8224 -17253 -8179
rect -17123 -8224 -17074 -8179
rect -18164 -8289 -18134 -8267
rect -18068 -8289 -18038 -8267
rect -17972 -8289 -17942 -8267
rect -17880 -8289 -17850 -8267
rect -17388 -8289 -17358 -8264
rect -17296 -8267 -17074 -8224
rect -17296 -8289 -17266 -8267
rect -17200 -8289 -17170 -8267
rect -17104 -8289 -17074 -8267
rect -17008 -8187 -16786 -8159
rect -17008 -8232 -16970 -8187
rect -16840 -8232 -16786 -8187
rect -17008 -8267 -16786 -8232
rect -17008 -8289 -16978 -8267
rect -16912 -8289 -16882 -8267
rect -16816 -8289 -16786 -8267
rect -16720 -8267 -16498 -8089
rect -16720 -8289 -16690 -8267
rect -16624 -8289 -16594 -8267
rect -16528 -8289 -16498 -8267
rect -16432 -7987 -16118 -7830
rect -15862 -7917 -15513 -7830
rect -16432 -8042 -16400 -7987
rect -16335 -8042 -16118 -7987
rect -16432 -8267 -16118 -8042
rect -16051 -7932 -15513 -7917
rect -15449 -7858 -15227 -7829
rect -15449 -7903 -15419 -7858
rect -15289 -7903 -15227 -7858
rect -15449 -7922 -15227 -7903
rect -15161 -7830 -15131 -7799
rect -15065 -7830 -15035 -7799
rect -14969 -7830 -14939 -7799
rect -15161 -7863 -14939 -7830
rect -15161 -7908 -15088 -7863
rect -14958 -7908 -14939 -7863
rect -15161 -7923 -14939 -7908
rect -14873 -7830 -14843 -7799
rect -14777 -7830 -14747 -7799
rect -14681 -7830 -14651 -7799
rect -14589 -7830 -14559 -7799
rect -14097 -7830 -14067 -7799
rect -14005 -7830 -13975 -7799
rect -13909 -7830 -13879 -7799
rect -13813 -7830 -13783 -7799
rect -13717 -7829 -13687 -7799
rect -13621 -7829 -13591 -7799
rect -13525 -7829 -13495 -7799
rect -16051 -8072 -16006 -7932
rect -15933 -7980 -15513 -7932
rect -15933 -8072 -14939 -7980
rect -16051 -8089 -14939 -8072
rect -15862 -8264 -15786 -8089
rect -15737 -8179 -15515 -8154
rect -15737 -8224 -15694 -8179
rect -15564 -8224 -15515 -8179
rect -16432 -8289 -16402 -8267
rect -16336 -8289 -16306 -8267
rect -16240 -8289 -16210 -8267
rect -16148 -8289 -16118 -8267
rect -15829 -8289 -15799 -8264
rect -15737 -8267 -15515 -8224
rect -15737 -8289 -15707 -8267
rect -15641 -8289 -15611 -8267
rect -15545 -8289 -15515 -8267
rect -15449 -8187 -15227 -8159
rect -15449 -8232 -15411 -8187
rect -15281 -8232 -15227 -8187
rect -15449 -8267 -15227 -8232
rect -15449 -8289 -15419 -8267
rect -15353 -8289 -15323 -8267
rect -15257 -8289 -15227 -8267
rect -15161 -8267 -14939 -8089
rect -15161 -8289 -15131 -8267
rect -15065 -8289 -15035 -8267
rect -14969 -8289 -14939 -8267
rect -14873 -7987 -14559 -7830
rect -14873 -8042 -14841 -7987
rect -14776 -8042 -14559 -7987
rect -14873 -8267 -14559 -8042
rect -14291 -7887 -13781 -7830
rect -14291 -7997 -14272 -7887
rect -14225 -7980 -13781 -7887
rect -13717 -7858 -13495 -7829
rect -13717 -7903 -13687 -7858
rect -13557 -7903 -13495 -7858
rect -13717 -7922 -13495 -7903
rect -13429 -7830 -13399 -7799
rect -13333 -7830 -13303 -7799
rect -13237 -7830 -13207 -7799
rect -13429 -7863 -13207 -7830
rect -13429 -7908 -13356 -7863
rect -13226 -7908 -13207 -7863
rect -13429 -7923 -13207 -7908
rect -13141 -7830 -13111 -7799
rect -13045 -7830 -13015 -7799
rect -12949 -7830 -12919 -7799
rect -12857 -7830 -12827 -7799
rect -12538 -7830 -12508 -7799
rect -12446 -7830 -12416 -7799
rect -12350 -7830 -12320 -7799
rect -12254 -7830 -12224 -7799
rect -12158 -7829 -12128 -7799
rect -12062 -7829 -12032 -7799
rect -11966 -7829 -11936 -7799
rect -14225 -7997 -13207 -7980
rect -14291 -8089 -13207 -7997
rect -14130 -8264 -14054 -8089
rect -14005 -8179 -13783 -8154
rect -14005 -8224 -13962 -8179
rect -13832 -8224 -13783 -8179
rect -14873 -8289 -14843 -8267
rect -14777 -8289 -14747 -8267
rect -14681 -8289 -14651 -8267
rect -14589 -8289 -14559 -8267
rect -14097 -8289 -14067 -8264
rect -14005 -8267 -13783 -8224
rect -14005 -8289 -13975 -8267
rect -13909 -8289 -13879 -8267
rect -13813 -8289 -13783 -8267
rect -13717 -8187 -13495 -8159
rect -13717 -8232 -13679 -8187
rect -13549 -8232 -13495 -8187
rect -13717 -8267 -13495 -8232
rect -13717 -8289 -13687 -8267
rect -13621 -8289 -13591 -8267
rect -13525 -8289 -13495 -8267
rect -13429 -8267 -13207 -8089
rect -13429 -8289 -13399 -8267
rect -13333 -8289 -13303 -8267
rect -13237 -8289 -13207 -8267
rect -13141 -7987 -12827 -7830
rect -12571 -7917 -12222 -7830
rect -13141 -8042 -13109 -7987
rect -13044 -8042 -12827 -7987
rect -13141 -8267 -12827 -8042
rect -12760 -7932 -12222 -7917
rect -12158 -7858 -11936 -7829
rect -12158 -7903 -12128 -7858
rect -11998 -7903 -11936 -7858
rect -12158 -7922 -11936 -7903
rect -11870 -7830 -11840 -7799
rect -11774 -7830 -11744 -7799
rect -11678 -7830 -11648 -7799
rect -11870 -7863 -11648 -7830
rect -11870 -7908 -11797 -7863
rect -11667 -7908 -11648 -7863
rect -11870 -7923 -11648 -7908
rect -11582 -7830 -11552 -7799
rect -11486 -7830 -11456 -7799
rect -11390 -7830 -11360 -7799
rect -11298 -7830 -11268 -7799
rect -10806 -7830 -10776 -7799
rect -10714 -7830 -10684 -7799
rect -10618 -7830 -10588 -7799
rect -10522 -7830 -10492 -7799
rect -10426 -7829 -10396 -7799
rect -10330 -7829 -10300 -7799
rect -10234 -7829 -10204 -7799
rect -12760 -8072 -12715 -7932
rect -12642 -7980 -12222 -7932
rect -12642 -8072 -11648 -7980
rect -12760 -8089 -11648 -8072
rect -12571 -8264 -12495 -8089
rect -12446 -8179 -12224 -8154
rect -12446 -8224 -12403 -8179
rect -12273 -8224 -12224 -8179
rect -13141 -8289 -13111 -8267
rect -13045 -8289 -13015 -8267
rect -12949 -8289 -12919 -8267
rect -12857 -8289 -12827 -8267
rect -12538 -8289 -12508 -8264
rect -12446 -8267 -12224 -8224
rect -12446 -8289 -12416 -8267
rect -12350 -8289 -12320 -8267
rect -12254 -8289 -12224 -8267
rect -12158 -8187 -11936 -8159
rect -12158 -8232 -12120 -8187
rect -11990 -8232 -11936 -8187
rect -12158 -8267 -11936 -8232
rect -12158 -8289 -12128 -8267
rect -12062 -8289 -12032 -8267
rect -11966 -8289 -11936 -8267
rect -11870 -8267 -11648 -8089
rect -11870 -8289 -11840 -8267
rect -11774 -8289 -11744 -8267
rect -11678 -8289 -11648 -8267
rect -11582 -7987 -11268 -7830
rect -11582 -8042 -11550 -7987
rect -11485 -8042 -11268 -7987
rect -11582 -8267 -11268 -8042
rect -11000 -7887 -10490 -7830
rect -11000 -7997 -10981 -7887
rect -10934 -7980 -10490 -7887
rect -10426 -7858 -10204 -7829
rect -10426 -7903 -10396 -7858
rect -10266 -7903 -10204 -7858
rect -10426 -7922 -10204 -7903
rect -10138 -7830 -10108 -7799
rect -10042 -7830 -10012 -7799
rect -9946 -7830 -9916 -7799
rect -10138 -7863 -9916 -7830
rect -10138 -7908 -10065 -7863
rect -9935 -7908 -9916 -7863
rect -10138 -7923 -9916 -7908
rect -9850 -7830 -9820 -7799
rect -9754 -7830 -9724 -7799
rect -9658 -7830 -9628 -7799
rect -9566 -7830 -9536 -7799
rect -9247 -7830 -9217 -7799
rect -9155 -7830 -9125 -7799
rect -9059 -7830 -9029 -7799
rect -8963 -7830 -8933 -7799
rect -8867 -7829 -8837 -7799
rect -8771 -7829 -8741 -7799
rect -8675 -7829 -8645 -7799
rect -10934 -7997 -9916 -7980
rect -11000 -8089 -9916 -7997
rect -10839 -8264 -10763 -8089
rect -10714 -8179 -10492 -8154
rect -10714 -8224 -10671 -8179
rect -10541 -8224 -10492 -8179
rect -11582 -8289 -11552 -8267
rect -11486 -8289 -11456 -8267
rect -11390 -8289 -11360 -8267
rect -11298 -8289 -11268 -8267
rect -10806 -8289 -10776 -8264
rect -10714 -8267 -10492 -8224
rect -10714 -8289 -10684 -8267
rect -10618 -8289 -10588 -8267
rect -10522 -8289 -10492 -8267
rect -10426 -8187 -10204 -8159
rect -10426 -8232 -10388 -8187
rect -10258 -8232 -10204 -8187
rect -10426 -8267 -10204 -8232
rect -10426 -8289 -10396 -8267
rect -10330 -8289 -10300 -8267
rect -10234 -8289 -10204 -8267
rect -10138 -8267 -9916 -8089
rect -10138 -8289 -10108 -8267
rect -10042 -8289 -10012 -8267
rect -9946 -8289 -9916 -8267
rect -9850 -7987 -9536 -7830
rect -9280 -7917 -8931 -7830
rect -9850 -8042 -9818 -7987
rect -9753 -8042 -9536 -7987
rect -9850 -8267 -9536 -8042
rect -9469 -7932 -8931 -7917
rect -8867 -7858 -8645 -7829
rect -8867 -7903 -8837 -7858
rect -8707 -7903 -8645 -7858
rect -8867 -7922 -8645 -7903
rect -8579 -7830 -8549 -7799
rect -8483 -7830 -8453 -7799
rect -8387 -7830 -8357 -7799
rect -8579 -7863 -8357 -7830
rect -8579 -7908 -8506 -7863
rect -8376 -7908 -8357 -7863
rect -8579 -7923 -8357 -7908
rect -8291 -7830 -8261 -7799
rect -8195 -7830 -8165 -7799
rect -8099 -7830 -8069 -7799
rect -8007 -7830 -7977 -7799
rect -9469 -8072 -9424 -7932
rect -9351 -7980 -8931 -7932
rect -9351 -8072 -8357 -7980
rect -9469 -8089 -8357 -8072
rect -9280 -8264 -9204 -8089
rect -9155 -8179 -8933 -8154
rect -9155 -8224 -9112 -8179
rect -8982 -8224 -8933 -8179
rect -9850 -8289 -9820 -8267
rect -9754 -8289 -9724 -8267
rect -9658 -8289 -9628 -8267
rect -9566 -8289 -9536 -8267
rect -9247 -8289 -9217 -8264
rect -9155 -8267 -8933 -8224
rect -9155 -8289 -9125 -8267
rect -9059 -8289 -9029 -8267
rect -8963 -8289 -8933 -8267
rect -8867 -8187 -8645 -8159
rect -8867 -8232 -8829 -8187
rect -8699 -8232 -8645 -8187
rect -8867 -8267 -8645 -8232
rect -8867 -8289 -8837 -8267
rect -8771 -8289 -8741 -8267
rect -8675 -8289 -8645 -8267
rect -8579 -8267 -8357 -8089
rect -8579 -8289 -8549 -8267
rect -8483 -8289 -8453 -8267
rect -8387 -8289 -8357 -8267
rect -8291 -7987 -7977 -7830
rect -8291 -8042 -8259 -7987
rect -8194 -8042 -7977 -7987
rect -8291 -8267 -7977 -8042
rect 11164 -7394 11194 -7368
rect 11260 -7394 11290 -7368
rect 11356 -7394 11386 -7368
rect 11452 -7394 11482 -7368
rect 7422 -8227 7452 -8194
rect -8291 -8289 -8261 -8267
rect -8195 -8289 -8165 -8267
rect -8099 -8289 -8069 -8267
rect -8007 -8289 -7977 -8267
rect 7238 -8257 7452 -8227
rect -20679 -8445 -20649 -8419
rect -20587 -8445 -20557 -8419
rect -20491 -8445 -20461 -8419
rect -20395 -8445 -20365 -8419
rect -20299 -8445 -20269 -8419
rect -20203 -8445 -20173 -8419
rect -20107 -8445 -20077 -8419
rect -20011 -8445 -19981 -8419
rect -19915 -8445 -19885 -8419
rect -19819 -8445 -19789 -8419
rect -19723 -8445 -19693 -8419
rect -19627 -8445 -19597 -8419
rect -19531 -8445 -19501 -8419
rect -19439 -8445 -19409 -8419
rect -19120 -8445 -19090 -8419
rect -19028 -8445 -18998 -8419
rect -18932 -8445 -18902 -8419
rect -18836 -8445 -18806 -8419
rect -18740 -8445 -18710 -8419
rect -18644 -8445 -18614 -8419
rect -18548 -8445 -18518 -8419
rect -18452 -8445 -18422 -8419
rect -18356 -8445 -18326 -8419
rect -18260 -8445 -18230 -8419
rect -18164 -8445 -18134 -8419
rect -18068 -8445 -18038 -8419
rect -17972 -8445 -17942 -8419
rect -17880 -8445 -17850 -8419
rect -17388 -8445 -17358 -8419
rect -17296 -8445 -17266 -8419
rect -17200 -8445 -17170 -8419
rect -17104 -8445 -17074 -8419
rect -17008 -8445 -16978 -8419
rect -16912 -8445 -16882 -8419
rect -16816 -8445 -16786 -8419
rect -16720 -8445 -16690 -8419
rect -16624 -8445 -16594 -8419
rect -16528 -8445 -16498 -8419
rect -16432 -8445 -16402 -8419
rect -16336 -8445 -16306 -8419
rect -16240 -8445 -16210 -8419
rect -16148 -8445 -16118 -8419
rect -15829 -8445 -15799 -8419
rect -15737 -8445 -15707 -8419
rect -15641 -8445 -15611 -8419
rect -15545 -8445 -15515 -8419
rect -15449 -8445 -15419 -8419
rect -15353 -8445 -15323 -8419
rect -15257 -8445 -15227 -8419
rect -15161 -8445 -15131 -8419
rect -15065 -8445 -15035 -8419
rect -14969 -8445 -14939 -8419
rect -14873 -8445 -14843 -8419
rect -14777 -8445 -14747 -8419
rect -14681 -8445 -14651 -8419
rect -14589 -8445 -14559 -8419
rect -14097 -8445 -14067 -8419
rect -14005 -8445 -13975 -8419
rect -13909 -8445 -13879 -8419
rect -13813 -8445 -13783 -8419
rect -13717 -8445 -13687 -8419
rect -13621 -8445 -13591 -8419
rect -13525 -8445 -13495 -8419
rect -13429 -8445 -13399 -8419
rect -13333 -8445 -13303 -8419
rect -13237 -8445 -13207 -8419
rect -13141 -8445 -13111 -8419
rect -13045 -8445 -13015 -8419
rect -12949 -8445 -12919 -8419
rect -12857 -8445 -12827 -8419
rect -12538 -8445 -12508 -8419
rect -12446 -8445 -12416 -8419
rect -12350 -8445 -12320 -8419
rect -12254 -8445 -12224 -8419
rect -12158 -8445 -12128 -8419
rect -12062 -8445 -12032 -8419
rect -11966 -8445 -11936 -8419
rect -11870 -8445 -11840 -8419
rect -11774 -8445 -11744 -8419
rect -11678 -8445 -11648 -8419
rect -11582 -8445 -11552 -8419
rect -11486 -8445 -11456 -8419
rect -11390 -8445 -11360 -8419
rect -11298 -8445 -11268 -8419
rect -10806 -8445 -10776 -8419
rect -10714 -8445 -10684 -8419
rect -10618 -8445 -10588 -8419
rect -10522 -8445 -10492 -8419
rect -10426 -8445 -10396 -8419
rect -10330 -8445 -10300 -8419
rect -10234 -8445 -10204 -8419
rect -10138 -8445 -10108 -8419
rect -10042 -8445 -10012 -8419
rect -9946 -8445 -9916 -8419
rect -9850 -8445 -9820 -8419
rect -9754 -8445 -9724 -8419
rect -9658 -8445 -9628 -8419
rect -9566 -8445 -9536 -8419
rect -9247 -8445 -9217 -8419
rect -9155 -8445 -9125 -8419
rect -9059 -8445 -9029 -8419
rect -8963 -8445 -8933 -8419
rect -8867 -8445 -8837 -8419
rect -8771 -8445 -8741 -8419
rect -8675 -8445 -8645 -8419
rect -8579 -8445 -8549 -8419
rect -8483 -8445 -8453 -8419
rect -8387 -8445 -8357 -8419
rect -8291 -8445 -8261 -8419
rect -8195 -8445 -8165 -8419
rect -8099 -8445 -8069 -8419
rect -8007 -8445 -7977 -8419
rect 7238 -8504 7268 -8257
rect 7518 -8299 7548 -8194
rect 7614 -8217 7644 -8194
rect 7374 -8437 7548 -8299
rect 7182 -8520 7326 -8504
rect 7182 -8554 7198 -8520
rect 7232 -8554 7326 -8520
rect 7182 -8570 7326 -8554
rect 7374 -8520 7518 -8437
rect 7590 -8479 7644 -8217
rect 7710 -8344 7740 -8194
rect 8370 -8227 8400 -8194
rect 8186 -8257 8400 -8227
rect 7710 -8374 7848 -8344
rect 7584 -8504 7644 -8479
rect 7758 -8504 7848 -8374
rect 8186 -8504 8216 -8257
rect 8466 -8299 8496 -8194
rect 8562 -8217 8592 -8194
rect 8322 -8437 8496 -8299
rect 7374 -8554 7390 -8520
rect 7424 -8554 7518 -8520
rect 7374 -8570 7518 -8554
rect 7566 -8520 7710 -8504
rect 7566 -8554 7582 -8520
rect 7616 -8554 7710 -8520
rect 7566 -8570 7710 -8554
rect 7758 -8520 7902 -8504
rect 7758 -8554 7774 -8520
rect 7808 -8554 7902 -8520
rect 7758 -8570 7902 -8554
rect 8130 -8520 8274 -8504
rect 8130 -8554 8146 -8520
rect 8180 -8554 8274 -8520
rect 8130 -8570 8274 -8554
rect 8322 -8520 8466 -8437
rect 8538 -8479 8592 -8217
rect 8658 -8344 8688 -8194
rect 9306 -8227 9336 -8194
rect 9122 -8257 9336 -8227
rect 8658 -8374 8796 -8344
rect 8532 -8504 8592 -8479
rect 8706 -8504 8796 -8374
rect 9122 -8504 9152 -8257
rect 9402 -8299 9432 -8194
rect 9498 -8217 9528 -8194
rect 9258 -8437 9432 -8299
rect 8322 -8554 8338 -8520
rect 8372 -8554 8466 -8520
rect 8322 -8570 8466 -8554
rect 8514 -8520 8658 -8504
rect 8514 -8554 8530 -8520
rect 8564 -8554 8658 -8520
rect 8514 -8570 8658 -8554
rect 8706 -8520 8850 -8504
rect 8706 -8554 8722 -8520
rect 8756 -8554 8850 -8520
rect 8706 -8570 8850 -8554
rect 9066 -8520 9210 -8504
rect 9066 -8554 9082 -8520
rect 9116 -8554 9210 -8520
rect 9066 -8570 9210 -8554
rect 9258 -8520 9402 -8437
rect 9474 -8479 9528 -8217
rect 9594 -8344 9624 -8194
rect 10237 -8226 10267 -8193
rect 10053 -8256 10267 -8226
rect 9594 -8374 9732 -8344
rect 9468 -8504 9528 -8479
rect 9642 -8504 9732 -8374
rect 10053 -8503 10083 -8256
rect 10333 -8298 10363 -8193
rect 10429 -8216 10459 -8193
rect 10189 -8436 10363 -8298
rect 9258 -8554 9274 -8520
rect 9308 -8554 9402 -8520
rect 9258 -8570 9402 -8554
rect 9450 -8520 9594 -8504
rect 9450 -8554 9466 -8520
rect 9500 -8554 9594 -8520
rect 9450 -8570 9594 -8554
rect 9642 -8520 9786 -8504
rect 9642 -8554 9658 -8520
rect 9692 -8554 9786 -8520
rect 9642 -8570 9786 -8554
rect 9997 -8519 10141 -8503
rect 9997 -8553 10013 -8519
rect 10047 -8553 10141 -8519
rect 9997 -8569 10141 -8553
rect 10189 -8519 10333 -8436
rect 10405 -8478 10459 -8216
rect 10525 -8343 10555 -8193
rect 12219 -7436 12249 -7300
rect 12315 -7229 12345 -7203
rect 12411 -7229 12441 -7203
rect 12507 -7229 12537 -7203
rect 12603 -7229 12633 -7203
rect 12699 -7229 12729 -7203
rect 12315 -7300 12729 -7229
rect 12315 -7342 12345 -7300
rect 12826 -7337 12842 -7111
rect 12876 -7113 12892 -7111
rect 12876 -7143 12923 -7113
rect 13137 -7143 13163 -7113
rect 12876 -7209 12892 -7143
rect 12876 -7239 12923 -7209
rect 13137 -7239 13163 -7209
rect 12876 -7305 12892 -7239
rect 12876 -7335 12923 -7305
rect 13137 -7335 13163 -7305
rect 12876 -7337 12892 -7335
rect 12297 -7358 12363 -7342
rect 12826 -7353 12892 -7337
rect 12297 -7392 12313 -7358
rect 12347 -7392 12363 -7358
rect 12297 -7408 12363 -7392
rect 12315 -7436 12345 -7408
rect 12826 -7557 12893 -7541
rect 12826 -7591 12842 -7557
rect 12876 -7559 12893 -7557
rect 12876 -7589 12923 -7559
rect 13123 -7589 13149 -7559
rect 12876 -7591 12893 -7589
rect 12826 -7607 12893 -7591
rect 12219 -7662 12249 -7636
rect 12315 -7662 12345 -7636
rect 11164 -8227 11194 -8194
rect 10980 -8257 11194 -8227
rect 10525 -8373 10663 -8343
rect 10399 -8503 10459 -8478
rect 10573 -8503 10663 -8373
rect 10189 -8553 10205 -8519
rect 10239 -8553 10333 -8519
rect 10189 -8569 10333 -8553
rect 10381 -8519 10525 -8503
rect 10381 -8553 10397 -8519
rect 10431 -8553 10525 -8519
rect 10381 -8569 10525 -8553
rect 10573 -8519 10717 -8503
rect 10980 -8504 11010 -8257
rect 11260 -8299 11290 -8194
rect 11356 -8217 11386 -8194
rect 11116 -8437 11290 -8299
rect 10573 -8553 10589 -8519
rect 10623 -8553 10717 -8519
rect 10573 -8569 10717 -8553
rect 7200 -8601 7230 -8570
rect 7296 -8601 7326 -8570
rect 7392 -8601 7422 -8570
rect 7488 -8601 7518 -8570
rect 7584 -8601 7614 -8570
rect 7680 -8601 7710 -8570
rect 7776 -8601 7806 -8570
rect 7872 -8601 7902 -8570
rect 8148 -8601 8178 -8570
rect 8244 -8601 8274 -8570
rect 8340 -8601 8370 -8570
rect 8436 -8601 8466 -8570
rect 8532 -8601 8562 -8570
rect 8628 -8601 8658 -8570
rect 8724 -8601 8754 -8570
rect 8820 -8601 8850 -8570
rect 9084 -8601 9114 -8570
rect 9180 -8601 9210 -8570
rect 9276 -8601 9306 -8570
rect 9372 -8601 9402 -8570
rect 9468 -8601 9498 -8570
rect 9564 -8601 9594 -8570
rect 9660 -8601 9690 -8570
rect 9756 -8601 9786 -8570
rect 10015 -8600 10045 -8569
rect 10111 -8600 10141 -8569
rect 10207 -8600 10237 -8569
rect 10303 -8600 10333 -8569
rect 10399 -8600 10429 -8569
rect 10495 -8600 10525 -8569
rect 10591 -8600 10621 -8569
rect 10687 -8600 10717 -8569
rect 10924 -8520 11068 -8504
rect 10924 -8554 10940 -8520
rect 10974 -8554 11068 -8520
rect 10924 -8570 11068 -8554
rect 11116 -8520 11260 -8437
rect 11332 -8479 11386 -8217
rect 11452 -8344 11482 -8194
rect 11452 -8374 11590 -8344
rect 11326 -8504 11386 -8479
rect 11500 -8504 11590 -8374
rect 11116 -8554 11132 -8520
rect 11166 -8554 11260 -8520
rect 11116 -8570 11260 -8554
rect 11308 -8520 11452 -8504
rect 11308 -8554 11324 -8520
rect 11358 -8554 11452 -8520
rect 11308 -8570 11452 -8554
rect 11500 -8520 11644 -8504
rect 11500 -8554 11516 -8520
rect 11550 -8554 11644 -8520
rect 11500 -8570 11644 -8554
rect -23680 -8736 -23614 -8720
rect -24334 -8782 -24304 -8751
rect -24238 -8782 -24208 -8751
rect -24142 -8782 -24112 -8751
rect -24046 -8782 -24016 -8751
rect -23950 -8782 -23920 -8751
rect -23854 -8782 -23824 -8751
rect -23680 -8962 -23664 -8736
rect -23630 -8738 -23614 -8736
rect -21943 -8736 -21877 -8720
rect -23630 -8768 -23583 -8738
rect -23369 -8768 -23343 -8738
rect -23630 -8834 -23614 -8768
rect -22598 -8782 -22568 -8751
rect -22502 -8782 -22472 -8751
rect -22406 -8782 -22376 -8751
rect -22310 -8782 -22280 -8751
rect -22214 -8782 -22184 -8751
rect -22118 -8782 -22088 -8751
rect -23630 -8864 -23583 -8834
rect -23369 -8864 -23343 -8834
rect -23630 -8930 -23614 -8864
rect -23630 -8960 -23583 -8930
rect -23369 -8960 -23343 -8930
rect -23630 -8962 -23614 -8960
rect -23680 -8978 -23614 -8962
rect -24334 -9022 -24304 -8996
rect -24238 -9022 -24208 -8996
rect -24142 -9022 -24112 -8996
rect -24335 -9043 -24112 -9022
rect -24335 -9078 -24318 -9043
rect -24284 -9052 -24112 -9043
rect -24046 -9022 -24016 -8996
rect -23950 -9022 -23920 -8996
rect -23854 -9022 -23824 -8996
rect -21943 -8962 -21927 -8736
rect -21893 -8738 -21877 -8736
rect -21893 -8768 -21846 -8738
rect -21632 -8768 -21606 -8738
rect -21893 -8834 -21877 -8768
rect -21893 -8864 -21846 -8834
rect -21632 -8864 -21606 -8834
rect -21893 -8930 -21877 -8864
rect -21893 -8960 -21846 -8930
rect -21632 -8960 -21606 -8930
rect -20468 -8950 -20438 -8919
rect -20372 -8950 -20342 -8919
rect -20276 -8950 -20246 -8919
rect -20180 -8950 -20150 -8919
rect -20084 -8950 -20054 -8919
rect -19988 -8950 -19958 -8919
rect -19359 -8950 -19329 -8919
rect -19263 -8950 -19233 -8919
rect -19167 -8950 -19137 -8919
rect -19071 -8950 -19041 -8919
rect -18975 -8950 -18945 -8919
rect -18879 -8950 -18849 -8919
rect -18477 -8950 -18447 -8919
rect -18381 -8950 -18351 -8919
rect -18285 -8950 -18255 -8919
rect -18189 -8950 -18159 -8919
rect -18093 -8950 -18063 -8919
rect -17997 -8950 -17967 -8919
rect -17177 -8950 -17147 -8919
rect -17081 -8950 -17051 -8919
rect -16985 -8950 -16955 -8919
rect -16889 -8950 -16859 -8919
rect -16793 -8950 -16763 -8919
rect -16697 -8950 -16667 -8919
rect -16068 -8950 -16038 -8919
rect -15972 -8950 -15942 -8919
rect -15876 -8950 -15846 -8919
rect -15780 -8950 -15750 -8919
rect -15684 -8950 -15654 -8919
rect -15588 -8950 -15558 -8919
rect -15186 -8950 -15156 -8919
rect -15090 -8950 -15060 -8919
rect -14994 -8950 -14964 -8919
rect -14898 -8950 -14868 -8919
rect -14802 -8950 -14772 -8919
rect -14706 -8950 -14676 -8919
rect -13886 -8950 -13856 -8919
rect -13790 -8950 -13760 -8919
rect -13694 -8950 -13664 -8919
rect -13598 -8950 -13568 -8919
rect -13502 -8950 -13472 -8919
rect -13406 -8950 -13376 -8919
rect -12777 -8950 -12747 -8919
rect -12681 -8950 -12651 -8919
rect -12585 -8950 -12555 -8919
rect -12489 -8950 -12459 -8919
rect -12393 -8950 -12363 -8919
rect -12297 -8950 -12267 -8919
rect -11895 -8950 -11865 -8919
rect -11799 -8950 -11769 -8919
rect -11703 -8950 -11673 -8919
rect -11607 -8950 -11577 -8919
rect -11511 -8950 -11481 -8919
rect -11415 -8950 -11385 -8919
rect -10595 -8950 -10565 -8919
rect -10499 -8950 -10469 -8919
rect -10403 -8950 -10373 -8919
rect -10307 -8950 -10277 -8919
rect -10211 -8950 -10181 -8919
rect -10115 -8950 -10085 -8919
rect -9486 -8950 -9456 -8919
rect -9390 -8950 -9360 -8919
rect -9294 -8950 -9264 -8919
rect -9198 -8950 -9168 -8919
rect -9102 -8950 -9072 -8919
rect -9006 -8950 -8976 -8919
rect -8604 -8950 -8574 -8919
rect -8508 -8950 -8478 -8919
rect -8412 -8950 -8382 -8919
rect -8316 -8950 -8286 -8919
rect -8220 -8950 -8190 -8919
rect -8124 -8950 -8094 -8919
rect 10942 -8601 10972 -8570
rect 11038 -8601 11068 -8570
rect 11134 -8601 11164 -8570
rect 11230 -8601 11260 -8570
rect 11326 -8601 11356 -8570
rect 11422 -8601 11452 -8570
rect 11518 -8601 11548 -8570
rect 11614 -8601 11644 -8570
rect 7200 -8949 7230 -8923
rect 7296 -8949 7326 -8923
rect 7392 -8949 7422 -8923
rect 7488 -8949 7518 -8923
rect 7584 -8949 7614 -8923
rect 7680 -8949 7710 -8923
rect 7776 -8949 7806 -8923
rect 7872 -8949 7902 -8923
rect 8148 -8949 8178 -8923
rect 8244 -8949 8274 -8923
rect 8340 -8949 8370 -8923
rect 8436 -8949 8466 -8923
rect 8532 -8949 8562 -8923
rect 8628 -8949 8658 -8923
rect 8724 -8949 8754 -8923
rect 8820 -8949 8850 -8923
rect 9084 -8949 9114 -8923
rect 9180 -8949 9210 -8923
rect 9276 -8949 9306 -8923
rect 9372 -8949 9402 -8923
rect 9468 -8949 9498 -8923
rect 9564 -8949 9594 -8923
rect 9660 -8949 9690 -8923
rect 9756 -8949 9786 -8923
rect 10015 -8948 10045 -8922
rect 10111 -8948 10141 -8922
rect 10207 -8948 10237 -8922
rect 10303 -8948 10333 -8922
rect 10399 -8948 10429 -8922
rect 10495 -8948 10525 -8922
rect 10591 -8948 10621 -8922
rect 10687 -8948 10717 -8922
rect 10942 -8949 10972 -8923
rect 11038 -8949 11068 -8923
rect 11134 -8949 11164 -8923
rect 11230 -8949 11260 -8923
rect 11326 -8949 11356 -8923
rect 11422 -8949 11452 -8923
rect 11518 -8949 11548 -8923
rect 11614 -8949 11644 -8923
rect -21893 -8962 -21877 -8960
rect -21943 -8978 -21877 -8962
rect -22598 -9022 -22568 -8996
rect -22502 -9022 -22472 -8996
rect -22406 -9022 -22376 -8996
rect -24046 -9043 -23824 -9022
rect -24284 -9078 -24268 -9052
rect -24335 -9089 -24268 -9078
rect -24046 -9078 -24029 -9043
rect -23995 -9052 -23824 -9043
rect -22599 -9043 -22376 -9022
rect -23995 -9078 -23979 -9052
rect -24046 -9089 -23979 -9078
rect -22599 -9078 -22582 -9043
rect -22548 -9052 -22376 -9043
rect -22310 -9022 -22280 -8996
rect -22214 -9022 -22184 -8996
rect -22118 -9022 -22088 -8996
rect -22310 -9043 -22088 -9022
rect -22548 -9078 -22532 -9052
rect -22599 -9089 -22532 -9078
rect -22310 -9078 -22293 -9043
rect -22259 -9052 -22088 -9043
rect -22259 -9078 -22243 -9052
rect -22310 -9089 -22243 -9078
rect -24335 -9284 -24292 -9089
rect -24250 -9167 -24184 -9151
rect -24250 -9202 -24234 -9167
rect -24200 -9188 -24184 -9167
rect -23680 -9182 -23613 -9166
rect -24200 -9202 -24162 -9188
rect -24250 -9218 -24162 -9202
rect -23762 -9218 -23736 -9188
rect -23680 -9216 -23664 -9182
rect -23630 -9184 -23613 -9182
rect -23630 -9214 -23583 -9184
rect -23383 -9214 -23357 -9184
rect -23630 -9216 -23613 -9214
rect -23680 -9232 -23613 -9216
rect -22599 -9284 -22556 -9089
rect -22514 -9167 -22448 -9151
rect -22514 -9202 -22498 -9167
rect -22464 -9188 -22448 -9167
rect -21943 -9182 -21876 -9166
rect -22464 -9202 -22426 -9188
rect -22514 -9218 -22426 -9202
rect -22026 -9218 -22000 -9188
rect -21943 -9216 -21927 -9182
rect -21893 -9184 -21876 -9182
rect -21893 -9214 -21846 -9184
rect -21646 -9214 -21620 -9184
rect -20468 -9190 -20438 -9164
rect -20372 -9190 -20342 -9164
rect -20276 -9190 -20246 -9164
rect -20469 -9211 -20246 -9190
rect -21893 -9216 -21876 -9214
rect -21943 -9232 -21876 -9216
rect -20469 -9246 -20452 -9211
rect -20418 -9220 -20246 -9211
rect -20180 -9190 -20150 -9164
rect -20084 -9190 -20054 -9164
rect -19988 -9190 -19958 -9164
rect -19359 -9190 -19329 -9164
rect -19263 -9190 -19233 -9164
rect -19167 -9190 -19137 -9164
rect -20180 -9211 -19958 -9190
rect -20418 -9246 -20402 -9220
rect -20469 -9257 -20402 -9246
rect -20180 -9246 -20163 -9211
rect -20129 -9220 -19958 -9211
rect -19360 -9211 -19137 -9190
rect -20129 -9246 -20113 -9220
rect -20180 -9257 -20113 -9246
rect -19360 -9246 -19343 -9211
rect -19309 -9220 -19137 -9211
rect -19071 -9190 -19041 -9164
rect -18975 -9190 -18945 -9164
rect -18879 -9190 -18849 -9164
rect -18477 -9190 -18447 -9164
rect -18381 -9190 -18351 -9164
rect -18285 -9190 -18255 -9164
rect -19071 -9211 -18849 -9190
rect -19309 -9246 -19293 -9220
rect -19360 -9257 -19293 -9246
rect -19071 -9246 -19054 -9211
rect -19020 -9220 -18849 -9211
rect -18478 -9211 -18255 -9190
rect -19020 -9246 -19004 -9220
rect -19071 -9257 -19004 -9246
rect -18478 -9246 -18461 -9211
rect -18427 -9220 -18255 -9211
rect -18189 -9190 -18159 -9164
rect -18093 -9190 -18063 -9164
rect -17997 -9190 -17967 -9164
rect -17177 -9190 -17147 -9164
rect -17081 -9190 -17051 -9164
rect -16985 -9190 -16955 -9164
rect -18189 -9211 -17967 -9190
rect -18427 -9246 -18411 -9220
rect -18478 -9257 -18411 -9246
rect -18189 -9246 -18172 -9211
rect -18138 -9220 -17967 -9211
rect -17178 -9211 -16955 -9190
rect -18138 -9246 -18122 -9220
rect -18189 -9257 -18122 -9246
rect -17178 -9246 -17161 -9211
rect -17127 -9220 -16955 -9211
rect -16889 -9190 -16859 -9164
rect -16793 -9190 -16763 -9164
rect -16697 -9190 -16667 -9164
rect -16068 -9190 -16038 -9164
rect -15972 -9190 -15942 -9164
rect -15876 -9190 -15846 -9164
rect -16889 -9211 -16667 -9190
rect -17127 -9246 -17111 -9220
rect -17178 -9257 -17111 -9246
rect -16889 -9246 -16872 -9211
rect -16838 -9220 -16667 -9211
rect -16069 -9211 -15846 -9190
rect -16838 -9246 -16822 -9220
rect -16889 -9257 -16822 -9246
rect -16069 -9246 -16052 -9211
rect -16018 -9220 -15846 -9211
rect -15780 -9190 -15750 -9164
rect -15684 -9190 -15654 -9164
rect -15588 -9190 -15558 -9164
rect -15186 -9190 -15156 -9164
rect -15090 -9190 -15060 -9164
rect -14994 -9190 -14964 -9164
rect -15780 -9211 -15558 -9190
rect -16018 -9246 -16002 -9220
rect -16069 -9257 -16002 -9246
rect -15780 -9246 -15763 -9211
rect -15729 -9220 -15558 -9211
rect -15187 -9211 -14964 -9190
rect -15729 -9246 -15713 -9220
rect -15780 -9257 -15713 -9246
rect -15187 -9246 -15170 -9211
rect -15136 -9220 -14964 -9211
rect -14898 -9190 -14868 -9164
rect -14802 -9190 -14772 -9164
rect -14706 -9190 -14676 -9164
rect -13886 -9190 -13856 -9164
rect -13790 -9190 -13760 -9164
rect -13694 -9190 -13664 -9164
rect -14898 -9211 -14676 -9190
rect -15136 -9246 -15120 -9220
rect -15187 -9257 -15120 -9246
rect -14898 -9246 -14881 -9211
rect -14847 -9220 -14676 -9211
rect -13887 -9211 -13664 -9190
rect -14847 -9246 -14831 -9220
rect -14898 -9257 -14831 -9246
rect -13887 -9246 -13870 -9211
rect -13836 -9220 -13664 -9211
rect -13598 -9190 -13568 -9164
rect -13502 -9190 -13472 -9164
rect -13406 -9190 -13376 -9164
rect -12777 -9190 -12747 -9164
rect -12681 -9190 -12651 -9164
rect -12585 -9190 -12555 -9164
rect -13598 -9211 -13376 -9190
rect -13836 -9246 -13820 -9220
rect -13887 -9257 -13820 -9246
rect -13598 -9246 -13581 -9211
rect -13547 -9220 -13376 -9211
rect -12778 -9211 -12555 -9190
rect -13547 -9246 -13531 -9220
rect -13598 -9257 -13531 -9246
rect -12778 -9246 -12761 -9211
rect -12727 -9220 -12555 -9211
rect -12489 -9190 -12459 -9164
rect -12393 -9190 -12363 -9164
rect -12297 -9190 -12267 -9164
rect -11895 -9190 -11865 -9164
rect -11799 -9190 -11769 -9164
rect -11703 -9190 -11673 -9164
rect -12489 -9211 -12267 -9190
rect -12727 -9246 -12711 -9220
rect -12778 -9257 -12711 -9246
rect -12489 -9246 -12472 -9211
rect -12438 -9220 -12267 -9211
rect -11896 -9211 -11673 -9190
rect -12438 -9246 -12422 -9220
rect -12489 -9257 -12422 -9246
rect -11896 -9246 -11879 -9211
rect -11845 -9220 -11673 -9211
rect -11607 -9190 -11577 -9164
rect -11511 -9190 -11481 -9164
rect -11415 -9190 -11385 -9164
rect -10595 -9190 -10565 -9164
rect -10499 -9190 -10469 -9164
rect -10403 -9190 -10373 -9164
rect -11607 -9211 -11385 -9190
rect -11845 -9246 -11829 -9220
rect -11896 -9257 -11829 -9246
rect -11607 -9246 -11590 -9211
rect -11556 -9220 -11385 -9211
rect -10596 -9211 -10373 -9190
rect -11556 -9246 -11540 -9220
rect -11607 -9257 -11540 -9246
rect -10596 -9246 -10579 -9211
rect -10545 -9220 -10373 -9211
rect -10307 -9190 -10277 -9164
rect -10211 -9190 -10181 -9164
rect -10115 -9190 -10085 -9164
rect -9486 -9190 -9456 -9164
rect -9390 -9190 -9360 -9164
rect -9294 -9190 -9264 -9164
rect -10307 -9211 -10085 -9190
rect -10545 -9246 -10529 -9220
rect -10596 -9257 -10529 -9246
rect -10307 -9246 -10290 -9211
rect -10256 -9220 -10085 -9211
rect -9487 -9211 -9264 -9190
rect -10256 -9246 -10240 -9220
rect -10307 -9257 -10240 -9246
rect -9487 -9246 -9470 -9211
rect -9436 -9220 -9264 -9211
rect -9198 -9190 -9168 -9164
rect -9102 -9190 -9072 -9164
rect -9006 -9190 -8976 -9164
rect -8604 -9190 -8574 -9164
rect -8508 -9190 -8478 -9164
rect -8412 -9190 -8382 -9164
rect -9198 -9211 -8976 -9190
rect -9436 -9246 -9420 -9220
rect -9487 -9257 -9420 -9246
rect -9198 -9246 -9181 -9211
rect -9147 -9220 -8976 -9211
rect -8605 -9211 -8382 -9190
rect -9147 -9246 -9131 -9220
rect -9198 -9257 -9131 -9246
rect -8605 -9246 -8588 -9211
rect -8554 -9220 -8382 -9211
rect -8316 -9190 -8286 -9164
rect -8220 -9190 -8190 -9164
rect -8124 -9190 -8094 -9164
rect -8316 -9211 -8094 -9190
rect -8554 -9246 -8538 -9220
rect -8605 -9257 -8538 -9246
rect -8316 -9246 -8299 -9211
rect -8265 -9220 -8094 -9211
rect -8265 -9246 -8249 -9220
rect -8316 -9257 -8249 -9246
rect -24335 -9300 -24162 -9284
rect -24335 -9335 -24234 -9300
rect -24200 -9314 -24162 -9300
rect -23762 -9314 -23736 -9284
rect -22599 -9300 -22426 -9284
rect -24200 -9335 -24184 -9314
rect -24335 -9351 -24184 -9335
rect -22599 -9335 -22498 -9300
rect -22464 -9314 -22426 -9300
rect -22026 -9314 -22000 -9284
rect -22464 -9335 -22448 -9314
rect -22599 -9351 -22448 -9335
rect -20469 -9452 -20426 -9257
rect -20384 -9335 -20318 -9319
rect -20384 -9370 -20368 -9335
rect -20334 -9356 -20318 -9335
rect -20334 -9370 -20296 -9356
rect -20384 -9386 -20296 -9370
rect -19896 -9386 -19870 -9356
rect -19360 -9452 -19317 -9257
rect -19275 -9335 -19209 -9319
rect -19275 -9370 -19259 -9335
rect -19225 -9356 -19209 -9335
rect -19225 -9370 -19187 -9356
rect -19275 -9386 -19187 -9370
rect -18787 -9386 -18761 -9356
rect -18478 -9452 -18435 -9257
rect -18393 -9335 -18327 -9319
rect -18393 -9370 -18377 -9335
rect -18343 -9356 -18327 -9335
rect -18343 -9370 -18305 -9356
rect -18393 -9386 -18305 -9370
rect -17905 -9386 -17879 -9356
rect -17178 -9452 -17135 -9257
rect -17093 -9335 -17027 -9319
rect -17093 -9370 -17077 -9335
rect -17043 -9356 -17027 -9335
rect -17043 -9370 -17005 -9356
rect -17093 -9386 -17005 -9370
rect -16605 -9386 -16579 -9356
rect -16069 -9452 -16026 -9257
rect -15984 -9335 -15918 -9319
rect -15984 -9370 -15968 -9335
rect -15934 -9356 -15918 -9335
rect -15934 -9370 -15896 -9356
rect -15984 -9386 -15896 -9370
rect -15496 -9386 -15470 -9356
rect -15187 -9452 -15144 -9257
rect -15102 -9335 -15036 -9319
rect -15102 -9370 -15086 -9335
rect -15052 -9356 -15036 -9335
rect -15052 -9370 -15014 -9356
rect -15102 -9386 -15014 -9370
rect -14614 -9386 -14588 -9356
rect -13887 -9452 -13844 -9257
rect -13802 -9335 -13736 -9319
rect -13802 -9370 -13786 -9335
rect -13752 -9356 -13736 -9335
rect -13752 -9370 -13714 -9356
rect -13802 -9386 -13714 -9370
rect -13314 -9386 -13288 -9356
rect -12778 -9452 -12735 -9257
rect -12693 -9335 -12627 -9319
rect -12693 -9370 -12677 -9335
rect -12643 -9356 -12627 -9335
rect -12643 -9370 -12605 -9356
rect -12693 -9386 -12605 -9370
rect -12205 -9386 -12179 -9356
rect -11896 -9452 -11853 -9257
rect -11811 -9335 -11745 -9319
rect -11811 -9370 -11795 -9335
rect -11761 -9356 -11745 -9335
rect -11761 -9370 -11723 -9356
rect -11811 -9386 -11723 -9370
rect -11323 -9386 -11297 -9356
rect -10596 -9452 -10553 -9257
rect -10511 -9335 -10445 -9319
rect -10511 -9370 -10495 -9335
rect -10461 -9356 -10445 -9335
rect -10461 -9370 -10423 -9356
rect -10511 -9386 -10423 -9370
rect -10023 -9386 -9997 -9356
rect -9487 -9452 -9444 -9257
rect -9402 -9335 -9336 -9319
rect -9402 -9370 -9386 -9335
rect -9352 -9356 -9336 -9335
rect -9352 -9370 -9314 -9356
rect -9402 -9386 -9314 -9370
rect -8914 -9386 -8888 -9356
rect -8605 -9452 -8562 -9257
rect -8520 -9335 -8454 -9319
rect -8520 -9370 -8504 -9335
rect -8470 -9356 -8454 -9335
rect -8470 -9370 -8432 -9356
rect -8520 -9386 -8432 -9370
rect -8032 -9386 -8006 -9356
rect -20469 -9468 -20296 -9452
rect -20469 -9503 -20368 -9468
rect -20334 -9482 -20296 -9468
rect -19896 -9482 -19870 -9452
rect -19360 -9468 -19187 -9452
rect -20334 -9503 -20318 -9482
rect -20469 -9519 -20318 -9503
rect -19360 -9503 -19259 -9468
rect -19225 -9482 -19187 -9468
rect -18787 -9482 -18761 -9452
rect -18478 -9468 -18305 -9452
rect -19225 -9503 -19209 -9482
rect -19360 -9519 -19209 -9503
rect -18478 -9503 -18377 -9468
rect -18343 -9482 -18305 -9468
rect -17905 -9482 -17879 -9452
rect -17178 -9468 -17005 -9452
rect -18343 -9503 -18327 -9482
rect -18478 -9519 -18327 -9503
rect -17178 -9503 -17077 -9468
rect -17043 -9482 -17005 -9468
rect -16605 -9482 -16579 -9452
rect -16069 -9468 -15896 -9452
rect -17043 -9503 -17027 -9482
rect -17178 -9519 -17027 -9503
rect -16069 -9503 -15968 -9468
rect -15934 -9482 -15896 -9468
rect -15496 -9482 -15470 -9452
rect -15187 -9468 -15014 -9452
rect -15934 -9503 -15918 -9482
rect -16069 -9519 -15918 -9503
rect -15187 -9503 -15086 -9468
rect -15052 -9482 -15014 -9468
rect -14614 -9482 -14588 -9452
rect -13887 -9468 -13714 -9452
rect -15052 -9503 -15036 -9482
rect -15187 -9519 -15036 -9503
rect -13887 -9503 -13786 -9468
rect -13752 -9482 -13714 -9468
rect -13314 -9482 -13288 -9452
rect -12778 -9468 -12605 -9452
rect -13752 -9503 -13736 -9482
rect -13887 -9519 -13736 -9503
rect -12778 -9503 -12677 -9468
rect -12643 -9482 -12605 -9468
rect -12205 -9482 -12179 -9452
rect -11896 -9468 -11723 -9452
rect -12643 -9503 -12627 -9482
rect -12778 -9519 -12627 -9503
rect -11896 -9503 -11795 -9468
rect -11761 -9482 -11723 -9468
rect -11323 -9482 -11297 -9452
rect -10596 -9468 -10423 -9452
rect -11761 -9503 -11745 -9482
rect -11896 -9519 -11745 -9503
rect -10596 -9503 -10495 -9468
rect -10461 -9482 -10423 -9468
rect -10023 -9482 -9997 -9452
rect -9487 -9468 -9314 -9452
rect -10461 -9503 -10445 -9482
rect -10596 -9519 -10445 -9503
rect -9487 -9503 -9386 -9468
rect -9352 -9482 -9314 -9468
rect -8914 -9482 -8888 -9452
rect -8605 -9468 -8432 -9452
rect -9352 -9503 -9336 -9482
rect -9487 -9519 -9336 -9503
rect -8605 -9503 -8504 -9468
rect -8470 -9482 -8432 -9468
rect -8032 -9482 -8006 -9452
rect -8470 -9503 -8454 -9482
rect -8605 -9519 -8454 -9503
rect 5561 -9721 5627 -9705
rect 5561 -9947 5577 -9721
rect 5611 -9723 5627 -9721
rect 6001 -9721 6067 -9705
rect 5611 -9753 5658 -9723
rect 5872 -9753 5898 -9723
rect 5611 -9819 5627 -9753
rect 5611 -9849 5658 -9819
rect 5872 -9849 5898 -9819
rect 5611 -9915 5627 -9849
rect 5611 -9945 5658 -9915
rect 5872 -9945 5898 -9915
rect 5611 -9947 5627 -9945
rect 5561 -9963 5627 -9947
rect 6001 -9947 6017 -9721
rect 6051 -9723 6067 -9721
rect 6441 -9721 6507 -9705
rect 6051 -9753 6098 -9723
rect 6312 -9753 6338 -9723
rect 6051 -9819 6067 -9753
rect 6051 -9849 6098 -9819
rect 6312 -9849 6338 -9819
rect 6051 -9915 6067 -9849
rect 6051 -9945 6098 -9915
rect 6312 -9945 6338 -9915
rect 6051 -9947 6067 -9945
rect 6001 -9963 6067 -9947
rect 6441 -9947 6457 -9721
rect 6491 -9723 6507 -9721
rect 6491 -9753 6538 -9723
rect 6752 -9753 6778 -9723
rect 6491 -9819 6507 -9753
rect 6491 -9849 6538 -9819
rect 6752 -9849 6778 -9819
rect 6491 -9915 6507 -9849
rect 6491 -9945 6538 -9915
rect 6752 -9945 6778 -9915
rect 6491 -9947 6507 -9945
rect 6441 -9963 6507 -9947
rect 5561 -10167 5628 -10151
rect 5561 -10201 5577 -10167
rect 5611 -10169 5628 -10167
rect 6001 -10167 6068 -10151
rect 5611 -10199 5658 -10169
rect 5858 -10199 5884 -10169
rect 5611 -10201 5628 -10199
rect 5561 -10217 5628 -10201
rect 6001 -10201 6017 -10167
rect 6051 -10169 6068 -10167
rect 6441 -10167 6508 -10151
rect 6051 -10199 6098 -10169
rect 6298 -10199 6324 -10169
rect 6051 -10201 6068 -10199
rect 6001 -10217 6068 -10201
rect 6441 -10201 6457 -10167
rect 6491 -10169 6508 -10167
rect 6491 -10199 6538 -10169
rect 6738 -10199 6764 -10169
rect 6491 -10201 6508 -10199
rect 6441 -10217 6508 -10201
rect 7200 -10365 7230 -10339
rect 7296 -10365 7326 -10339
rect 7392 -10365 7422 -10339
rect 7488 -10365 7518 -10339
rect 7584 -10365 7614 -10339
rect 7680 -10365 7710 -10339
rect 7776 -10365 7806 -10339
rect 7872 -10365 7902 -10339
rect 8148 -10365 8178 -10339
rect 8244 -10365 8274 -10339
rect 8340 -10365 8370 -10339
rect 8436 -10365 8466 -10339
rect 8532 -10365 8562 -10339
rect 8628 -10365 8658 -10339
rect 8724 -10365 8754 -10339
rect 8820 -10365 8850 -10339
rect 9084 -10365 9114 -10339
rect 9180 -10365 9210 -10339
rect 9276 -10365 9306 -10339
rect 9372 -10365 9402 -10339
rect 9468 -10365 9498 -10339
rect 9564 -10365 9594 -10339
rect 9660 -10365 9690 -10339
rect 9756 -10365 9786 -10339
rect 10015 -10365 10045 -10339
rect 10111 -10365 10141 -10339
rect 10207 -10365 10237 -10339
rect 10303 -10365 10333 -10339
rect 10399 -10365 10429 -10339
rect 10495 -10365 10525 -10339
rect 10591 -10365 10621 -10339
rect 10687 -10365 10717 -10339
rect 10942 -10365 10972 -10339
rect 11038 -10365 11068 -10339
rect 11134 -10365 11164 -10339
rect 11230 -10365 11260 -10339
rect 11326 -10365 11356 -10339
rect 11422 -10365 11452 -10339
rect 11518 -10365 11548 -10339
rect 11614 -10365 11644 -10339
rect -20679 -10513 -20649 -10487
rect -20587 -10513 -20557 -10482
rect -20491 -10513 -20461 -10482
rect -20395 -10513 -20365 -10482
rect -20299 -10513 -20269 -10482
rect -20203 -10513 -20173 -10482
rect -20107 -10513 -20077 -10482
rect -20011 -10513 -19981 -10482
rect -19915 -10513 -19885 -10482
rect -19819 -10513 -19789 -10482
rect -19723 -10513 -19693 -10482
rect -19627 -10513 -19597 -10482
rect -19531 -10513 -19501 -10482
rect -19439 -10513 -19409 -10487
rect -19120 -10513 -19090 -10487
rect -19028 -10513 -18998 -10482
rect -18932 -10513 -18902 -10482
rect -18836 -10513 -18806 -10482
rect -18740 -10513 -18710 -10482
rect -18644 -10513 -18614 -10482
rect -18548 -10513 -18518 -10482
rect -18452 -10513 -18422 -10482
rect -18356 -10513 -18326 -10482
rect -18260 -10513 -18230 -10482
rect -18164 -10513 -18134 -10482
rect -18068 -10513 -18038 -10482
rect -17972 -10513 -17942 -10482
rect -17880 -10513 -17850 -10487
rect -17388 -10513 -17358 -10487
rect -17296 -10513 -17266 -10482
rect -17200 -10513 -17170 -10482
rect -17104 -10513 -17074 -10482
rect -17008 -10513 -16978 -10482
rect -16912 -10513 -16882 -10482
rect -16816 -10513 -16786 -10482
rect -16720 -10513 -16690 -10482
rect -16624 -10513 -16594 -10482
rect -16528 -10513 -16498 -10482
rect -16432 -10513 -16402 -10482
rect -16336 -10513 -16306 -10482
rect -16240 -10513 -16210 -10482
rect -16148 -10513 -16118 -10487
rect -15829 -10513 -15799 -10487
rect -15737 -10513 -15707 -10482
rect -15641 -10513 -15611 -10482
rect -15545 -10513 -15515 -10482
rect -15449 -10513 -15419 -10482
rect -15353 -10513 -15323 -10482
rect -15257 -10513 -15227 -10482
rect -15161 -10513 -15131 -10482
rect -15065 -10513 -15035 -10482
rect -14969 -10513 -14939 -10482
rect -14873 -10513 -14843 -10482
rect -14777 -10513 -14747 -10482
rect -14681 -10513 -14651 -10482
rect -14589 -10513 -14559 -10487
rect -14097 -10513 -14067 -10487
rect -14005 -10513 -13975 -10482
rect -13909 -10513 -13879 -10482
rect -13813 -10513 -13783 -10482
rect -13717 -10513 -13687 -10482
rect -13621 -10513 -13591 -10482
rect -13525 -10513 -13495 -10482
rect -13429 -10513 -13399 -10482
rect -13333 -10513 -13303 -10482
rect -13237 -10513 -13207 -10482
rect -13141 -10513 -13111 -10482
rect -13045 -10513 -13015 -10482
rect -12949 -10513 -12919 -10482
rect -12857 -10513 -12827 -10487
rect -12538 -10513 -12508 -10487
rect -12446 -10513 -12416 -10482
rect -12350 -10513 -12320 -10482
rect -12254 -10513 -12224 -10482
rect -12158 -10513 -12128 -10482
rect -12062 -10513 -12032 -10482
rect -11966 -10513 -11936 -10482
rect -11870 -10513 -11840 -10482
rect -11774 -10513 -11744 -10482
rect -11678 -10513 -11648 -10482
rect -11582 -10513 -11552 -10482
rect -11486 -10513 -11456 -10482
rect -11390 -10513 -11360 -10482
rect -11298 -10513 -11268 -10487
rect -10806 -10513 -10776 -10487
rect -10714 -10513 -10684 -10482
rect -10618 -10513 -10588 -10482
rect -10522 -10513 -10492 -10482
rect -10426 -10513 -10396 -10482
rect -10330 -10513 -10300 -10482
rect -10234 -10513 -10204 -10482
rect -10138 -10513 -10108 -10482
rect -10042 -10513 -10012 -10482
rect -9946 -10513 -9916 -10482
rect -9850 -10513 -9820 -10482
rect -9754 -10513 -9724 -10482
rect -9658 -10513 -9628 -10482
rect -9566 -10513 -9536 -10487
rect -9247 -10513 -9217 -10487
rect -9155 -10513 -9125 -10482
rect -9059 -10513 -9029 -10482
rect -8963 -10513 -8933 -10482
rect -8867 -10513 -8837 -10482
rect -8771 -10513 -8741 -10482
rect -8675 -10513 -8645 -10482
rect -8579 -10513 -8549 -10482
rect -8483 -10513 -8453 -10482
rect -8387 -10513 -8357 -10482
rect -8291 -10513 -8261 -10482
rect -8195 -10513 -8165 -10482
rect -8099 -10513 -8069 -10482
rect -8007 -10513 -7977 -10487
rect -23680 -10708 -23614 -10692
rect -24334 -10754 -24304 -10723
rect -24238 -10754 -24208 -10723
rect -24142 -10754 -24112 -10723
rect -24046 -10754 -24016 -10723
rect -23950 -10754 -23920 -10723
rect -23854 -10754 -23824 -10723
rect -23680 -10934 -23664 -10708
rect -23630 -10710 -23614 -10708
rect -21947 -10708 -21881 -10692
rect -23630 -10740 -23583 -10710
rect -23369 -10740 -23343 -10710
rect -23630 -10806 -23614 -10740
rect -22597 -10754 -22567 -10723
rect -22501 -10754 -22471 -10723
rect -22405 -10754 -22375 -10723
rect -22309 -10754 -22279 -10723
rect -22213 -10754 -22183 -10723
rect -22117 -10754 -22087 -10723
rect -23630 -10836 -23583 -10806
rect -23369 -10836 -23343 -10806
rect -23630 -10902 -23614 -10836
rect -23630 -10932 -23583 -10902
rect -23369 -10932 -23343 -10902
rect -23630 -10934 -23614 -10932
rect -23680 -10950 -23614 -10934
rect -24334 -10994 -24304 -10968
rect -24238 -10994 -24208 -10968
rect -24142 -10994 -24112 -10968
rect -24335 -11015 -24112 -10994
rect -24335 -11050 -24318 -11015
rect -24284 -11024 -24112 -11015
rect -24046 -10994 -24016 -10968
rect -23950 -10994 -23920 -10968
rect -23854 -10994 -23824 -10968
rect -21947 -10934 -21931 -10708
rect -21897 -10710 -21881 -10708
rect -21897 -10740 -21850 -10710
rect -21636 -10740 -21610 -10710
rect -21897 -10806 -21881 -10740
rect -21897 -10836 -21850 -10806
rect -21636 -10836 -21610 -10806
rect -21897 -10902 -21881 -10836
rect -21897 -10932 -21850 -10902
rect -21636 -10932 -21610 -10902
rect -21897 -10934 -21881 -10932
rect -21947 -10950 -21881 -10934
rect -22597 -10994 -22567 -10968
rect -22501 -10994 -22471 -10968
rect -22405 -10994 -22375 -10968
rect -24046 -11015 -23824 -10994
rect -24284 -11050 -24268 -11024
rect -24335 -11061 -24268 -11050
rect -24046 -11050 -24029 -11015
rect -23995 -11024 -23824 -11015
rect -22598 -11015 -22375 -10994
rect -23995 -11050 -23979 -11024
rect -24046 -11061 -23979 -11050
rect -22598 -11050 -22581 -11015
rect -22547 -11024 -22375 -11015
rect -22309 -10994 -22279 -10968
rect -22213 -10994 -22183 -10968
rect -22117 -10994 -22087 -10968
rect -22309 -11015 -22087 -10994
rect -22547 -11050 -22531 -11024
rect -22598 -11061 -22531 -11050
rect -22309 -11050 -22292 -11015
rect -22258 -11024 -22087 -11015
rect -22258 -11050 -22242 -11024
rect -22309 -11061 -22242 -11050
rect -24335 -11256 -24292 -11061
rect -24250 -11139 -24184 -11123
rect -24250 -11174 -24234 -11139
rect -24200 -11160 -24184 -11139
rect -23680 -11154 -23613 -11138
rect -24200 -11174 -24162 -11160
rect -24250 -11190 -24162 -11174
rect -23762 -11190 -23736 -11160
rect -23680 -11188 -23664 -11154
rect -23630 -11156 -23613 -11154
rect -23630 -11186 -23583 -11156
rect -23383 -11186 -23357 -11156
rect -23630 -11188 -23613 -11186
rect -23680 -11204 -23613 -11188
rect -22598 -11256 -22555 -11061
rect 7200 -10718 7230 -10687
rect 7296 -10718 7326 -10687
rect 7392 -10718 7422 -10687
rect 7488 -10718 7518 -10687
rect 7584 -10718 7614 -10687
rect 7680 -10718 7710 -10687
rect 7776 -10718 7806 -10687
rect 7872 -10718 7902 -10687
rect 8148 -10718 8178 -10687
rect 8244 -10718 8274 -10687
rect 8340 -10718 8370 -10687
rect 8436 -10718 8466 -10687
rect 8532 -10718 8562 -10687
rect 8628 -10718 8658 -10687
rect 8724 -10718 8754 -10687
rect 8820 -10718 8850 -10687
rect 9084 -10718 9114 -10687
rect 9180 -10718 9210 -10687
rect 9276 -10718 9306 -10687
rect 9372 -10718 9402 -10687
rect 9468 -10718 9498 -10687
rect 9564 -10718 9594 -10687
rect 9660 -10718 9690 -10687
rect 9756 -10718 9786 -10687
rect 10015 -10718 10045 -10687
rect 10111 -10718 10141 -10687
rect 10207 -10718 10237 -10687
rect 10303 -10718 10333 -10687
rect 10399 -10718 10429 -10687
rect 10495 -10718 10525 -10687
rect 10591 -10718 10621 -10687
rect 10687 -10718 10717 -10687
rect 10942 -10718 10972 -10687
rect 11038 -10718 11068 -10687
rect 11134 -10718 11164 -10687
rect 11230 -10718 11260 -10687
rect 11326 -10718 11356 -10687
rect 11422 -10718 11452 -10687
rect 11518 -10718 11548 -10687
rect 11614 -10718 11644 -10687
rect 7182 -10734 7326 -10718
rect 7182 -10768 7198 -10734
rect 7232 -10768 7326 -10734
rect 7182 -10784 7326 -10768
rect 7374 -10734 7518 -10718
rect 7374 -10768 7390 -10734
rect 7424 -10768 7518 -10734
rect 7238 -11031 7268 -10784
rect 7374 -10851 7518 -10768
rect 7566 -10734 7710 -10718
rect 7566 -10768 7582 -10734
rect 7616 -10768 7710 -10734
rect 7566 -10784 7710 -10768
rect 7758 -10734 7902 -10718
rect 7758 -10768 7774 -10734
rect 7808 -10768 7902 -10734
rect 7758 -10784 7902 -10768
rect 8130 -10734 8274 -10718
rect 8130 -10768 8146 -10734
rect 8180 -10768 8274 -10734
rect 8130 -10784 8274 -10768
rect 8322 -10734 8466 -10718
rect 8322 -10768 8338 -10734
rect 8372 -10768 8466 -10734
rect 7584 -10809 7644 -10784
rect 7374 -10989 7548 -10851
rect 7238 -11061 7452 -11031
rect -20679 -11094 -20649 -11063
rect -20587 -11094 -20557 -11063
rect -20491 -11094 -20461 -11063
rect -20395 -11094 -20365 -11063
rect -20299 -11093 -20269 -11063
rect -20203 -11093 -20173 -11063
rect -20107 -11093 -20077 -11063
rect -22513 -11139 -22447 -11123
rect -22513 -11174 -22497 -11139
rect -22463 -11160 -22447 -11139
rect -21947 -11154 -21880 -11138
rect -22463 -11174 -22425 -11160
rect -22513 -11190 -22425 -11174
rect -22025 -11190 -21999 -11160
rect -21947 -11188 -21931 -11154
rect -21897 -11156 -21880 -11154
rect -20873 -11151 -20363 -11094
rect -21897 -11186 -21850 -11156
rect -21650 -11186 -21624 -11156
rect -21897 -11188 -21880 -11186
rect -21947 -11204 -21880 -11188
rect -24335 -11272 -24162 -11256
rect -24335 -11307 -24234 -11272
rect -24200 -11286 -24162 -11272
rect -23762 -11286 -23736 -11256
rect -22598 -11272 -22425 -11256
rect -24200 -11307 -24184 -11286
rect -24335 -11323 -24184 -11307
rect -22598 -11307 -22497 -11272
rect -22463 -11286 -22425 -11272
rect -22025 -11286 -21999 -11256
rect -20873 -11261 -20854 -11151
rect -20807 -11244 -20363 -11151
rect -20299 -11122 -20077 -11093
rect -20299 -11167 -20269 -11122
rect -20139 -11167 -20077 -11122
rect -20299 -11186 -20077 -11167
rect -20011 -11094 -19981 -11063
rect -19915 -11094 -19885 -11063
rect -19819 -11094 -19789 -11063
rect -20011 -11127 -19789 -11094
rect -20011 -11172 -19938 -11127
rect -19808 -11172 -19789 -11127
rect -20011 -11187 -19789 -11172
rect -19723 -11094 -19693 -11063
rect -19627 -11094 -19597 -11063
rect -19531 -11094 -19501 -11063
rect -19439 -11094 -19409 -11063
rect -19120 -11094 -19090 -11063
rect -19028 -11094 -18998 -11063
rect -18932 -11094 -18902 -11063
rect -18836 -11094 -18806 -11063
rect -18740 -11093 -18710 -11063
rect -18644 -11093 -18614 -11063
rect -18548 -11093 -18518 -11063
rect -20807 -11261 -19789 -11244
rect -22463 -11307 -22447 -11286
rect -22598 -11323 -22447 -11307
rect -20873 -11353 -19789 -11261
rect -20712 -11528 -20636 -11353
rect -20587 -11443 -20365 -11418
rect -20587 -11488 -20544 -11443
rect -20414 -11488 -20365 -11443
rect -20679 -11553 -20649 -11528
rect -20587 -11531 -20365 -11488
rect -20587 -11553 -20557 -11531
rect -20491 -11553 -20461 -11531
rect -20395 -11553 -20365 -11531
rect -20299 -11451 -20077 -11423
rect -20299 -11496 -20261 -11451
rect -20131 -11496 -20077 -11451
rect -20299 -11531 -20077 -11496
rect -20299 -11553 -20269 -11531
rect -20203 -11553 -20173 -11531
rect -20107 -11553 -20077 -11531
rect -20011 -11531 -19789 -11353
rect -20011 -11553 -19981 -11531
rect -19915 -11553 -19885 -11531
rect -19819 -11553 -19789 -11531
rect -19723 -11251 -19409 -11094
rect -19153 -11181 -18804 -11094
rect -19723 -11306 -19691 -11251
rect -19626 -11306 -19409 -11251
rect -19723 -11531 -19409 -11306
rect -19342 -11196 -18804 -11181
rect -18740 -11122 -18518 -11093
rect -18740 -11167 -18710 -11122
rect -18580 -11167 -18518 -11122
rect -18740 -11186 -18518 -11167
rect -18452 -11094 -18422 -11063
rect -18356 -11094 -18326 -11063
rect -18260 -11094 -18230 -11063
rect -18452 -11127 -18230 -11094
rect -18452 -11172 -18379 -11127
rect -18249 -11172 -18230 -11127
rect -18452 -11187 -18230 -11172
rect -18164 -11094 -18134 -11063
rect -18068 -11094 -18038 -11063
rect -17972 -11094 -17942 -11063
rect -17880 -11094 -17850 -11063
rect -17388 -11094 -17358 -11063
rect -17296 -11094 -17266 -11063
rect -17200 -11094 -17170 -11063
rect -17104 -11094 -17074 -11063
rect -17008 -11093 -16978 -11063
rect -16912 -11093 -16882 -11063
rect -16816 -11093 -16786 -11063
rect -19342 -11336 -19297 -11196
rect -19224 -11244 -18804 -11196
rect -19224 -11336 -18230 -11244
rect -19342 -11353 -18230 -11336
rect -19153 -11528 -19077 -11353
rect -19028 -11443 -18806 -11418
rect -19028 -11488 -18985 -11443
rect -18855 -11488 -18806 -11443
rect -19723 -11553 -19693 -11531
rect -19627 -11553 -19597 -11531
rect -19531 -11553 -19501 -11531
rect -19439 -11553 -19409 -11531
rect -19120 -11553 -19090 -11528
rect -19028 -11531 -18806 -11488
rect -19028 -11553 -18998 -11531
rect -18932 -11553 -18902 -11531
rect -18836 -11553 -18806 -11531
rect -18740 -11451 -18518 -11423
rect -18740 -11496 -18702 -11451
rect -18572 -11496 -18518 -11451
rect -18740 -11531 -18518 -11496
rect -18740 -11553 -18710 -11531
rect -18644 -11553 -18614 -11531
rect -18548 -11553 -18518 -11531
rect -18452 -11531 -18230 -11353
rect -18452 -11553 -18422 -11531
rect -18356 -11553 -18326 -11531
rect -18260 -11553 -18230 -11531
rect -18164 -11251 -17850 -11094
rect -18164 -11306 -18132 -11251
rect -18067 -11306 -17850 -11251
rect -18164 -11531 -17850 -11306
rect -17582 -11151 -17072 -11094
rect -17582 -11261 -17563 -11151
rect -17516 -11244 -17072 -11151
rect -17008 -11122 -16786 -11093
rect -17008 -11167 -16978 -11122
rect -16848 -11167 -16786 -11122
rect -17008 -11186 -16786 -11167
rect -16720 -11094 -16690 -11063
rect -16624 -11094 -16594 -11063
rect -16528 -11094 -16498 -11063
rect -16720 -11127 -16498 -11094
rect -16720 -11172 -16647 -11127
rect -16517 -11172 -16498 -11127
rect -16720 -11187 -16498 -11172
rect -16432 -11094 -16402 -11063
rect -16336 -11094 -16306 -11063
rect -16240 -11094 -16210 -11063
rect -16148 -11094 -16118 -11063
rect -15829 -11094 -15799 -11063
rect -15737 -11094 -15707 -11063
rect -15641 -11094 -15611 -11063
rect -15545 -11094 -15515 -11063
rect -15449 -11093 -15419 -11063
rect -15353 -11093 -15323 -11063
rect -15257 -11093 -15227 -11063
rect -17516 -11261 -16498 -11244
rect -17582 -11353 -16498 -11261
rect -17421 -11528 -17345 -11353
rect -17296 -11443 -17074 -11418
rect -17296 -11488 -17253 -11443
rect -17123 -11488 -17074 -11443
rect -18164 -11553 -18134 -11531
rect -18068 -11553 -18038 -11531
rect -17972 -11553 -17942 -11531
rect -17880 -11553 -17850 -11531
rect -17388 -11553 -17358 -11528
rect -17296 -11531 -17074 -11488
rect -17296 -11553 -17266 -11531
rect -17200 -11553 -17170 -11531
rect -17104 -11553 -17074 -11531
rect -17008 -11451 -16786 -11423
rect -17008 -11496 -16970 -11451
rect -16840 -11496 -16786 -11451
rect -17008 -11531 -16786 -11496
rect -17008 -11553 -16978 -11531
rect -16912 -11553 -16882 -11531
rect -16816 -11553 -16786 -11531
rect -16720 -11531 -16498 -11353
rect -16720 -11553 -16690 -11531
rect -16624 -11553 -16594 -11531
rect -16528 -11553 -16498 -11531
rect -16432 -11251 -16118 -11094
rect -15862 -11181 -15513 -11094
rect -16432 -11306 -16400 -11251
rect -16335 -11306 -16118 -11251
rect -16432 -11531 -16118 -11306
rect -16051 -11196 -15513 -11181
rect -15449 -11122 -15227 -11093
rect -15449 -11167 -15419 -11122
rect -15289 -11167 -15227 -11122
rect -15449 -11186 -15227 -11167
rect -15161 -11094 -15131 -11063
rect -15065 -11094 -15035 -11063
rect -14969 -11094 -14939 -11063
rect -15161 -11127 -14939 -11094
rect -15161 -11172 -15088 -11127
rect -14958 -11172 -14939 -11127
rect -15161 -11187 -14939 -11172
rect -14873 -11094 -14843 -11063
rect -14777 -11094 -14747 -11063
rect -14681 -11094 -14651 -11063
rect -14589 -11094 -14559 -11063
rect -14097 -11094 -14067 -11063
rect -14005 -11094 -13975 -11063
rect -13909 -11094 -13879 -11063
rect -13813 -11094 -13783 -11063
rect -13717 -11093 -13687 -11063
rect -13621 -11093 -13591 -11063
rect -13525 -11093 -13495 -11063
rect -16051 -11336 -16006 -11196
rect -15933 -11244 -15513 -11196
rect -15933 -11336 -14939 -11244
rect -16051 -11353 -14939 -11336
rect -15862 -11528 -15786 -11353
rect -15737 -11443 -15515 -11418
rect -15737 -11488 -15694 -11443
rect -15564 -11488 -15515 -11443
rect -16432 -11553 -16402 -11531
rect -16336 -11553 -16306 -11531
rect -16240 -11553 -16210 -11531
rect -16148 -11553 -16118 -11531
rect -15829 -11553 -15799 -11528
rect -15737 -11531 -15515 -11488
rect -15737 -11553 -15707 -11531
rect -15641 -11553 -15611 -11531
rect -15545 -11553 -15515 -11531
rect -15449 -11451 -15227 -11423
rect -15449 -11496 -15411 -11451
rect -15281 -11496 -15227 -11451
rect -15449 -11531 -15227 -11496
rect -15449 -11553 -15419 -11531
rect -15353 -11553 -15323 -11531
rect -15257 -11553 -15227 -11531
rect -15161 -11531 -14939 -11353
rect -15161 -11553 -15131 -11531
rect -15065 -11553 -15035 -11531
rect -14969 -11553 -14939 -11531
rect -14873 -11251 -14559 -11094
rect -14873 -11306 -14841 -11251
rect -14776 -11306 -14559 -11251
rect -14873 -11531 -14559 -11306
rect -14291 -11151 -13781 -11094
rect -14291 -11261 -14272 -11151
rect -14225 -11244 -13781 -11151
rect -13717 -11122 -13495 -11093
rect -13717 -11167 -13687 -11122
rect -13557 -11167 -13495 -11122
rect -13717 -11186 -13495 -11167
rect -13429 -11094 -13399 -11063
rect -13333 -11094 -13303 -11063
rect -13237 -11094 -13207 -11063
rect -13429 -11127 -13207 -11094
rect -13429 -11172 -13356 -11127
rect -13226 -11172 -13207 -11127
rect -13429 -11187 -13207 -11172
rect -13141 -11094 -13111 -11063
rect -13045 -11094 -13015 -11063
rect -12949 -11094 -12919 -11063
rect -12857 -11094 -12827 -11063
rect -12538 -11094 -12508 -11063
rect -12446 -11094 -12416 -11063
rect -12350 -11094 -12320 -11063
rect -12254 -11094 -12224 -11063
rect -12158 -11093 -12128 -11063
rect -12062 -11093 -12032 -11063
rect -11966 -11093 -11936 -11063
rect -14225 -11261 -13207 -11244
rect -14291 -11353 -13207 -11261
rect -14130 -11528 -14054 -11353
rect -14005 -11443 -13783 -11418
rect -14005 -11488 -13962 -11443
rect -13832 -11488 -13783 -11443
rect -14873 -11553 -14843 -11531
rect -14777 -11553 -14747 -11531
rect -14681 -11553 -14651 -11531
rect -14589 -11553 -14559 -11531
rect -14097 -11553 -14067 -11528
rect -14005 -11531 -13783 -11488
rect -14005 -11553 -13975 -11531
rect -13909 -11553 -13879 -11531
rect -13813 -11553 -13783 -11531
rect -13717 -11451 -13495 -11423
rect -13717 -11496 -13679 -11451
rect -13549 -11496 -13495 -11451
rect -13717 -11531 -13495 -11496
rect -13717 -11553 -13687 -11531
rect -13621 -11553 -13591 -11531
rect -13525 -11553 -13495 -11531
rect -13429 -11531 -13207 -11353
rect -13429 -11553 -13399 -11531
rect -13333 -11553 -13303 -11531
rect -13237 -11553 -13207 -11531
rect -13141 -11251 -12827 -11094
rect -12571 -11181 -12222 -11094
rect -13141 -11306 -13109 -11251
rect -13044 -11306 -12827 -11251
rect -13141 -11531 -12827 -11306
rect -12760 -11196 -12222 -11181
rect -12158 -11122 -11936 -11093
rect -12158 -11167 -12128 -11122
rect -11998 -11167 -11936 -11122
rect -12158 -11186 -11936 -11167
rect -11870 -11094 -11840 -11063
rect -11774 -11094 -11744 -11063
rect -11678 -11094 -11648 -11063
rect -11870 -11127 -11648 -11094
rect -11870 -11172 -11797 -11127
rect -11667 -11172 -11648 -11127
rect -11870 -11187 -11648 -11172
rect -11582 -11094 -11552 -11063
rect -11486 -11094 -11456 -11063
rect -11390 -11094 -11360 -11063
rect -11298 -11094 -11268 -11063
rect -10806 -11094 -10776 -11063
rect -10714 -11094 -10684 -11063
rect -10618 -11094 -10588 -11063
rect -10522 -11094 -10492 -11063
rect -10426 -11093 -10396 -11063
rect -10330 -11093 -10300 -11063
rect -10234 -11093 -10204 -11063
rect -12760 -11336 -12715 -11196
rect -12642 -11244 -12222 -11196
rect -12642 -11336 -11648 -11244
rect -12760 -11353 -11648 -11336
rect -12571 -11528 -12495 -11353
rect -12446 -11443 -12224 -11418
rect -12446 -11488 -12403 -11443
rect -12273 -11488 -12224 -11443
rect -13141 -11553 -13111 -11531
rect -13045 -11553 -13015 -11531
rect -12949 -11553 -12919 -11531
rect -12857 -11553 -12827 -11531
rect -12538 -11553 -12508 -11528
rect -12446 -11531 -12224 -11488
rect -12446 -11553 -12416 -11531
rect -12350 -11553 -12320 -11531
rect -12254 -11553 -12224 -11531
rect -12158 -11451 -11936 -11423
rect -12158 -11496 -12120 -11451
rect -11990 -11496 -11936 -11451
rect -12158 -11531 -11936 -11496
rect -12158 -11553 -12128 -11531
rect -12062 -11553 -12032 -11531
rect -11966 -11553 -11936 -11531
rect -11870 -11531 -11648 -11353
rect -11870 -11553 -11840 -11531
rect -11774 -11553 -11744 -11531
rect -11678 -11553 -11648 -11531
rect -11582 -11251 -11268 -11094
rect -11582 -11306 -11550 -11251
rect -11485 -11306 -11268 -11251
rect -11582 -11531 -11268 -11306
rect -11000 -11151 -10490 -11094
rect -11000 -11261 -10981 -11151
rect -10934 -11244 -10490 -11151
rect -10426 -11122 -10204 -11093
rect -10426 -11167 -10396 -11122
rect -10266 -11167 -10204 -11122
rect -10426 -11186 -10204 -11167
rect -10138 -11094 -10108 -11063
rect -10042 -11094 -10012 -11063
rect -9946 -11094 -9916 -11063
rect -10138 -11127 -9916 -11094
rect -10138 -11172 -10065 -11127
rect -9935 -11172 -9916 -11127
rect -10138 -11187 -9916 -11172
rect -9850 -11094 -9820 -11063
rect -9754 -11094 -9724 -11063
rect -9658 -11094 -9628 -11063
rect -9566 -11094 -9536 -11063
rect -9247 -11094 -9217 -11063
rect -9155 -11094 -9125 -11063
rect -9059 -11094 -9029 -11063
rect -8963 -11094 -8933 -11063
rect -8867 -11093 -8837 -11063
rect -8771 -11093 -8741 -11063
rect -8675 -11093 -8645 -11063
rect -10934 -11261 -9916 -11244
rect -11000 -11353 -9916 -11261
rect -10839 -11528 -10763 -11353
rect -10714 -11443 -10492 -11418
rect -10714 -11488 -10671 -11443
rect -10541 -11488 -10492 -11443
rect -11582 -11553 -11552 -11531
rect -11486 -11553 -11456 -11531
rect -11390 -11553 -11360 -11531
rect -11298 -11553 -11268 -11531
rect -10806 -11553 -10776 -11528
rect -10714 -11531 -10492 -11488
rect -10714 -11553 -10684 -11531
rect -10618 -11553 -10588 -11531
rect -10522 -11553 -10492 -11531
rect -10426 -11451 -10204 -11423
rect -10426 -11496 -10388 -11451
rect -10258 -11496 -10204 -11451
rect -10426 -11531 -10204 -11496
rect -10426 -11553 -10396 -11531
rect -10330 -11553 -10300 -11531
rect -10234 -11553 -10204 -11531
rect -10138 -11531 -9916 -11353
rect -10138 -11553 -10108 -11531
rect -10042 -11553 -10012 -11531
rect -9946 -11553 -9916 -11531
rect -9850 -11251 -9536 -11094
rect -9280 -11181 -8931 -11094
rect -9850 -11306 -9818 -11251
rect -9753 -11306 -9536 -11251
rect -9850 -11531 -9536 -11306
rect -9469 -11196 -8931 -11181
rect -8867 -11122 -8645 -11093
rect -8867 -11167 -8837 -11122
rect -8707 -11167 -8645 -11122
rect -8867 -11186 -8645 -11167
rect -8579 -11094 -8549 -11063
rect -8483 -11094 -8453 -11063
rect -8387 -11094 -8357 -11063
rect -8579 -11127 -8357 -11094
rect -8579 -11172 -8506 -11127
rect -8376 -11172 -8357 -11127
rect -8579 -11187 -8357 -11172
rect -8291 -11094 -8261 -11063
rect -8195 -11094 -8165 -11063
rect -8099 -11094 -8069 -11063
rect -8007 -11094 -7977 -11063
rect 7422 -11094 7452 -11061
rect 7518 -11094 7548 -10989
rect 7590 -11071 7644 -10809
rect 7758 -10914 7848 -10784
rect 7614 -11094 7644 -11071
rect 7710 -10944 7848 -10914
rect 7710 -11094 7740 -10944
rect 8186 -11031 8216 -10784
rect 8322 -10851 8466 -10768
rect 8514 -10734 8658 -10718
rect 8514 -10768 8530 -10734
rect 8564 -10768 8658 -10734
rect 8514 -10784 8658 -10768
rect 8706 -10734 8850 -10718
rect 8706 -10768 8722 -10734
rect 8756 -10768 8850 -10734
rect 8706 -10784 8850 -10768
rect 9066 -10734 9210 -10718
rect 9066 -10768 9082 -10734
rect 9116 -10768 9210 -10734
rect 9066 -10784 9210 -10768
rect 9258 -10734 9402 -10718
rect 9258 -10768 9274 -10734
rect 9308 -10768 9402 -10734
rect 8532 -10809 8592 -10784
rect 8322 -10989 8496 -10851
rect 8186 -11061 8400 -11031
rect 8370 -11094 8400 -11061
rect 8466 -11094 8496 -10989
rect 8538 -11071 8592 -10809
rect 8706 -10914 8796 -10784
rect 8562 -11094 8592 -11071
rect 8658 -10944 8796 -10914
rect 8658 -11094 8688 -10944
rect 9122 -11031 9152 -10784
rect 9258 -10851 9402 -10768
rect 9450 -10734 9594 -10718
rect 9450 -10768 9466 -10734
rect 9500 -10768 9594 -10734
rect 9450 -10784 9594 -10768
rect 9642 -10734 9786 -10718
rect 9642 -10768 9658 -10734
rect 9692 -10768 9786 -10734
rect 9642 -10784 9786 -10768
rect 9997 -10734 10141 -10718
rect 9997 -10768 10013 -10734
rect 10047 -10768 10141 -10734
rect 9997 -10784 10141 -10768
rect 10189 -10734 10333 -10718
rect 10189 -10768 10205 -10734
rect 10239 -10768 10333 -10734
rect 9468 -10809 9528 -10784
rect 9258 -10989 9432 -10851
rect 9122 -11061 9336 -11031
rect 9306 -11094 9336 -11061
rect 9402 -11094 9432 -10989
rect 9474 -11071 9528 -10809
rect 9642 -10914 9732 -10784
rect 9498 -11094 9528 -11071
rect 9594 -10944 9732 -10914
rect 9594 -11094 9624 -10944
rect 10053 -11031 10083 -10784
rect 10189 -10851 10333 -10768
rect 10381 -10734 10525 -10718
rect 10381 -10768 10397 -10734
rect 10431 -10768 10525 -10734
rect 10381 -10784 10525 -10768
rect 10573 -10734 10717 -10718
rect 10573 -10768 10589 -10734
rect 10623 -10768 10717 -10734
rect 10573 -10784 10717 -10768
rect 10924 -10734 11068 -10718
rect 10924 -10768 10940 -10734
rect 10974 -10768 11068 -10734
rect 10924 -10784 11068 -10768
rect 11116 -10734 11260 -10718
rect 11116 -10768 11132 -10734
rect 11166 -10768 11260 -10734
rect 10399 -10809 10459 -10784
rect 10189 -10989 10363 -10851
rect 10053 -11061 10267 -11031
rect 10237 -11094 10267 -11061
rect 10333 -11094 10363 -10989
rect 10405 -11071 10459 -10809
rect 10573 -10914 10663 -10784
rect 10429 -11094 10459 -11071
rect 10525 -10944 10663 -10914
rect 10525 -11094 10555 -10944
rect 10980 -11031 11010 -10784
rect 11116 -10851 11260 -10768
rect 11308 -10734 11452 -10718
rect 11308 -10768 11324 -10734
rect 11358 -10768 11452 -10734
rect 11308 -10784 11452 -10768
rect 11500 -10734 11644 -10718
rect 11500 -10768 11516 -10734
rect 11550 -10768 11644 -10734
rect 11500 -10784 11644 -10768
rect 11326 -10809 11386 -10784
rect 11116 -10989 11290 -10851
rect 10980 -11061 11194 -11031
rect 11164 -11094 11194 -11061
rect 11260 -11094 11290 -10989
rect 11332 -11071 11386 -10809
rect 11500 -10914 11590 -10784
rect 11356 -11094 11386 -11071
rect 11452 -10944 11590 -10914
rect 11452 -11094 11482 -10944
rect -9469 -11336 -9424 -11196
rect -9351 -11244 -8931 -11196
rect -9351 -11336 -8357 -11244
rect -9469 -11353 -8357 -11336
rect -9280 -11528 -9204 -11353
rect -9155 -11443 -8933 -11418
rect -9155 -11488 -9112 -11443
rect -8982 -11488 -8933 -11443
rect -9850 -11553 -9820 -11531
rect -9754 -11553 -9724 -11531
rect -9658 -11553 -9628 -11531
rect -9566 -11553 -9536 -11531
rect -9247 -11553 -9217 -11528
rect -9155 -11531 -8933 -11488
rect -9155 -11553 -9125 -11531
rect -9059 -11553 -9029 -11531
rect -8963 -11553 -8933 -11531
rect -8867 -11451 -8645 -11423
rect -8867 -11496 -8829 -11451
rect -8699 -11496 -8645 -11451
rect -8867 -11531 -8645 -11496
rect -8867 -11553 -8837 -11531
rect -8771 -11553 -8741 -11531
rect -8675 -11553 -8645 -11531
rect -8579 -11531 -8357 -11353
rect -8579 -11553 -8549 -11531
rect -8483 -11553 -8453 -11531
rect -8387 -11553 -8357 -11531
rect -8291 -11251 -7977 -11094
rect -8291 -11306 -8259 -11251
rect -8194 -11306 -7977 -11251
rect -8291 -11531 -7977 -11306
rect -8291 -11553 -8261 -11531
rect -8195 -11553 -8165 -11531
rect -8099 -11553 -8069 -11531
rect -8007 -11553 -7977 -11531
rect -20679 -11709 -20649 -11683
rect -20587 -11709 -20557 -11683
rect -20491 -11709 -20461 -11683
rect -20395 -11709 -20365 -11683
rect -20299 -11709 -20269 -11683
rect -20203 -11709 -20173 -11683
rect -20107 -11709 -20077 -11683
rect -20011 -11709 -19981 -11683
rect -19915 -11709 -19885 -11683
rect -19819 -11709 -19789 -11683
rect -19723 -11709 -19693 -11683
rect -19627 -11709 -19597 -11683
rect -19531 -11709 -19501 -11683
rect -19439 -11709 -19409 -11683
rect -19120 -11709 -19090 -11683
rect -19028 -11709 -18998 -11683
rect -18932 -11709 -18902 -11683
rect -18836 -11709 -18806 -11683
rect -18740 -11709 -18710 -11683
rect -18644 -11709 -18614 -11683
rect -18548 -11709 -18518 -11683
rect -18452 -11709 -18422 -11683
rect -18356 -11709 -18326 -11683
rect -18260 -11709 -18230 -11683
rect -18164 -11709 -18134 -11683
rect -18068 -11709 -18038 -11683
rect -17972 -11709 -17942 -11683
rect -17880 -11709 -17850 -11683
rect -17388 -11709 -17358 -11683
rect -17296 -11709 -17266 -11683
rect -17200 -11709 -17170 -11683
rect -17104 -11709 -17074 -11683
rect -17008 -11709 -16978 -11683
rect -16912 -11709 -16882 -11683
rect -16816 -11709 -16786 -11683
rect -16720 -11709 -16690 -11683
rect -16624 -11709 -16594 -11683
rect -16528 -11709 -16498 -11683
rect -16432 -11709 -16402 -11683
rect -16336 -11709 -16306 -11683
rect -16240 -11709 -16210 -11683
rect -16148 -11709 -16118 -11683
rect -15829 -11709 -15799 -11683
rect -15737 -11709 -15707 -11683
rect -15641 -11709 -15611 -11683
rect -15545 -11709 -15515 -11683
rect -15449 -11709 -15419 -11683
rect -15353 -11709 -15323 -11683
rect -15257 -11709 -15227 -11683
rect -15161 -11709 -15131 -11683
rect -15065 -11709 -15035 -11683
rect -14969 -11709 -14939 -11683
rect -14873 -11709 -14843 -11683
rect -14777 -11709 -14747 -11683
rect -14681 -11709 -14651 -11683
rect -14589 -11709 -14559 -11683
rect -14097 -11709 -14067 -11683
rect -14005 -11709 -13975 -11683
rect -13909 -11709 -13879 -11683
rect -13813 -11709 -13783 -11683
rect -13717 -11709 -13687 -11683
rect -13621 -11709 -13591 -11683
rect -13525 -11709 -13495 -11683
rect -13429 -11709 -13399 -11683
rect -13333 -11709 -13303 -11683
rect -13237 -11709 -13207 -11683
rect -13141 -11709 -13111 -11683
rect -13045 -11709 -13015 -11683
rect -12949 -11709 -12919 -11683
rect -12857 -11709 -12827 -11683
rect -12538 -11709 -12508 -11683
rect -12446 -11709 -12416 -11683
rect -12350 -11709 -12320 -11683
rect -12254 -11709 -12224 -11683
rect -12158 -11709 -12128 -11683
rect -12062 -11709 -12032 -11683
rect -11966 -11709 -11936 -11683
rect -11870 -11709 -11840 -11683
rect -11774 -11709 -11744 -11683
rect -11678 -11709 -11648 -11683
rect -11582 -11709 -11552 -11683
rect -11486 -11709 -11456 -11683
rect -11390 -11709 -11360 -11683
rect -11298 -11709 -11268 -11683
rect -10806 -11709 -10776 -11683
rect -10714 -11709 -10684 -11683
rect -10618 -11709 -10588 -11683
rect -10522 -11709 -10492 -11683
rect -10426 -11709 -10396 -11683
rect -10330 -11709 -10300 -11683
rect -10234 -11709 -10204 -11683
rect -10138 -11709 -10108 -11683
rect -10042 -11709 -10012 -11683
rect -9946 -11709 -9916 -11683
rect -9850 -11709 -9820 -11683
rect -9754 -11709 -9724 -11683
rect -9658 -11709 -9628 -11683
rect -9566 -11709 -9536 -11683
rect -9247 -11709 -9217 -11683
rect -9155 -11709 -9125 -11683
rect -9059 -11709 -9029 -11683
rect -8963 -11709 -8933 -11683
rect -8867 -11709 -8837 -11683
rect -8771 -11709 -8741 -11683
rect -8675 -11709 -8645 -11683
rect -8579 -11709 -8549 -11683
rect -8483 -11709 -8453 -11683
rect -8387 -11709 -8357 -11683
rect -8291 -11709 -8261 -11683
rect -8195 -11709 -8165 -11683
rect -8099 -11709 -8069 -11683
rect -8007 -11709 -7977 -11683
rect 11835 -11575 11865 -11549
rect 11931 -11575 11961 -11549
rect 12027 -11575 12057 -11549
rect 12123 -11575 12153 -11549
rect 12219 -11575 12249 -11549
rect 12315 -11575 12345 -11549
rect 12411 -11575 12441 -11549
rect 12507 -11575 12537 -11549
rect 12603 -11575 12633 -11549
rect 12699 -11575 12729 -11549
rect 12826 -11739 12892 -11723
rect 11835 -11857 11865 -11831
rect 11931 -11857 11961 -11831
rect 12027 -11857 12057 -11831
rect 12123 -11857 12153 -11831
rect 12219 -11857 12249 -11831
rect 11835 -11881 12249 -11857
rect -23680 -12000 -23614 -11984
rect -24334 -12046 -24304 -12015
rect -24238 -12046 -24208 -12015
rect -24142 -12046 -24112 -12015
rect -24046 -12046 -24016 -12015
rect -23950 -12046 -23920 -12015
rect -23854 -12046 -23824 -12015
rect -23680 -12226 -23664 -12000
rect -23630 -12002 -23614 -12000
rect 7422 -11920 7452 -11894
rect 7518 -11920 7548 -11894
rect 7614 -11920 7644 -11894
rect 7710 -11920 7740 -11894
rect 8370 -11920 8400 -11894
rect 8466 -11920 8496 -11894
rect 8562 -11920 8592 -11894
rect 8658 -11920 8688 -11894
rect 9306 -11920 9336 -11894
rect 9402 -11920 9432 -11894
rect 9498 -11920 9528 -11894
rect 9594 -11920 9624 -11894
rect 10237 -11920 10267 -11894
rect 10333 -11920 10363 -11894
rect 10429 -11920 10459 -11894
rect 10525 -11920 10555 -11894
rect 11164 -11920 11194 -11894
rect 11260 -11920 11290 -11894
rect 11356 -11920 11386 -11894
rect 11452 -11920 11482 -11894
rect 11835 -11915 12170 -11881
rect 12204 -11915 12249 -11881
rect 11835 -11928 12249 -11915
rect -21951 -12000 -21885 -11984
rect -23630 -12032 -23583 -12002
rect -23369 -12032 -23343 -12002
rect -23630 -12098 -23614 -12032
rect -22597 -12046 -22567 -12015
rect -22501 -12046 -22471 -12015
rect -22405 -12046 -22375 -12015
rect -22309 -12046 -22279 -12015
rect -22213 -12046 -22183 -12015
rect -22117 -12046 -22087 -12015
rect -23630 -12128 -23583 -12098
rect -23369 -12128 -23343 -12098
rect -23630 -12194 -23614 -12128
rect -23630 -12224 -23583 -12194
rect -23369 -12224 -23343 -12194
rect -23630 -12226 -23614 -12224
rect -23680 -12242 -23614 -12226
rect -24334 -12286 -24304 -12260
rect -24238 -12286 -24208 -12260
rect -24142 -12286 -24112 -12260
rect -24335 -12307 -24112 -12286
rect -24335 -12342 -24318 -12307
rect -24284 -12316 -24112 -12307
rect -24046 -12286 -24016 -12260
rect -23950 -12286 -23920 -12260
rect -23854 -12286 -23824 -12260
rect -21951 -12226 -21935 -12000
rect -21901 -12002 -21885 -12000
rect -21901 -12032 -21854 -12002
rect -21640 -12032 -21614 -12002
rect 7422 -12022 7452 -11996
rect 7518 -12022 7548 -11996
rect 7614 -12022 7644 -11996
rect 7710 -12022 7740 -11996
rect 8370 -12022 8400 -11996
rect 8466 -12022 8496 -11996
rect 8562 -12022 8592 -11996
rect 8658 -12022 8688 -11996
rect 9306 -12022 9336 -11996
rect 9402 -12022 9432 -11996
rect 9498 -12022 9528 -11996
rect 9594 -12022 9624 -11996
rect 10237 -12021 10267 -11995
rect 10333 -12021 10363 -11995
rect 10429 -12021 10459 -11995
rect 10525 -12021 10555 -11995
rect -21901 -12098 -21885 -12032
rect -21901 -12128 -21854 -12098
rect -21640 -12128 -21614 -12098
rect -21901 -12194 -21885 -12128
rect -21901 -12224 -21854 -12194
rect -21640 -12224 -21614 -12194
rect -20468 -12214 -20438 -12183
rect -20372 -12214 -20342 -12183
rect -20276 -12214 -20246 -12183
rect -20180 -12214 -20150 -12183
rect -20084 -12214 -20054 -12183
rect -19988 -12214 -19958 -12183
rect -19359 -12214 -19329 -12183
rect -19263 -12214 -19233 -12183
rect -19167 -12214 -19137 -12183
rect -19071 -12214 -19041 -12183
rect -18975 -12214 -18945 -12183
rect -18879 -12214 -18849 -12183
rect -18477 -12214 -18447 -12183
rect -18381 -12214 -18351 -12183
rect -18285 -12214 -18255 -12183
rect -18189 -12214 -18159 -12183
rect -18093 -12214 -18063 -12183
rect -17997 -12214 -17967 -12183
rect -17177 -12214 -17147 -12183
rect -17081 -12214 -17051 -12183
rect -16985 -12214 -16955 -12183
rect -16889 -12214 -16859 -12183
rect -16793 -12214 -16763 -12183
rect -16697 -12214 -16667 -12183
rect -16068 -12214 -16038 -12183
rect -15972 -12214 -15942 -12183
rect -15876 -12214 -15846 -12183
rect -15780 -12214 -15750 -12183
rect -15684 -12214 -15654 -12183
rect -15588 -12214 -15558 -12183
rect -15186 -12214 -15156 -12183
rect -15090 -12214 -15060 -12183
rect -14994 -12214 -14964 -12183
rect -14898 -12214 -14868 -12183
rect -14802 -12214 -14772 -12183
rect -14706 -12214 -14676 -12183
rect -13886 -12214 -13856 -12183
rect -13790 -12214 -13760 -12183
rect -13694 -12214 -13664 -12183
rect -13598 -12214 -13568 -12183
rect -13502 -12214 -13472 -12183
rect -13406 -12214 -13376 -12183
rect -12777 -12214 -12747 -12183
rect -12681 -12214 -12651 -12183
rect -12585 -12214 -12555 -12183
rect -12489 -12214 -12459 -12183
rect -12393 -12214 -12363 -12183
rect -12297 -12214 -12267 -12183
rect -11895 -12214 -11865 -12183
rect -11799 -12214 -11769 -12183
rect -11703 -12214 -11673 -12183
rect -11607 -12214 -11577 -12183
rect -11511 -12214 -11481 -12183
rect -11415 -12214 -11385 -12183
rect -10595 -12214 -10565 -12183
rect -10499 -12214 -10469 -12183
rect -10403 -12214 -10373 -12183
rect -10307 -12214 -10277 -12183
rect -10211 -12214 -10181 -12183
rect -10115 -12214 -10085 -12183
rect -9486 -12214 -9456 -12183
rect -9390 -12214 -9360 -12183
rect -9294 -12214 -9264 -12183
rect -9198 -12214 -9168 -12183
rect -9102 -12214 -9072 -12183
rect -9006 -12214 -8976 -12183
rect -8604 -12214 -8574 -12183
rect -8508 -12214 -8478 -12183
rect -8412 -12214 -8382 -12183
rect -8316 -12214 -8286 -12183
rect -8220 -12214 -8190 -12183
rect -8124 -12214 -8094 -12183
rect -21901 -12226 -21885 -12224
rect -21951 -12242 -21885 -12226
rect -22597 -12286 -22567 -12260
rect -22501 -12286 -22471 -12260
rect -22405 -12286 -22375 -12260
rect -24046 -12307 -23824 -12286
rect -24284 -12342 -24268 -12316
rect -24335 -12353 -24268 -12342
rect -24046 -12342 -24029 -12307
rect -23995 -12316 -23824 -12307
rect -22598 -12307 -22375 -12286
rect -23995 -12342 -23979 -12316
rect -24046 -12353 -23979 -12342
rect -22598 -12342 -22581 -12307
rect -22547 -12316 -22375 -12307
rect -22309 -12286 -22279 -12260
rect -22213 -12286 -22183 -12260
rect -22117 -12286 -22087 -12260
rect -22309 -12307 -22087 -12286
rect -22547 -12342 -22531 -12316
rect -22598 -12353 -22531 -12342
rect -22309 -12342 -22292 -12307
rect -22258 -12316 -22087 -12307
rect -22258 -12342 -22242 -12316
rect -22309 -12353 -22242 -12342
rect -24335 -12548 -24292 -12353
rect -24250 -12431 -24184 -12415
rect -24250 -12466 -24234 -12431
rect -24200 -12452 -24184 -12431
rect -23680 -12446 -23613 -12430
rect -24200 -12466 -24162 -12452
rect -24250 -12482 -24162 -12466
rect -23762 -12482 -23736 -12452
rect -23680 -12480 -23664 -12446
rect -23630 -12448 -23613 -12446
rect -23630 -12478 -23583 -12448
rect -23383 -12478 -23357 -12448
rect -23630 -12480 -23613 -12478
rect -23680 -12496 -23613 -12480
rect -22598 -12548 -22555 -12353
rect -22513 -12431 -22447 -12415
rect -22513 -12466 -22497 -12431
rect -22463 -12452 -22447 -12431
rect -21951 -12446 -21884 -12430
rect -22463 -12466 -22425 -12452
rect -22513 -12482 -22425 -12466
rect -22025 -12482 -21999 -12452
rect -21951 -12480 -21935 -12446
rect -21901 -12448 -21884 -12446
rect -21901 -12478 -21854 -12448
rect -21654 -12478 -21628 -12448
rect -20468 -12454 -20438 -12428
rect -20372 -12454 -20342 -12428
rect -20276 -12454 -20246 -12428
rect -20469 -12475 -20246 -12454
rect -21901 -12480 -21884 -12478
rect -21951 -12496 -21884 -12480
rect -20469 -12510 -20452 -12475
rect -20418 -12484 -20246 -12475
rect -20180 -12454 -20150 -12428
rect -20084 -12454 -20054 -12428
rect -19988 -12454 -19958 -12428
rect -19359 -12454 -19329 -12428
rect -19263 -12454 -19233 -12428
rect -19167 -12454 -19137 -12428
rect -20180 -12475 -19958 -12454
rect -20418 -12510 -20402 -12484
rect -20469 -12521 -20402 -12510
rect -20180 -12510 -20163 -12475
rect -20129 -12484 -19958 -12475
rect -19360 -12475 -19137 -12454
rect -20129 -12510 -20113 -12484
rect -20180 -12521 -20113 -12510
rect -19360 -12510 -19343 -12475
rect -19309 -12484 -19137 -12475
rect -19071 -12454 -19041 -12428
rect -18975 -12454 -18945 -12428
rect -18879 -12454 -18849 -12428
rect -18477 -12454 -18447 -12428
rect -18381 -12454 -18351 -12428
rect -18285 -12454 -18255 -12428
rect -19071 -12475 -18849 -12454
rect -19309 -12510 -19293 -12484
rect -19360 -12521 -19293 -12510
rect -19071 -12510 -19054 -12475
rect -19020 -12484 -18849 -12475
rect -18478 -12475 -18255 -12454
rect -19020 -12510 -19004 -12484
rect -19071 -12521 -19004 -12510
rect -18478 -12510 -18461 -12475
rect -18427 -12484 -18255 -12475
rect -18189 -12454 -18159 -12428
rect -18093 -12454 -18063 -12428
rect -17997 -12454 -17967 -12428
rect -17177 -12454 -17147 -12428
rect -17081 -12454 -17051 -12428
rect -16985 -12454 -16955 -12428
rect -18189 -12475 -17967 -12454
rect -18427 -12510 -18411 -12484
rect -18478 -12521 -18411 -12510
rect -18189 -12510 -18172 -12475
rect -18138 -12484 -17967 -12475
rect -17178 -12475 -16955 -12454
rect -18138 -12510 -18122 -12484
rect -18189 -12521 -18122 -12510
rect -17178 -12510 -17161 -12475
rect -17127 -12484 -16955 -12475
rect -16889 -12454 -16859 -12428
rect -16793 -12454 -16763 -12428
rect -16697 -12454 -16667 -12428
rect -16068 -12454 -16038 -12428
rect -15972 -12454 -15942 -12428
rect -15876 -12454 -15846 -12428
rect -16889 -12475 -16667 -12454
rect -17127 -12510 -17111 -12484
rect -17178 -12521 -17111 -12510
rect -16889 -12510 -16872 -12475
rect -16838 -12484 -16667 -12475
rect -16069 -12475 -15846 -12454
rect -16838 -12510 -16822 -12484
rect -16889 -12521 -16822 -12510
rect -16069 -12510 -16052 -12475
rect -16018 -12484 -15846 -12475
rect -15780 -12454 -15750 -12428
rect -15684 -12454 -15654 -12428
rect -15588 -12454 -15558 -12428
rect -15186 -12454 -15156 -12428
rect -15090 -12454 -15060 -12428
rect -14994 -12454 -14964 -12428
rect -15780 -12475 -15558 -12454
rect -16018 -12510 -16002 -12484
rect -16069 -12521 -16002 -12510
rect -15780 -12510 -15763 -12475
rect -15729 -12484 -15558 -12475
rect -15187 -12475 -14964 -12454
rect -15729 -12510 -15713 -12484
rect -15780 -12521 -15713 -12510
rect -15187 -12510 -15170 -12475
rect -15136 -12484 -14964 -12475
rect -14898 -12454 -14868 -12428
rect -14802 -12454 -14772 -12428
rect -14706 -12454 -14676 -12428
rect -13886 -12454 -13856 -12428
rect -13790 -12454 -13760 -12428
rect -13694 -12454 -13664 -12428
rect -14898 -12475 -14676 -12454
rect -15136 -12510 -15120 -12484
rect -15187 -12521 -15120 -12510
rect -14898 -12510 -14881 -12475
rect -14847 -12484 -14676 -12475
rect -13887 -12475 -13664 -12454
rect -14847 -12510 -14831 -12484
rect -14898 -12521 -14831 -12510
rect -13887 -12510 -13870 -12475
rect -13836 -12484 -13664 -12475
rect -13598 -12454 -13568 -12428
rect -13502 -12454 -13472 -12428
rect -13406 -12454 -13376 -12428
rect -12777 -12454 -12747 -12428
rect -12681 -12454 -12651 -12428
rect -12585 -12454 -12555 -12428
rect -13598 -12475 -13376 -12454
rect -13836 -12510 -13820 -12484
rect -13887 -12521 -13820 -12510
rect -13598 -12510 -13581 -12475
rect -13547 -12484 -13376 -12475
rect -12778 -12475 -12555 -12454
rect -13547 -12510 -13531 -12484
rect -13598 -12521 -13531 -12510
rect -12778 -12510 -12761 -12475
rect -12727 -12484 -12555 -12475
rect -12489 -12454 -12459 -12428
rect -12393 -12454 -12363 -12428
rect -12297 -12454 -12267 -12428
rect -11895 -12454 -11865 -12428
rect -11799 -12454 -11769 -12428
rect -11703 -12454 -11673 -12428
rect -12489 -12475 -12267 -12454
rect -12727 -12510 -12711 -12484
rect -12778 -12521 -12711 -12510
rect -12489 -12510 -12472 -12475
rect -12438 -12484 -12267 -12475
rect -11896 -12475 -11673 -12454
rect -12438 -12510 -12422 -12484
rect -12489 -12521 -12422 -12510
rect -11896 -12510 -11879 -12475
rect -11845 -12484 -11673 -12475
rect -11607 -12454 -11577 -12428
rect -11511 -12454 -11481 -12428
rect -11415 -12454 -11385 -12428
rect -10595 -12454 -10565 -12428
rect -10499 -12454 -10469 -12428
rect -10403 -12454 -10373 -12428
rect -11607 -12475 -11385 -12454
rect -11845 -12510 -11829 -12484
rect -11896 -12521 -11829 -12510
rect -11607 -12510 -11590 -12475
rect -11556 -12484 -11385 -12475
rect -10596 -12475 -10373 -12454
rect -11556 -12510 -11540 -12484
rect -11607 -12521 -11540 -12510
rect -10596 -12510 -10579 -12475
rect -10545 -12484 -10373 -12475
rect -10307 -12454 -10277 -12428
rect -10211 -12454 -10181 -12428
rect -10115 -12454 -10085 -12428
rect -9486 -12454 -9456 -12428
rect -9390 -12454 -9360 -12428
rect -9294 -12454 -9264 -12428
rect -10307 -12475 -10085 -12454
rect -10545 -12510 -10529 -12484
rect -10596 -12521 -10529 -12510
rect -10307 -12510 -10290 -12475
rect -10256 -12484 -10085 -12475
rect -9487 -12475 -9264 -12454
rect -10256 -12510 -10240 -12484
rect -10307 -12521 -10240 -12510
rect -9487 -12510 -9470 -12475
rect -9436 -12484 -9264 -12475
rect -9198 -12454 -9168 -12428
rect -9102 -12454 -9072 -12428
rect -9006 -12454 -8976 -12428
rect -8604 -12454 -8574 -12428
rect -8508 -12454 -8478 -12428
rect -8412 -12454 -8382 -12428
rect -9198 -12475 -8976 -12454
rect -9436 -12510 -9420 -12484
rect -9487 -12521 -9420 -12510
rect -9198 -12510 -9181 -12475
rect -9147 -12484 -8976 -12475
rect -8605 -12475 -8382 -12454
rect -9147 -12510 -9131 -12484
rect -9198 -12521 -9131 -12510
rect -8605 -12510 -8588 -12475
rect -8554 -12484 -8382 -12475
rect -8316 -12454 -8286 -12428
rect -8220 -12454 -8190 -12428
rect -8124 -12454 -8094 -12428
rect -8316 -12475 -8094 -12454
rect -8554 -12510 -8538 -12484
rect -8605 -12521 -8538 -12510
rect -8316 -12510 -8299 -12475
rect -8265 -12484 -8094 -12475
rect -8265 -12510 -8249 -12484
rect -8316 -12521 -8249 -12510
rect -24335 -12564 -24162 -12548
rect -24335 -12599 -24234 -12564
rect -24200 -12578 -24162 -12564
rect -23762 -12578 -23736 -12548
rect -22598 -12564 -22425 -12548
rect -24200 -12599 -24184 -12578
rect -24335 -12615 -24184 -12599
rect -22598 -12599 -22497 -12564
rect -22463 -12578 -22425 -12564
rect -22025 -12578 -21999 -12548
rect -22463 -12599 -22447 -12578
rect -22598 -12615 -22447 -12599
rect -20469 -12716 -20426 -12521
rect -20384 -12599 -20318 -12583
rect -20384 -12634 -20368 -12599
rect -20334 -12620 -20318 -12599
rect -20334 -12634 -20296 -12620
rect -20384 -12650 -20296 -12634
rect -19896 -12650 -19870 -12620
rect -19360 -12716 -19317 -12521
rect -19275 -12599 -19209 -12583
rect -19275 -12634 -19259 -12599
rect -19225 -12620 -19209 -12599
rect -19225 -12634 -19187 -12620
rect -19275 -12650 -19187 -12634
rect -18787 -12650 -18761 -12620
rect -18478 -12716 -18435 -12521
rect -18393 -12599 -18327 -12583
rect -18393 -12634 -18377 -12599
rect -18343 -12620 -18327 -12599
rect -18343 -12634 -18305 -12620
rect -18393 -12650 -18305 -12634
rect -17905 -12650 -17879 -12620
rect -17178 -12716 -17135 -12521
rect -17093 -12599 -17027 -12583
rect -17093 -12634 -17077 -12599
rect -17043 -12620 -17027 -12599
rect -17043 -12634 -17005 -12620
rect -17093 -12650 -17005 -12634
rect -16605 -12650 -16579 -12620
rect -16069 -12716 -16026 -12521
rect -15984 -12599 -15918 -12583
rect -15984 -12634 -15968 -12599
rect -15934 -12620 -15918 -12599
rect -15934 -12634 -15896 -12620
rect -15984 -12650 -15896 -12634
rect -15496 -12650 -15470 -12620
rect -15187 -12716 -15144 -12521
rect -15102 -12599 -15036 -12583
rect -15102 -12634 -15086 -12599
rect -15052 -12620 -15036 -12599
rect -15052 -12634 -15014 -12620
rect -15102 -12650 -15014 -12634
rect -14614 -12650 -14588 -12620
rect -13887 -12716 -13844 -12521
rect -13802 -12599 -13736 -12583
rect -13802 -12634 -13786 -12599
rect -13752 -12620 -13736 -12599
rect -13752 -12634 -13714 -12620
rect -13802 -12650 -13714 -12634
rect -13314 -12650 -13288 -12620
rect -12778 -12716 -12735 -12521
rect -12693 -12599 -12627 -12583
rect -12693 -12634 -12677 -12599
rect -12643 -12620 -12627 -12599
rect -12643 -12634 -12605 -12620
rect -12693 -12650 -12605 -12634
rect -12205 -12650 -12179 -12620
rect -11896 -12716 -11853 -12521
rect -11811 -12599 -11745 -12583
rect -11811 -12634 -11795 -12599
rect -11761 -12620 -11745 -12599
rect -11761 -12634 -11723 -12620
rect -11811 -12650 -11723 -12634
rect -11323 -12650 -11297 -12620
rect -10596 -12716 -10553 -12521
rect -10511 -12599 -10445 -12583
rect -10511 -12634 -10495 -12599
rect -10461 -12620 -10445 -12599
rect -10461 -12634 -10423 -12620
rect -10511 -12650 -10423 -12634
rect -10023 -12650 -9997 -12620
rect -9487 -12716 -9444 -12521
rect -9402 -12599 -9336 -12583
rect -9402 -12634 -9386 -12599
rect -9352 -12620 -9336 -12599
rect -9352 -12634 -9314 -12620
rect -9402 -12650 -9314 -12634
rect -8914 -12650 -8888 -12620
rect -8605 -12716 -8562 -12521
rect -8520 -12599 -8454 -12583
rect -8520 -12634 -8504 -12599
rect -8470 -12620 -8454 -12599
rect -8470 -12634 -8432 -12620
rect -8520 -12650 -8432 -12634
rect -8032 -12650 -8006 -12620
rect -20469 -12732 -20296 -12716
rect -20469 -12767 -20368 -12732
rect -20334 -12746 -20296 -12732
rect -19896 -12746 -19870 -12716
rect -19360 -12732 -19187 -12716
rect -20334 -12767 -20318 -12746
rect -20469 -12783 -20318 -12767
rect -19360 -12767 -19259 -12732
rect -19225 -12746 -19187 -12732
rect -18787 -12746 -18761 -12716
rect -18478 -12732 -18305 -12716
rect -19225 -12767 -19209 -12746
rect -19360 -12783 -19209 -12767
rect -18478 -12767 -18377 -12732
rect -18343 -12746 -18305 -12732
rect -17905 -12746 -17879 -12716
rect -17178 -12732 -17005 -12716
rect -18343 -12767 -18327 -12746
rect -18478 -12783 -18327 -12767
rect -17178 -12767 -17077 -12732
rect -17043 -12746 -17005 -12732
rect -16605 -12746 -16579 -12716
rect -16069 -12732 -15896 -12716
rect -17043 -12767 -17027 -12746
rect -17178 -12783 -17027 -12767
rect -16069 -12767 -15968 -12732
rect -15934 -12746 -15896 -12732
rect -15496 -12746 -15470 -12716
rect -15187 -12732 -15014 -12716
rect -15934 -12767 -15918 -12746
rect -16069 -12783 -15918 -12767
rect -15187 -12767 -15086 -12732
rect -15052 -12746 -15014 -12732
rect -14614 -12746 -14588 -12716
rect -13887 -12732 -13714 -12716
rect -15052 -12767 -15036 -12746
rect -15187 -12783 -15036 -12767
rect -13887 -12767 -13786 -12732
rect -13752 -12746 -13714 -12732
rect -13314 -12746 -13288 -12716
rect -12778 -12732 -12605 -12716
rect -13752 -12767 -13736 -12746
rect -13887 -12783 -13736 -12767
rect -12778 -12767 -12677 -12732
rect -12643 -12746 -12605 -12732
rect -12205 -12746 -12179 -12716
rect -11896 -12732 -11723 -12716
rect -12643 -12767 -12627 -12746
rect -12778 -12783 -12627 -12767
rect -11896 -12767 -11795 -12732
rect -11761 -12746 -11723 -12732
rect -11323 -12746 -11297 -12716
rect -10596 -12732 -10423 -12716
rect -11761 -12767 -11745 -12746
rect -11896 -12783 -11745 -12767
rect -10596 -12767 -10495 -12732
rect -10461 -12746 -10423 -12732
rect -10023 -12746 -9997 -12716
rect -9487 -12732 -9314 -12716
rect -10461 -12767 -10445 -12746
rect -10596 -12783 -10445 -12767
rect -9487 -12767 -9386 -12732
rect -9352 -12746 -9314 -12732
rect -8914 -12746 -8888 -12716
rect -8605 -12732 -8432 -12716
rect -9352 -12767 -9336 -12746
rect -9487 -12783 -9336 -12767
rect -8605 -12767 -8504 -12732
rect -8470 -12746 -8432 -12732
rect -8032 -12746 -8006 -12716
rect -8470 -12767 -8454 -12746
rect -8605 -12783 -8454 -12767
rect 11164 -12022 11194 -11996
rect 11260 -12022 11290 -11996
rect 11356 -12022 11386 -11996
rect 11452 -12022 11482 -11996
rect 7422 -12855 7452 -12822
rect 7238 -12885 7452 -12855
rect 7238 -13132 7268 -12885
rect 7518 -12927 7548 -12822
rect 7614 -12845 7644 -12822
rect 7374 -13065 7548 -12927
rect 7182 -13148 7326 -13132
rect 7182 -13182 7198 -13148
rect 7232 -13182 7326 -13148
rect 7182 -13198 7326 -13182
rect 7374 -13148 7518 -13065
rect 7590 -13107 7644 -12845
rect 7710 -12972 7740 -12822
rect 8370 -12855 8400 -12822
rect 8186 -12885 8400 -12855
rect 7710 -13002 7848 -12972
rect 7584 -13132 7644 -13107
rect 7758 -13132 7848 -13002
rect 8186 -13132 8216 -12885
rect 8466 -12927 8496 -12822
rect 8562 -12845 8592 -12822
rect 8322 -13065 8496 -12927
rect 7374 -13182 7390 -13148
rect 7424 -13182 7518 -13148
rect 7374 -13198 7518 -13182
rect 7566 -13148 7710 -13132
rect 7566 -13182 7582 -13148
rect 7616 -13182 7710 -13148
rect 7566 -13198 7710 -13182
rect 7758 -13148 7902 -13132
rect 7758 -13182 7774 -13148
rect 7808 -13182 7902 -13148
rect 7758 -13198 7902 -13182
rect 8130 -13148 8274 -13132
rect 8130 -13182 8146 -13148
rect 8180 -13182 8274 -13148
rect 8130 -13198 8274 -13182
rect 8322 -13148 8466 -13065
rect 8538 -13107 8592 -12845
rect 8658 -12972 8688 -12822
rect 9306 -12855 9336 -12822
rect 9122 -12885 9336 -12855
rect 8658 -13002 8796 -12972
rect 8532 -13132 8592 -13107
rect 8706 -13132 8796 -13002
rect 9122 -13132 9152 -12885
rect 9402 -12927 9432 -12822
rect 9498 -12845 9528 -12822
rect 9258 -13065 9432 -12927
rect 8322 -13182 8338 -13148
rect 8372 -13182 8466 -13148
rect 8322 -13198 8466 -13182
rect 8514 -13148 8658 -13132
rect 8514 -13182 8530 -13148
rect 8564 -13182 8658 -13148
rect 8514 -13198 8658 -13182
rect 8706 -13148 8850 -13132
rect 8706 -13182 8722 -13148
rect 8756 -13182 8850 -13148
rect 8706 -13198 8850 -13182
rect 9066 -13148 9210 -13132
rect 9066 -13182 9082 -13148
rect 9116 -13182 9210 -13148
rect 9066 -13198 9210 -13182
rect 9258 -13148 9402 -13065
rect 9474 -13107 9528 -12845
rect 9594 -12972 9624 -12822
rect 10237 -12854 10267 -12821
rect 10053 -12884 10267 -12854
rect 9594 -13002 9732 -12972
rect 9468 -13132 9528 -13107
rect 9642 -13132 9732 -13002
rect 10053 -13131 10083 -12884
rect 10333 -12926 10363 -12821
rect 10429 -12844 10459 -12821
rect 10189 -13064 10363 -12926
rect 9258 -13182 9274 -13148
rect 9308 -13182 9402 -13148
rect 9258 -13198 9402 -13182
rect 9450 -13148 9594 -13132
rect 9450 -13182 9466 -13148
rect 9500 -13182 9594 -13148
rect 9450 -13198 9594 -13182
rect 9642 -13148 9786 -13132
rect 9642 -13182 9658 -13148
rect 9692 -13182 9786 -13148
rect 9642 -13198 9786 -13182
rect 9997 -13147 10141 -13131
rect 9997 -13181 10013 -13147
rect 10047 -13181 10141 -13147
rect 9997 -13197 10141 -13181
rect 10189 -13147 10333 -13064
rect 10405 -13106 10459 -12844
rect 10525 -12971 10555 -12821
rect 12219 -12064 12249 -11928
rect 12315 -11857 12345 -11831
rect 12411 -11857 12441 -11831
rect 12507 -11857 12537 -11831
rect 12603 -11857 12633 -11831
rect 12699 -11857 12729 -11831
rect 12315 -11928 12729 -11857
rect 12315 -11970 12345 -11928
rect 12826 -11965 12842 -11739
rect 12876 -11741 12892 -11739
rect 12876 -11771 12923 -11741
rect 13137 -11771 13163 -11741
rect 12876 -11837 12892 -11771
rect 12876 -11867 12923 -11837
rect 13137 -11867 13163 -11837
rect 12876 -11933 12892 -11867
rect 12876 -11963 12923 -11933
rect 13137 -11963 13163 -11933
rect 12876 -11965 12892 -11963
rect 12297 -11986 12363 -11970
rect 12826 -11981 12892 -11965
rect 12297 -12020 12313 -11986
rect 12347 -12020 12363 -11986
rect 12297 -12036 12363 -12020
rect 12315 -12064 12345 -12036
rect 12826 -12185 12893 -12169
rect 12826 -12219 12842 -12185
rect 12876 -12187 12893 -12185
rect 12876 -12217 12923 -12187
rect 13123 -12217 13149 -12187
rect 12876 -12219 12893 -12217
rect 12826 -12235 12893 -12219
rect 12219 -12290 12249 -12264
rect 12315 -12290 12345 -12264
rect 11164 -12855 11194 -12822
rect 10980 -12885 11194 -12855
rect 10525 -13001 10663 -12971
rect 10399 -13131 10459 -13106
rect 10573 -13131 10663 -13001
rect 10189 -13181 10205 -13147
rect 10239 -13181 10333 -13147
rect 10189 -13197 10333 -13181
rect 10381 -13147 10525 -13131
rect 10381 -13181 10397 -13147
rect 10431 -13181 10525 -13147
rect 10381 -13197 10525 -13181
rect 10573 -13147 10717 -13131
rect 10980 -13132 11010 -12885
rect 11260 -12927 11290 -12822
rect 11356 -12845 11386 -12822
rect 11116 -13065 11290 -12927
rect 10573 -13181 10589 -13147
rect 10623 -13181 10717 -13147
rect 10573 -13197 10717 -13181
rect 7200 -13229 7230 -13198
rect 7296 -13229 7326 -13198
rect 7392 -13229 7422 -13198
rect 7488 -13229 7518 -13198
rect 7584 -13229 7614 -13198
rect 7680 -13229 7710 -13198
rect 7776 -13229 7806 -13198
rect 7872 -13229 7902 -13198
rect 8148 -13229 8178 -13198
rect 8244 -13229 8274 -13198
rect 8340 -13229 8370 -13198
rect 8436 -13229 8466 -13198
rect 8532 -13229 8562 -13198
rect 8628 -13229 8658 -13198
rect 8724 -13229 8754 -13198
rect 8820 -13229 8850 -13198
rect 9084 -13229 9114 -13198
rect 9180 -13229 9210 -13198
rect 9276 -13229 9306 -13198
rect 9372 -13229 9402 -13198
rect 9468 -13229 9498 -13198
rect 9564 -13229 9594 -13198
rect 9660 -13229 9690 -13198
rect 9756 -13229 9786 -13198
rect 10015 -13228 10045 -13197
rect 10111 -13228 10141 -13197
rect 10207 -13228 10237 -13197
rect 10303 -13228 10333 -13197
rect 10399 -13228 10429 -13197
rect 10495 -13228 10525 -13197
rect 10591 -13228 10621 -13197
rect 10687 -13228 10717 -13197
rect 10924 -13148 11068 -13132
rect 10924 -13182 10940 -13148
rect 10974 -13182 11068 -13148
rect 10924 -13198 11068 -13182
rect 11116 -13148 11260 -13065
rect 11332 -13107 11386 -12845
rect 11452 -12972 11482 -12822
rect 11452 -13002 11590 -12972
rect 11326 -13132 11386 -13107
rect 11500 -13132 11590 -13002
rect 11116 -13182 11132 -13148
rect 11166 -13182 11260 -13148
rect 11116 -13198 11260 -13182
rect 11308 -13148 11452 -13132
rect 11308 -13182 11324 -13148
rect 11358 -13182 11452 -13148
rect 11308 -13198 11452 -13182
rect 11500 -13148 11644 -13132
rect 11500 -13182 11516 -13148
rect 11550 -13182 11644 -13148
rect 11500 -13198 11644 -13182
rect 10942 -13229 10972 -13198
rect 11038 -13229 11068 -13198
rect 11134 -13229 11164 -13198
rect 11230 -13229 11260 -13198
rect 11326 -13229 11356 -13198
rect 11422 -13229 11452 -13198
rect 11518 -13229 11548 -13198
rect 11614 -13229 11644 -13198
rect 7200 -13577 7230 -13551
rect 7296 -13577 7326 -13551
rect 7392 -13577 7422 -13551
rect 7488 -13577 7518 -13551
rect 7584 -13577 7614 -13551
rect 7680 -13577 7710 -13551
rect 7776 -13577 7806 -13551
rect 7872 -13577 7902 -13551
rect 8148 -13577 8178 -13551
rect 8244 -13577 8274 -13551
rect 8340 -13577 8370 -13551
rect 8436 -13577 8466 -13551
rect 8532 -13577 8562 -13551
rect 8628 -13577 8658 -13551
rect 8724 -13577 8754 -13551
rect 8820 -13577 8850 -13551
rect 9084 -13577 9114 -13551
rect 9180 -13577 9210 -13551
rect 9276 -13577 9306 -13551
rect 9372 -13577 9402 -13551
rect 9468 -13577 9498 -13551
rect 9564 -13577 9594 -13551
rect 9660 -13577 9690 -13551
rect 9756 -13577 9786 -13551
rect 10015 -13576 10045 -13550
rect 10111 -13576 10141 -13550
rect 10207 -13576 10237 -13550
rect 10303 -13576 10333 -13550
rect 10399 -13576 10429 -13550
rect 10495 -13576 10525 -13550
rect 10591 -13576 10621 -13550
rect 10687 -13576 10717 -13550
rect 10942 -13577 10972 -13551
rect 11038 -13577 11068 -13551
rect 11134 -13577 11164 -13551
rect 11230 -13577 11260 -13551
rect 11326 -13577 11356 -13551
rect 11422 -13577 11452 -13551
rect 11518 -13577 11548 -13551
rect 11614 -13577 11644 -13551
rect -2050 -13818 -2020 -13792
rect -1954 -13818 -1924 -13792
rect -1858 -13818 -1828 -13792
rect -1604 -13832 -1574 -13806
rect -2050 -14063 -2020 -14032
rect -1954 -14063 -1924 -14032
rect -1858 -14063 -1828 -14032
rect -1604 -14062 -1574 -14032
rect -2068 -14079 -1810 -14063
rect -4784 -14122 -4526 -14106
rect -12342 -14181 -12316 -14151
rect -11766 -14181 -11276 -14151
rect -11146 -14181 -11120 -14151
rect -4784 -14156 -4768 -14122
rect -4542 -14156 -4526 -14122
rect -4784 -14172 -4526 -14156
rect -4338 -14122 -4272 -14106
rect -4338 -14156 -4322 -14122
rect -4288 -14156 -4272 -14122
rect -2068 -14113 -2052 -14079
rect -1826 -14113 -1810 -14079
rect -2068 -14129 -1810 -14113
rect -1622 -14079 -1556 -14062
rect -1622 -14113 -1606 -14079
rect -1572 -14113 -1556 -14079
rect -1622 -14129 -1556 -14113
rect -17703 -14591 -17677 -14561
rect -17421 -14591 -17324 -14561
rect -17395 -14657 -17324 -14591
rect -17703 -14687 -17677 -14657
rect -17421 -14687 -17324 -14657
rect -17395 -14753 -17324 -14687
rect -17703 -14783 -17677 -14753
rect -17421 -14783 -17324 -14753
rect -17395 -14849 -17324 -14783
rect -17703 -14879 -17677 -14849
rect -17421 -14879 -17324 -14849
rect -24043 -14916 -24013 -14890
rect -23947 -14916 -23917 -14890
rect -24480 -15008 -24449 -14978
rect -24235 -15008 -24179 -14978
rect -24209 -15074 -24179 -15008
rect -24480 -15104 -24449 -15074
rect -24235 -15104 -24179 -15074
rect -24209 -15133 -24179 -15104
rect -24209 -15149 -24142 -15133
rect -24209 -15170 -24188 -15149
rect -24480 -15200 -24449 -15170
rect -24235 -15183 -24188 -15170
rect -24153 -15183 -24142 -15149
rect -24235 -15200 -24142 -15183
rect -24480 -15296 -24449 -15266
rect -24235 -15296 -24179 -15266
rect -24209 -15362 -24179 -15296
rect -17395 -14945 -17324 -14879
rect -17282 -14943 -17216 -14927
rect -17282 -14945 -17266 -14943
rect -17703 -14975 -17677 -14945
rect -17421 -14975 -17266 -14945
rect -17282 -14977 -17266 -14975
rect -17232 -14945 -17216 -14943
rect -17232 -14975 -17188 -14945
rect -16988 -14975 -16962 -14945
rect -17232 -14977 -17216 -14975
rect -17282 -14993 -17216 -14977
rect -17703 -15071 -17677 -15041
rect -17421 -15071 -17188 -15041
rect -16988 -15071 -16962 -15041
rect -24043 -15338 -24013 -15316
rect -24480 -15392 -24449 -15362
rect -24235 -15392 -24179 -15362
rect -24209 -15422 -24179 -15392
rect -24080 -15354 -24013 -15338
rect -24080 -15388 -24064 -15354
rect -24029 -15388 -24013 -15354
rect -24080 -15404 -24013 -15388
rect -23947 -15338 -23917 -15316
rect -23947 -15354 -23880 -15338
rect -23947 -15388 -23931 -15354
rect -23896 -15388 -23880 -15354
rect -24209 -15438 -24142 -15422
rect -24209 -15458 -24188 -15438
rect -24480 -15488 -24449 -15458
rect -24235 -15472 -24188 -15458
rect -24153 -15446 -24142 -15438
rect -23947 -15446 -23880 -15388
rect -24153 -15472 -23880 -15446
rect -24235 -15488 -23880 -15472
rect -24209 -15489 -23880 -15488
rect -17395 -15086 -17324 -15071
rect -17395 -15120 -17371 -15086
rect -17337 -15120 -17324 -15086
rect -17395 -15137 -17324 -15120
rect -17703 -15167 -17677 -15137
rect -17421 -15167 -17324 -15137
rect -17395 -15233 -17324 -15167
rect -17703 -15263 -17677 -15233
rect -17421 -15263 -17324 -15233
rect -17395 -15329 -17324 -15263
rect -17703 -15359 -17677 -15329
rect -17421 -15359 -17324 -15329
rect -17395 -15425 -17324 -15359
rect -11735 -14243 -11298 -14181
rect -4766 -14203 -4736 -14172
rect -4670 -14203 -4640 -14172
rect -4574 -14203 -4544 -14172
rect -4338 -14173 -4272 -14156
rect -4320 -14203 -4290 -14173
rect -2050 -14197 -2020 -14171
rect -1954 -14197 -1924 -14171
rect -1858 -14197 -1828 -14171
rect -12347 -14273 -12316 -14243
rect -11766 -14273 -11276 -14243
rect -11146 -14273 -11120 -14243
rect -11735 -14339 -11298 -14273
rect -12347 -14369 -12316 -14339
rect -11766 -14368 -11276 -14339
rect -11766 -14369 -11578 -14368
rect -11735 -14433 -11578 -14369
rect -11523 -14369 -11276 -14368
rect -11146 -14369 -11120 -14339
rect -11523 -14433 -11298 -14369
rect -11735 -14435 -11298 -14433
rect -12347 -14465 -12316 -14435
rect -11766 -14465 -11276 -14435
rect -11146 -14465 -11120 -14435
rect -12347 -14561 -12316 -14531
rect -11766 -14550 -11642 -14531
rect -11766 -14561 -11702 -14550
rect -11735 -14627 -11702 -14561
rect -12347 -14657 -12316 -14627
rect -11766 -14657 -11702 -14627
rect -11735 -14680 -11702 -14657
rect -11657 -14680 -11642 -14550
rect -11735 -14723 -11642 -14680
rect -12347 -14753 -12316 -14723
rect -11766 -14753 -11642 -14723
rect -11585 -14561 -11276 -14531
rect -11146 -14561 -11120 -14531
rect -11585 -14627 -11298 -14561
rect -11585 -14657 -11276 -14627
rect -11146 -14657 -11120 -14627
rect -11585 -14723 -11298 -14657
rect -11585 -14753 -11276 -14723
rect -11146 -14753 -11120 -14723
rect -12347 -14849 -12316 -14819
rect -11766 -14849 -11643 -14819
rect -11736 -14881 -11643 -14849
rect -11736 -14915 -11707 -14881
rect -12347 -14945 -12316 -14915
rect -11766 -14945 -11707 -14915
rect -11736 -15011 -11707 -14945
rect -11662 -15011 -11643 -14881
rect -12347 -15041 -12316 -15011
rect -11766 -15041 -11643 -15011
rect -11585 -15105 -11476 -14753
rect -11406 -14849 -11276 -14819
rect -11146 -14849 -11120 -14819
rect -11406 -14873 -11298 -14849
rect -11406 -15003 -11378 -14873
rect -11333 -14915 -11298 -14873
rect -11333 -14945 -11276 -14915
rect -11146 -14945 -11120 -14915
rect -11333 -15003 -11298 -14945
rect -11406 -15011 -11298 -15003
rect -11406 -15041 -11276 -15011
rect -11146 -15041 -11120 -15011
rect -11735 -15107 -11476 -15105
rect -12347 -15137 -12316 -15107
rect -11766 -15137 -11476 -15107
rect -11735 -15203 -11476 -15137
rect -12347 -15233 -12316 -15203
rect -11766 -15233 -11476 -15203
rect -11735 -15299 -11476 -15233
rect -12347 -15329 -12316 -15299
rect -11766 -15329 -11476 -15299
rect -11411 -15137 -11276 -15107
rect -11146 -15137 -11120 -15107
rect -11411 -15156 -11298 -15137
rect -11411 -15286 -11386 -15156
rect -11341 -15203 -11298 -15156
rect -11341 -15233 -11276 -15203
rect -11146 -15233 -11120 -15203
rect -11341 -15286 -11298 -15233
rect -11411 -15299 -11298 -15286
rect -11411 -15329 -11276 -15299
rect -11146 -15329 -11120 -15299
rect -11735 -15378 -11476 -15329
rect -11735 -15391 -11301 -15378
rect -4766 -14443 -4736 -14417
rect -4670 -14443 -4640 -14417
rect -4574 -14443 -4544 -14417
rect -4320 -14429 -4290 -14403
rect -1604 -14211 -1574 -14185
rect 5561 -14249 5627 -14233
rect -2050 -14442 -2020 -14411
rect -1954 -14442 -1924 -14411
rect -1858 -14442 -1828 -14411
rect -1604 -14441 -1574 -14411
rect -2068 -14458 -1810 -14442
rect -2068 -14492 -2052 -14458
rect -1826 -14492 -1810 -14458
rect -2068 -14508 -1810 -14492
rect -1622 -14458 -1556 -14441
rect -1622 -14492 -1606 -14458
rect -1572 -14492 -1556 -14458
rect 5561 -14475 5577 -14249
rect 5611 -14251 5627 -14249
rect 6001 -14249 6067 -14233
rect 5611 -14281 5658 -14251
rect 5872 -14281 5898 -14251
rect 5611 -14347 5627 -14281
rect 5611 -14377 5658 -14347
rect 5872 -14377 5898 -14347
rect 5611 -14443 5627 -14377
rect 5611 -14473 5658 -14443
rect 5872 -14473 5898 -14443
rect 5611 -14475 5627 -14473
rect 5561 -14491 5627 -14475
rect -1622 -14508 -1556 -14492
rect 6001 -14475 6017 -14249
rect 6051 -14251 6067 -14249
rect 6441 -14249 6507 -14233
rect 6051 -14281 6098 -14251
rect 6312 -14281 6338 -14251
rect 6051 -14347 6067 -14281
rect 6051 -14377 6098 -14347
rect 6312 -14377 6338 -14347
rect 6051 -14443 6067 -14377
rect 6051 -14473 6098 -14443
rect 6312 -14473 6338 -14443
rect 6051 -14475 6067 -14473
rect 6001 -14491 6067 -14475
rect 6441 -14475 6457 -14249
rect 6491 -14251 6507 -14249
rect 6491 -14281 6538 -14251
rect 6752 -14281 6778 -14251
rect 6491 -14347 6507 -14281
rect 6491 -14377 6538 -14347
rect 6752 -14377 6778 -14347
rect 6491 -14443 6507 -14377
rect 6491 -14473 6538 -14443
rect 6752 -14473 6778 -14443
rect 6491 -14475 6507 -14473
rect 6441 -14491 6507 -14475
rect -4784 -14562 -4526 -14546
rect -4784 -14596 -4768 -14562
rect -4542 -14596 -4526 -14562
rect -4784 -14612 -4526 -14596
rect -4338 -14562 -4272 -14546
rect -4338 -14596 -4322 -14562
rect -4288 -14596 -4272 -14562
rect -4766 -14643 -4736 -14612
rect -4670 -14643 -4640 -14612
rect -4574 -14643 -4544 -14612
rect -4338 -14613 -4272 -14596
rect -4320 -14643 -4290 -14613
rect -2050 -14637 -2020 -14611
rect -1954 -14637 -1924 -14611
rect -1858 -14637 -1828 -14611
rect -4766 -14883 -4736 -14857
rect -4670 -14883 -4640 -14857
rect -4574 -14883 -4544 -14857
rect -4320 -14869 -4290 -14843
rect -1604 -14651 -1574 -14625
rect 5561 -14695 5628 -14679
rect 5561 -14729 5577 -14695
rect 5611 -14697 5628 -14695
rect 6001 -14695 6068 -14679
rect 5611 -14727 5658 -14697
rect 5858 -14727 5884 -14697
rect 5611 -14729 5628 -14727
rect 5561 -14745 5628 -14729
rect 6001 -14729 6017 -14695
rect 6051 -14697 6068 -14695
rect 6441 -14695 6508 -14679
rect 6051 -14727 6098 -14697
rect 6298 -14727 6324 -14697
rect 6051 -14729 6068 -14727
rect 6001 -14745 6068 -14729
rect 6441 -14729 6457 -14695
rect 6491 -14697 6508 -14695
rect 6491 -14727 6538 -14697
rect 6738 -14727 6764 -14697
rect 6491 -14729 6508 -14727
rect 6441 -14745 6508 -14729
rect -2050 -14882 -2020 -14851
rect -1954 -14882 -1924 -14851
rect -1858 -14882 -1828 -14851
rect -1604 -14881 -1574 -14851
rect -2068 -14898 -1810 -14882
rect -4784 -14941 -4526 -14925
rect -4784 -14975 -4768 -14941
rect -4542 -14975 -4526 -14941
rect -4784 -14991 -4526 -14975
rect -4338 -14941 -4272 -14925
rect -4338 -14975 -4322 -14941
rect -4288 -14975 -4272 -14941
rect -2068 -14932 -2052 -14898
rect -1826 -14932 -1810 -14898
rect -2068 -14948 -1810 -14932
rect -1622 -14898 -1556 -14881
rect 7200 -14893 7230 -14867
rect 7296 -14893 7326 -14867
rect 7392 -14893 7422 -14867
rect 7488 -14893 7518 -14867
rect 7584 -14893 7614 -14867
rect 7680 -14893 7710 -14867
rect 7776 -14893 7806 -14867
rect 7872 -14893 7902 -14867
rect 8148 -14893 8178 -14867
rect 8244 -14893 8274 -14867
rect 8340 -14893 8370 -14867
rect 8436 -14893 8466 -14867
rect 8532 -14893 8562 -14867
rect 8628 -14893 8658 -14867
rect 8724 -14893 8754 -14867
rect 8820 -14893 8850 -14867
rect 9084 -14893 9114 -14867
rect 9180 -14893 9210 -14867
rect 9276 -14893 9306 -14867
rect 9372 -14893 9402 -14867
rect 9468 -14893 9498 -14867
rect 9564 -14893 9594 -14867
rect 9660 -14893 9690 -14867
rect 9756 -14893 9786 -14867
rect 10015 -14893 10045 -14867
rect 10111 -14893 10141 -14867
rect 10207 -14893 10237 -14867
rect 10303 -14893 10333 -14867
rect 10399 -14893 10429 -14867
rect 10495 -14893 10525 -14867
rect 10591 -14893 10621 -14867
rect 10687 -14893 10717 -14867
rect 10942 -14893 10972 -14867
rect 11038 -14893 11068 -14867
rect 11134 -14893 11164 -14867
rect 11230 -14893 11260 -14867
rect 11326 -14893 11356 -14867
rect 11422 -14893 11452 -14867
rect 11518 -14893 11548 -14867
rect 11614 -14893 11644 -14867
rect -1622 -14932 -1606 -14898
rect -1572 -14932 -1556 -14898
rect -1622 -14948 -1556 -14932
rect -4766 -15022 -4736 -14991
rect -4670 -15022 -4640 -14991
rect -4574 -15022 -4544 -14991
rect -4338 -14992 -4272 -14975
rect -4320 -15022 -4290 -14992
rect -2050 -15016 -2020 -14990
rect -1954 -15016 -1924 -14990
rect -1858 -15016 -1828 -14990
rect -4766 -15262 -4736 -15236
rect -4670 -15262 -4640 -15236
rect -4574 -15262 -4544 -15236
rect -4320 -15248 -4290 -15222
rect -1604 -15030 -1574 -15004
rect -2050 -15261 -2020 -15230
rect -1954 -15261 -1924 -15230
rect -1858 -15261 -1828 -15230
rect -1604 -15260 -1574 -15230
rect 7200 -15246 7230 -15215
rect 7296 -15246 7326 -15215
rect 7392 -15246 7422 -15215
rect 7488 -15246 7518 -15215
rect 7584 -15246 7614 -15215
rect 7680 -15246 7710 -15215
rect 7776 -15246 7806 -15215
rect 7872 -15246 7902 -15215
rect 8148 -15246 8178 -15215
rect 8244 -15246 8274 -15215
rect 8340 -15246 8370 -15215
rect 8436 -15246 8466 -15215
rect 8532 -15246 8562 -15215
rect 8628 -15246 8658 -15215
rect 8724 -15246 8754 -15215
rect 8820 -15246 8850 -15215
rect 9084 -15246 9114 -15215
rect 9180 -15246 9210 -15215
rect 9276 -15246 9306 -15215
rect 9372 -15246 9402 -15215
rect 9468 -15246 9498 -15215
rect 9564 -15246 9594 -15215
rect 9660 -15246 9690 -15215
rect 9756 -15246 9786 -15215
rect 10015 -15246 10045 -15215
rect 10111 -15246 10141 -15215
rect 10207 -15246 10237 -15215
rect 10303 -15246 10333 -15215
rect 10399 -15246 10429 -15215
rect 10495 -15246 10525 -15215
rect 10591 -15246 10621 -15215
rect 10687 -15246 10717 -15215
rect 10942 -15246 10972 -15215
rect 11038 -15246 11068 -15215
rect 11134 -15246 11164 -15215
rect 11230 -15246 11260 -15215
rect 11326 -15246 11356 -15215
rect 11422 -15246 11452 -15215
rect 11518 -15246 11548 -15215
rect 11614 -15246 11644 -15215
rect -2068 -15277 -1810 -15261
rect -2068 -15311 -2052 -15277
rect -1826 -15311 -1810 -15277
rect -8117 -15346 -8087 -15320
rect -8021 -15346 -7991 -15320
rect -7925 -15346 -7895 -15320
rect -2068 -15327 -1810 -15311
rect -1622 -15277 -1556 -15260
rect -1622 -15311 -1606 -15277
rect -1572 -15311 -1556 -15277
rect -1622 -15327 -1556 -15311
rect 7182 -15262 7326 -15246
rect 7182 -15296 7198 -15262
rect 7232 -15296 7326 -15262
rect 7182 -15312 7326 -15296
rect 7374 -15262 7518 -15246
rect 7374 -15296 7390 -15262
rect 7424 -15296 7518 -15262
rect -12342 -15421 -12316 -15391
rect -11766 -15421 -11276 -15391
rect -11146 -15421 -11120 -15391
rect -17703 -15455 -17677 -15425
rect -17421 -15455 -17324 -15425
rect -11735 -15454 -11301 -15421
rect -11585 -15515 -11476 -15454
rect -11579 -15604 -11481 -15515
rect -7671 -15360 -7641 -15334
rect -4784 -15381 -4526 -15365
rect -4784 -15415 -4768 -15381
rect -4542 -15415 -4526 -15381
rect -4784 -15431 -4526 -15415
rect -4338 -15381 -4272 -15365
rect -4338 -15415 -4322 -15381
rect -4288 -15415 -4272 -15381
rect -4766 -15462 -4736 -15431
rect -4670 -15462 -4640 -15431
rect -4574 -15462 -4544 -15431
rect -4338 -15432 -4272 -15415
rect -4320 -15462 -4290 -15432
rect -2050 -15456 -2020 -15430
rect -1954 -15456 -1924 -15430
rect -1858 -15456 -1828 -15430
rect -8117 -15591 -8087 -15560
rect -8021 -15591 -7991 -15560
rect -7925 -15591 -7895 -15560
rect -7671 -15590 -7641 -15560
rect -11579 -15658 -11557 -15604
rect -11503 -15658 -11481 -15604
rect -8135 -15607 -7877 -15591
rect -8135 -15641 -8119 -15607
rect -7893 -15641 -7877 -15607
rect -8135 -15657 -7877 -15641
rect -7689 -15607 -7623 -15590
rect -7689 -15641 -7673 -15607
rect -7639 -15641 -7623 -15607
rect -7689 -15657 -7623 -15641
rect -11579 -15674 -11481 -15658
rect -4766 -15702 -4736 -15676
rect -4670 -15702 -4640 -15676
rect -4574 -15702 -4544 -15676
rect -4320 -15688 -4290 -15662
rect -1604 -15470 -1574 -15444
rect 7238 -15559 7268 -15312
rect 7374 -15379 7518 -15296
rect 7566 -15262 7710 -15246
rect 7566 -15296 7582 -15262
rect 7616 -15296 7710 -15262
rect 7566 -15312 7710 -15296
rect 7758 -15262 7902 -15246
rect 7758 -15296 7774 -15262
rect 7808 -15296 7902 -15262
rect 7758 -15312 7902 -15296
rect 8130 -15262 8274 -15246
rect 8130 -15296 8146 -15262
rect 8180 -15296 8274 -15262
rect 8130 -15312 8274 -15296
rect 8322 -15262 8466 -15246
rect 8322 -15296 8338 -15262
rect 8372 -15296 8466 -15262
rect 7584 -15337 7644 -15312
rect 7374 -15517 7548 -15379
rect 7238 -15589 7452 -15559
rect 7422 -15622 7452 -15589
rect 7518 -15622 7548 -15517
rect 7590 -15599 7644 -15337
rect 7758 -15442 7848 -15312
rect 7614 -15622 7644 -15599
rect 7710 -15472 7848 -15442
rect 7710 -15622 7740 -15472
rect 8186 -15559 8216 -15312
rect 8322 -15379 8466 -15296
rect 8514 -15262 8658 -15246
rect 8514 -15296 8530 -15262
rect 8564 -15296 8658 -15262
rect 8514 -15312 8658 -15296
rect 8706 -15262 8850 -15246
rect 8706 -15296 8722 -15262
rect 8756 -15296 8850 -15262
rect 8706 -15312 8850 -15296
rect 9066 -15262 9210 -15246
rect 9066 -15296 9082 -15262
rect 9116 -15296 9210 -15262
rect 9066 -15312 9210 -15296
rect 9258 -15262 9402 -15246
rect 9258 -15296 9274 -15262
rect 9308 -15296 9402 -15262
rect 8532 -15337 8592 -15312
rect 8322 -15517 8496 -15379
rect 8186 -15589 8400 -15559
rect 8370 -15622 8400 -15589
rect 8466 -15622 8496 -15517
rect 8538 -15599 8592 -15337
rect 8706 -15442 8796 -15312
rect 8562 -15622 8592 -15599
rect 8658 -15472 8796 -15442
rect 8658 -15622 8688 -15472
rect 9122 -15559 9152 -15312
rect 9258 -15379 9402 -15296
rect 9450 -15262 9594 -15246
rect 9450 -15296 9466 -15262
rect 9500 -15296 9594 -15262
rect 9450 -15312 9594 -15296
rect 9642 -15262 9786 -15246
rect 9642 -15296 9658 -15262
rect 9692 -15296 9786 -15262
rect 9642 -15312 9786 -15296
rect 9997 -15262 10141 -15246
rect 9997 -15296 10013 -15262
rect 10047 -15296 10141 -15262
rect 9997 -15312 10141 -15296
rect 10189 -15262 10333 -15246
rect 10189 -15296 10205 -15262
rect 10239 -15296 10333 -15262
rect 9468 -15337 9528 -15312
rect 9258 -15517 9432 -15379
rect 9122 -15589 9336 -15559
rect 9306 -15622 9336 -15589
rect 9402 -15622 9432 -15517
rect 9474 -15599 9528 -15337
rect 9642 -15442 9732 -15312
rect 9498 -15622 9528 -15599
rect 9594 -15472 9732 -15442
rect 9594 -15622 9624 -15472
rect 10053 -15559 10083 -15312
rect 10189 -15379 10333 -15296
rect 10381 -15262 10525 -15246
rect 10381 -15296 10397 -15262
rect 10431 -15296 10525 -15262
rect 10381 -15312 10525 -15296
rect 10573 -15262 10717 -15246
rect 10573 -15296 10589 -15262
rect 10623 -15296 10717 -15262
rect 10573 -15312 10717 -15296
rect 10924 -15262 11068 -15246
rect 10924 -15296 10940 -15262
rect 10974 -15296 11068 -15262
rect 10924 -15312 11068 -15296
rect 11116 -15262 11260 -15246
rect 11116 -15296 11132 -15262
rect 11166 -15296 11260 -15262
rect 10399 -15337 10459 -15312
rect 10189 -15517 10363 -15379
rect 10053 -15589 10267 -15559
rect 10237 -15622 10267 -15589
rect 10333 -15622 10363 -15517
rect 10405 -15599 10459 -15337
rect 10573 -15442 10663 -15312
rect 10429 -15622 10459 -15599
rect 10525 -15472 10663 -15442
rect 10525 -15622 10555 -15472
rect 10980 -15559 11010 -15312
rect 11116 -15379 11260 -15296
rect 11308 -15262 11452 -15246
rect 11308 -15296 11324 -15262
rect 11358 -15296 11452 -15262
rect 11308 -15312 11452 -15296
rect 11500 -15262 11644 -15246
rect 11500 -15296 11516 -15262
rect 11550 -15296 11644 -15262
rect 11500 -15312 11644 -15296
rect 11326 -15337 11386 -15312
rect 11116 -15517 11290 -15379
rect 10980 -15589 11194 -15559
rect 11164 -15622 11194 -15589
rect 11260 -15622 11290 -15517
rect 11332 -15599 11386 -15337
rect 11500 -15442 11590 -15312
rect 11356 -15622 11386 -15599
rect 11452 -15472 11590 -15442
rect 11452 -15622 11482 -15472
rect -2050 -15701 -2020 -15670
rect -1954 -15701 -1924 -15670
rect -1858 -15701 -1828 -15670
rect -1604 -15700 -1574 -15670
rect -2068 -15717 -1810 -15701
rect -4784 -15760 -4526 -15744
rect -4784 -15794 -4768 -15760
rect -4542 -15794 -4526 -15760
rect -4784 -15810 -4526 -15794
rect -4338 -15760 -4272 -15744
rect -4338 -15794 -4322 -15760
rect -4288 -15794 -4272 -15760
rect -2068 -15751 -2052 -15717
rect -1826 -15751 -1810 -15717
rect -2068 -15767 -1810 -15751
rect -1622 -15717 -1556 -15700
rect -1622 -15751 -1606 -15717
rect -1572 -15751 -1556 -15717
rect -1622 -15767 -1556 -15751
rect -8116 -15846 -8086 -15820
rect -8020 -15846 -7990 -15820
rect -7924 -15846 -7894 -15820
rect -17703 -15991 -17677 -15961
rect -17421 -15991 -17324 -15961
rect -17395 -16057 -17324 -15991
rect -24042 -16101 -24012 -16075
rect -23946 -16101 -23916 -16075
rect -17703 -16087 -17677 -16057
rect -17421 -16087 -17324 -16057
rect -7670 -15860 -7640 -15834
rect -4766 -15841 -4736 -15810
rect -4670 -15841 -4640 -15810
rect -4574 -15841 -4544 -15810
rect -4338 -15811 -4272 -15794
rect -4320 -15841 -4290 -15811
rect -2050 -15835 -2020 -15809
rect -1954 -15835 -1924 -15809
rect -1858 -15835 -1828 -15809
rect -24479 -16193 -24448 -16163
rect -24234 -16193 -24178 -16163
rect -24208 -16259 -24178 -16193
rect -24479 -16289 -24448 -16259
rect -24234 -16289 -24178 -16259
rect -24208 -16318 -24178 -16289
rect -24208 -16334 -24141 -16318
rect -24208 -16355 -24187 -16334
rect -24479 -16385 -24448 -16355
rect -24234 -16368 -24187 -16355
rect -24152 -16368 -24141 -16334
rect -24234 -16385 -24141 -16368
rect -24479 -16481 -24448 -16451
rect -24234 -16481 -24178 -16451
rect -24208 -16547 -24178 -16481
rect -17395 -16153 -17324 -16087
rect -8116 -16091 -8086 -16060
rect -8020 -16091 -7990 -16060
rect -7924 -16091 -7894 -16060
rect -7670 -16090 -7640 -16060
rect -4766 -16081 -4736 -16055
rect -4670 -16081 -4640 -16055
rect -4574 -16081 -4544 -16055
rect -4320 -16067 -4290 -16041
rect -1604 -15849 -1574 -15823
rect -2050 -16080 -2020 -16049
rect -1954 -16080 -1924 -16049
rect -1858 -16080 -1828 -16049
rect -1604 -16079 -1574 -16049
rect -17703 -16183 -17677 -16153
rect -17421 -16183 -17324 -16153
rect -8134 -16107 -7876 -16091
rect -8134 -16141 -8118 -16107
rect -7892 -16141 -7876 -16107
rect -8134 -16157 -7876 -16141
rect -7688 -16107 -7622 -16090
rect -7688 -16141 -7672 -16107
rect -7638 -16141 -7622 -16107
rect -7688 -16157 -7622 -16141
rect -2068 -16096 -1810 -16080
rect -2068 -16130 -2052 -16096
rect -1826 -16130 -1810 -16096
rect -2068 -16146 -1810 -16130
rect -1622 -16096 -1556 -16079
rect -1622 -16130 -1606 -16096
rect -1572 -16130 -1556 -16096
rect -1622 -16146 -1556 -16130
rect -17395 -16249 -17324 -16183
rect -17703 -16279 -17677 -16249
rect -17421 -16279 -17324 -16249
rect -4784 -16200 -4526 -16184
rect -4784 -16234 -4768 -16200
rect -4542 -16234 -4526 -16200
rect -4784 -16250 -4526 -16234
rect -4338 -16200 -4272 -16184
rect -4338 -16234 -4322 -16200
rect -4288 -16234 -4272 -16200
rect -17395 -16345 -17324 -16279
rect -4766 -16281 -4736 -16250
rect -4670 -16281 -4640 -16250
rect -4574 -16281 -4544 -16250
rect -4338 -16251 -4272 -16234
rect -4320 -16281 -4290 -16251
rect -2050 -16275 -2020 -16249
rect -1954 -16275 -1924 -16249
rect -1858 -16275 -1828 -16249
rect -17282 -16343 -17216 -16327
rect -17282 -16345 -17266 -16343
rect -17703 -16375 -17677 -16345
rect -17421 -16375 -17266 -16345
rect -17282 -16377 -17266 -16375
rect -17232 -16345 -17216 -16343
rect -17232 -16375 -17188 -16345
rect -16988 -16375 -16962 -16345
rect -17232 -16377 -17216 -16375
rect -17282 -16393 -17216 -16377
rect -17703 -16471 -17677 -16441
rect -17421 -16471 -17188 -16441
rect -16988 -16471 -16962 -16441
rect -24042 -16523 -24012 -16501
rect -24479 -16577 -24448 -16547
rect -24234 -16577 -24178 -16547
rect -24208 -16607 -24178 -16577
rect -24079 -16539 -24012 -16523
rect -24079 -16573 -24063 -16539
rect -24028 -16573 -24012 -16539
rect -24079 -16589 -24012 -16573
rect -23946 -16523 -23916 -16501
rect -23946 -16539 -23879 -16523
rect -23946 -16573 -23930 -16539
rect -23895 -16573 -23879 -16539
rect -24208 -16623 -24141 -16607
rect -24208 -16643 -24187 -16623
rect -24479 -16673 -24448 -16643
rect -24234 -16657 -24187 -16643
rect -24152 -16631 -24141 -16623
rect -23946 -16631 -23879 -16573
rect -24152 -16657 -23879 -16631
rect -24234 -16673 -23879 -16657
rect -24208 -16674 -23879 -16673
rect -17395 -16486 -17324 -16471
rect -17395 -16520 -17371 -16486
rect -17337 -16520 -17324 -16486
rect -17395 -16537 -17324 -16520
rect -8117 -16326 -8087 -16300
rect -8021 -16326 -7991 -16300
rect -7925 -16326 -7895 -16300
rect -17703 -16567 -17677 -16537
rect -17421 -16567 -17324 -16537
rect -7671 -16340 -7641 -16314
rect -4766 -16521 -4736 -16495
rect -4670 -16521 -4640 -16495
rect -4574 -16521 -4544 -16495
rect -4320 -16507 -4290 -16481
rect -1604 -16289 -1574 -16263
rect 11835 -16103 11865 -16077
rect 11931 -16103 11961 -16077
rect 12027 -16103 12057 -16077
rect 12123 -16103 12153 -16077
rect 12219 -16103 12249 -16077
rect 12315 -16103 12345 -16077
rect 12411 -16103 12441 -16077
rect 12507 -16103 12537 -16077
rect 12603 -16103 12633 -16077
rect 12699 -16103 12729 -16077
rect 12826 -16267 12892 -16251
rect 11835 -16385 11865 -16359
rect 11931 -16385 11961 -16359
rect 12027 -16385 12057 -16359
rect 12123 -16385 12153 -16359
rect 12219 -16385 12249 -16359
rect 11835 -16409 12249 -16385
rect 7422 -16448 7452 -16422
rect 7518 -16448 7548 -16422
rect 7614 -16448 7644 -16422
rect 7710 -16448 7740 -16422
rect 8370 -16448 8400 -16422
rect 8466 -16448 8496 -16422
rect 8562 -16448 8592 -16422
rect 8658 -16448 8688 -16422
rect 9306 -16448 9336 -16422
rect 9402 -16448 9432 -16422
rect 9498 -16448 9528 -16422
rect 9594 -16448 9624 -16422
rect 10237 -16448 10267 -16422
rect 10333 -16448 10363 -16422
rect 10429 -16448 10459 -16422
rect 10525 -16448 10555 -16422
rect 11164 -16448 11194 -16422
rect 11260 -16448 11290 -16422
rect 11356 -16448 11386 -16422
rect 11452 -16448 11482 -16422
rect 11835 -16443 12170 -16409
rect 12204 -16443 12249 -16409
rect 11835 -16456 12249 -16443
rect -2050 -16520 -2020 -16489
rect -1954 -16520 -1924 -16489
rect -1858 -16520 -1828 -16489
rect -1604 -16519 -1574 -16489
rect -2068 -16536 -1810 -16520
rect -17395 -16633 -17324 -16567
rect -8117 -16571 -8087 -16540
rect -8021 -16571 -7991 -16540
rect -7925 -16571 -7895 -16540
rect -7671 -16570 -7641 -16540
rect -17703 -16663 -17677 -16633
rect -17421 -16663 -17324 -16633
rect -8135 -16587 -7877 -16571
rect -8135 -16621 -8119 -16587
rect -7893 -16621 -7877 -16587
rect -8135 -16637 -7877 -16621
rect -7689 -16587 -7623 -16570
rect -7689 -16621 -7673 -16587
rect -7639 -16621 -7623 -16587
rect -7689 -16637 -7623 -16621
rect -4784 -16579 -4526 -16563
rect -4784 -16613 -4768 -16579
rect -4542 -16613 -4526 -16579
rect -4784 -16629 -4526 -16613
rect -4338 -16579 -4272 -16563
rect -4338 -16613 -4322 -16579
rect -4288 -16613 -4272 -16579
rect -2068 -16570 -2052 -16536
rect -1826 -16570 -1810 -16536
rect -2068 -16586 -1810 -16570
rect -1622 -16536 -1556 -16519
rect -1622 -16570 -1606 -16536
rect -1572 -16570 -1556 -16536
rect 7422 -16550 7452 -16524
rect 7518 -16550 7548 -16524
rect 7614 -16550 7644 -16524
rect 7710 -16550 7740 -16524
rect 8370 -16550 8400 -16524
rect 8466 -16550 8496 -16524
rect 8562 -16550 8592 -16524
rect 8658 -16550 8688 -16524
rect 9306 -16550 9336 -16524
rect 9402 -16550 9432 -16524
rect 9498 -16550 9528 -16524
rect 9594 -16550 9624 -16524
rect 10237 -16549 10267 -16523
rect 10333 -16549 10363 -16523
rect 10429 -16549 10459 -16523
rect 10525 -16549 10555 -16523
rect -1622 -16586 -1556 -16570
rect -4766 -16660 -4736 -16629
rect -4670 -16660 -4640 -16629
rect -4574 -16660 -4544 -16629
rect -4338 -16630 -4272 -16613
rect -4320 -16660 -4290 -16630
rect -2050 -16654 -2020 -16628
rect -1954 -16654 -1924 -16628
rect -1858 -16654 -1828 -16628
rect -17395 -16729 -17324 -16663
rect -17703 -16759 -17677 -16729
rect -17421 -16759 -17324 -16729
rect -17395 -16825 -17324 -16759
rect -17703 -16855 -17677 -16825
rect -17421 -16855 -17324 -16825
rect -8117 -16826 -8087 -16800
rect -8021 -16826 -7991 -16800
rect -7925 -16826 -7895 -16800
rect -12340 -16997 -12314 -16967
rect -11764 -16997 -11274 -16967
rect -11144 -16997 -11118 -16967
rect -24037 -17314 -24007 -17288
rect -23941 -17314 -23911 -17288
rect -24474 -17406 -24443 -17376
rect -24229 -17406 -24173 -17376
rect -24203 -17472 -24173 -17406
rect -24474 -17502 -24443 -17472
rect -24229 -17502 -24173 -17472
rect -24203 -17531 -24173 -17502
rect -24203 -17547 -24136 -17531
rect -24203 -17568 -24182 -17547
rect -24474 -17598 -24443 -17568
rect -24229 -17581 -24182 -17568
rect -24147 -17581 -24136 -17547
rect -24229 -17598 -24136 -17581
rect -24474 -17694 -24443 -17664
rect -24229 -17694 -24173 -17664
rect -24203 -17760 -24173 -17694
rect -17703 -17391 -17677 -17361
rect -17421 -17391 -17324 -17361
rect -17395 -17457 -17324 -17391
rect -17703 -17487 -17677 -17457
rect -17421 -17487 -17324 -17457
rect -17395 -17553 -17324 -17487
rect -17703 -17583 -17677 -17553
rect -17421 -17583 -17324 -17553
rect -17395 -17649 -17324 -17583
rect -17703 -17679 -17677 -17649
rect -17421 -17679 -17324 -17649
rect -24037 -17736 -24007 -17714
rect -24474 -17790 -24443 -17760
rect -24229 -17790 -24173 -17760
rect -24203 -17820 -24173 -17790
rect -24074 -17752 -24007 -17736
rect -24074 -17786 -24058 -17752
rect -24023 -17786 -24007 -17752
rect -24074 -17802 -24007 -17786
rect -23941 -17736 -23911 -17714
rect -23941 -17752 -23874 -17736
rect -17395 -17745 -17324 -17679
rect -17282 -17743 -17216 -17727
rect -17282 -17745 -17266 -17743
rect -23941 -17786 -23925 -17752
rect -23890 -17786 -23874 -17752
rect -17703 -17775 -17677 -17745
rect -17421 -17775 -17266 -17745
rect -24203 -17836 -24136 -17820
rect -24203 -17856 -24182 -17836
rect -24474 -17886 -24443 -17856
rect -24229 -17870 -24182 -17856
rect -24147 -17844 -24136 -17836
rect -23941 -17844 -23874 -17786
rect -17282 -17777 -17266 -17775
rect -17232 -17745 -17216 -17743
rect -17232 -17775 -17188 -17745
rect -16988 -17775 -16962 -17745
rect -17232 -17777 -17216 -17775
rect -17282 -17793 -17216 -17777
rect -24147 -17870 -23874 -17844
rect -24229 -17886 -23874 -17870
rect -17703 -17871 -17677 -17841
rect -17421 -17871 -17188 -17841
rect -16988 -17871 -16962 -17841
rect -24203 -17887 -23874 -17886
rect -21556 -18034 -21526 -18008
rect -21460 -18034 -21430 -18008
rect -21364 -18034 -21334 -18008
rect -21110 -18048 -21080 -18022
rect -21556 -18279 -21526 -18248
rect -21460 -18279 -21430 -18248
rect -21364 -18279 -21334 -18248
rect -21110 -18278 -21080 -18248
rect -21574 -18295 -21316 -18279
rect -21574 -18329 -21558 -18295
rect -21332 -18329 -21316 -18295
rect -21574 -18345 -21316 -18329
rect -21128 -18295 -21062 -18278
rect -21128 -18329 -21112 -18295
rect -21078 -18329 -21062 -18295
rect -17395 -17886 -17324 -17871
rect -17395 -17920 -17371 -17886
rect -17337 -17920 -17324 -17886
rect -17395 -17937 -17324 -17920
rect -15965 -17905 -15935 -17879
rect -15869 -17905 -15839 -17879
rect -15773 -17905 -15743 -17879
rect -17703 -17967 -17677 -17937
rect -17421 -17967 -17324 -17937
rect -17395 -18033 -17324 -17967
rect -17703 -18063 -17677 -18033
rect -17421 -18063 -17324 -18033
rect -17395 -18129 -17324 -18063
rect -15519 -17919 -15489 -17893
rect -17703 -18159 -17677 -18129
rect -17421 -18159 -17324 -18129
rect -15965 -18150 -15935 -18119
rect -15869 -18150 -15839 -18119
rect -15773 -18150 -15743 -18119
rect -15519 -18149 -15489 -18119
rect -17395 -18225 -17324 -18159
rect -15983 -18166 -15725 -18150
rect -15983 -18200 -15967 -18166
rect -15741 -18200 -15725 -18166
rect -15983 -18216 -15725 -18200
rect -15537 -18166 -15471 -18149
rect -15537 -18200 -15521 -18166
rect -15487 -18200 -15471 -18166
rect -15537 -18216 -15471 -18200
rect -11733 -17059 -11296 -16997
rect -12345 -17089 -12314 -17059
rect -11764 -17089 -11274 -17059
rect -11144 -17089 -11118 -17059
rect -11733 -17155 -11296 -17089
rect -12345 -17185 -12314 -17155
rect -11764 -17184 -11274 -17155
rect -11764 -17185 -11576 -17184
rect -11733 -17249 -11576 -17185
rect -11521 -17185 -11274 -17184
rect -11144 -17185 -11118 -17155
rect -11521 -17249 -11296 -17185
rect -11733 -17251 -11296 -17249
rect -12345 -17281 -12314 -17251
rect -11764 -17281 -11274 -17251
rect -11144 -17281 -11118 -17251
rect -12345 -17377 -12314 -17347
rect -11764 -17366 -11640 -17347
rect -11764 -17377 -11700 -17366
rect -11733 -17443 -11700 -17377
rect -12345 -17473 -12314 -17443
rect -11764 -17473 -11700 -17443
rect -11733 -17496 -11700 -17473
rect -11655 -17496 -11640 -17366
rect -11733 -17539 -11640 -17496
rect -12345 -17569 -12314 -17539
rect -11764 -17569 -11640 -17539
rect -11583 -17377 -11274 -17347
rect -11144 -17377 -11118 -17347
rect -11583 -17443 -11296 -17377
rect -11583 -17473 -11274 -17443
rect -11144 -17473 -11118 -17443
rect -11583 -17539 -11296 -17473
rect -11583 -17569 -11274 -17539
rect -11144 -17569 -11118 -17539
rect -12345 -17665 -12314 -17635
rect -11764 -17665 -11641 -17635
rect -11734 -17697 -11641 -17665
rect -11734 -17731 -11705 -17697
rect -12345 -17761 -12314 -17731
rect -11764 -17761 -11705 -17731
rect -11734 -17827 -11705 -17761
rect -11660 -17827 -11641 -17697
rect -12345 -17857 -12314 -17827
rect -11764 -17857 -11641 -17827
rect -11583 -17921 -11474 -17569
rect -11404 -17665 -11274 -17635
rect -11144 -17665 -11118 -17635
rect -11404 -17689 -11296 -17665
rect -11404 -17819 -11376 -17689
rect -11331 -17731 -11296 -17689
rect -11331 -17761 -11274 -17731
rect -11144 -17761 -11118 -17731
rect -11331 -17819 -11296 -17761
rect -11404 -17827 -11296 -17819
rect -11404 -17857 -11274 -17827
rect -11144 -17857 -11118 -17827
rect -11733 -17923 -11474 -17921
rect -12345 -17953 -12314 -17923
rect -11764 -17953 -11474 -17923
rect -11733 -18019 -11474 -17953
rect -12345 -18049 -12314 -18019
rect -11764 -18049 -11474 -18019
rect -11733 -18115 -11474 -18049
rect -12345 -18145 -12314 -18115
rect -11764 -18145 -11474 -18115
rect -11409 -17953 -11274 -17923
rect -11144 -17953 -11118 -17923
rect -11409 -17972 -11296 -17953
rect -11409 -18102 -11384 -17972
rect -11339 -18019 -11296 -17972
rect -11339 -18049 -11274 -18019
rect -11144 -18049 -11118 -18019
rect -11339 -18102 -11296 -18049
rect -11409 -18115 -11296 -18102
rect -11409 -18145 -11274 -18115
rect -11144 -18145 -11118 -18115
rect -11733 -18194 -11474 -18145
rect -11733 -18207 -11299 -18194
rect -7671 -16840 -7641 -16814
rect -4766 -16900 -4736 -16874
rect -4670 -16900 -4640 -16874
rect -4574 -16900 -4544 -16874
rect -4320 -16886 -4290 -16860
rect -1604 -16668 -1574 -16642
rect -2050 -16899 -2020 -16868
rect -1954 -16899 -1924 -16868
rect -1858 -16899 -1828 -16868
rect -1604 -16898 -1574 -16868
rect -2068 -16915 -1810 -16899
rect -2068 -16949 -2052 -16915
rect -1826 -16949 -1810 -16915
rect -2068 -16965 -1810 -16949
rect -1622 -16915 -1556 -16898
rect -1622 -16949 -1606 -16915
rect -1572 -16949 -1556 -16915
rect -1622 -16965 -1556 -16949
rect -4784 -17019 -4526 -17003
rect -8117 -17071 -8087 -17040
rect -8021 -17071 -7991 -17040
rect -7925 -17071 -7895 -17040
rect -7671 -17070 -7641 -17040
rect -4784 -17053 -4768 -17019
rect -4542 -17053 -4526 -17019
rect -4784 -17069 -4526 -17053
rect -4338 -17019 -4272 -17003
rect -4338 -17053 -4322 -17019
rect -4288 -17053 -4272 -17019
rect -8135 -17087 -7877 -17071
rect -8135 -17121 -8119 -17087
rect -7893 -17121 -7877 -17087
rect -8135 -17137 -7877 -17121
rect -7689 -17087 -7623 -17070
rect -7689 -17121 -7673 -17087
rect -7639 -17121 -7623 -17087
rect -4766 -17100 -4736 -17069
rect -4670 -17100 -4640 -17069
rect -4574 -17100 -4544 -17069
rect -4338 -17070 -4272 -17053
rect -4320 -17100 -4290 -17070
rect -2050 -17094 -2020 -17068
rect -1954 -17094 -1924 -17068
rect -1858 -17094 -1828 -17068
rect -7689 -17137 -7623 -17121
rect -8117 -17306 -8087 -17280
rect -8021 -17306 -7991 -17280
rect -7925 -17306 -7895 -17280
rect -7671 -17320 -7641 -17294
rect -4766 -17340 -4736 -17314
rect -4670 -17340 -4640 -17314
rect -4574 -17340 -4544 -17314
rect -4320 -17326 -4290 -17300
rect -1604 -17108 -1574 -17082
rect -2050 -17339 -2020 -17308
rect -1954 -17339 -1924 -17308
rect -1858 -17339 -1828 -17308
rect -1604 -17338 -1574 -17308
rect -2068 -17355 -1810 -17339
rect -4784 -17398 -4526 -17382
rect -4784 -17432 -4768 -17398
rect -4542 -17432 -4526 -17398
rect -4784 -17448 -4526 -17432
rect -4338 -17398 -4272 -17382
rect -4338 -17432 -4322 -17398
rect -4288 -17432 -4272 -17398
rect -2068 -17389 -2052 -17355
rect -1826 -17389 -1810 -17355
rect -2068 -17405 -1810 -17389
rect -1622 -17355 -1556 -17338
rect 11164 -16550 11194 -16524
rect 11260 -16550 11290 -16524
rect 11356 -16550 11386 -16524
rect 11452 -16550 11482 -16524
rect -1622 -17389 -1606 -17355
rect -1572 -17389 -1556 -17355
rect 7422 -17383 7452 -17350
rect -1622 -17405 -1556 -17389
rect -4766 -17479 -4736 -17448
rect -4670 -17479 -4640 -17448
rect -4574 -17479 -4544 -17448
rect -4338 -17449 -4272 -17432
rect 7238 -17413 7452 -17383
rect -4320 -17479 -4290 -17449
rect -2050 -17473 -2020 -17447
rect -1954 -17473 -1924 -17447
rect -1858 -17473 -1828 -17447
rect -8117 -17551 -8087 -17520
rect -8021 -17551 -7991 -17520
rect -7925 -17551 -7895 -17520
rect -7671 -17550 -7641 -17520
rect -8135 -17567 -7877 -17551
rect -8135 -17601 -8119 -17567
rect -7893 -17601 -7877 -17567
rect -8135 -17617 -7877 -17601
rect -7689 -17567 -7623 -17550
rect -7689 -17601 -7673 -17567
rect -7639 -17601 -7623 -17567
rect -7689 -17617 -7623 -17601
rect -4766 -17719 -4736 -17693
rect -4670 -17719 -4640 -17693
rect -4574 -17719 -4544 -17693
rect -4320 -17705 -4290 -17679
rect -1604 -17487 -1574 -17461
rect 7238 -17660 7268 -17413
rect 7518 -17455 7548 -17350
rect 7614 -17373 7644 -17350
rect 7374 -17593 7548 -17455
rect 7182 -17676 7326 -17660
rect -2050 -17718 -2020 -17687
rect -1954 -17718 -1924 -17687
rect -1858 -17718 -1828 -17687
rect -1604 -17717 -1574 -17687
rect 7182 -17710 7198 -17676
rect 7232 -17710 7326 -17676
rect -2068 -17734 -1810 -17718
rect -8117 -17766 -8087 -17740
rect -8021 -17766 -7991 -17740
rect -7925 -17766 -7895 -17740
rect -7671 -17780 -7641 -17754
rect -2068 -17768 -2052 -17734
rect -1826 -17768 -1810 -17734
rect -2068 -17784 -1810 -17768
rect -1622 -17734 -1556 -17717
rect 7182 -17726 7326 -17710
rect 7374 -17676 7518 -17593
rect 7590 -17635 7644 -17373
rect 7710 -17500 7740 -17350
rect 8370 -17383 8400 -17350
rect 8186 -17413 8400 -17383
rect 7710 -17530 7848 -17500
rect 7584 -17660 7644 -17635
rect 7758 -17660 7848 -17530
rect 8186 -17660 8216 -17413
rect 8466 -17455 8496 -17350
rect 8562 -17373 8592 -17350
rect 8322 -17593 8496 -17455
rect 7374 -17710 7390 -17676
rect 7424 -17710 7518 -17676
rect 7374 -17726 7518 -17710
rect 7566 -17676 7710 -17660
rect 7566 -17710 7582 -17676
rect 7616 -17710 7710 -17676
rect 7566 -17726 7710 -17710
rect 7758 -17676 7902 -17660
rect 7758 -17710 7774 -17676
rect 7808 -17710 7902 -17676
rect 7758 -17726 7902 -17710
rect 8130 -17676 8274 -17660
rect 8130 -17710 8146 -17676
rect 8180 -17710 8274 -17676
rect 8130 -17726 8274 -17710
rect 8322 -17676 8466 -17593
rect 8538 -17635 8592 -17373
rect 8658 -17500 8688 -17350
rect 9306 -17383 9336 -17350
rect 9122 -17413 9336 -17383
rect 8658 -17530 8796 -17500
rect 8532 -17660 8592 -17635
rect 8706 -17660 8796 -17530
rect 9122 -17660 9152 -17413
rect 9402 -17455 9432 -17350
rect 9498 -17373 9528 -17350
rect 9258 -17593 9432 -17455
rect 8322 -17710 8338 -17676
rect 8372 -17710 8466 -17676
rect 8322 -17726 8466 -17710
rect 8514 -17676 8658 -17660
rect 8514 -17710 8530 -17676
rect 8564 -17710 8658 -17676
rect 8514 -17726 8658 -17710
rect 8706 -17676 8850 -17660
rect 8706 -17710 8722 -17676
rect 8756 -17710 8850 -17676
rect 8706 -17726 8850 -17710
rect 9066 -17676 9210 -17660
rect 9066 -17710 9082 -17676
rect 9116 -17710 9210 -17676
rect 9066 -17726 9210 -17710
rect 9258 -17676 9402 -17593
rect 9474 -17635 9528 -17373
rect 9594 -17500 9624 -17350
rect 10237 -17382 10267 -17349
rect 10053 -17412 10267 -17382
rect 9594 -17530 9732 -17500
rect 9468 -17660 9528 -17635
rect 9642 -17660 9732 -17530
rect 10053 -17659 10083 -17412
rect 10333 -17454 10363 -17349
rect 10429 -17372 10459 -17349
rect 10189 -17592 10363 -17454
rect 9258 -17710 9274 -17676
rect 9308 -17710 9402 -17676
rect 9258 -17726 9402 -17710
rect 9450 -17676 9594 -17660
rect 9450 -17710 9466 -17676
rect 9500 -17710 9594 -17676
rect 9450 -17726 9594 -17710
rect 9642 -17676 9786 -17660
rect 9642 -17710 9658 -17676
rect 9692 -17710 9786 -17676
rect 9642 -17726 9786 -17710
rect 9997 -17675 10141 -17659
rect 9997 -17709 10013 -17675
rect 10047 -17709 10141 -17675
rect 9997 -17725 10141 -17709
rect 10189 -17675 10333 -17592
rect 10405 -17634 10459 -17372
rect 10525 -17499 10555 -17349
rect 12219 -16592 12249 -16456
rect 12315 -16385 12345 -16359
rect 12411 -16385 12441 -16359
rect 12507 -16385 12537 -16359
rect 12603 -16385 12633 -16359
rect 12699 -16385 12729 -16359
rect 12315 -16456 12729 -16385
rect 12315 -16498 12345 -16456
rect 12826 -16493 12842 -16267
rect 12876 -16269 12892 -16267
rect 12876 -16299 12923 -16269
rect 13137 -16299 13163 -16269
rect 12876 -16365 12892 -16299
rect 12876 -16395 12923 -16365
rect 13137 -16395 13163 -16365
rect 12876 -16461 12892 -16395
rect 12876 -16491 12923 -16461
rect 13137 -16491 13163 -16461
rect 12876 -16493 12892 -16491
rect 12297 -16514 12363 -16498
rect 12826 -16509 12892 -16493
rect 12297 -16548 12313 -16514
rect 12347 -16548 12363 -16514
rect 12297 -16564 12363 -16548
rect 12315 -16592 12345 -16564
rect 12826 -16713 12893 -16697
rect 12826 -16747 12842 -16713
rect 12876 -16715 12893 -16713
rect 12876 -16745 12923 -16715
rect 13123 -16745 13149 -16715
rect 12876 -16747 12893 -16745
rect 12826 -16763 12893 -16747
rect 12219 -16818 12249 -16792
rect 12315 -16818 12345 -16792
rect 16209 -17049 16239 -17023
rect 16305 -17049 16335 -17023
rect 16401 -17049 16431 -17023
rect 16497 -17049 16527 -17023
rect 16209 -17264 16239 -17249
rect 16017 -17294 16239 -17264
rect 11164 -17383 11194 -17350
rect 10980 -17413 11194 -17383
rect 10525 -17529 10663 -17499
rect 10399 -17659 10459 -17634
rect 10573 -17659 10663 -17529
rect 10189 -17709 10205 -17675
rect 10239 -17709 10333 -17675
rect 10189 -17725 10333 -17709
rect 10381 -17675 10525 -17659
rect 10381 -17709 10397 -17675
rect 10431 -17709 10525 -17675
rect 10381 -17725 10525 -17709
rect 10573 -17675 10717 -17659
rect 10980 -17660 11010 -17413
rect 11260 -17455 11290 -17350
rect 11356 -17373 11386 -17350
rect 11116 -17593 11290 -17455
rect 10573 -17709 10589 -17675
rect 10623 -17709 10717 -17675
rect 10573 -17725 10717 -17709
rect -1622 -17768 -1606 -17734
rect -1572 -17768 -1556 -17734
rect 7200 -17757 7230 -17726
rect 7296 -17757 7326 -17726
rect 7392 -17757 7422 -17726
rect 7488 -17757 7518 -17726
rect 7584 -17757 7614 -17726
rect 7680 -17757 7710 -17726
rect 7776 -17757 7806 -17726
rect 7872 -17757 7902 -17726
rect 8148 -17757 8178 -17726
rect 8244 -17757 8274 -17726
rect 8340 -17757 8370 -17726
rect 8436 -17757 8466 -17726
rect 8532 -17757 8562 -17726
rect 8628 -17757 8658 -17726
rect 8724 -17757 8754 -17726
rect 8820 -17757 8850 -17726
rect 9084 -17757 9114 -17726
rect 9180 -17757 9210 -17726
rect 9276 -17757 9306 -17726
rect 9372 -17757 9402 -17726
rect 9468 -17757 9498 -17726
rect 9564 -17757 9594 -17726
rect 9660 -17757 9690 -17726
rect 9756 -17757 9786 -17726
rect 10015 -17756 10045 -17725
rect 10111 -17756 10141 -17725
rect 10207 -17756 10237 -17725
rect 10303 -17756 10333 -17725
rect 10399 -17756 10429 -17725
rect 10495 -17756 10525 -17725
rect 10591 -17756 10621 -17725
rect 10687 -17756 10717 -17725
rect 10924 -17676 11068 -17660
rect 10924 -17710 10940 -17676
rect 10974 -17710 11068 -17676
rect 10924 -17726 11068 -17710
rect 11116 -17676 11260 -17593
rect 11332 -17635 11386 -17373
rect 11452 -17500 11482 -17350
rect 11452 -17530 11590 -17500
rect 11326 -17660 11386 -17635
rect 11500 -17660 11590 -17530
rect 16017 -17570 16047 -17294
rect 16305 -17570 16335 -17249
rect 15981 -17586 16047 -17570
rect 15981 -17611 15997 -17586
rect 15825 -17620 15997 -17611
rect 16031 -17620 16047 -17586
rect 16269 -17586 16335 -17570
rect 16269 -17611 16285 -17586
rect 15825 -17641 16047 -17620
rect 11116 -17710 11132 -17676
rect 11166 -17710 11260 -17676
rect 11116 -17726 11260 -17710
rect 11308 -17676 11452 -17660
rect 11308 -17710 11324 -17676
rect 11358 -17710 11452 -17676
rect 11308 -17726 11452 -17710
rect 11500 -17676 11644 -17660
rect 15825 -17667 15855 -17641
rect 15921 -17667 15951 -17641
rect 16017 -17667 16047 -17641
rect 16113 -17620 16285 -17611
rect 16319 -17620 16335 -17586
rect 16113 -17641 16335 -17620
rect 16113 -17667 16143 -17641
rect 16209 -17667 16239 -17641
rect 16305 -17667 16335 -17641
rect 16401 -17570 16431 -17249
rect 16497 -17287 16527 -17249
rect 16497 -17304 16719 -17287
rect 16497 -17317 16669 -17304
rect 16653 -17338 16669 -17317
rect 16703 -17338 16719 -17304
rect 16653 -17354 16719 -17338
rect 16401 -17586 16467 -17570
rect 16401 -17620 16417 -17586
rect 16451 -17611 16467 -17586
rect 16689 -17611 16719 -17354
rect 16451 -17620 16623 -17611
rect 16401 -17641 16623 -17620
rect 16401 -17667 16431 -17641
rect 16497 -17667 16527 -17641
rect 16593 -17667 16623 -17641
rect 16689 -17641 16911 -17611
rect 16689 -17667 16719 -17641
rect 16785 -17667 16815 -17641
rect 16881 -17667 16911 -17641
rect 11500 -17710 11516 -17676
rect 11550 -17710 11644 -17676
rect 11500 -17726 11644 -17710
rect -1622 -17784 -1556 -17768
rect -4784 -17838 -4526 -17822
rect -4784 -17872 -4768 -17838
rect -4542 -17872 -4526 -17838
rect -4784 -17888 -4526 -17872
rect -4338 -17838 -4272 -17822
rect -4338 -17872 -4322 -17838
rect -4288 -17872 -4272 -17838
rect -4766 -17919 -4736 -17888
rect -4670 -17919 -4640 -17888
rect -4574 -17919 -4544 -17888
rect -4338 -17889 -4272 -17872
rect -4320 -17919 -4290 -17889
rect -2050 -17913 -2020 -17887
rect -1954 -17913 -1924 -17887
rect -1858 -17913 -1828 -17887
rect -8117 -18011 -8087 -17980
rect -8021 -18011 -7991 -17980
rect -7925 -18011 -7895 -17980
rect -7671 -18010 -7641 -17980
rect -8135 -18027 -7877 -18011
rect -8135 -18061 -8119 -18027
rect -7893 -18061 -7877 -18027
rect -8135 -18077 -7877 -18061
rect -7689 -18027 -7623 -18010
rect -7689 -18061 -7673 -18027
rect -7639 -18061 -7623 -18027
rect -7689 -18077 -7623 -18061
rect -4766 -18159 -4736 -18133
rect -4670 -18159 -4640 -18133
rect -4574 -18159 -4544 -18133
rect -4320 -18145 -4290 -18119
rect -1604 -17927 -1574 -17901
rect 10942 -17757 10972 -17726
rect 11038 -17757 11068 -17726
rect 11134 -17757 11164 -17726
rect 11230 -17757 11260 -17726
rect 11326 -17757 11356 -17726
rect 11422 -17757 11452 -17726
rect 11518 -17757 11548 -17726
rect 11614 -17757 11644 -17726
rect 7200 -18105 7230 -18079
rect 7296 -18105 7326 -18079
rect 7392 -18105 7422 -18079
rect 7488 -18105 7518 -18079
rect 7584 -18105 7614 -18079
rect 7680 -18105 7710 -18079
rect 7776 -18105 7806 -18079
rect 7872 -18105 7902 -18079
rect 8148 -18105 8178 -18079
rect 8244 -18105 8274 -18079
rect 8340 -18105 8370 -18079
rect 8436 -18105 8466 -18079
rect 8532 -18105 8562 -18079
rect 8628 -18105 8658 -18079
rect 8724 -18105 8754 -18079
rect 8820 -18105 8850 -18079
rect 9084 -18105 9114 -18079
rect 9180 -18105 9210 -18079
rect 9276 -18105 9306 -18079
rect 9372 -18105 9402 -18079
rect 9468 -18105 9498 -18079
rect 9564 -18105 9594 -18079
rect 9660 -18105 9690 -18079
rect 9756 -18105 9786 -18079
rect 10015 -18104 10045 -18078
rect 10111 -18104 10141 -18078
rect 10207 -18104 10237 -18078
rect 10303 -18104 10333 -18078
rect 10399 -18104 10429 -18078
rect 10495 -18104 10525 -18078
rect 10591 -18104 10621 -18078
rect 10687 -18104 10717 -18078
rect 10942 -18105 10972 -18079
rect 11038 -18105 11068 -18079
rect 11134 -18105 11164 -18079
rect 11230 -18105 11260 -18079
rect 11326 -18105 11356 -18079
rect 11422 -18105 11452 -18079
rect 11518 -18105 11548 -18079
rect 11614 -18105 11644 -18079
rect -2050 -18158 -2020 -18127
rect -1954 -18158 -1924 -18127
rect -1858 -18158 -1828 -18127
rect -1604 -18157 -1574 -18127
rect -2068 -18174 -1810 -18158
rect -17703 -18255 -17677 -18225
rect -17421 -18255 -17324 -18225
rect -12340 -18237 -12314 -18207
rect -11764 -18237 -11274 -18207
rect -11144 -18237 -11118 -18207
rect -8131 -18226 -8101 -18200
rect -8035 -18226 -8005 -18200
rect -7939 -18226 -7909 -18200
rect -11733 -18270 -11299 -18237
rect -21128 -18345 -21062 -18329
rect -11583 -18331 -11474 -18270
rect -15964 -18405 -15934 -18379
rect -15868 -18405 -15838 -18379
rect -15772 -18405 -15742 -18379
rect -24022 -18433 -23992 -18407
rect -23926 -18433 -23896 -18407
rect -24459 -18525 -24428 -18495
rect -24214 -18525 -24158 -18495
rect -24188 -18591 -24158 -18525
rect -24459 -18621 -24428 -18591
rect -24214 -18621 -24158 -18591
rect -24188 -18650 -24158 -18621
rect -24188 -18666 -24121 -18650
rect -24188 -18687 -24167 -18666
rect -24459 -18717 -24428 -18687
rect -24214 -18700 -24167 -18687
rect -24132 -18700 -24121 -18666
rect -24214 -18717 -24121 -18700
rect -24459 -18813 -24428 -18783
rect -24214 -18813 -24158 -18783
rect -24188 -18879 -24158 -18813
rect -21555 -18534 -21525 -18508
rect -21459 -18534 -21429 -18508
rect -21363 -18534 -21333 -18508
rect -21109 -18548 -21079 -18522
rect -15518 -18419 -15488 -18393
rect -11577 -18413 -11479 -18331
rect -11577 -18467 -11555 -18413
rect -11501 -18467 -11479 -18413
rect -7685 -18240 -7655 -18214
rect -4784 -18217 -4526 -18201
rect -4784 -18251 -4768 -18217
rect -4542 -18251 -4526 -18217
rect -4784 -18267 -4526 -18251
rect -4338 -18217 -4272 -18201
rect -4338 -18251 -4322 -18217
rect -4288 -18251 -4272 -18217
rect -2068 -18208 -2052 -18174
rect -1826 -18208 -1810 -18174
rect -2068 -18224 -1810 -18208
rect -1622 -18174 -1556 -18157
rect -1622 -18208 -1606 -18174
rect -1572 -18208 -1556 -18174
rect -1622 -18224 -1556 -18208
rect -4766 -18298 -4736 -18267
rect -4670 -18298 -4640 -18267
rect -4574 -18298 -4544 -18267
rect -4338 -18268 -4272 -18251
rect -4320 -18298 -4290 -18268
rect -2050 -18292 -2020 -18266
rect -1954 -18292 -1924 -18266
rect -1858 -18292 -1828 -18266
rect -11577 -18483 -11479 -18467
rect -8131 -18471 -8101 -18440
rect -8035 -18471 -8005 -18440
rect -7939 -18471 -7909 -18440
rect -7685 -18470 -7655 -18440
rect -8149 -18487 -7891 -18471
rect -8149 -18521 -8133 -18487
rect -7907 -18521 -7891 -18487
rect -8149 -18537 -7891 -18521
rect -7703 -18487 -7637 -18470
rect -7703 -18521 -7687 -18487
rect -7653 -18521 -7637 -18487
rect -7703 -18537 -7637 -18521
rect -4766 -18538 -4736 -18512
rect -4670 -18538 -4640 -18512
rect -4574 -18538 -4544 -18512
rect -4320 -18524 -4290 -18498
rect -1604 -18306 -1574 -18280
rect -2050 -18537 -2020 -18506
rect -1954 -18537 -1924 -18506
rect -1858 -18537 -1828 -18506
rect -1604 -18536 -1574 -18506
rect 17356 -18275 17386 -18244
rect 17452 -18275 17482 -18244
rect 17548 -18275 17578 -18244
rect 17644 -18275 17674 -18244
rect 17740 -18275 17770 -18244
rect 17836 -18275 17866 -18244
rect 17999 -18307 18065 -18291
rect 17356 -18515 17386 -18489
rect 17452 -18515 17482 -18489
rect 17548 -18515 17578 -18489
rect -2068 -18553 -1810 -18537
rect -2068 -18587 -2052 -18553
rect -1826 -18587 -1810 -18553
rect -2068 -18603 -1810 -18587
rect -1622 -18553 -1556 -18536
rect -1622 -18587 -1606 -18553
rect -1572 -18587 -1556 -18553
rect -1622 -18603 -1556 -18587
rect -15964 -18650 -15934 -18619
rect -15868 -18650 -15838 -18619
rect -15772 -18650 -15742 -18619
rect -15518 -18649 -15488 -18619
rect -15982 -18666 -15724 -18650
rect -15982 -18700 -15966 -18666
rect -15740 -18700 -15724 -18666
rect -15982 -18716 -15724 -18700
rect -15536 -18666 -15470 -18649
rect -15536 -18700 -15520 -18666
rect -15486 -18700 -15470 -18666
rect -4784 -18657 -4526 -18641
rect -15536 -18716 -15470 -18700
rect -8129 -18706 -8099 -18680
rect -8033 -18706 -8003 -18680
rect -7937 -18706 -7907 -18680
rect -4784 -18691 -4768 -18657
rect -4542 -18691 -4526 -18657
rect -21555 -18779 -21525 -18748
rect -21459 -18779 -21429 -18748
rect -21363 -18779 -21333 -18748
rect -21109 -18778 -21079 -18748
rect -21573 -18795 -21315 -18779
rect -21573 -18829 -21557 -18795
rect -21331 -18829 -21315 -18795
rect -24022 -18855 -23992 -18833
rect -24459 -18909 -24428 -18879
rect -24214 -18909 -24158 -18879
rect -24188 -18939 -24158 -18909
rect -24059 -18871 -23992 -18855
rect -24059 -18905 -24043 -18871
rect -24008 -18905 -23992 -18871
rect -24059 -18921 -23992 -18905
rect -23926 -18855 -23896 -18833
rect -21573 -18845 -21315 -18829
rect -21127 -18795 -21061 -18778
rect -17703 -18791 -17677 -18761
rect -17421 -18791 -17324 -18761
rect -21127 -18829 -21111 -18795
rect -21077 -18829 -21061 -18795
rect -21127 -18845 -21061 -18829
rect -23926 -18871 -23859 -18855
rect -17395 -18857 -17324 -18791
rect -23926 -18905 -23910 -18871
rect -23875 -18905 -23859 -18871
rect -17703 -18887 -17677 -18857
rect -17421 -18887 -17324 -18857
rect -15965 -18885 -15935 -18859
rect -15869 -18885 -15839 -18859
rect -15773 -18885 -15743 -18859
rect -24188 -18955 -24121 -18939
rect -24188 -18975 -24167 -18955
rect -24459 -19005 -24428 -18975
rect -24214 -18989 -24167 -18975
rect -24132 -18963 -24121 -18955
rect -23926 -18963 -23859 -18905
rect -17395 -18953 -17324 -18887
rect -24132 -18989 -23859 -18963
rect -17703 -18983 -17677 -18953
rect -17421 -18983 -17324 -18953
rect -24214 -19005 -23859 -18989
rect -24188 -19006 -23859 -19005
rect -21556 -19014 -21526 -18988
rect -21460 -19014 -21430 -18988
rect -21364 -19014 -21334 -18988
rect -21110 -19028 -21080 -19002
rect -17395 -19049 -17324 -18983
rect -17703 -19079 -17677 -19049
rect -17421 -19079 -17324 -19049
rect -17395 -19145 -17324 -19079
rect -17282 -19143 -17216 -19127
rect -17282 -19145 -17266 -19143
rect -17703 -19175 -17677 -19145
rect -17421 -19175 -17266 -19145
rect -17282 -19177 -17266 -19175
rect -17232 -19145 -17216 -19143
rect -15519 -18899 -15489 -18873
rect -7683 -18720 -7653 -18694
rect -4784 -18707 -4526 -18691
rect -4338 -18657 -4272 -18641
rect 15825 -18549 15855 -18523
rect 15921 -18549 15951 -18523
rect 16017 -18549 16047 -18523
rect 16113 -18549 16143 -18523
rect 16209 -18549 16239 -18523
rect 16305 -18549 16335 -18523
rect 16401 -18549 16431 -18523
rect 16497 -18549 16527 -18523
rect 16593 -18549 16623 -18523
rect 16689 -18549 16719 -18523
rect 16785 -18549 16815 -18523
rect 16881 -18549 16911 -18523
rect 17355 -18536 17578 -18515
rect 17355 -18571 17372 -18536
rect 17406 -18545 17578 -18536
rect 17644 -18515 17674 -18489
rect 17740 -18515 17770 -18489
rect 17836 -18515 17866 -18489
rect 17644 -18536 17866 -18515
rect 17406 -18571 17422 -18545
rect 17355 -18582 17422 -18571
rect 17644 -18571 17661 -18536
rect 17695 -18545 17866 -18536
rect 17999 -18533 18015 -18307
rect 18049 -18309 18065 -18307
rect 18049 -18339 18096 -18309
rect 18310 -18339 18336 -18309
rect 18049 -18405 18065 -18339
rect 18049 -18435 18096 -18405
rect 18310 -18435 18336 -18405
rect 18049 -18501 18065 -18435
rect 18049 -18531 18096 -18501
rect 18310 -18531 18336 -18501
rect 18049 -18533 18065 -18531
rect 17695 -18571 17711 -18545
rect 17999 -18549 18065 -18533
rect 17644 -18582 17711 -18571
rect 15825 -18649 15855 -18623
rect 15921 -18649 15951 -18623
rect 16017 -18649 16047 -18623
rect 16113 -18649 16143 -18623
rect 16209 -18649 16239 -18623
rect 16305 -18649 16335 -18623
rect 16401 -18649 16431 -18623
rect 16497 -18649 16527 -18623
rect 16593 -18649 16623 -18623
rect 16689 -18649 16719 -18623
rect 16785 -18649 16815 -18623
rect 16881 -18649 16911 -18623
rect -4338 -18691 -4322 -18657
rect -4288 -18691 -4272 -18657
rect -4766 -18738 -4736 -18707
rect -4670 -18738 -4640 -18707
rect -4574 -18738 -4544 -18707
rect -4338 -18708 -4272 -18691
rect -4320 -18738 -4290 -18708
rect -2050 -18732 -2020 -18706
rect -1954 -18732 -1924 -18706
rect -1858 -18732 -1828 -18706
rect -8129 -18951 -8099 -18920
rect -8033 -18951 -8003 -18920
rect -7937 -18951 -7907 -18920
rect -7683 -18950 -7653 -18920
rect -8147 -18967 -7889 -18951
rect -8147 -19001 -8131 -18967
rect -7905 -19001 -7889 -18967
rect -8147 -19017 -7889 -19001
rect -7701 -18967 -7635 -18950
rect -7701 -19001 -7685 -18967
rect -7651 -19001 -7635 -18967
rect -4766 -18978 -4736 -18952
rect -4670 -18978 -4640 -18952
rect -4574 -18978 -4544 -18952
rect -4320 -18964 -4290 -18938
rect -1604 -18746 -1574 -18720
rect 5561 -18777 5627 -18761
rect -2050 -18977 -2020 -18946
rect -1954 -18977 -1924 -18946
rect -1858 -18977 -1828 -18946
rect -1604 -18976 -1574 -18946
rect -7701 -19017 -7635 -19001
rect -2068 -18993 -1810 -18977
rect -4784 -19036 -4526 -19020
rect -4784 -19070 -4768 -19036
rect -4542 -19070 -4526 -19036
rect -4784 -19086 -4526 -19070
rect -4338 -19036 -4272 -19020
rect -4338 -19070 -4322 -19036
rect -4288 -19070 -4272 -19036
rect -2068 -19027 -2052 -18993
rect -1826 -19027 -1810 -18993
rect -2068 -19043 -1810 -19027
rect -1622 -18993 -1556 -18976
rect -1622 -19027 -1606 -18993
rect -1572 -19027 -1556 -18993
rect 5561 -19003 5577 -18777
rect 5611 -18779 5627 -18777
rect 6001 -18777 6067 -18761
rect 5611 -18809 5658 -18779
rect 5872 -18809 5898 -18779
rect 5611 -18875 5627 -18809
rect 5611 -18905 5658 -18875
rect 5872 -18905 5898 -18875
rect 5611 -18971 5627 -18905
rect 5611 -19001 5658 -18971
rect 5872 -19001 5898 -18971
rect 5611 -19003 5627 -19001
rect 5561 -19019 5627 -19003
rect -1622 -19043 -1556 -19027
rect 6001 -19003 6017 -18777
rect 6051 -18779 6067 -18777
rect 6441 -18777 6507 -18761
rect 6051 -18809 6098 -18779
rect 6312 -18809 6338 -18779
rect 6051 -18875 6067 -18809
rect 6051 -18905 6098 -18875
rect 6312 -18905 6338 -18875
rect 6051 -18971 6067 -18905
rect 6051 -19001 6098 -18971
rect 6312 -19001 6338 -18971
rect 6051 -19003 6067 -19001
rect 6001 -19019 6067 -19003
rect 6441 -19003 6457 -18777
rect 6491 -18779 6507 -18777
rect 6491 -18809 6538 -18779
rect 6752 -18809 6778 -18779
rect 6491 -18875 6507 -18809
rect 6491 -18905 6538 -18875
rect 6752 -18905 6778 -18875
rect 6491 -18971 6507 -18905
rect 6491 -19001 6538 -18971
rect 6752 -19001 6778 -18971
rect 6491 -19003 6507 -19001
rect 6441 -19019 6507 -19003
rect -17232 -19175 -17188 -19145
rect -16988 -19175 -16962 -19145
rect -17232 -19177 -17216 -19175
rect -17282 -19193 -17216 -19177
rect -21556 -19259 -21526 -19228
rect -21460 -19259 -21430 -19228
rect -21364 -19259 -21334 -19228
rect -21110 -19258 -21080 -19228
rect -21574 -19275 -21316 -19259
rect -21574 -19309 -21558 -19275
rect -21332 -19309 -21316 -19275
rect -21574 -19325 -21316 -19309
rect -21128 -19275 -21062 -19258
rect -17703 -19271 -17677 -19241
rect -17421 -19271 -17188 -19241
rect -16988 -19271 -16962 -19241
rect -21128 -19309 -21112 -19275
rect -21078 -19309 -21062 -19275
rect -21128 -19325 -21062 -19309
rect -21556 -19514 -21526 -19488
rect -21460 -19514 -21430 -19488
rect -21364 -19514 -21334 -19488
rect -24020 -19627 -23990 -19601
rect -23924 -19627 -23894 -19601
rect -24457 -19719 -24426 -19689
rect -24212 -19719 -24156 -19689
rect -24186 -19785 -24156 -19719
rect -24457 -19815 -24426 -19785
rect -24212 -19815 -24156 -19785
rect -24186 -19844 -24156 -19815
rect -24186 -19860 -24119 -19844
rect -24186 -19881 -24165 -19860
rect -24457 -19911 -24426 -19881
rect -24212 -19894 -24165 -19881
rect -24130 -19894 -24119 -19860
rect -24212 -19911 -24119 -19894
rect -24457 -20007 -24426 -19977
rect -24212 -20007 -24156 -19977
rect -24186 -20073 -24156 -20007
rect -21110 -19528 -21080 -19502
rect -17395 -19286 -17324 -19271
rect -17395 -19320 -17371 -19286
rect -17337 -19320 -17324 -19286
rect -17395 -19337 -17324 -19320
rect -15965 -19130 -15935 -19099
rect -15869 -19130 -15839 -19099
rect -15773 -19130 -15743 -19099
rect -15519 -19129 -15489 -19099
rect -4766 -19117 -4736 -19086
rect -4670 -19117 -4640 -19086
rect -4574 -19117 -4544 -19086
rect -4338 -19087 -4272 -19070
rect -4320 -19117 -4290 -19087
rect -2050 -19111 -2020 -19085
rect -1954 -19111 -1924 -19085
rect -1858 -19111 -1828 -19085
rect -15983 -19146 -15725 -19130
rect -15983 -19180 -15967 -19146
rect -15741 -19180 -15725 -19146
rect -15983 -19196 -15725 -19180
rect -15537 -19146 -15471 -19129
rect -15537 -19180 -15521 -19146
rect -15487 -19180 -15471 -19146
rect -15537 -19196 -15471 -19180
rect -17703 -19367 -17677 -19337
rect -17421 -19367 -17324 -19337
rect -4766 -19357 -4736 -19331
rect -4670 -19357 -4640 -19331
rect -4574 -19357 -4544 -19331
rect -4320 -19343 -4290 -19317
rect -1604 -19125 -1574 -19099
rect 5561 -19223 5628 -19207
rect 5561 -19257 5577 -19223
rect 5611 -19225 5628 -19223
rect 6001 -19223 6068 -19207
rect 5611 -19255 5658 -19225
rect 5858 -19255 5884 -19225
rect 5611 -19257 5628 -19255
rect 5561 -19273 5628 -19257
rect 6001 -19257 6017 -19223
rect 6051 -19225 6068 -19223
rect 6441 -19223 6508 -19207
rect 6051 -19255 6098 -19225
rect 6298 -19255 6324 -19225
rect 6051 -19257 6068 -19255
rect 6001 -19273 6068 -19257
rect 6441 -19257 6457 -19223
rect 6491 -19225 6508 -19223
rect 6491 -19255 6538 -19225
rect 6738 -19255 6764 -19225
rect 6491 -19257 6508 -19255
rect 6441 -19273 6508 -19257
rect -2050 -19356 -2020 -19325
rect -1954 -19356 -1924 -19325
rect -1858 -19356 -1828 -19325
rect -1604 -19355 -1574 -19325
rect -17395 -19433 -17324 -19367
rect -15965 -19385 -15935 -19359
rect -15869 -19385 -15839 -19359
rect -15773 -19385 -15743 -19359
rect -2068 -19372 -1810 -19356
rect -17703 -19463 -17677 -19433
rect -17421 -19463 -17324 -19433
rect -17395 -19529 -17324 -19463
rect -17703 -19559 -17677 -19529
rect -17421 -19559 -17324 -19529
rect -17395 -19625 -17324 -19559
rect -15519 -19399 -15489 -19373
rect -2068 -19406 -2052 -19372
rect -1826 -19406 -1810 -19372
rect -2068 -19422 -1810 -19406
rect -1622 -19372 -1556 -19355
rect -1622 -19406 -1606 -19372
rect -1572 -19406 -1556 -19372
rect -1622 -19422 -1556 -19406
rect 7200 -19421 7230 -19395
rect 7296 -19421 7326 -19395
rect 7392 -19421 7422 -19395
rect 7488 -19421 7518 -19395
rect 7584 -19421 7614 -19395
rect 7680 -19421 7710 -19395
rect 7776 -19421 7806 -19395
rect 7872 -19421 7902 -19395
rect 8148 -19421 8178 -19395
rect 8244 -19421 8274 -19395
rect 8340 -19421 8370 -19395
rect 8436 -19421 8466 -19395
rect 8532 -19421 8562 -19395
rect 8628 -19421 8658 -19395
rect 8724 -19421 8754 -19395
rect 8820 -19421 8850 -19395
rect 9084 -19421 9114 -19395
rect 9180 -19421 9210 -19395
rect 9276 -19421 9306 -19395
rect 9372 -19421 9402 -19395
rect 9468 -19421 9498 -19395
rect 9564 -19421 9594 -19395
rect 9660 -19421 9690 -19395
rect 9756 -19421 9786 -19395
rect 10015 -19421 10045 -19395
rect 10111 -19421 10141 -19395
rect 10207 -19421 10237 -19395
rect 10303 -19421 10333 -19395
rect 10399 -19421 10429 -19395
rect 10495 -19421 10525 -19395
rect 10591 -19421 10621 -19395
rect 10687 -19421 10717 -19395
rect 10942 -19421 10972 -19395
rect 11038 -19421 11068 -19395
rect 11134 -19421 11164 -19395
rect 11230 -19421 11260 -19395
rect 11326 -19421 11356 -19395
rect 11422 -19421 11452 -19395
rect 11518 -19421 11548 -19395
rect 11614 -19421 11644 -19395
rect -4784 -19476 -4526 -19460
rect -4784 -19510 -4768 -19476
rect -4542 -19510 -4526 -19476
rect -4784 -19526 -4526 -19510
rect -4338 -19476 -4272 -19460
rect -4338 -19510 -4322 -19476
rect -4288 -19510 -4272 -19476
rect -4766 -19557 -4736 -19526
rect -4670 -19557 -4640 -19526
rect -4574 -19557 -4544 -19526
rect -4338 -19527 -4272 -19510
rect -4320 -19557 -4290 -19527
rect -2050 -19551 -2020 -19525
rect -1954 -19551 -1924 -19525
rect -1858 -19551 -1828 -19525
rect -17703 -19655 -17677 -19625
rect -17421 -19655 -17324 -19625
rect -15965 -19630 -15935 -19599
rect -15869 -19630 -15839 -19599
rect -15773 -19630 -15743 -19599
rect -15519 -19629 -15489 -19599
rect -15983 -19646 -15725 -19630
rect -15983 -19680 -15967 -19646
rect -15741 -19680 -15725 -19646
rect -15983 -19696 -15725 -19680
rect -15537 -19646 -15471 -19629
rect -15537 -19680 -15521 -19646
rect -15487 -19680 -15471 -19646
rect -15537 -19696 -15471 -19680
rect -21556 -19759 -21526 -19728
rect -21460 -19759 -21430 -19728
rect -21364 -19759 -21334 -19728
rect -21110 -19758 -21080 -19728
rect -21574 -19775 -21316 -19759
rect -21574 -19809 -21558 -19775
rect -21332 -19809 -21316 -19775
rect -21574 -19825 -21316 -19809
rect -21128 -19775 -21062 -19758
rect -21128 -19809 -21112 -19775
rect -21078 -19809 -21062 -19775
rect -4766 -19797 -4736 -19771
rect -4670 -19797 -4640 -19771
rect -4574 -19797 -4544 -19771
rect -4320 -19783 -4290 -19757
rect -1604 -19565 -1574 -19539
rect 17355 -18777 17398 -18582
rect 17440 -18660 17506 -18644
rect 17440 -18695 17456 -18660
rect 17490 -18681 17506 -18660
rect 17490 -18695 17528 -18681
rect 17440 -18711 17528 -18695
rect 17928 -18711 17954 -18681
rect 17999 -18753 18066 -18737
rect 17355 -18793 17528 -18777
rect 17355 -18828 17456 -18793
rect 17490 -18807 17528 -18793
rect 17928 -18807 17954 -18777
rect 17999 -18787 18015 -18753
rect 18049 -18755 18066 -18753
rect 18049 -18785 18096 -18755
rect 18296 -18785 18322 -18755
rect 18049 -18787 18066 -18785
rect 17999 -18803 18066 -18787
rect 17490 -18828 17506 -18807
rect 17355 -18844 17506 -18828
rect 15825 -19531 15855 -19505
rect 15921 -19531 15951 -19505
rect 16017 -19531 16047 -19505
rect 15825 -19552 16047 -19531
rect 15825 -19561 15997 -19552
rect 15981 -19586 15997 -19561
rect 16031 -19586 16047 -19552
rect 16113 -19531 16143 -19505
rect 16209 -19531 16239 -19505
rect 16305 -19531 16335 -19505
rect 16113 -19552 16335 -19531
rect 16113 -19561 16285 -19552
rect 15981 -19602 16047 -19586
rect 16269 -19586 16285 -19561
rect 16319 -19586 16335 -19552
rect 16269 -19602 16335 -19586
rect -2050 -19796 -2020 -19765
rect -1954 -19796 -1924 -19765
rect -1858 -19796 -1828 -19765
rect -1604 -19795 -1574 -19765
rect 7200 -19774 7230 -19743
rect 7296 -19774 7326 -19743
rect 7392 -19774 7422 -19743
rect 7488 -19774 7518 -19743
rect 7584 -19774 7614 -19743
rect 7680 -19774 7710 -19743
rect 7776 -19774 7806 -19743
rect 7872 -19774 7902 -19743
rect 8148 -19774 8178 -19743
rect 8244 -19774 8274 -19743
rect 8340 -19774 8370 -19743
rect 8436 -19774 8466 -19743
rect 8532 -19774 8562 -19743
rect 8628 -19774 8658 -19743
rect 8724 -19774 8754 -19743
rect 8820 -19774 8850 -19743
rect 9084 -19774 9114 -19743
rect 9180 -19774 9210 -19743
rect 9276 -19774 9306 -19743
rect 9372 -19774 9402 -19743
rect 9468 -19774 9498 -19743
rect 9564 -19774 9594 -19743
rect 9660 -19774 9690 -19743
rect 9756 -19774 9786 -19743
rect 10015 -19774 10045 -19743
rect 10111 -19774 10141 -19743
rect 10207 -19774 10237 -19743
rect 10303 -19774 10333 -19743
rect 10399 -19774 10429 -19743
rect 10495 -19774 10525 -19743
rect 10591 -19774 10621 -19743
rect 10687 -19774 10717 -19743
rect 10942 -19774 10972 -19743
rect 11038 -19774 11068 -19743
rect 11134 -19774 11164 -19743
rect 11230 -19774 11260 -19743
rect 11326 -19774 11356 -19743
rect 11422 -19774 11452 -19743
rect 11518 -19774 11548 -19743
rect 11614 -19774 11644 -19743
rect 7182 -19790 7326 -19774
rect -21128 -19825 -21062 -19809
rect -2068 -19812 -1810 -19796
rect -15965 -19865 -15935 -19839
rect -15869 -19865 -15839 -19839
rect -15773 -19865 -15743 -19839
rect -21556 -19994 -21526 -19968
rect -21460 -19994 -21430 -19968
rect -21364 -19994 -21334 -19968
rect -24020 -20049 -23990 -20027
rect -24457 -20103 -24426 -20073
rect -24212 -20103 -24156 -20073
rect -24186 -20133 -24156 -20103
rect -24057 -20065 -23990 -20049
rect -24057 -20099 -24041 -20065
rect -24006 -20099 -23990 -20065
rect -24057 -20115 -23990 -20099
rect -23924 -20049 -23894 -20027
rect -23924 -20065 -23857 -20049
rect -23924 -20099 -23908 -20065
rect -23873 -20099 -23857 -20065
rect -24186 -20149 -24119 -20133
rect -24186 -20169 -24165 -20149
rect -24457 -20199 -24426 -20169
rect -24212 -20183 -24165 -20169
rect -24130 -20157 -24119 -20149
rect -23924 -20157 -23857 -20099
rect -24130 -20183 -23857 -20157
rect -24212 -20199 -23857 -20183
rect -24186 -20200 -23857 -20199
rect -21110 -20008 -21080 -19982
rect -15519 -19879 -15489 -19853
rect -4784 -19855 -4526 -19839
rect -4784 -19889 -4768 -19855
rect -4542 -19889 -4526 -19855
rect -4784 -19905 -4526 -19889
rect -4338 -19855 -4272 -19839
rect -4338 -19889 -4322 -19855
rect -4288 -19889 -4272 -19855
rect -2068 -19846 -2052 -19812
rect -1826 -19846 -1810 -19812
rect -2068 -19862 -1810 -19846
rect -1622 -19812 -1556 -19795
rect -1622 -19846 -1606 -19812
rect -1572 -19846 -1556 -19812
rect 7182 -19824 7198 -19790
rect 7232 -19824 7326 -19790
rect 7182 -19840 7326 -19824
rect 7374 -19790 7518 -19774
rect 7374 -19824 7390 -19790
rect 7424 -19824 7518 -19790
rect -1622 -19862 -1556 -19846
rect -12340 -19954 -12314 -19924
rect -11764 -19954 -11274 -19924
rect -11144 -19954 -11118 -19924
rect -4766 -19936 -4736 -19905
rect -4670 -19936 -4640 -19905
rect -4574 -19936 -4544 -19905
rect -4338 -19906 -4272 -19889
rect -4320 -19936 -4290 -19906
rect -2050 -19930 -2020 -19904
rect -1954 -19930 -1924 -19904
rect -1858 -19930 -1828 -19904
rect -15965 -20110 -15935 -20079
rect -15869 -20110 -15839 -20079
rect -15773 -20110 -15743 -20079
rect -15519 -20109 -15489 -20079
rect -15983 -20126 -15725 -20110
rect -15983 -20160 -15967 -20126
rect -15741 -20160 -15725 -20126
rect -17703 -20191 -17677 -20161
rect -17421 -20191 -17324 -20161
rect -15983 -20176 -15725 -20160
rect -15537 -20126 -15471 -20109
rect -15537 -20160 -15521 -20126
rect -15487 -20160 -15471 -20126
rect -15537 -20176 -15471 -20160
rect -21556 -20239 -21526 -20208
rect -21460 -20239 -21430 -20208
rect -21364 -20239 -21334 -20208
rect -21110 -20238 -21080 -20208
rect -21574 -20255 -21316 -20239
rect -21574 -20289 -21558 -20255
rect -21332 -20289 -21316 -20255
rect -21574 -20305 -21316 -20289
rect -21128 -20255 -21062 -20238
rect -21128 -20289 -21112 -20255
rect -21078 -20289 -21062 -20255
rect -17395 -20257 -17324 -20191
rect -17703 -20287 -17677 -20257
rect -17421 -20287 -17324 -20257
rect -21128 -20305 -21062 -20289
rect -17395 -20353 -17324 -20287
rect -15965 -20325 -15935 -20299
rect -15869 -20325 -15839 -20299
rect -15773 -20325 -15743 -20299
rect -17703 -20383 -17677 -20353
rect -17421 -20383 -17324 -20353
rect -21556 -20454 -21526 -20428
rect -21460 -20454 -21430 -20428
rect -21364 -20454 -21334 -20428
rect -21110 -20468 -21080 -20442
rect -17395 -20449 -17324 -20383
rect -17703 -20479 -17677 -20449
rect -17421 -20479 -17324 -20449
rect -17395 -20545 -17324 -20479
rect -17282 -20543 -17216 -20527
rect -17282 -20545 -17266 -20543
rect -17703 -20575 -17677 -20545
rect -17421 -20575 -17266 -20545
rect -17282 -20577 -17266 -20575
rect -17232 -20545 -17216 -20543
rect -17232 -20575 -17188 -20545
rect -16988 -20575 -16962 -20545
rect -17232 -20577 -17216 -20575
rect -17282 -20593 -17216 -20577
rect -21556 -20699 -21526 -20668
rect -21460 -20699 -21430 -20668
rect -21364 -20699 -21334 -20668
rect -21110 -20698 -21080 -20668
rect -17703 -20671 -17677 -20641
rect -17421 -20671 -17188 -20641
rect -16988 -20671 -16962 -20641
rect -21574 -20715 -21316 -20699
rect -21574 -20749 -21558 -20715
rect -21332 -20749 -21316 -20715
rect -21574 -20765 -21316 -20749
rect -21128 -20715 -21062 -20698
rect -21128 -20749 -21112 -20715
rect -21078 -20749 -21062 -20715
rect -21128 -20765 -21062 -20749
rect -23989 -20827 -23959 -20801
rect -23893 -20827 -23863 -20801
rect -24426 -20919 -24395 -20889
rect -24181 -20919 -24125 -20889
rect -24155 -20985 -24125 -20919
rect -24426 -21015 -24395 -20985
rect -24181 -21015 -24125 -20985
rect -24155 -21044 -24125 -21015
rect -24155 -21060 -24088 -21044
rect -24155 -21081 -24134 -21060
rect -24426 -21111 -24395 -21081
rect -24181 -21094 -24134 -21081
rect -24099 -21094 -24088 -21060
rect -24181 -21111 -24088 -21094
rect -24426 -21207 -24395 -21177
rect -24181 -21207 -24125 -21177
rect -24155 -21273 -24125 -21207
rect -21570 -20914 -21540 -20888
rect -21474 -20914 -21444 -20888
rect -21378 -20914 -21348 -20888
rect -21124 -20928 -21094 -20902
rect -17395 -20686 -17324 -20671
rect -17395 -20720 -17371 -20686
rect -17337 -20720 -17324 -20686
rect -17395 -20737 -17324 -20720
rect -15519 -20339 -15489 -20313
rect -15965 -20570 -15935 -20539
rect -15869 -20570 -15839 -20539
rect -15773 -20570 -15743 -20539
rect -15519 -20569 -15489 -20539
rect -15983 -20586 -15725 -20570
rect -15983 -20620 -15967 -20586
rect -15741 -20620 -15725 -20586
rect -15983 -20636 -15725 -20620
rect -15537 -20586 -15471 -20569
rect -15537 -20620 -15521 -20586
rect -15487 -20620 -15471 -20586
rect -15537 -20636 -15471 -20620
rect -17703 -20767 -17677 -20737
rect -17421 -20767 -17324 -20737
rect -17395 -20833 -17324 -20767
rect -15979 -20785 -15949 -20759
rect -15883 -20785 -15853 -20759
rect -15787 -20785 -15757 -20759
rect -17703 -20863 -17677 -20833
rect -17421 -20863 -17324 -20833
rect -17395 -20929 -17324 -20863
rect -17703 -20959 -17677 -20929
rect -17421 -20959 -17324 -20929
rect -17395 -21025 -17324 -20959
rect -15533 -20799 -15503 -20773
rect -17703 -21055 -17677 -21025
rect -17421 -21055 -17324 -21025
rect -15979 -21030 -15949 -20999
rect -15883 -21030 -15853 -20999
rect -15787 -21030 -15757 -20999
rect -15533 -21029 -15503 -20999
rect -15997 -21046 -15739 -21030
rect -15997 -21080 -15981 -21046
rect -15755 -21080 -15739 -21046
rect -15997 -21096 -15739 -21080
rect -15551 -21046 -15485 -21029
rect -15551 -21080 -15535 -21046
rect -15501 -21080 -15485 -21046
rect -15551 -21096 -15485 -21080
rect -11733 -20016 -11296 -19954
rect -12345 -20046 -12314 -20016
rect -11764 -20046 -11274 -20016
rect -11144 -20046 -11118 -20016
rect -11733 -20112 -11296 -20046
rect -12345 -20142 -12314 -20112
rect -11764 -20141 -11274 -20112
rect -11764 -20142 -11576 -20141
rect -11733 -20206 -11576 -20142
rect -11521 -20142 -11274 -20141
rect -11144 -20142 -11118 -20112
rect -11521 -20206 -11296 -20142
rect -11733 -20208 -11296 -20206
rect -12345 -20238 -12314 -20208
rect -11764 -20238 -11274 -20208
rect -11144 -20238 -11118 -20208
rect -12345 -20334 -12314 -20304
rect -11764 -20323 -11640 -20304
rect -11764 -20334 -11700 -20323
rect -11733 -20400 -11700 -20334
rect -12345 -20430 -12314 -20400
rect -11764 -20430 -11700 -20400
rect -11733 -20453 -11700 -20430
rect -11655 -20453 -11640 -20323
rect -11733 -20496 -11640 -20453
rect -12345 -20526 -12314 -20496
rect -11764 -20526 -11640 -20496
rect -11583 -20334 -11274 -20304
rect -11144 -20334 -11118 -20304
rect -11583 -20400 -11296 -20334
rect -11583 -20430 -11274 -20400
rect -11144 -20430 -11118 -20400
rect -11583 -20496 -11296 -20430
rect -11583 -20526 -11274 -20496
rect -11144 -20526 -11118 -20496
rect -12345 -20622 -12314 -20592
rect -11764 -20622 -11641 -20592
rect -11734 -20654 -11641 -20622
rect -11734 -20688 -11705 -20654
rect -12345 -20718 -12314 -20688
rect -11764 -20718 -11705 -20688
rect -11734 -20784 -11705 -20718
rect -11660 -20784 -11641 -20654
rect -12345 -20814 -12314 -20784
rect -11764 -20814 -11641 -20784
rect -11583 -20878 -11474 -20526
rect -11404 -20622 -11274 -20592
rect -11144 -20622 -11118 -20592
rect -11404 -20646 -11296 -20622
rect -11404 -20776 -11376 -20646
rect -11331 -20688 -11296 -20646
rect -11331 -20718 -11274 -20688
rect -11144 -20718 -11118 -20688
rect -11331 -20776 -11296 -20718
rect -11404 -20784 -11296 -20776
rect -11404 -20814 -11274 -20784
rect -11144 -20814 -11118 -20784
rect -11733 -20880 -11474 -20878
rect -12345 -20910 -12314 -20880
rect -11764 -20910 -11474 -20880
rect -11733 -20976 -11474 -20910
rect -12345 -21006 -12314 -20976
rect -11764 -21006 -11474 -20976
rect -11733 -21072 -11474 -21006
rect -12345 -21102 -12314 -21072
rect -11764 -21102 -11474 -21072
rect -11409 -20910 -11274 -20880
rect -11144 -20910 -11118 -20880
rect -11409 -20929 -11296 -20910
rect -11409 -21059 -11384 -20929
rect -11339 -20976 -11296 -20929
rect -11339 -21006 -11274 -20976
rect -11144 -21006 -11118 -20976
rect -11339 -21059 -11296 -21006
rect -11409 -21072 -11296 -21059
rect -11409 -21102 -11274 -21072
rect -11144 -21102 -11118 -21072
rect -21570 -21159 -21540 -21128
rect -21474 -21159 -21444 -21128
rect -21378 -21159 -21348 -21128
rect -21124 -21158 -21094 -21128
rect -21588 -21175 -21330 -21159
rect -21588 -21209 -21572 -21175
rect -21346 -21209 -21330 -21175
rect -21588 -21225 -21330 -21209
rect -21142 -21175 -21076 -21158
rect -11733 -21151 -11474 -21102
rect -11733 -21164 -11299 -21151
rect -4766 -20176 -4736 -20150
rect -4670 -20176 -4640 -20150
rect -4574 -20176 -4544 -20150
rect -4320 -20162 -4290 -20136
rect -1604 -19944 -1574 -19918
rect 7238 -20087 7268 -19840
rect 7374 -19907 7518 -19824
rect 7566 -19790 7710 -19774
rect 7566 -19824 7582 -19790
rect 7616 -19824 7710 -19790
rect 7566 -19840 7710 -19824
rect 7758 -19790 7902 -19774
rect 7758 -19824 7774 -19790
rect 7808 -19824 7902 -19790
rect 7758 -19840 7902 -19824
rect 8130 -19790 8274 -19774
rect 8130 -19824 8146 -19790
rect 8180 -19824 8274 -19790
rect 8130 -19840 8274 -19824
rect 8322 -19790 8466 -19774
rect 8322 -19824 8338 -19790
rect 8372 -19824 8466 -19790
rect 7584 -19865 7644 -19840
rect 7374 -20045 7548 -19907
rect 7238 -20117 7452 -20087
rect -2050 -20175 -2020 -20144
rect -1954 -20175 -1924 -20144
rect -1858 -20175 -1828 -20144
rect -1604 -20174 -1574 -20144
rect 7422 -20150 7452 -20117
rect 7518 -20150 7548 -20045
rect 7590 -20127 7644 -19865
rect 7758 -19970 7848 -19840
rect 7614 -20150 7644 -20127
rect 7710 -20000 7848 -19970
rect 7710 -20150 7740 -20000
rect 8186 -20087 8216 -19840
rect 8322 -19907 8466 -19824
rect 8514 -19790 8658 -19774
rect 8514 -19824 8530 -19790
rect 8564 -19824 8658 -19790
rect 8514 -19840 8658 -19824
rect 8706 -19790 8850 -19774
rect 8706 -19824 8722 -19790
rect 8756 -19824 8850 -19790
rect 8706 -19840 8850 -19824
rect 9066 -19790 9210 -19774
rect 9066 -19824 9082 -19790
rect 9116 -19824 9210 -19790
rect 9066 -19840 9210 -19824
rect 9258 -19790 9402 -19774
rect 9258 -19824 9274 -19790
rect 9308 -19824 9402 -19790
rect 8532 -19865 8592 -19840
rect 8322 -20045 8496 -19907
rect 8186 -20117 8400 -20087
rect 8370 -20150 8400 -20117
rect 8466 -20150 8496 -20045
rect 8538 -20127 8592 -19865
rect 8706 -19970 8796 -19840
rect 8562 -20150 8592 -20127
rect 8658 -20000 8796 -19970
rect 8658 -20150 8688 -20000
rect 9122 -20087 9152 -19840
rect 9258 -19907 9402 -19824
rect 9450 -19790 9594 -19774
rect 9450 -19824 9466 -19790
rect 9500 -19824 9594 -19790
rect 9450 -19840 9594 -19824
rect 9642 -19790 9786 -19774
rect 9642 -19824 9658 -19790
rect 9692 -19824 9786 -19790
rect 9642 -19840 9786 -19824
rect 9997 -19790 10141 -19774
rect 9997 -19824 10013 -19790
rect 10047 -19824 10141 -19790
rect 9997 -19840 10141 -19824
rect 10189 -19790 10333 -19774
rect 10189 -19824 10205 -19790
rect 10239 -19824 10333 -19790
rect 9468 -19865 9528 -19840
rect 9258 -20045 9432 -19907
rect 9122 -20117 9336 -20087
rect 9306 -20150 9336 -20117
rect 9402 -20150 9432 -20045
rect 9474 -20127 9528 -19865
rect 9642 -19970 9732 -19840
rect 9498 -20150 9528 -20127
rect 9594 -20000 9732 -19970
rect 9594 -20150 9624 -20000
rect 10053 -20087 10083 -19840
rect 10189 -19907 10333 -19824
rect 10381 -19790 10525 -19774
rect 10381 -19824 10397 -19790
rect 10431 -19824 10525 -19790
rect 10381 -19840 10525 -19824
rect 10573 -19790 10717 -19774
rect 10573 -19824 10589 -19790
rect 10623 -19824 10717 -19790
rect 10573 -19840 10717 -19824
rect 10924 -19790 11068 -19774
rect 10924 -19824 10940 -19790
rect 10974 -19824 11068 -19790
rect 10924 -19840 11068 -19824
rect 11116 -19790 11260 -19774
rect 11116 -19824 11132 -19790
rect 11166 -19824 11260 -19790
rect 10399 -19865 10459 -19840
rect 10189 -20045 10363 -19907
rect 10053 -20117 10267 -20087
rect 10237 -20150 10267 -20117
rect 10333 -20150 10363 -20045
rect 10405 -20127 10459 -19865
rect 10573 -19970 10663 -19840
rect 10429 -20150 10459 -20127
rect 10525 -20000 10663 -19970
rect 10525 -20150 10555 -20000
rect 10980 -20087 11010 -19840
rect 11116 -19907 11260 -19824
rect 11308 -19790 11452 -19774
rect 11308 -19824 11324 -19790
rect 11358 -19824 11452 -19790
rect 11308 -19840 11452 -19824
rect 11500 -19790 11644 -19774
rect 11500 -19824 11516 -19790
rect 11550 -19824 11644 -19790
rect 11500 -19840 11644 -19824
rect 11326 -19865 11386 -19840
rect 11116 -20045 11290 -19907
rect 10980 -20117 11194 -20087
rect 11164 -20150 11194 -20117
rect 11260 -20150 11290 -20045
rect 11332 -20127 11386 -19865
rect 11500 -19970 11590 -19840
rect 16017 -19878 16047 -19602
rect 16017 -19908 16239 -19878
rect 16209 -19923 16239 -19908
rect 16305 -19923 16335 -19602
rect 16401 -19531 16431 -19505
rect 16497 -19531 16527 -19505
rect 16593 -19531 16623 -19505
rect 16401 -19552 16623 -19531
rect 16401 -19586 16417 -19552
rect 16451 -19561 16623 -19552
rect 16689 -19531 16719 -19505
rect 16785 -19531 16815 -19505
rect 16881 -19531 16911 -19505
rect 16689 -19561 16911 -19531
rect 16451 -19586 16467 -19561
rect 16401 -19602 16467 -19586
rect 16401 -19923 16431 -19602
rect 16689 -19818 16719 -19561
rect 16653 -19834 16719 -19818
rect 16653 -19855 16669 -19834
rect 16497 -19868 16669 -19855
rect 16703 -19868 16719 -19834
rect 16497 -19885 16719 -19868
rect 16497 -19923 16527 -19885
rect 11356 -20150 11386 -20127
rect 11452 -20000 11590 -19970
rect 11452 -20150 11482 -20000
rect 16209 -20149 16239 -20123
rect 16305 -20149 16335 -20123
rect 16401 -20149 16431 -20123
rect 16497 -20149 16527 -20123
rect -2068 -20191 -1810 -20175
rect -2068 -20225 -2052 -20191
rect -1826 -20225 -1810 -20191
rect -2068 -20241 -1810 -20225
rect -1622 -20191 -1556 -20174
rect -1622 -20225 -1606 -20191
rect -1572 -20225 -1556 -20191
rect -1622 -20241 -1556 -20225
rect -4784 -20295 -4526 -20279
rect -4784 -20329 -4768 -20295
rect -4542 -20329 -4526 -20295
rect -4784 -20345 -4526 -20329
rect -4338 -20295 -4272 -20279
rect -4338 -20329 -4322 -20295
rect -4288 -20329 -4272 -20295
rect -4766 -20376 -4736 -20345
rect -4670 -20376 -4640 -20345
rect -4574 -20376 -4544 -20345
rect -4338 -20346 -4272 -20329
rect -4320 -20376 -4290 -20346
rect -2050 -20370 -2020 -20344
rect -1954 -20370 -1924 -20344
rect -1858 -20370 -1828 -20344
rect -4766 -20616 -4736 -20590
rect -4670 -20616 -4640 -20590
rect -4574 -20616 -4544 -20590
rect -4320 -20602 -4290 -20576
rect -1604 -20384 -1574 -20358
rect -2050 -20615 -2020 -20584
rect -1954 -20615 -1924 -20584
rect -1858 -20615 -1828 -20584
rect -1604 -20614 -1574 -20584
rect -2068 -20631 -1810 -20615
rect -4784 -20674 -4526 -20658
rect -4784 -20708 -4768 -20674
rect -4542 -20708 -4526 -20674
rect -4784 -20724 -4526 -20708
rect -4338 -20674 -4272 -20658
rect -4338 -20708 -4322 -20674
rect -4288 -20708 -4272 -20674
rect -2068 -20665 -2052 -20631
rect -1826 -20665 -1810 -20631
rect -2068 -20681 -1810 -20665
rect -1622 -20631 -1556 -20614
rect -1622 -20665 -1606 -20631
rect -1572 -20665 -1556 -20631
rect -1622 -20681 -1556 -20665
rect -4766 -20755 -4736 -20724
rect -4670 -20755 -4640 -20724
rect -4574 -20755 -4544 -20724
rect -4338 -20725 -4272 -20708
rect -4320 -20755 -4290 -20725
rect 11835 -20631 11865 -20605
rect 11931 -20631 11961 -20605
rect 12027 -20631 12057 -20605
rect 12123 -20631 12153 -20605
rect 12219 -20631 12249 -20605
rect 12315 -20631 12345 -20605
rect 12411 -20631 12441 -20605
rect 12507 -20631 12537 -20605
rect 12603 -20631 12633 -20605
rect 12699 -20631 12729 -20605
rect 12826 -20795 12892 -20779
rect 11835 -20913 11865 -20887
rect 11931 -20913 11961 -20887
rect 12027 -20913 12057 -20887
rect 12123 -20913 12153 -20887
rect 12219 -20913 12249 -20887
rect 11835 -20937 12249 -20913
rect -4766 -20995 -4736 -20969
rect -4670 -20995 -4640 -20969
rect -4574 -20995 -4544 -20969
rect -4320 -20981 -4290 -20955
rect 7422 -20976 7452 -20950
rect 7518 -20976 7548 -20950
rect 7614 -20976 7644 -20950
rect 7710 -20976 7740 -20950
rect 8370 -20976 8400 -20950
rect 8466 -20976 8496 -20950
rect 8562 -20976 8592 -20950
rect 8658 -20976 8688 -20950
rect 9306 -20976 9336 -20950
rect 9402 -20976 9432 -20950
rect 9498 -20976 9528 -20950
rect 9594 -20976 9624 -20950
rect 10237 -20976 10267 -20950
rect 10333 -20976 10363 -20950
rect 10429 -20976 10459 -20950
rect 10525 -20976 10555 -20950
rect 11164 -20976 11194 -20950
rect 11260 -20976 11290 -20950
rect 11356 -20976 11386 -20950
rect 11452 -20976 11482 -20950
rect 11835 -20971 12170 -20937
rect 12204 -20971 12249 -20937
rect 11835 -20984 12249 -20971
rect 7422 -21078 7452 -21052
rect 7518 -21078 7548 -21052
rect 7614 -21078 7644 -21052
rect 7710 -21078 7740 -21052
rect 8370 -21078 8400 -21052
rect 8466 -21078 8496 -21052
rect 8562 -21078 8592 -21052
rect 8658 -21078 8688 -21052
rect 9306 -21078 9336 -21052
rect 9402 -21078 9432 -21052
rect 9498 -21078 9528 -21052
rect 9594 -21078 9624 -21052
rect 10237 -21077 10267 -21051
rect 10333 -21077 10363 -21051
rect 10429 -21077 10459 -21051
rect 10525 -21077 10555 -21051
rect -21142 -21209 -21126 -21175
rect -21092 -21209 -21076 -21175
rect -12340 -21194 -12314 -21164
rect -11764 -21194 -11274 -21164
rect -11144 -21194 -11118 -21164
rect -21142 -21225 -21076 -21209
rect -23989 -21249 -23959 -21227
rect -24426 -21303 -24395 -21273
rect -24181 -21303 -24125 -21273
rect -24155 -21333 -24125 -21303
rect -24026 -21265 -23959 -21249
rect -24026 -21299 -24010 -21265
rect -23975 -21299 -23959 -21265
rect -24026 -21315 -23959 -21299
rect -23893 -21249 -23863 -21227
rect -23893 -21265 -23826 -21249
rect -15977 -21265 -15947 -21239
rect -15881 -21265 -15851 -21239
rect -15785 -21265 -15755 -21239
rect -11733 -21227 -11299 -21194
rect -23893 -21299 -23877 -21265
rect -23842 -21299 -23826 -21265
rect -24155 -21349 -24088 -21333
rect -24155 -21369 -24134 -21349
rect -24426 -21399 -24395 -21369
rect -24181 -21383 -24134 -21369
rect -24099 -21357 -24088 -21349
rect -23893 -21357 -23826 -21299
rect -24099 -21383 -23826 -21357
rect -24181 -21399 -23826 -21383
rect -21568 -21394 -21538 -21368
rect -21472 -21394 -21442 -21368
rect -21376 -21394 -21346 -21368
rect -24155 -21400 -23826 -21399
rect -21122 -21408 -21092 -21382
rect -15531 -21279 -15501 -21253
rect -11583 -21288 -11474 -21227
rect -11571 -21389 -11485 -21288
rect -11571 -21431 -11549 -21389
rect -11507 -21431 -11485 -21389
rect -11571 -21447 -11485 -21431
rect -15977 -21510 -15947 -21479
rect -15881 -21510 -15851 -21479
rect -15785 -21510 -15755 -21479
rect -15531 -21509 -15501 -21479
rect -15995 -21526 -15737 -21510
rect -15995 -21560 -15979 -21526
rect -15753 -21560 -15737 -21526
rect -17703 -21591 -17677 -21561
rect -17421 -21591 -17324 -21561
rect -15995 -21576 -15737 -21560
rect -15549 -21526 -15483 -21509
rect -15549 -21560 -15533 -21526
rect -15499 -21560 -15483 -21526
rect -15549 -21576 -15483 -21560
rect -21568 -21639 -21538 -21608
rect -21472 -21639 -21442 -21608
rect -21376 -21639 -21346 -21608
rect -21122 -21638 -21092 -21608
rect -21586 -21655 -21328 -21639
rect -21586 -21689 -21570 -21655
rect -21344 -21689 -21328 -21655
rect -21586 -21705 -21328 -21689
rect -21140 -21655 -21074 -21638
rect -21140 -21689 -21124 -21655
rect -21090 -21689 -21074 -21655
rect -17395 -21657 -17324 -21591
rect -17703 -21687 -17677 -21657
rect -17421 -21687 -17324 -21657
rect -21140 -21705 -21074 -21689
rect -17395 -21753 -17324 -21687
rect -17703 -21783 -17677 -21753
rect -17421 -21783 -17324 -21753
rect -17395 -21849 -17324 -21783
rect -17703 -21879 -17677 -21849
rect -17421 -21879 -17324 -21849
rect 11164 -21078 11194 -21052
rect 11260 -21078 11290 -21052
rect 11356 -21078 11386 -21052
rect 11452 -21078 11482 -21052
rect -17395 -21945 -17324 -21879
rect -17282 -21943 -17216 -21927
rect -17282 -21945 -17266 -21943
rect -17703 -21975 -17677 -21945
rect -17421 -21975 -17266 -21945
rect -17282 -21977 -17266 -21975
rect -17232 -21945 -17216 -21943
rect -17232 -21975 -17188 -21945
rect -16988 -21975 -16962 -21945
rect -17232 -21977 -17216 -21975
rect -17282 -21993 -17216 -21977
rect -17703 -22071 -17677 -22041
rect -17421 -22071 -17188 -22041
rect -16988 -22071 -16962 -22041
rect -23990 -22130 -23960 -22104
rect -23894 -22130 -23864 -22104
rect -24427 -22222 -24396 -22192
rect -24182 -22222 -24126 -22192
rect -24156 -22288 -24126 -22222
rect -24427 -22318 -24396 -22288
rect -24182 -22318 -24126 -22288
rect -24156 -22347 -24126 -22318
rect -24156 -22363 -24089 -22347
rect -24156 -22384 -24135 -22363
rect -24427 -22414 -24396 -22384
rect -24182 -22397 -24135 -22384
rect -24100 -22397 -24089 -22363
rect -24182 -22414 -24089 -22397
rect -24427 -22510 -24396 -22480
rect -24182 -22510 -24126 -22480
rect -24156 -22576 -24126 -22510
rect -17395 -22086 -17324 -22071
rect -17395 -22120 -17371 -22086
rect -17337 -22120 -17324 -22086
rect -17395 -22137 -17324 -22120
rect 7422 -21911 7452 -21878
rect 7238 -21941 7452 -21911
rect -17703 -22167 -17677 -22137
rect -17421 -22167 -17324 -22137
rect -17395 -22233 -17324 -22167
rect 7238 -22188 7268 -21941
rect 7518 -21983 7548 -21878
rect 7614 -21901 7644 -21878
rect 7374 -22121 7548 -21983
rect -17703 -22263 -17677 -22233
rect -17421 -22263 -17324 -22233
rect 7182 -22204 7326 -22188
rect 7182 -22238 7198 -22204
rect 7232 -22238 7326 -22204
rect 7182 -22254 7326 -22238
rect 7374 -22204 7518 -22121
rect 7590 -22163 7644 -21901
rect 7710 -22028 7740 -21878
rect 8370 -21911 8400 -21878
rect 8186 -21941 8400 -21911
rect 7710 -22058 7848 -22028
rect 7584 -22188 7644 -22163
rect 7758 -22188 7848 -22058
rect 8186 -22188 8216 -21941
rect 8466 -21983 8496 -21878
rect 8562 -21901 8592 -21878
rect 8322 -22121 8496 -21983
rect 7374 -22238 7390 -22204
rect 7424 -22238 7518 -22204
rect 7374 -22254 7518 -22238
rect 7566 -22204 7710 -22188
rect 7566 -22238 7582 -22204
rect 7616 -22238 7710 -22204
rect 7566 -22254 7710 -22238
rect 7758 -22204 7902 -22188
rect 7758 -22238 7774 -22204
rect 7808 -22238 7902 -22204
rect 7758 -22254 7902 -22238
rect 8130 -22204 8274 -22188
rect 8130 -22238 8146 -22204
rect 8180 -22238 8274 -22204
rect 8130 -22254 8274 -22238
rect 8322 -22204 8466 -22121
rect 8538 -22163 8592 -21901
rect 8658 -22028 8688 -21878
rect 9306 -21911 9336 -21878
rect 9122 -21941 9336 -21911
rect 8658 -22058 8796 -22028
rect 8532 -22188 8592 -22163
rect 8706 -22188 8796 -22058
rect 9122 -22188 9152 -21941
rect 9402 -21983 9432 -21878
rect 9498 -21901 9528 -21878
rect 9258 -22121 9432 -21983
rect 8322 -22238 8338 -22204
rect 8372 -22238 8466 -22204
rect 8322 -22254 8466 -22238
rect 8514 -22204 8658 -22188
rect 8514 -22238 8530 -22204
rect 8564 -22238 8658 -22204
rect 8514 -22254 8658 -22238
rect 8706 -22204 8850 -22188
rect 8706 -22238 8722 -22204
rect 8756 -22238 8850 -22204
rect 8706 -22254 8850 -22238
rect 9066 -22204 9210 -22188
rect 9066 -22238 9082 -22204
rect 9116 -22238 9210 -22204
rect 9066 -22254 9210 -22238
rect 9258 -22204 9402 -22121
rect 9474 -22163 9528 -21901
rect 9594 -22028 9624 -21878
rect 10237 -21910 10267 -21877
rect 10053 -21940 10267 -21910
rect 9594 -22058 9732 -22028
rect 9468 -22188 9528 -22163
rect 9642 -22188 9732 -22058
rect 10053 -22187 10083 -21940
rect 10333 -21982 10363 -21877
rect 10429 -21900 10459 -21877
rect 10189 -22120 10363 -21982
rect 9258 -22238 9274 -22204
rect 9308 -22238 9402 -22204
rect 9258 -22254 9402 -22238
rect 9450 -22204 9594 -22188
rect 9450 -22238 9466 -22204
rect 9500 -22238 9594 -22204
rect 9450 -22254 9594 -22238
rect 9642 -22204 9786 -22188
rect 9642 -22238 9658 -22204
rect 9692 -22238 9786 -22204
rect 9642 -22254 9786 -22238
rect 9997 -22203 10141 -22187
rect 9997 -22237 10013 -22203
rect 10047 -22237 10141 -22203
rect 9997 -22253 10141 -22237
rect 10189 -22203 10333 -22120
rect 10405 -22162 10459 -21900
rect 10525 -22027 10555 -21877
rect 12219 -21120 12249 -20984
rect 12315 -20913 12345 -20887
rect 12411 -20913 12441 -20887
rect 12507 -20913 12537 -20887
rect 12603 -20913 12633 -20887
rect 12699 -20913 12729 -20887
rect 12315 -20984 12729 -20913
rect 12315 -21026 12345 -20984
rect 12826 -21021 12842 -20795
rect 12876 -20797 12892 -20795
rect 12876 -20827 12923 -20797
rect 13137 -20827 13163 -20797
rect 12876 -20893 12892 -20827
rect 12876 -20923 12923 -20893
rect 13137 -20923 13163 -20893
rect 12876 -20989 12892 -20923
rect 12876 -21019 12923 -20989
rect 13137 -21019 13163 -20989
rect 12876 -21021 12892 -21019
rect 12297 -21042 12363 -21026
rect 12826 -21037 12892 -21021
rect 12297 -21076 12313 -21042
rect 12347 -21076 12363 -21042
rect 12297 -21092 12363 -21076
rect 12315 -21120 12345 -21092
rect 12826 -21241 12893 -21225
rect 12826 -21275 12842 -21241
rect 12876 -21243 12893 -21241
rect 12876 -21273 12923 -21243
rect 13123 -21273 13149 -21243
rect 12876 -21275 12893 -21273
rect 12826 -21291 12893 -21275
rect 12219 -21346 12249 -21320
rect 12315 -21346 12345 -21320
rect 11164 -21911 11194 -21878
rect 10980 -21941 11194 -21911
rect 10525 -22057 10663 -22027
rect 10399 -22187 10459 -22162
rect 10573 -22187 10663 -22057
rect 10189 -22237 10205 -22203
rect 10239 -22237 10333 -22203
rect 10189 -22253 10333 -22237
rect 10381 -22203 10525 -22187
rect 10381 -22237 10397 -22203
rect 10431 -22237 10525 -22203
rect 10381 -22253 10525 -22237
rect 10573 -22203 10717 -22187
rect 10980 -22188 11010 -21941
rect 11260 -21983 11290 -21878
rect 11356 -21901 11386 -21878
rect 11116 -22121 11290 -21983
rect 10573 -22237 10589 -22203
rect 10623 -22237 10717 -22203
rect 10573 -22253 10717 -22237
rect -17395 -22329 -17324 -22263
rect 7200 -22285 7230 -22254
rect 7296 -22285 7326 -22254
rect 7392 -22285 7422 -22254
rect 7488 -22285 7518 -22254
rect 7584 -22285 7614 -22254
rect 7680 -22285 7710 -22254
rect 7776 -22285 7806 -22254
rect 7872 -22285 7902 -22254
rect 8148 -22285 8178 -22254
rect 8244 -22285 8274 -22254
rect 8340 -22285 8370 -22254
rect 8436 -22285 8466 -22254
rect 8532 -22285 8562 -22254
rect 8628 -22285 8658 -22254
rect 8724 -22285 8754 -22254
rect 8820 -22285 8850 -22254
rect 9084 -22285 9114 -22254
rect 9180 -22285 9210 -22254
rect 9276 -22285 9306 -22254
rect 9372 -22285 9402 -22254
rect 9468 -22285 9498 -22254
rect 9564 -22285 9594 -22254
rect 9660 -22285 9690 -22254
rect 9756 -22285 9786 -22254
rect 10015 -22284 10045 -22253
rect 10111 -22284 10141 -22253
rect 10207 -22284 10237 -22253
rect 10303 -22284 10333 -22253
rect 10399 -22284 10429 -22253
rect 10495 -22284 10525 -22253
rect 10591 -22284 10621 -22253
rect 10687 -22284 10717 -22253
rect 10924 -22204 11068 -22188
rect 10924 -22238 10940 -22204
rect 10974 -22238 11068 -22204
rect 10924 -22254 11068 -22238
rect 11116 -22204 11260 -22121
rect 11332 -22163 11386 -21901
rect 11452 -22028 11482 -21878
rect 11452 -22058 11590 -22028
rect 11326 -22188 11386 -22163
rect 11500 -22188 11590 -22058
rect 11116 -22238 11132 -22204
rect 11166 -22238 11260 -22204
rect 11116 -22254 11260 -22238
rect 11308 -22204 11452 -22188
rect 11308 -22238 11324 -22204
rect 11358 -22238 11452 -22204
rect 11308 -22254 11452 -22238
rect 11500 -22204 11644 -22188
rect 11500 -22238 11516 -22204
rect 11550 -22238 11644 -22204
rect 11500 -22254 11644 -22238
rect -17703 -22359 -17677 -22329
rect -17421 -22359 -17324 -22329
rect -17395 -22425 -17324 -22359
rect -17703 -22455 -17677 -22425
rect -17421 -22455 -17324 -22425
rect -23990 -22552 -23960 -22530
rect -24427 -22606 -24396 -22576
rect -24182 -22606 -24126 -22576
rect -24156 -22636 -24126 -22606
rect -24027 -22568 -23960 -22552
rect -24027 -22602 -24011 -22568
rect -23976 -22602 -23960 -22568
rect -24027 -22618 -23960 -22602
rect -23894 -22552 -23864 -22530
rect -12340 -22533 -12314 -22503
rect -11764 -22533 -11274 -22503
rect -11144 -22533 -11118 -22503
rect -23894 -22568 -23827 -22552
rect -23894 -22602 -23878 -22568
rect -23843 -22602 -23827 -22568
rect -24156 -22652 -24089 -22636
rect -24156 -22672 -24135 -22652
rect -24427 -22702 -24396 -22672
rect -24182 -22686 -24135 -22672
rect -24100 -22660 -24089 -22652
rect -23894 -22660 -23827 -22602
rect -24100 -22686 -23827 -22660
rect -24182 -22702 -23827 -22686
rect -24156 -22703 -23827 -22702
rect -17703 -22991 -17677 -22961
rect -17421 -22991 -17324 -22961
rect -17395 -23057 -17324 -22991
rect -17703 -23087 -17677 -23057
rect -17421 -23087 -17324 -23057
rect -17395 -23153 -17324 -23087
rect -17703 -23183 -17677 -23153
rect -17421 -23183 -17324 -23153
rect -17395 -23249 -17324 -23183
rect -17703 -23279 -17677 -23249
rect -17421 -23279 -17324 -23249
rect -17395 -23345 -17324 -23279
rect -17282 -23343 -17216 -23327
rect -17282 -23345 -17266 -23343
rect -17703 -23375 -17677 -23345
rect -17421 -23375 -17266 -23345
rect -23990 -23439 -23960 -23413
rect -23894 -23439 -23864 -23413
rect -17282 -23377 -17266 -23375
rect -17232 -23345 -17216 -23343
rect -17232 -23375 -17188 -23345
rect -16988 -23375 -16962 -23345
rect -17232 -23377 -17216 -23375
rect -17282 -23393 -17216 -23377
rect -24427 -23531 -24396 -23501
rect -24182 -23531 -24126 -23501
rect -24156 -23597 -24126 -23531
rect -24427 -23627 -24396 -23597
rect -24182 -23627 -24126 -23597
rect -24156 -23656 -24126 -23627
rect -24156 -23672 -24089 -23656
rect -24156 -23693 -24135 -23672
rect -24427 -23723 -24396 -23693
rect -24182 -23706 -24135 -23693
rect -24100 -23706 -24089 -23672
rect -24182 -23723 -24089 -23706
rect -24427 -23819 -24396 -23789
rect -24182 -23819 -24126 -23789
rect -24156 -23885 -24126 -23819
rect -17703 -23471 -17677 -23441
rect -17421 -23471 -17188 -23441
rect -16988 -23471 -16962 -23441
rect -23990 -23861 -23960 -23839
rect -24427 -23915 -24396 -23885
rect -24182 -23915 -24126 -23885
rect -24156 -23945 -24126 -23915
rect -24027 -23877 -23960 -23861
rect -24027 -23911 -24011 -23877
rect -23976 -23911 -23960 -23877
rect -24027 -23927 -23960 -23911
rect -23894 -23861 -23864 -23839
rect -23894 -23877 -23827 -23861
rect -23894 -23911 -23878 -23877
rect -23843 -23911 -23827 -23877
rect -17395 -23486 -17324 -23471
rect -17395 -23520 -17371 -23486
rect -17337 -23520 -17324 -23486
rect -17395 -23537 -17324 -23520
rect -17703 -23567 -17677 -23537
rect -17421 -23567 -17324 -23537
rect -17395 -23633 -17324 -23567
rect -17703 -23663 -17677 -23633
rect -17421 -23663 -17324 -23633
rect -17395 -23729 -17324 -23663
rect -17703 -23759 -17677 -23729
rect -17421 -23759 -17324 -23729
rect -11733 -22595 -11296 -22533
rect -12345 -22625 -12314 -22595
rect -11764 -22625 -11274 -22595
rect -11144 -22625 -11118 -22595
rect -11733 -22691 -11296 -22625
rect -12345 -22721 -12314 -22691
rect -11764 -22720 -11274 -22691
rect -11764 -22721 -11576 -22720
rect -11733 -22785 -11576 -22721
rect -11521 -22721 -11274 -22720
rect -11144 -22721 -11118 -22691
rect -11521 -22785 -11296 -22721
rect -11733 -22787 -11296 -22785
rect -12345 -22817 -12314 -22787
rect -11764 -22817 -11274 -22787
rect -11144 -22817 -11118 -22787
rect -12345 -22913 -12314 -22883
rect -11764 -22902 -11640 -22883
rect -11764 -22913 -11700 -22902
rect -11733 -22979 -11700 -22913
rect -12345 -23009 -12314 -22979
rect -11764 -23009 -11700 -22979
rect -11733 -23032 -11700 -23009
rect -11655 -23032 -11640 -22902
rect -11733 -23075 -11640 -23032
rect -12345 -23105 -12314 -23075
rect -11764 -23105 -11640 -23075
rect -11583 -22913 -11274 -22883
rect -11144 -22913 -11118 -22883
rect -11583 -22979 -11296 -22913
rect -11583 -23009 -11274 -22979
rect -11144 -23009 -11118 -22979
rect -11583 -23075 -11296 -23009
rect -11583 -23105 -11274 -23075
rect -11144 -23105 -11118 -23075
rect -12345 -23201 -12314 -23171
rect -11764 -23201 -11641 -23171
rect -11734 -23233 -11641 -23201
rect -11734 -23267 -11705 -23233
rect -12345 -23297 -12314 -23267
rect -11764 -23297 -11705 -23267
rect -11734 -23363 -11705 -23297
rect -11660 -23363 -11641 -23233
rect -12345 -23393 -12314 -23363
rect -11764 -23393 -11641 -23363
rect -11583 -23457 -11474 -23105
rect -11404 -23201 -11274 -23171
rect -11144 -23201 -11118 -23171
rect -11404 -23225 -11296 -23201
rect -11404 -23355 -11376 -23225
rect -11331 -23267 -11296 -23225
rect -11331 -23297 -11274 -23267
rect -11144 -23297 -11118 -23267
rect -11331 -23355 -11296 -23297
rect -11404 -23363 -11296 -23355
rect -11404 -23393 -11274 -23363
rect -11144 -23393 -11118 -23363
rect -11733 -23459 -11474 -23457
rect -12345 -23489 -12314 -23459
rect -11764 -23489 -11474 -23459
rect -11733 -23555 -11474 -23489
rect -12345 -23585 -12314 -23555
rect -11764 -23585 -11474 -23555
rect -11733 -23651 -11474 -23585
rect -12345 -23681 -12314 -23651
rect -11764 -23681 -11474 -23651
rect -11409 -23489 -11274 -23459
rect -11144 -23489 -11118 -23459
rect -11409 -23508 -11296 -23489
rect -11409 -23638 -11384 -23508
rect -11339 -23555 -11296 -23508
rect -11339 -23585 -11274 -23555
rect -11144 -23585 -11118 -23555
rect -11339 -23638 -11296 -23585
rect -11409 -23651 -11296 -23638
rect -11409 -23681 -11274 -23651
rect -11144 -23681 -11118 -23651
rect -11733 -23730 -11474 -23681
rect -11733 -23743 -11299 -23730
rect 10942 -22285 10972 -22254
rect 11038 -22285 11068 -22254
rect 11134 -22285 11164 -22254
rect 11230 -22285 11260 -22254
rect 11326 -22285 11356 -22254
rect 11422 -22285 11452 -22254
rect 11518 -22285 11548 -22254
rect 11614 -22285 11644 -22254
rect 7200 -22633 7230 -22607
rect 7296 -22633 7326 -22607
rect 7392 -22633 7422 -22607
rect 7488 -22633 7518 -22607
rect 7584 -22633 7614 -22607
rect 7680 -22633 7710 -22607
rect 7776 -22633 7806 -22607
rect 7872 -22633 7902 -22607
rect 8148 -22633 8178 -22607
rect 8244 -22633 8274 -22607
rect 8340 -22633 8370 -22607
rect 8436 -22633 8466 -22607
rect 8532 -22633 8562 -22607
rect 8628 -22633 8658 -22607
rect 8724 -22633 8754 -22607
rect 8820 -22633 8850 -22607
rect 9084 -22633 9114 -22607
rect 9180 -22633 9210 -22607
rect 9276 -22633 9306 -22607
rect 9372 -22633 9402 -22607
rect 9468 -22633 9498 -22607
rect 9564 -22633 9594 -22607
rect 9660 -22633 9690 -22607
rect 9756 -22633 9786 -22607
rect 10015 -22632 10045 -22606
rect 10111 -22632 10141 -22606
rect 10207 -22632 10237 -22606
rect 10303 -22632 10333 -22606
rect 10399 -22632 10429 -22606
rect 10495 -22632 10525 -22606
rect 10591 -22632 10621 -22606
rect 10687 -22632 10717 -22606
rect 10942 -22633 10972 -22607
rect 11038 -22633 11068 -22607
rect 11134 -22633 11164 -22607
rect 11230 -22633 11260 -22607
rect 11326 -22633 11356 -22607
rect 11422 -22633 11452 -22607
rect 11518 -22633 11548 -22607
rect 11614 -22633 11644 -22607
rect 5561 -23305 5627 -23289
rect 5561 -23531 5577 -23305
rect 5611 -23307 5627 -23305
rect 6001 -23305 6067 -23289
rect 5611 -23337 5658 -23307
rect 5872 -23337 5898 -23307
rect 5611 -23403 5627 -23337
rect 5611 -23433 5658 -23403
rect 5872 -23433 5898 -23403
rect 5611 -23499 5627 -23433
rect 5611 -23529 5658 -23499
rect 5872 -23529 5898 -23499
rect 5611 -23531 5627 -23529
rect 5561 -23547 5627 -23531
rect 6001 -23531 6017 -23305
rect 6051 -23307 6067 -23305
rect 6441 -23305 6507 -23289
rect 6051 -23337 6098 -23307
rect 6312 -23337 6338 -23307
rect 6051 -23403 6067 -23337
rect 6051 -23433 6098 -23403
rect 6312 -23433 6338 -23403
rect 6051 -23499 6067 -23433
rect 6051 -23529 6098 -23499
rect 6312 -23529 6338 -23499
rect 6051 -23531 6067 -23529
rect 6001 -23547 6067 -23531
rect 6441 -23531 6457 -23305
rect 6491 -23307 6507 -23305
rect 6491 -23337 6538 -23307
rect 6752 -23337 6778 -23307
rect 6491 -23403 6507 -23337
rect 6491 -23433 6538 -23403
rect 6752 -23433 6778 -23403
rect 6491 -23499 6507 -23433
rect 6491 -23529 6538 -23499
rect 6752 -23529 6778 -23499
rect 6491 -23531 6507 -23529
rect 6441 -23547 6507 -23531
rect -17395 -23825 -17324 -23759
rect -12340 -23773 -12314 -23743
rect -11764 -23773 -11274 -23743
rect -11144 -23773 -11118 -23743
rect 5561 -23751 5628 -23735
rect -17703 -23855 -17677 -23825
rect -17421 -23855 -17324 -23825
rect -11733 -23806 -11299 -23773
rect -11583 -23867 -11474 -23806
rect 5561 -23785 5577 -23751
rect 5611 -23753 5628 -23751
rect 6001 -23751 6068 -23735
rect 5611 -23783 5658 -23753
rect 5858 -23783 5884 -23753
rect 5611 -23785 5628 -23783
rect 5561 -23801 5628 -23785
rect 6001 -23785 6017 -23751
rect 6051 -23753 6068 -23751
rect 6441 -23751 6508 -23735
rect 6051 -23783 6098 -23753
rect 6298 -23783 6324 -23753
rect 6051 -23785 6068 -23783
rect 6001 -23801 6068 -23785
rect 6441 -23785 6457 -23751
rect 6491 -23753 6508 -23751
rect 6491 -23783 6538 -23753
rect 6738 -23783 6764 -23753
rect 6491 -23785 6508 -23783
rect 6441 -23801 6508 -23785
rect -24156 -23961 -24089 -23945
rect -24156 -23981 -24135 -23961
rect -24427 -24011 -24396 -23981
rect -24182 -23995 -24135 -23981
rect -24100 -23969 -24089 -23961
rect -23894 -23969 -23827 -23911
rect -24100 -23995 -23827 -23969
rect -24182 -24011 -23827 -23995
rect -24156 -24012 -23827 -24011
rect -11575 -23970 -11482 -23867
rect 7200 -23949 7230 -23923
rect 7296 -23949 7326 -23923
rect 7392 -23949 7422 -23923
rect 7488 -23949 7518 -23923
rect 7584 -23949 7614 -23923
rect 7680 -23949 7710 -23923
rect 7776 -23949 7806 -23923
rect 7872 -23949 7902 -23923
rect 8148 -23949 8178 -23923
rect 8244 -23949 8274 -23923
rect 8340 -23949 8370 -23923
rect 8436 -23949 8466 -23923
rect 8532 -23949 8562 -23923
rect 8628 -23949 8658 -23923
rect 8724 -23949 8754 -23923
rect 8820 -23949 8850 -23923
rect 9084 -23949 9114 -23923
rect 9180 -23949 9210 -23923
rect 9276 -23949 9306 -23923
rect 9372 -23949 9402 -23923
rect 9468 -23949 9498 -23923
rect 9564 -23949 9594 -23923
rect 9660 -23949 9690 -23923
rect 9756 -23949 9786 -23923
rect 10015 -23949 10045 -23923
rect 10111 -23949 10141 -23923
rect 10207 -23949 10237 -23923
rect 10303 -23949 10333 -23923
rect 10399 -23949 10429 -23923
rect 10495 -23949 10525 -23923
rect 10591 -23949 10621 -23923
rect 10687 -23949 10717 -23923
rect 10942 -23949 10972 -23923
rect 11038 -23949 11068 -23923
rect 11134 -23949 11164 -23923
rect 11230 -23949 11260 -23923
rect 11326 -23949 11356 -23923
rect 11422 -23949 11452 -23923
rect 11518 -23949 11548 -23923
rect 11614 -23949 11644 -23923
rect -11575 -24019 -11553 -23970
rect -11504 -24019 -11482 -23970
rect -11575 -24035 -11482 -24019
rect 7200 -24302 7230 -24271
rect 7296 -24302 7326 -24271
rect 7392 -24302 7422 -24271
rect 7488 -24302 7518 -24271
rect 7584 -24302 7614 -24271
rect 7680 -24302 7710 -24271
rect 7776 -24302 7806 -24271
rect 7872 -24302 7902 -24271
rect 8148 -24302 8178 -24271
rect 8244 -24302 8274 -24271
rect 8340 -24302 8370 -24271
rect 8436 -24302 8466 -24271
rect 8532 -24302 8562 -24271
rect 8628 -24302 8658 -24271
rect 8724 -24302 8754 -24271
rect 8820 -24302 8850 -24271
rect 9084 -24302 9114 -24271
rect 9180 -24302 9210 -24271
rect 9276 -24302 9306 -24271
rect 9372 -24302 9402 -24271
rect 9468 -24302 9498 -24271
rect 9564 -24302 9594 -24271
rect 9660 -24302 9690 -24271
rect 9756 -24302 9786 -24271
rect 10015 -24302 10045 -24271
rect 10111 -24302 10141 -24271
rect 10207 -24302 10237 -24271
rect 10303 -24302 10333 -24271
rect 10399 -24302 10429 -24271
rect 10495 -24302 10525 -24271
rect 10591 -24302 10621 -24271
rect 10687 -24302 10717 -24271
rect 10942 -24302 10972 -24271
rect 11038 -24302 11068 -24271
rect 11134 -24302 11164 -24271
rect 11230 -24302 11260 -24271
rect 11326 -24302 11356 -24271
rect 11422 -24302 11452 -24271
rect 11518 -24302 11548 -24271
rect 11614 -24302 11644 -24271
rect 7182 -24318 7326 -24302
rect 7182 -24352 7198 -24318
rect 7232 -24352 7326 -24318
rect -17703 -24391 -17677 -24361
rect -17421 -24391 -17324 -24361
rect 7182 -24368 7326 -24352
rect 7374 -24318 7518 -24302
rect 7374 -24352 7390 -24318
rect 7424 -24352 7518 -24318
rect -17395 -24457 -17324 -24391
rect -17703 -24487 -17677 -24457
rect -17421 -24487 -17324 -24457
rect -17395 -24553 -17324 -24487
rect -17703 -24583 -17677 -24553
rect -17421 -24583 -17324 -24553
rect -17395 -24649 -17324 -24583
rect 7238 -24615 7268 -24368
rect 7374 -24435 7518 -24352
rect 7566 -24318 7710 -24302
rect 7566 -24352 7582 -24318
rect 7616 -24352 7710 -24318
rect 7566 -24368 7710 -24352
rect 7758 -24318 7902 -24302
rect 7758 -24352 7774 -24318
rect 7808 -24352 7902 -24318
rect 7758 -24368 7902 -24352
rect 8130 -24318 8274 -24302
rect 8130 -24352 8146 -24318
rect 8180 -24352 8274 -24318
rect 8130 -24368 8274 -24352
rect 8322 -24318 8466 -24302
rect 8322 -24352 8338 -24318
rect 8372 -24352 8466 -24318
rect 7584 -24393 7644 -24368
rect 7374 -24573 7548 -24435
rect 7238 -24645 7452 -24615
rect -17703 -24679 -17677 -24649
rect -17421 -24679 -17324 -24649
rect 7422 -24678 7452 -24645
rect 7518 -24678 7548 -24573
rect 7590 -24655 7644 -24393
rect 7758 -24498 7848 -24368
rect 7614 -24678 7644 -24655
rect 7710 -24528 7848 -24498
rect 7710 -24678 7740 -24528
rect 8186 -24615 8216 -24368
rect 8322 -24435 8466 -24352
rect 8514 -24318 8658 -24302
rect 8514 -24352 8530 -24318
rect 8564 -24352 8658 -24318
rect 8514 -24368 8658 -24352
rect 8706 -24318 8850 -24302
rect 8706 -24352 8722 -24318
rect 8756 -24352 8850 -24318
rect 8706 -24368 8850 -24352
rect 9066 -24318 9210 -24302
rect 9066 -24352 9082 -24318
rect 9116 -24352 9210 -24318
rect 9066 -24368 9210 -24352
rect 9258 -24318 9402 -24302
rect 9258 -24352 9274 -24318
rect 9308 -24352 9402 -24318
rect 8532 -24393 8592 -24368
rect 8322 -24573 8496 -24435
rect 8186 -24645 8400 -24615
rect 8370 -24678 8400 -24645
rect 8466 -24678 8496 -24573
rect 8538 -24655 8592 -24393
rect 8706 -24498 8796 -24368
rect 8562 -24678 8592 -24655
rect 8658 -24528 8796 -24498
rect 8658 -24678 8688 -24528
rect 9122 -24615 9152 -24368
rect 9258 -24435 9402 -24352
rect 9450 -24318 9594 -24302
rect 9450 -24352 9466 -24318
rect 9500 -24352 9594 -24318
rect 9450 -24368 9594 -24352
rect 9642 -24318 9786 -24302
rect 9642 -24352 9658 -24318
rect 9692 -24352 9786 -24318
rect 9642 -24368 9786 -24352
rect 9997 -24318 10141 -24302
rect 9997 -24352 10013 -24318
rect 10047 -24352 10141 -24318
rect 9997 -24368 10141 -24352
rect 10189 -24318 10333 -24302
rect 10189 -24352 10205 -24318
rect 10239 -24352 10333 -24318
rect 9468 -24393 9528 -24368
rect 9258 -24573 9432 -24435
rect 9122 -24645 9336 -24615
rect 9306 -24678 9336 -24645
rect 9402 -24678 9432 -24573
rect 9474 -24655 9528 -24393
rect 9642 -24498 9732 -24368
rect 9498 -24678 9528 -24655
rect 9594 -24528 9732 -24498
rect 9594 -24678 9624 -24528
rect 10053 -24615 10083 -24368
rect 10189 -24435 10333 -24352
rect 10381 -24318 10525 -24302
rect 10381 -24352 10397 -24318
rect 10431 -24352 10525 -24318
rect 10381 -24368 10525 -24352
rect 10573 -24318 10717 -24302
rect 10573 -24352 10589 -24318
rect 10623 -24352 10717 -24318
rect 10573 -24368 10717 -24352
rect 10924 -24318 11068 -24302
rect 10924 -24352 10940 -24318
rect 10974 -24352 11068 -24318
rect 10924 -24368 11068 -24352
rect 11116 -24318 11260 -24302
rect 11116 -24352 11132 -24318
rect 11166 -24352 11260 -24318
rect 10399 -24393 10459 -24368
rect 10189 -24573 10363 -24435
rect 10053 -24645 10267 -24615
rect 10237 -24678 10267 -24645
rect 10333 -24678 10363 -24573
rect 10405 -24655 10459 -24393
rect 10573 -24498 10663 -24368
rect 10429 -24678 10459 -24655
rect 10525 -24528 10663 -24498
rect 10525 -24678 10555 -24528
rect 10980 -24615 11010 -24368
rect 11116 -24435 11260 -24352
rect 11308 -24318 11452 -24302
rect 11308 -24352 11324 -24318
rect 11358 -24352 11452 -24318
rect 11308 -24368 11452 -24352
rect 11500 -24318 11644 -24302
rect 11500 -24352 11516 -24318
rect 11550 -24352 11644 -24318
rect 11500 -24368 11644 -24352
rect 11326 -24393 11386 -24368
rect 11116 -24573 11290 -24435
rect 10980 -24645 11194 -24615
rect 11164 -24678 11194 -24645
rect 11260 -24678 11290 -24573
rect 11332 -24655 11386 -24393
rect 11500 -24498 11590 -24368
rect 11356 -24678 11386 -24655
rect 11452 -24528 11590 -24498
rect 11452 -24678 11482 -24528
rect -17395 -24745 -17324 -24679
rect -17282 -24743 -17216 -24727
rect -17282 -24745 -17266 -24743
rect -17703 -24775 -17677 -24745
rect -17421 -24775 -17266 -24745
rect -17282 -24777 -17266 -24775
rect -17232 -24745 -17216 -24743
rect -17232 -24775 -17188 -24745
rect -16988 -24775 -16962 -24745
rect -17232 -24777 -17216 -24775
rect -17282 -24793 -17216 -24777
rect -17703 -24871 -17677 -24841
rect -17421 -24871 -17188 -24841
rect -16988 -24871 -16962 -24841
rect -17395 -24886 -17324 -24871
rect -17395 -24920 -17371 -24886
rect -17337 -24920 -17324 -24886
rect -17395 -24937 -17324 -24920
rect -17703 -24967 -17677 -24937
rect -17421 -24967 -17324 -24937
rect -17395 -25033 -17324 -24967
rect -17703 -25063 -17677 -25033
rect -17421 -25063 -17324 -25033
rect -17395 -25129 -17324 -25063
rect -17703 -25159 -17677 -25129
rect -17421 -25159 -17324 -25129
rect -17395 -25225 -17324 -25159
rect -17703 -25255 -17677 -25225
rect -17421 -25255 -17324 -25225
rect -12340 -25301 -12314 -25271
rect -11764 -25301 -11274 -25271
rect -11144 -25301 -11118 -25271
rect -11733 -25363 -11296 -25301
rect -12345 -25393 -12314 -25363
rect -11764 -25393 -11274 -25363
rect -11144 -25393 -11118 -25363
rect -11733 -25459 -11296 -25393
rect -12345 -25489 -12314 -25459
rect -11764 -25488 -11274 -25459
rect -11764 -25489 -11576 -25488
rect -11733 -25553 -11576 -25489
rect -11521 -25489 -11274 -25488
rect -11144 -25489 -11118 -25459
rect -11521 -25553 -11296 -25489
rect -11733 -25555 -11296 -25553
rect -12345 -25585 -12314 -25555
rect -11764 -25585 -11274 -25555
rect -11144 -25585 -11118 -25555
rect -12345 -25681 -12314 -25651
rect -11764 -25670 -11640 -25651
rect -11764 -25681 -11700 -25670
rect -11733 -25747 -11700 -25681
rect -12345 -25777 -12314 -25747
rect -11764 -25777 -11700 -25747
rect -11733 -25800 -11700 -25777
rect -11655 -25800 -11640 -25670
rect -11733 -25843 -11640 -25800
rect -12345 -25873 -12314 -25843
rect -11764 -25873 -11640 -25843
rect -11583 -25681 -11274 -25651
rect -11144 -25681 -11118 -25651
rect -11583 -25747 -11296 -25681
rect -11583 -25777 -11274 -25747
rect -11144 -25777 -11118 -25747
rect -11583 -25843 -11296 -25777
rect -11583 -25873 -11274 -25843
rect -11144 -25873 -11118 -25843
rect -12345 -25969 -12314 -25939
rect -11764 -25969 -11641 -25939
rect -11734 -26001 -11641 -25969
rect -11734 -26035 -11705 -26001
rect -12345 -26065 -12314 -26035
rect -11764 -26065 -11705 -26035
rect -11734 -26131 -11705 -26065
rect -11660 -26131 -11641 -26001
rect -12345 -26161 -12314 -26131
rect -11764 -26161 -11641 -26131
rect -11583 -26225 -11474 -25873
rect -11404 -25969 -11274 -25939
rect -11144 -25969 -11118 -25939
rect -11404 -25993 -11296 -25969
rect -11404 -26123 -11376 -25993
rect -11331 -26035 -11296 -25993
rect -11331 -26065 -11274 -26035
rect -11144 -26065 -11118 -26035
rect -11331 -26123 -11296 -26065
rect -11404 -26131 -11296 -26123
rect -11404 -26161 -11274 -26131
rect -11144 -26161 -11118 -26131
rect -11733 -26227 -11474 -26225
rect -12345 -26257 -12314 -26227
rect -11764 -26257 -11474 -26227
rect -11733 -26323 -11474 -26257
rect -12345 -26353 -12314 -26323
rect -11764 -26353 -11474 -26323
rect -11733 -26419 -11474 -26353
rect -12345 -26449 -12314 -26419
rect -11764 -26449 -11474 -26419
rect -11409 -26257 -11274 -26227
rect -11144 -26257 -11118 -26227
rect -11409 -26276 -11296 -26257
rect -11409 -26406 -11384 -26276
rect -11339 -26323 -11296 -26276
rect -11339 -26353 -11274 -26323
rect -11144 -26353 -11118 -26323
rect -11339 -26406 -11296 -26353
rect -11409 -26419 -11296 -26406
rect -11409 -26449 -11274 -26419
rect -11144 -26449 -11118 -26419
rect -11733 -26498 -11474 -26449
rect -11733 -26511 -11299 -26498
rect 11835 -25159 11865 -25133
rect 11931 -25159 11961 -25133
rect 12027 -25159 12057 -25133
rect 12123 -25159 12153 -25133
rect 12219 -25159 12249 -25133
rect 12315 -25159 12345 -25133
rect 12411 -25159 12441 -25133
rect 12507 -25159 12537 -25133
rect 12603 -25159 12633 -25133
rect 12699 -25159 12729 -25133
rect 12826 -25323 12892 -25307
rect 11835 -25441 11865 -25415
rect 11931 -25441 11961 -25415
rect 12027 -25441 12057 -25415
rect 12123 -25441 12153 -25415
rect 12219 -25441 12249 -25415
rect 11835 -25465 12249 -25441
rect 7422 -25504 7452 -25478
rect 7518 -25504 7548 -25478
rect 7614 -25504 7644 -25478
rect 7710 -25504 7740 -25478
rect 8370 -25504 8400 -25478
rect 8466 -25504 8496 -25478
rect 8562 -25504 8592 -25478
rect 8658 -25504 8688 -25478
rect 9306 -25504 9336 -25478
rect 9402 -25504 9432 -25478
rect 9498 -25504 9528 -25478
rect 9594 -25504 9624 -25478
rect 10237 -25504 10267 -25478
rect 10333 -25504 10363 -25478
rect 10429 -25504 10459 -25478
rect 10525 -25504 10555 -25478
rect 11164 -25504 11194 -25478
rect 11260 -25504 11290 -25478
rect 11356 -25504 11386 -25478
rect 11452 -25504 11482 -25478
rect 11835 -25499 12170 -25465
rect 12204 -25499 12249 -25465
rect 11835 -25512 12249 -25499
rect 7422 -25606 7452 -25580
rect 7518 -25606 7548 -25580
rect 7614 -25606 7644 -25580
rect 7710 -25606 7740 -25580
rect 8370 -25606 8400 -25580
rect 8466 -25606 8496 -25580
rect 8562 -25606 8592 -25580
rect 8658 -25606 8688 -25580
rect 9306 -25606 9336 -25580
rect 9402 -25606 9432 -25580
rect 9498 -25606 9528 -25580
rect 9594 -25606 9624 -25580
rect 10237 -25605 10267 -25579
rect 10333 -25605 10363 -25579
rect 10429 -25605 10459 -25579
rect 10525 -25605 10555 -25579
rect 11164 -25606 11194 -25580
rect 11260 -25606 11290 -25580
rect 11356 -25606 11386 -25580
rect 11452 -25606 11482 -25580
rect 7422 -26439 7452 -26406
rect 7238 -26469 7452 -26439
rect -12340 -26541 -12314 -26511
rect -11764 -26541 -11274 -26511
rect -11144 -26541 -11118 -26511
rect -11733 -26574 -11299 -26541
rect -11583 -26635 -11474 -26574
rect -11576 -26758 -11480 -26635
rect 7238 -26716 7268 -26469
rect 7518 -26511 7548 -26406
rect 7614 -26429 7644 -26406
rect 7374 -26649 7548 -26511
rect -11576 -26810 -11554 -26758
rect -11502 -26810 -11480 -26758
rect 7182 -26732 7326 -26716
rect 7182 -26766 7198 -26732
rect 7232 -26766 7326 -26732
rect 7182 -26782 7326 -26766
rect 7374 -26732 7518 -26649
rect 7590 -26691 7644 -26429
rect 7710 -26556 7740 -26406
rect 8370 -26439 8400 -26406
rect 8186 -26469 8400 -26439
rect 7710 -26586 7848 -26556
rect 7584 -26716 7644 -26691
rect 7758 -26716 7848 -26586
rect 8186 -26716 8216 -26469
rect 8466 -26511 8496 -26406
rect 8562 -26429 8592 -26406
rect 8322 -26649 8496 -26511
rect 7374 -26766 7390 -26732
rect 7424 -26766 7518 -26732
rect 7374 -26782 7518 -26766
rect 7566 -26732 7710 -26716
rect 7566 -26766 7582 -26732
rect 7616 -26766 7710 -26732
rect 7566 -26782 7710 -26766
rect 7758 -26732 7902 -26716
rect 7758 -26766 7774 -26732
rect 7808 -26766 7902 -26732
rect 7758 -26782 7902 -26766
rect 8130 -26732 8274 -26716
rect 8130 -26766 8146 -26732
rect 8180 -26766 8274 -26732
rect 8130 -26782 8274 -26766
rect 8322 -26732 8466 -26649
rect 8538 -26691 8592 -26429
rect 8658 -26556 8688 -26406
rect 9306 -26439 9336 -26406
rect 9122 -26469 9336 -26439
rect 8658 -26586 8796 -26556
rect 8532 -26716 8592 -26691
rect 8706 -26716 8796 -26586
rect 9122 -26716 9152 -26469
rect 9402 -26511 9432 -26406
rect 9498 -26429 9528 -26406
rect 9258 -26649 9432 -26511
rect 8322 -26766 8338 -26732
rect 8372 -26766 8466 -26732
rect 8322 -26782 8466 -26766
rect 8514 -26732 8658 -26716
rect 8514 -26766 8530 -26732
rect 8564 -26766 8658 -26732
rect 8514 -26782 8658 -26766
rect 8706 -26732 8850 -26716
rect 8706 -26766 8722 -26732
rect 8756 -26766 8850 -26732
rect 8706 -26782 8850 -26766
rect 9066 -26732 9210 -26716
rect 9066 -26766 9082 -26732
rect 9116 -26766 9210 -26732
rect 9066 -26782 9210 -26766
rect 9258 -26732 9402 -26649
rect 9474 -26691 9528 -26429
rect 9594 -26556 9624 -26406
rect 10237 -26438 10267 -26405
rect 10053 -26468 10267 -26438
rect 9594 -26586 9732 -26556
rect 9468 -26716 9528 -26691
rect 9642 -26716 9732 -26586
rect 10053 -26715 10083 -26468
rect 10333 -26510 10363 -26405
rect 10429 -26428 10459 -26405
rect 10189 -26648 10363 -26510
rect 9258 -26766 9274 -26732
rect 9308 -26766 9402 -26732
rect 9258 -26782 9402 -26766
rect 9450 -26732 9594 -26716
rect 9450 -26766 9466 -26732
rect 9500 -26766 9594 -26732
rect 9450 -26782 9594 -26766
rect 9642 -26732 9786 -26716
rect 9642 -26766 9658 -26732
rect 9692 -26766 9786 -26732
rect 9642 -26782 9786 -26766
rect 9997 -26731 10141 -26715
rect 9997 -26765 10013 -26731
rect 10047 -26765 10141 -26731
rect 9997 -26781 10141 -26765
rect 10189 -26731 10333 -26648
rect 10405 -26690 10459 -26428
rect 10525 -26555 10555 -26405
rect 12219 -25648 12249 -25512
rect 12315 -25441 12345 -25415
rect 12411 -25441 12441 -25415
rect 12507 -25441 12537 -25415
rect 12603 -25441 12633 -25415
rect 12699 -25441 12729 -25415
rect 12315 -25512 12729 -25441
rect 12315 -25554 12345 -25512
rect 12826 -25549 12842 -25323
rect 12876 -25325 12892 -25323
rect 12876 -25355 12923 -25325
rect 13137 -25355 13163 -25325
rect 12876 -25421 12892 -25355
rect 12876 -25451 12923 -25421
rect 13137 -25451 13163 -25421
rect 12876 -25517 12892 -25451
rect 12876 -25547 12923 -25517
rect 13137 -25547 13163 -25517
rect 12876 -25549 12892 -25547
rect 12297 -25570 12363 -25554
rect 12826 -25565 12892 -25549
rect 12297 -25604 12313 -25570
rect 12347 -25604 12363 -25570
rect 12297 -25620 12363 -25604
rect 12315 -25648 12345 -25620
rect 12826 -25769 12893 -25753
rect 12826 -25803 12842 -25769
rect 12876 -25771 12893 -25769
rect 12876 -25801 12923 -25771
rect 13123 -25801 13149 -25771
rect 12876 -25803 12893 -25801
rect 12826 -25819 12893 -25803
rect 12219 -25874 12249 -25848
rect 12315 -25874 12345 -25848
rect 11164 -26439 11194 -26406
rect 10980 -26469 11194 -26439
rect 10525 -26585 10663 -26555
rect 10399 -26715 10459 -26690
rect 10573 -26715 10663 -26585
rect 10189 -26765 10205 -26731
rect 10239 -26765 10333 -26731
rect 10189 -26781 10333 -26765
rect 10381 -26731 10525 -26715
rect 10381 -26765 10397 -26731
rect 10431 -26765 10525 -26731
rect 10381 -26781 10525 -26765
rect 10573 -26731 10717 -26715
rect 10980 -26716 11010 -26469
rect 11260 -26511 11290 -26406
rect 11356 -26429 11386 -26406
rect 11116 -26649 11290 -26511
rect 10573 -26765 10589 -26731
rect 10623 -26765 10717 -26731
rect 10573 -26781 10717 -26765
rect -11576 -26832 -11480 -26810
rect 7200 -26813 7230 -26782
rect 7296 -26813 7326 -26782
rect 7392 -26813 7422 -26782
rect 7488 -26813 7518 -26782
rect 7584 -26813 7614 -26782
rect 7680 -26813 7710 -26782
rect 7776 -26813 7806 -26782
rect 7872 -26813 7902 -26782
rect 8148 -26813 8178 -26782
rect 8244 -26813 8274 -26782
rect 8340 -26813 8370 -26782
rect 8436 -26813 8466 -26782
rect 8532 -26813 8562 -26782
rect 8628 -26813 8658 -26782
rect 8724 -26813 8754 -26782
rect 8820 -26813 8850 -26782
rect 9084 -26813 9114 -26782
rect 9180 -26813 9210 -26782
rect 9276 -26813 9306 -26782
rect 9372 -26813 9402 -26782
rect 9468 -26813 9498 -26782
rect 9564 -26813 9594 -26782
rect 9660 -26813 9690 -26782
rect 9756 -26813 9786 -26782
rect 10015 -26812 10045 -26781
rect 10111 -26812 10141 -26781
rect 10207 -26812 10237 -26781
rect 10303 -26812 10333 -26781
rect 10399 -26812 10429 -26781
rect 10495 -26812 10525 -26781
rect 10591 -26812 10621 -26781
rect 10687 -26812 10717 -26781
rect 10924 -26732 11068 -26716
rect 10924 -26766 10940 -26732
rect 10974 -26766 11068 -26732
rect 10924 -26782 11068 -26766
rect 11116 -26732 11260 -26649
rect 11332 -26691 11386 -26429
rect 11452 -26556 11482 -26406
rect 11452 -26586 11590 -26556
rect 11326 -26716 11386 -26691
rect 11500 -26716 11590 -26586
rect 11116 -26766 11132 -26732
rect 11166 -26766 11260 -26732
rect 11116 -26782 11260 -26766
rect 11308 -26732 11452 -26716
rect 11308 -26766 11324 -26732
rect 11358 -26766 11452 -26732
rect 11308 -26782 11452 -26766
rect 11500 -26732 11644 -26716
rect 11500 -26766 11516 -26732
rect 11550 -26766 11644 -26732
rect 11500 -26782 11644 -26766
rect 10942 -26813 10972 -26782
rect 11038 -26813 11068 -26782
rect 11134 -26813 11164 -26782
rect 11230 -26813 11260 -26782
rect 11326 -26813 11356 -26782
rect 11422 -26813 11452 -26782
rect 11518 -26813 11548 -26782
rect 11614 -26813 11644 -26782
rect 7200 -27161 7230 -27135
rect 7296 -27161 7326 -27135
rect 7392 -27161 7422 -27135
rect 7488 -27161 7518 -27135
rect 7584 -27161 7614 -27135
rect 7680 -27161 7710 -27135
rect 7776 -27161 7806 -27135
rect 7872 -27161 7902 -27135
rect 8148 -27161 8178 -27135
rect 8244 -27161 8274 -27135
rect 8340 -27161 8370 -27135
rect 8436 -27161 8466 -27135
rect 8532 -27161 8562 -27135
rect 8628 -27161 8658 -27135
rect 8724 -27161 8754 -27135
rect 8820 -27161 8850 -27135
rect 9084 -27161 9114 -27135
rect 9180 -27161 9210 -27135
rect 9276 -27161 9306 -27135
rect 9372 -27161 9402 -27135
rect 9468 -27161 9498 -27135
rect 9564 -27161 9594 -27135
rect 9660 -27161 9690 -27135
rect 9756 -27161 9786 -27135
rect 10015 -27160 10045 -27134
rect 10111 -27160 10141 -27134
rect 10207 -27160 10237 -27134
rect 10303 -27160 10333 -27134
rect 10399 -27160 10429 -27134
rect 10495 -27160 10525 -27134
rect 10591 -27160 10621 -27134
rect 10687 -27160 10717 -27134
rect 10942 -27161 10972 -27135
rect 11038 -27161 11068 -27135
rect 11134 -27161 11164 -27135
rect 11230 -27161 11260 -27135
rect 11326 -27161 11356 -27135
rect 11422 -27161 11452 -27135
rect 11518 -27161 11548 -27135
rect 11614 -27161 11644 -27135
rect 5561 -27833 5627 -27817
rect -12340 -27934 -12314 -27904
rect -11764 -27934 -11274 -27904
rect -11144 -27934 -11118 -27904
rect -11733 -27996 -11296 -27934
rect -12345 -28026 -12314 -27996
rect -11764 -28026 -11274 -27996
rect -11144 -28026 -11118 -27996
rect -11733 -28092 -11296 -28026
rect -12345 -28122 -12314 -28092
rect -11764 -28121 -11274 -28092
rect -11764 -28122 -11576 -28121
rect -11733 -28186 -11576 -28122
rect -11521 -28122 -11274 -28121
rect -11144 -28122 -11118 -28092
rect -11521 -28186 -11296 -28122
rect -11733 -28188 -11296 -28186
rect -12345 -28218 -12314 -28188
rect -11764 -28218 -11274 -28188
rect -11144 -28218 -11118 -28188
rect -12345 -28314 -12314 -28284
rect -11764 -28303 -11640 -28284
rect -11764 -28314 -11700 -28303
rect -11733 -28380 -11700 -28314
rect -12345 -28410 -12314 -28380
rect -11764 -28410 -11700 -28380
rect -11733 -28433 -11700 -28410
rect -11655 -28433 -11640 -28303
rect -11733 -28476 -11640 -28433
rect -12345 -28506 -12314 -28476
rect -11764 -28506 -11640 -28476
rect -11583 -28314 -11274 -28284
rect -11144 -28314 -11118 -28284
rect -11583 -28380 -11296 -28314
rect -11583 -28410 -11274 -28380
rect -11144 -28410 -11118 -28380
rect -11583 -28476 -11296 -28410
rect -11583 -28506 -11274 -28476
rect -11144 -28506 -11118 -28476
rect -12345 -28602 -12314 -28572
rect -11764 -28602 -11641 -28572
rect -11734 -28634 -11641 -28602
rect -11734 -28668 -11705 -28634
rect -12345 -28698 -12314 -28668
rect -11764 -28698 -11705 -28668
rect -11734 -28764 -11705 -28698
rect -11660 -28764 -11641 -28634
rect -12345 -28794 -12314 -28764
rect -11764 -28794 -11641 -28764
rect -11583 -28858 -11474 -28506
rect -11404 -28602 -11274 -28572
rect -11144 -28602 -11118 -28572
rect -11404 -28626 -11296 -28602
rect -11404 -28756 -11376 -28626
rect -11331 -28668 -11296 -28626
rect -11331 -28698 -11274 -28668
rect -11144 -28698 -11118 -28668
rect -11331 -28756 -11296 -28698
rect -11404 -28764 -11296 -28756
rect -11404 -28794 -11274 -28764
rect -11144 -28794 -11118 -28764
rect -11733 -28860 -11474 -28858
rect -12345 -28890 -12314 -28860
rect -11764 -28890 -11474 -28860
rect -11733 -28956 -11474 -28890
rect -12345 -28986 -12314 -28956
rect -11764 -28986 -11474 -28956
rect -11733 -29052 -11474 -28986
rect -12345 -29082 -12314 -29052
rect -11764 -29082 -11474 -29052
rect -11409 -28890 -11274 -28860
rect -11144 -28890 -11118 -28860
rect -11409 -28909 -11296 -28890
rect -11409 -29039 -11384 -28909
rect -11339 -28956 -11296 -28909
rect -11339 -28986 -11274 -28956
rect -11144 -28986 -11118 -28956
rect -11339 -29039 -11296 -28986
rect -11409 -29052 -11296 -29039
rect -11409 -29082 -11274 -29052
rect -11144 -29082 -11118 -29052
rect -11733 -29131 -11474 -29082
rect -11733 -29144 -11299 -29131
rect 5561 -28059 5577 -27833
rect 5611 -27835 5627 -27833
rect 6001 -27833 6067 -27817
rect 5611 -27865 5658 -27835
rect 5872 -27865 5898 -27835
rect 5611 -27931 5627 -27865
rect 5611 -27961 5658 -27931
rect 5872 -27961 5898 -27931
rect 5611 -28027 5627 -27961
rect 5611 -28057 5658 -28027
rect 5872 -28057 5898 -28027
rect 5611 -28059 5627 -28057
rect 5561 -28075 5627 -28059
rect 6001 -28059 6017 -27833
rect 6051 -27835 6067 -27833
rect 6441 -27833 6507 -27817
rect 6051 -27865 6098 -27835
rect 6312 -27865 6338 -27835
rect 6051 -27931 6067 -27865
rect 6051 -27961 6098 -27931
rect 6312 -27961 6338 -27931
rect 6051 -28027 6067 -27961
rect 6051 -28057 6098 -28027
rect 6312 -28057 6338 -28027
rect 6051 -28059 6067 -28057
rect 6001 -28075 6067 -28059
rect 6441 -28059 6457 -27833
rect 6491 -27835 6507 -27833
rect 6491 -27865 6538 -27835
rect 6752 -27865 6778 -27835
rect 6491 -27931 6507 -27865
rect 6491 -27961 6538 -27931
rect 6752 -27961 6778 -27931
rect 6491 -28027 6507 -27961
rect 6491 -28057 6538 -28027
rect 6752 -28057 6778 -28027
rect 6491 -28059 6507 -28057
rect 6441 -28075 6507 -28059
rect 5561 -28279 5628 -28263
rect 5561 -28313 5577 -28279
rect 5611 -28281 5628 -28279
rect 6001 -28279 6068 -28263
rect 5611 -28311 5658 -28281
rect 5858 -28311 5884 -28281
rect 5611 -28313 5628 -28311
rect 5561 -28329 5628 -28313
rect 6001 -28313 6017 -28279
rect 6051 -28281 6068 -28279
rect 6441 -28279 6508 -28263
rect 6051 -28311 6098 -28281
rect 6298 -28311 6324 -28281
rect 6051 -28313 6068 -28311
rect 6001 -28329 6068 -28313
rect 6441 -28313 6457 -28279
rect 6491 -28281 6508 -28279
rect 6491 -28311 6538 -28281
rect 6738 -28311 6764 -28281
rect 6491 -28313 6508 -28311
rect 6441 -28329 6508 -28313
rect 7200 -28477 7230 -28451
rect 7296 -28477 7326 -28451
rect 7392 -28477 7422 -28451
rect 7488 -28477 7518 -28451
rect 7584 -28477 7614 -28451
rect 7680 -28477 7710 -28451
rect 7776 -28477 7806 -28451
rect 7872 -28477 7902 -28451
rect 8148 -28477 8178 -28451
rect 8244 -28477 8274 -28451
rect 8340 -28477 8370 -28451
rect 8436 -28477 8466 -28451
rect 8532 -28477 8562 -28451
rect 8628 -28477 8658 -28451
rect 8724 -28477 8754 -28451
rect 8820 -28477 8850 -28451
rect 9084 -28477 9114 -28451
rect 9180 -28477 9210 -28451
rect 9276 -28477 9306 -28451
rect 9372 -28477 9402 -28451
rect 9468 -28477 9498 -28451
rect 9564 -28477 9594 -28451
rect 9660 -28477 9690 -28451
rect 9756 -28477 9786 -28451
rect 10015 -28477 10045 -28451
rect 10111 -28477 10141 -28451
rect 10207 -28477 10237 -28451
rect 10303 -28477 10333 -28451
rect 10399 -28477 10429 -28451
rect 10495 -28477 10525 -28451
rect 10591 -28477 10621 -28451
rect 10687 -28477 10717 -28451
rect 10942 -28477 10972 -28451
rect 11038 -28477 11068 -28451
rect 11134 -28477 11164 -28451
rect 11230 -28477 11260 -28451
rect 11326 -28477 11356 -28451
rect 11422 -28477 11452 -28451
rect 11518 -28477 11548 -28451
rect 11614 -28477 11644 -28451
rect 7200 -28830 7230 -28799
rect 7296 -28830 7326 -28799
rect 7392 -28830 7422 -28799
rect 7488 -28830 7518 -28799
rect 7584 -28830 7614 -28799
rect 7680 -28830 7710 -28799
rect 7776 -28830 7806 -28799
rect 7872 -28830 7902 -28799
rect 8148 -28830 8178 -28799
rect 8244 -28830 8274 -28799
rect 8340 -28830 8370 -28799
rect 8436 -28830 8466 -28799
rect 8532 -28830 8562 -28799
rect 8628 -28830 8658 -28799
rect 8724 -28830 8754 -28799
rect 8820 -28830 8850 -28799
rect 9084 -28830 9114 -28799
rect 9180 -28830 9210 -28799
rect 9276 -28830 9306 -28799
rect 9372 -28830 9402 -28799
rect 9468 -28830 9498 -28799
rect 9564 -28830 9594 -28799
rect 9660 -28830 9690 -28799
rect 9756 -28830 9786 -28799
rect 10015 -28830 10045 -28799
rect 10111 -28830 10141 -28799
rect 10207 -28830 10237 -28799
rect 10303 -28830 10333 -28799
rect 10399 -28830 10429 -28799
rect 10495 -28830 10525 -28799
rect 10591 -28830 10621 -28799
rect 10687 -28830 10717 -28799
rect 10942 -28830 10972 -28799
rect 11038 -28830 11068 -28799
rect 11134 -28830 11164 -28799
rect 11230 -28830 11260 -28799
rect 11326 -28830 11356 -28799
rect 11422 -28830 11452 -28799
rect 11518 -28830 11548 -28799
rect 11614 -28830 11644 -28799
rect 7182 -28846 7326 -28830
rect 7182 -28880 7198 -28846
rect 7232 -28880 7326 -28846
rect 7182 -28896 7326 -28880
rect 7374 -28846 7518 -28830
rect 7374 -28880 7390 -28846
rect 7424 -28880 7518 -28846
rect 7238 -29143 7268 -28896
rect 7374 -28963 7518 -28880
rect 7566 -28846 7710 -28830
rect 7566 -28880 7582 -28846
rect 7616 -28880 7710 -28846
rect 7566 -28896 7710 -28880
rect 7758 -28846 7902 -28830
rect 7758 -28880 7774 -28846
rect 7808 -28880 7902 -28846
rect 7758 -28896 7902 -28880
rect 8130 -28846 8274 -28830
rect 8130 -28880 8146 -28846
rect 8180 -28880 8274 -28846
rect 8130 -28896 8274 -28880
rect 8322 -28846 8466 -28830
rect 8322 -28880 8338 -28846
rect 8372 -28880 8466 -28846
rect 7584 -28921 7644 -28896
rect 7374 -29101 7548 -28963
rect -12340 -29174 -12314 -29144
rect -11764 -29174 -11274 -29144
rect -11144 -29174 -11118 -29144
rect 7238 -29173 7452 -29143
rect -11733 -29207 -11299 -29174
rect -11583 -29268 -11474 -29207
rect 7422 -29206 7452 -29173
rect 7518 -29206 7548 -29101
rect 7590 -29183 7644 -28921
rect 7758 -29026 7848 -28896
rect 7614 -29206 7644 -29183
rect 7710 -29056 7848 -29026
rect 7710 -29206 7740 -29056
rect 8186 -29143 8216 -28896
rect 8322 -28963 8466 -28880
rect 8514 -28846 8658 -28830
rect 8514 -28880 8530 -28846
rect 8564 -28880 8658 -28846
rect 8514 -28896 8658 -28880
rect 8706 -28846 8850 -28830
rect 8706 -28880 8722 -28846
rect 8756 -28880 8850 -28846
rect 8706 -28896 8850 -28880
rect 9066 -28846 9210 -28830
rect 9066 -28880 9082 -28846
rect 9116 -28880 9210 -28846
rect 9066 -28896 9210 -28880
rect 9258 -28846 9402 -28830
rect 9258 -28880 9274 -28846
rect 9308 -28880 9402 -28846
rect 8532 -28921 8592 -28896
rect 8322 -29101 8496 -28963
rect 8186 -29173 8400 -29143
rect 8370 -29206 8400 -29173
rect 8466 -29206 8496 -29101
rect 8538 -29183 8592 -28921
rect 8706 -29026 8796 -28896
rect 8562 -29206 8592 -29183
rect 8658 -29056 8796 -29026
rect 8658 -29206 8688 -29056
rect 9122 -29143 9152 -28896
rect 9258 -28963 9402 -28880
rect 9450 -28846 9594 -28830
rect 9450 -28880 9466 -28846
rect 9500 -28880 9594 -28846
rect 9450 -28896 9594 -28880
rect 9642 -28846 9786 -28830
rect 9642 -28880 9658 -28846
rect 9692 -28880 9786 -28846
rect 9642 -28896 9786 -28880
rect 9997 -28846 10141 -28830
rect 9997 -28880 10013 -28846
rect 10047 -28880 10141 -28846
rect 9997 -28896 10141 -28880
rect 10189 -28846 10333 -28830
rect 10189 -28880 10205 -28846
rect 10239 -28880 10333 -28846
rect 9468 -28921 9528 -28896
rect 9258 -29101 9432 -28963
rect 9122 -29173 9336 -29143
rect 9306 -29206 9336 -29173
rect 9402 -29206 9432 -29101
rect 9474 -29183 9528 -28921
rect 9642 -29026 9732 -28896
rect 9498 -29206 9528 -29183
rect 9594 -29056 9732 -29026
rect 9594 -29206 9624 -29056
rect 10053 -29143 10083 -28896
rect 10189 -28963 10333 -28880
rect 10381 -28846 10525 -28830
rect 10381 -28880 10397 -28846
rect 10431 -28880 10525 -28846
rect 10381 -28896 10525 -28880
rect 10573 -28846 10717 -28830
rect 10573 -28880 10589 -28846
rect 10623 -28880 10717 -28846
rect 10573 -28896 10717 -28880
rect 10924 -28846 11068 -28830
rect 10924 -28880 10940 -28846
rect 10974 -28880 11068 -28846
rect 10924 -28896 11068 -28880
rect 11116 -28846 11260 -28830
rect 11116 -28880 11132 -28846
rect 11166 -28880 11260 -28846
rect 10399 -28921 10459 -28896
rect 10189 -29101 10363 -28963
rect 10053 -29173 10267 -29143
rect 10237 -29206 10267 -29173
rect 10333 -29206 10363 -29101
rect 10405 -29183 10459 -28921
rect 10573 -29026 10663 -28896
rect 10429 -29206 10459 -29183
rect 10525 -29056 10663 -29026
rect 10525 -29206 10555 -29056
rect 10980 -29143 11010 -28896
rect 11116 -28963 11260 -28880
rect 11308 -28846 11452 -28830
rect 11308 -28880 11324 -28846
rect 11358 -28880 11452 -28846
rect 11308 -28896 11452 -28880
rect 11500 -28846 11644 -28830
rect 11500 -28880 11516 -28846
rect 11550 -28880 11644 -28846
rect 11500 -28896 11644 -28880
rect 11326 -28921 11386 -28896
rect 11116 -29101 11290 -28963
rect 10980 -29173 11194 -29143
rect 11164 -29206 11194 -29173
rect 11260 -29206 11290 -29101
rect 11332 -29183 11386 -28921
rect 11500 -29026 11590 -28896
rect 11356 -29206 11386 -29183
rect 11452 -29056 11590 -29026
rect 11452 -29206 11482 -29056
rect -11575 -29395 -11482 -29268
rect -11575 -29443 -11552 -29395
rect -11504 -29443 -11482 -29395
rect -11575 -29465 -11482 -29443
rect 11835 -29687 11865 -29661
rect 11931 -29687 11961 -29661
rect 12027 -29687 12057 -29661
rect 12123 -29687 12153 -29661
rect 12219 -29687 12249 -29661
rect 12315 -29687 12345 -29661
rect 12411 -29687 12441 -29661
rect 12507 -29687 12537 -29661
rect 12603 -29687 12633 -29661
rect 12699 -29687 12729 -29661
rect 12826 -29851 12892 -29835
rect 11835 -29969 11865 -29943
rect 11931 -29969 11961 -29943
rect 12027 -29969 12057 -29943
rect 12123 -29969 12153 -29943
rect 12219 -29969 12249 -29943
rect 11835 -29993 12249 -29969
rect 7422 -30032 7452 -30006
rect 7518 -30032 7548 -30006
rect 7614 -30032 7644 -30006
rect 7710 -30032 7740 -30006
rect 8370 -30032 8400 -30006
rect 8466 -30032 8496 -30006
rect 8562 -30032 8592 -30006
rect 8658 -30032 8688 -30006
rect 9306 -30032 9336 -30006
rect 9402 -30032 9432 -30006
rect 9498 -30032 9528 -30006
rect 9594 -30032 9624 -30006
rect 10237 -30032 10267 -30006
rect 10333 -30032 10363 -30006
rect 10429 -30032 10459 -30006
rect 10525 -30032 10555 -30006
rect 11164 -30032 11194 -30006
rect 11260 -30032 11290 -30006
rect 11356 -30032 11386 -30006
rect 11452 -30032 11482 -30006
rect 11835 -30027 12170 -29993
rect 12204 -30027 12249 -29993
rect 11835 -30040 12249 -30027
rect 7422 -30134 7452 -30108
rect 7518 -30134 7548 -30108
rect 7614 -30134 7644 -30108
rect 7710 -30134 7740 -30108
rect 8370 -30134 8400 -30108
rect 8466 -30134 8496 -30108
rect 8562 -30134 8592 -30108
rect 8658 -30134 8688 -30108
rect 9306 -30134 9336 -30108
rect 9402 -30134 9432 -30108
rect 9498 -30134 9528 -30108
rect 9594 -30134 9624 -30108
rect 10237 -30133 10267 -30107
rect 10333 -30133 10363 -30107
rect 10429 -30133 10459 -30107
rect 10525 -30133 10555 -30107
rect -12340 -30543 -12314 -30513
rect -11764 -30543 -11274 -30513
rect -11144 -30543 -11118 -30513
rect -11733 -30605 -11296 -30543
rect -12345 -30635 -12314 -30605
rect -11764 -30635 -11274 -30605
rect -11144 -30635 -11118 -30605
rect -11733 -30701 -11296 -30635
rect -12345 -30731 -12314 -30701
rect -11764 -30730 -11274 -30701
rect -11764 -30731 -11576 -30730
rect -11733 -30795 -11576 -30731
rect -11521 -30731 -11274 -30730
rect -11144 -30731 -11118 -30701
rect -11521 -30795 -11296 -30731
rect -11733 -30797 -11296 -30795
rect -12345 -30827 -12314 -30797
rect -11764 -30827 -11274 -30797
rect -11144 -30827 -11118 -30797
rect -12345 -30923 -12314 -30893
rect -11764 -30912 -11640 -30893
rect -11764 -30923 -11700 -30912
rect -11733 -30989 -11700 -30923
rect -12345 -31019 -12314 -30989
rect -11764 -31019 -11700 -30989
rect -11733 -31042 -11700 -31019
rect -11655 -31042 -11640 -30912
rect -11733 -31085 -11640 -31042
rect -12345 -31115 -12314 -31085
rect -11764 -31115 -11640 -31085
rect -11583 -30923 -11274 -30893
rect -11144 -30923 -11118 -30893
rect -11583 -30989 -11296 -30923
rect -11583 -31019 -11274 -30989
rect -11144 -31019 -11118 -30989
rect -11583 -31085 -11296 -31019
rect -11583 -31115 -11274 -31085
rect -11144 -31115 -11118 -31085
rect -12345 -31211 -12314 -31181
rect -11764 -31211 -11641 -31181
rect -11734 -31243 -11641 -31211
rect -11734 -31277 -11705 -31243
rect -12345 -31307 -12314 -31277
rect -11764 -31307 -11705 -31277
rect -11734 -31373 -11705 -31307
rect -11660 -31373 -11641 -31243
rect -12345 -31403 -12314 -31373
rect -11764 -31403 -11641 -31373
rect -11583 -31467 -11474 -31115
rect -11404 -31211 -11274 -31181
rect -11144 -31211 -11118 -31181
rect -11404 -31235 -11296 -31211
rect -11404 -31365 -11376 -31235
rect -11331 -31277 -11296 -31235
rect -11331 -31307 -11274 -31277
rect -11144 -31307 -11118 -31277
rect -11331 -31365 -11296 -31307
rect -11404 -31373 -11296 -31365
rect -11404 -31403 -11274 -31373
rect -11144 -31403 -11118 -31373
rect -11733 -31469 -11474 -31467
rect -12345 -31499 -12314 -31469
rect -11764 -31499 -11474 -31469
rect -11733 -31565 -11474 -31499
rect -12345 -31595 -12314 -31565
rect -11764 -31595 -11474 -31565
rect -11733 -31661 -11474 -31595
rect -12345 -31691 -12314 -31661
rect -11764 -31691 -11474 -31661
rect -11409 -31499 -11274 -31469
rect -11144 -31499 -11118 -31469
rect -11409 -31518 -11296 -31499
rect -11409 -31648 -11384 -31518
rect -11339 -31565 -11296 -31518
rect -11339 -31595 -11274 -31565
rect -11144 -31595 -11118 -31565
rect -11339 -31648 -11296 -31595
rect -11409 -31661 -11296 -31648
rect -11409 -31691 -11274 -31661
rect -11144 -31691 -11118 -31661
rect -11733 -31740 -11474 -31691
rect -11733 -31753 -11299 -31740
rect 11164 -30134 11194 -30108
rect 11260 -30134 11290 -30108
rect 11356 -30134 11386 -30108
rect 11452 -30134 11482 -30108
rect 7422 -30967 7452 -30934
rect 7238 -30997 7452 -30967
rect 7238 -31244 7268 -30997
rect 7518 -31039 7548 -30934
rect 7614 -30957 7644 -30934
rect 7374 -31177 7548 -31039
rect 7182 -31260 7326 -31244
rect 7182 -31294 7198 -31260
rect 7232 -31294 7326 -31260
rect 7182 -31310 7326 -31294
rect 7374 -31260 7518 -31177
rect 7590 -31219 7644 -30957
rect 7710 -31084 7740 -30934
rect 8370 -30967 8400 -30934
rect 8186 -30997 8400 -30967
rect 7710 -31114 7848 -31084
rect 7584 -31244 7644 -31219
rect 7758 -31244 7848 -31114
rect 8186 -31244 8216 -30997
rect 8466 -31039 8496 -30934
rect 8562 -30957 8592 -30934
rect 8322 -31177 8496 -31039
rect 7374 -31294 7390 -31260
rect 7424 -31294 7518 -31260
rect 7374 -31310 7518 -31294
rect 7566 -31260 7710 -31244
rect 7566 -31294 7582 -31260
rect 7616 -31294 7710 -31260
rect 7566 -31310 7710 -31294
rect 7758 -31260 7902 -31244
rect 7758 -31294 7774 -31260
rect 7808 -31294 7902 -31260
rect 7758 -31310 7902 -31294
rect 8130 -31260 8274 -31244
rect 8130 -31294 8146 -31260
rect 8180 -31294 8274 -31260
rect 8130 -31310 8274 -31294
rect 8322 -31260 8466 -31177
rect 8538 -31219 8592 -30957
rect 8658 -31084 8688 -30934
rect 9306 -30967 9336 -30934
rect 9122 -30997 9336 -30967
rect 8658 -31114 8796 -31084
rect 8532 -31244 8592 -31219
rect 8706 -31244 8796 -31114
rect 9122 -31244 9152 -30997
rect 9402 -31039 9432 -30934
rect 9498 -30957 9528 -30934
rect 9258 -31177 9432 -31039
rect 8322 -31294 8338 -31260
rect 8372 -31294 8466 -31260
rect 8322 -31310 8466 -31294
rect 8514 -31260 8658 -31244
rect 8514 -31294 8530 -31260
rect 8564 -31294 8658 -31260
rect 8514 -31310 8658 -31294
rect 8706 -31260 8850 -31244
rect 8706 -31294 8722 -31260
rect 8756 -31294 8850 -31260
rect 8706 -31310 8850 -31294
rect 9066 -31260 9210 -31244
rect 9066 -31294 9082 -31260
rect 9116 -31294 9210 -31260
rect 9066 -31310 9210 -31294
rect 9258 -31260 9402 -31177
rect 9474 -31219 9528 -30957
rect 9594 -31084 9624 -30934
rect 10237 -30966 10267 -30933
rect 10053 -30996 10267 -30966
rect 9594 -31114 9732 -31084
rect 9468 -31244 9528 -31219
rect 9642 -31244 9732 -31114
rect 10053 -31243 10083 -30996
rect 10333 -31038 10363 -30933
rect 10429 -30956 10459 -30933
rect 10189 -31176 10363 -31038
rect 9258 -31294 9274 -31260
rect 9308 -31294 9402 -31260
rect 9258 -31310 9402 -31294
rect 9450 -31260 9594 -31244
rect 9450 -31294 9466 -31260
rect 9500 -31294 9594 -31260
rect 9450 -31310 9594 -31294
rect 9642 -31260 9786 -31244
rect 9642 -31294 9658 -31260
rect 9692 -31294 9786 -31260
rect 9642 -31310 9786 -31294
rect 9997 -31259 10141 -31243
rect 9997 -31293 10013 -31259
rect 10047 -31293 10141 -31259
rect 9997 -31309 10141 -31293
rect 10189 -31259 10333 -31176
rect 10405 -31218 10459 -30956
rect 10525 -31083 10555 -30933
rect 12219 -30176 12249 -30040
rect 12315 -29969 12345 -29943
rect 12411 -29969 12441 -29943
rect 12507 -29969 12537 -29943
rect 12603 -29969 12633 -29943
rect 12699 -29969 12729 -29943
rect 12315 -30040 12729 -29969
rect 12315 -30082 12345 -30040
rect 12826 -30077 12842 -29851
rect 12876 -29853 12892 -29851
rect 12876 -29883 12923 -29853
rect 13137 -29883 13163 -29853
rect 12876 -29949 12892 -29883
rect 12876 -29979 12923 -29949
rect 13137 -29979 13163 -29949
rect 12876 -30045 12892 -29979
rect 12876 -30075 12923 -30045
rect 13137 -30075 13163 -30045
rect 12876 -30077 12892 -30075
rect 12297 -30098 12363 -30082
rect 12826 -30093 12892 -30077
rect 12297 -30132 12313 -30098
rect 12347 -30132 12363 -30098
rect 12297 -30148 12363 -30132
rect 12315 -30176 12345 -30148
rect 12826 -30297 12893 -30281
rect 12826 -30331 12842 -30297
rect 12876 -30299 12893 -30297
rect 12876 -30329 12923 -30299
rect 13123 -30329 13149 -30299
rect 12876 -30331 12893 -30329
rect 12826 -30347 12893 -30331
rect 12219 -30402 12249 -30376
rect 12315 -30402 12345 -30376
rect 11164 -30967 11194 -30934
rect 10980 -30997 11194 -30967
rect 10525 -31113 10663 -31083
rect 10399 -31243 10459 -31218
rect 10573 -31243 10663 -31113
rect 10189 -31293 10205 -31259
rect 10239 -31293 10333 -31259
rect 10189 -31309 10333 -31293
rect 10381 -31259 10525 -31243
rect 10381 -31293 10397 -31259
rect 10431 -31293 10525 -31259
rect 10381 -31309 10525 -31293
rect 10573 -31259 10717 -31243
rect 10980 -31244 11010 -30997
rect 11260 -31039 11290 -30934
rect 11356 -30957 11386 -30934
rect 11116 -31177 11290 -31039
rect 10573 -31293 10589 -31259
rect 10623 -31293 10717 -31259
rect 10573 -31309 10717 -31293
rect 7200 -31341 7230 -31310
rect 7296 -31341 7326 -31310
rect 7392 -31341 7422 -31310
rect 7488 -31341 7518 -31310
rect 7584 -31341 7614 -31310
rect 7680 -31341 7710 -31310
rect 7776 -31341 7806 -31310
rect 7872 -31341 7902 -31310
rect 8148 -31341 8178 -31310
rect 8244 -31341 8274 -31310
rect 8340 -31341 8370 -31310
rect 8436 -31341 8466 -31310
rect 8532 -31341 8562 -31310
rect 8628 -31341 8658 -31310
rect 8724 -31341 8754 -31310
rect 8820 -31341 8850 -31310
rect 9084 -31341 9114 -31310
rect 9180 -31341 9210 -31310
rect 9276 -31341 9306 -31310
rect 9372 -31341 9402 -31310
rect 9468 -31341 9498 -31310
rect 9564 -31341 9594 -31310
rect 9660 -31341 9690 -31310
rect 9756 -31341 9786 -31310
rect 10015 -31340 10045 -31309
rect 10111 -31340 10141 -31309
rect 10207 -31340 10237 -31309
rect 10303 -31340 10333 -31309
rect 10399 -31340 10429 -31309
rect 10495 -31340 10525 -31309
rect 10591 -31340 10621 -31309
rect 10687 -31340 10717 -31309
rect 10924 -31260 11068 -31244
rect 10924 -31294 10940 -31260
rect 10974 -31294 11068 -31260
rect 10924 -31310 11068 -31294
rect 11116 -31260 11260 -31177
rect 11332 -31219 11386 -30957
rect 11452 -31084 11482 -30934
rect 11452 -31114 11590 -31084
rect 11326 -31244 11386 -31219
rect 11500 -31244 11590 -31114
rect 11116 -31294 11132 -31260
rect 11166 -31294 11260 -31260
rect 11116 -31310 11260 -31294
rect 11308 -31260 11452 -31244
rect 11308 -31294 11324 -31260
rect 11358 -31294 11452 -31260
rect 11308 -31310 11452 -31294
rect 11500 -31260 11644 -31244
rect 11500 -31294 11516 -31260
rect 11550 -31294 11644 -31260
rect 11500 -31310 11644 -31294
rect 10942 -31341 10972 -31310
rect 11038 -31341 11068 -31310
rect 11134 -31341 11164 -31310
rect 11230 -31341 11260 -31310
rect 11326 -31341 11356 -31310
rect 11422 -31341 11452 -31310
rect 11518 -31341 11548 -31310
rect 11614 -31341 11644 -31310
rect 7200 -31689 7230 -31663
rect 7296 -31689 7326 -31663
rect 7392 -31689 7422 -31663
rect 7488 -31689 7518 -31663
rect 7584 -31689 7614 -31663
rect 7680 -31689 7710 -31663
rect 7776 -31689 7806 -31663
rect 7872 -31689 7902 -31663
rect 8148 -31689 8178 -31663
rect 8244 -31689 8274 -31663
rect 8340 -31689 8370 -31663
rect 8436 -31689 8466 -31663
rect 8532 -31689 8562 -31663
rect 8628 -31689 8658 -31663
rect 8724 -31689 8754 -31663
rect 8820 -31689 8850 -31663
rect 9084 -31689 9114 -31663
rect 9180 -31689 9210 -31663
rect 9276 -31689 9306 -31663
rect 9372 -31689 9402 -31663
rect 9468 -31689 9498 -31663
rect 9564 -31689 9594 -31663
rect 9660 -31689 9690 -31663
rect 9756 -31689 9786 -31663
rect 10015 -31688 10045 -31662
rect 10111 -31688 10141 -31662
rect 10207 -31688 10237 -31662
rect 10303 -31688 10333 -31662
rect 10399 -31688 10429 -31662
rect 10495 -31688 10525 -31662
rect 10591 -31688 10621 -31662
rect 10687 -31688 10717 -31662
rect 10942 -31689 10972 -31663
rect 11038 -31689 11068 -31663
rect 11134 -31689 11164 -31663
rect 11230 -31689 11260 -31663
rect 11326 -31689 11356 -31663
rect 11422 -31689 11452 -31663
rect 11518 -31689 11548 -31663
rect 11614 -31689 11644 -31663
rect -12340 -31783 -12314 -31753
rect -11764 -31783 -11274 -31753
rect -11144 -31783 -11118 -31753
rect -11733 -31816 -11299 -31783
rect -11583 -31937 -11474 -31816
rect -11583 -31988 -11554 -31937
rect -11503 -31988 -11474 -31937
rect -11583 -32010 -11474 -31988
rect 5561 -32361 5627 -32345
rect 5561 -32587 5577 -32361
rect 5611 -32363 5627 -32361
rect 6001 -32361 6067 -32345
rect 5611 -32393 5658 -32363
rect 5872 -32393 5898 -32363
rect 5611 -32459 5627 -32393
rect 5611 -32489 5658 -32459
rect 5872 -32489 5898 -32459
rect 5611 -32555 5627 -32489
rect 5611 -32585 5658 -32555
rect 5872 -32585 5898 -32555
rect 5611 -32587 5627 -32585
rect 5561 -32603 5627 -32587
rect 6001 -32587 6017 -32361
rect 6051 -32363 6067 -32361
rect 6441 -32361 6507 -32345
rect 6051 -32393 6098 -32363
rect 6312 -32393 6338 -32363
rect 6051 -32459 6067 -32393
rect 6051 -32489 6098 -32459
rect 6312 -32489 6338 -32459
rect 6051 -32555 6067 -32489
rect 6051 -32585 6098 -32555
rect 6312 -32585 6338 -32555
rect 6051 -32587 6067 -32585
rect 6001 -32603 6067 -32587
rect 6441 -32587 6457 -32361
rect 6491 -32363 6507 -32361
rect 6491 -32393 6538 -32363
rect 6752 -32393 6778 -32363
rect 6491 -32459 6507 -32393
rect 6491 -32489 6538 -32459
rect 6752 -32489 6778 -32459
rect 6491 -32555 6507 -32489
rect 6491 -32585 6538 -32555
rect 6752 -32585 6778 -32555
rect 6491 -32587 6507 -32585
rect 6441 -32603 6507 -32587
rect 5561 -32807 5628 -32791
rect 5561 -32841 5577 -32807
rect 5611 -32809 5628 -32807
rect 6001 -32807 6068 -32791
rect 5611 -32839 5658 -32809
rect 5858 -32839 5884 -32809
rect 5611 -32841 5628 -32839
rect 5561 -32857 5628 -32841
rect 6001 -32841 6017 -32807
rect 6051 -32809 6068 -32807
rect 6441 -32807 6508 -32791
rect 6051 -32839 6098 -32809
rect 6298 -32839 6324 -32809
rect 6051 -32841 6068 -32839
rect 6001 -32857 6068 -32841
rect 6441 -32841 6457 -32807
rect 6491 -32809 6508 -32807
rect 6491 -32839 6538 -32809
rect 6738 -32839 6764 -32809
rect 6491 -32841 6508 -32839
rect 6441 -32857 6508 -32841
rect 7200 -33005 7230 -32979
rect 7296 -33005 7326 -32979
rect 7392 -33005 7422 -32979
rect 7488 -33005 7518 -32979
rect 7584 -33005 7614 -32979
rect 7680 -33005 7710 -32979
rect 7776 -33005 7806 -32979
rect 7872 -33005 7902 -32979
rect 8148 -33005 8178 -32979
rect 8244 -33005 8274 -32979
rect 8340 -33005 8370 -32979
rect 8436 -33005 8466 -32979
rect 8532 -33005 8562 -32979
rect 8628 -33005 8658 -32979
rect 8724 -33005 8754 -32979
rect 8820 -33005 8850 -32979
rect 9084 -33005 9114 -32979
rect 9180 -33005 9210 -32979
rect 9276 -33005 9306 -32979
rect 9372 -33005 9402 -32979
rect 9468 -33005 9498 -32979
rect 9564 -33005 9594 -32979
rect 9660 -33005 9690 -32979
rect 9756 -33005 9786 -32979
rect 10015 -33005 10045 -32979
rect 10111 -33005 10141 -32979
rect 10207 -33005 10237 -32979
rect 10303 -33005 10333 -32979
rect 10399 -33005 10429 -32979
rect 10495 -33005 10525 -32979
rect 10591 -33005 10621 -32979
rect 10687 -33005 10717 -32979
rect 10942 -33005 10972 -32979
rect 11038 -33005 11068 -32979
rect 11134 -33005 11164 -32979
rect 11230 -33005 11260 -32979
rect 11326 -33005 11356 -32979
rect 11422 -33005 11452 -32979
rect 11518 -33005 11548 -32979
rect 11614 -33005 11644 -32979
rect -12342 -33163 -12316 -33133
rect -11766 -33163 -11276 -33133
rect -11146 -33163 -11120 -33133
rect -11735 -33225 -11298 -33163
rect -12347 -33255 -12316 -33225
rect -11766 -33255 -11276 -33225
rect -11146 -33255 -11120 -33225
rect -11735 -33321 -11298 -33255
rect -12347 -33351 -12316 -33321
rect -11766 -33350 -11276 -33321
rect -11766 -33351 -11578 -33350
rect -11735 -33415 -11578 -33351
rect -11523 -33351 -11276 -33350
rect -11146 -33351 -11120 -33321
rect -11523 -33415 -11298 -33351
rect -11735 -33417 -11298 -33415
rect -12347 -33447 -12316 -33417
rect -11766 -33447 -11276 -33417
rect -11146 -33447 -11120 -33417
rect -12347 -33543 -12316 -33513
rect -11766 -33532 -11642 -33513
rect -11766 -33543 -11702 -33532
rect -11735 -33609 -11702 -33543
rect -12347 -33639 -12316 -33609
rect -11766 -33639 -11702 -33609
rect -11735 -33662 -11702 -33639
rect -11657 -33662 -11642 -33532
rect -11735 -33705 -11642 -33662
rect -12347 -33735 -12316 -33705
rect -11766 -33735 -11642 -33705
rect -11585 -33543 -11276 -33513
rect -11146 -33543 -11120 -33513
rect -11585 -33609 -11298 -33543
rect -11585 -33639 -11276 -33609
rect -11146 -33639 -11120 -33609
rect -11585 -33705 -11298 -33639
rect -11585 -33735 -11276 -33705
rect -11146 -33735 -11120 -33705
rect -12347 -33831 -12316 -33801
rect -11766 -33831 -11643 -33801
rect -11736 -33863 -11643 -33831
rect -11736 -33897 -11707 -33863
rect -12347 -33927 -12316 -33897
rect -11766 -33927 -11707 -33897
rect -11736 -33993 -11707 -33927
rect -11662 -33993 -11643 -33863
rect -12347 -34023 -12316 -33993
rect -11766 -34023 -11643 -33993
rect -11585 -34087 -11476 -33735
rect -11406 -33831 -11276 -33801
rect -11146 -33831 -11120 -33801
rect -11406 -33855 -11298 -33831
rect -11406 -33985 -11378 -33855
rect -11333 -33897 -11298 -33855
rect -11333 -33927 -11276 -33897
rect -11146 -33927 -11120 -33897
rect -11333 -33985 -11298 -33927
rect -11406 -33993 -11298 -33985
rect -11406 -34023 -11276 -33993
rect -11146 -34023 -11120 -33993
rect -11735 -34089 -11476 -34087
rect -12347 -34119 -12316 -34089
rect -11766 -34119 -11476 -34089
rect -11735 -34185 -11476 -34119
rect -12347 -34215 -12316 -34185
rect -11766 -34215 -11476 -34185
rect -11735 -34281 -11476 -34215
rect -12347 -34311 -12316 -34281
rect -11766 -34311 -11476 -34281
rect -11411 -34119 -11276 -34089
rect -11146 -34119 -11120 -34089
rect -11411 -34138 -11298 -34119
rect -11411 -34268 -11386 -34138
rect -11341 -34185 -11298 -34138
rect -11341 -34215 -11276 -34185
rect -11146 -34215 -11120 -34185
rect -11341 -34268 -11298 -34215
rect -11411 -34281 -11298 -34268
rect -11411 -34311 -11276 -34281
rect -11146 -34311 -11120 -34281
rect -11735 -34360 -11476 -34311
rect -11735 -34373 -11301 -34360
rect 7200 -33358 7230 -33327
rect 7296 -33358 7326 -33327
rect 7392 -33358 7422 -33327
rect 7488 -33358 7518 -33327
rect 7584 -33358 7614 -33327
rect 7680 -33358 7710 -33327
rect 7776 -33358 7806 -33327
rect 7872 -33358 7902 -33327
rect 8148 -33358 8178 -33327
rect 8244 -33358 8274 -33327
rect 8340 -33358 8370 -33327
rect 8436 -33358 8466 -33327
rect 8532 -33358 8562 -33327
rect 8628 -33358 8658 -33327
rect 8724 -33358 8754 -33327
rect 8820 -33358 8850 -33327
rect 9084 -33358 9114 -33327
rect 9180 -33358 9210 -33327
rect 9276 -33358 9306 -33327
rect 9372 -33358 9402 -33327
rect 9468 -33358 9498 -33327
rect 9564 -33358 9594 -33327
rect 9660 -33358 9690 -33327
rect 9756 -33358 9786 -33327
rect 10015 -33358 10045 -33327
rect 10111 -33358 10141 -33327
rect 10207 -33358 10237 -33327
rect 10303 -33358 10333 -33327
rect 10399 -33358 10429 -33327
rect 10495 -33358 10525 -33327
rect 10591 -33358 10621 -33327
rect 10687 -33358 10717 -33327
rect 10942 -33358 10972 -33327
rect 11038 -33358 11068 -33327
rect 11134 -33358 11164 -33327
rect 11230 -33358 11260 -33327
rect 11326 -33358 11356 -33327
rect 11422 -33358 11452 -33327
rect 11518 -33358 11548 -33327
rect 11614 -33358 11644 -33327
rect 7182 -33374 7326 -33358
rect 7182 -33408 7198 -33374
rect 7232 -33408 7326 -33374
rect 7182 -33424 7326 -33408
rect 7374 -33374 7518 -33358
rect 7374 -33408 7390 -33374
rect 7424 -33408 7518 -33374
rect 7238 -33671 7268 -33424
rect 7374 -33491 7518 -33408
rect 7566 -33374 7710 -33358
rect 7566 -33408 7582 -33374
rect 7616 -33408 7710 -33374
rect 7566 -33424 7710 -33408
rect 7758 -33374 7902 -33358
rect 7758 -33408 7774 -33374
rect 7808 -33408 7902 -33374
rect 7758 -33424 7902 -33408
rect 8130 -33374 8274 -33358
rect 8130 -33408 8146 -33374
rect 8180 -33408 8274 -33374
rect 8130 -33424 8274 -33408
rect 8322 -33374 8466 -33358
rect 8322 -33408 8338 -33374
rect 8372 -33408 8466 -33374
rect 7584 -33449 7644 -33424
rect 7374 -33629 7548 -33491
rect 7238 -33701 7452 -33671
rect 7422 -33734 7452 -33701
rect 7518 -33734 7548 -33629
rect 7590 -33711 7644 -33449
rect 7758 -33554 7848 -33424
rect 7614 -33734 7644 -33711
rect 7710 -33584 7848 -33554
rect 7710 -33734 7740 -33584
rect 8186 -33671 8216 -33424
rect 8322 -33491 8466 -33408
rect 8514 -33374 8658 -33358
rect 8514 -33408 8530 -33374
rect 8564 -33408 8658 -33374
rect 8514 -33424 8658 -33408
rect 8706 -33374 8850 -33358
rect 8706 -33408 8722 -33374
rect 8756 -33408 8850 -33374
rect 8706 -33424 8850 -33408
rect 9066 -33374 9210 -33358
rect 9066 -33408 9082 -33374
rect 9116 -33408 9210 -33374
rect 9066 -33424 9210 -33408
rect 9258 -33374 9402 -33358
rect 9258 -33408 9274 -33374
rect 9308 -33408 9402 -33374
rect 8532 -33449 8592 -33424
rect 8322 -33629 8496 -33491
rect 8186 -33701 8400 -33671
rect 8370 -33734 8400 -33701
rect 8466 -33734 8496 -33629
rect 8538 -33711 8592 -33449
rect 8706 -33554 8796 -33424
rect 8562 -33734 8592 -33711
rect 8658 -33584 8796 -33554
rect 8658 -33734 8688 -33584
rect 9122 -33671 9152 -33424
rect 9258 -33491 9402 -33408
rect 9450 -33374 9594 -33358
rect 9450 -33408 9466 -33374
rect 9500 -33408 9594 -33374
rect 9450 -33424 9594 -33408
rect 9642 -33374 9786 -33358
rect 9642 -33408 9658 -33374
rect 9692 -33408 9786 -33374
rect 9642 -33424 9786 -33408
rect 9997 -33374 10141 -33358
rect 9997 -33408 10013 -33374
rect 10047 -33408 10141 -33374
rect 9997 -33424 10141 -33408
rect 10189 -33374 10333 -33358
rect 10189 -33408 10205 -33374
rect 10239 -33408 10333 -33374
rect 9468 -33449 9528 -33424
rect 9258 -33629 9432 -33491
rect 9122 -33701 9336 -33671
rect 9306 -33734 9336 -33701
rect 9402 -33734 9432 -33629
rect 9474 -33711 9528 -33449
rect 9642 -33554 9732 -33424
rect 9498 -33734 9528 -33711
rect 9594 -33584 9732 -33554
rect 9594 -33734 9624 -33584
rect 10053 -33671 10083 -33424
rect 10189 -33491 10333 -33408
rect 10381 -33374 10525 -33358
rect 10381 -33408 10397 -33374
rect 10431 -33408 10525 -33374
rect 10381 -33424 10525 -33408
rect 10573 -33374 10717 -33358
rect 10573 -33408 10589 -33374
rect 10623 -33408 10717 -33374
rect 10573 -33424 10717 -33408
rect 10924 -33374 11068 -33358
rect 10924 -33408 10940 -33374
rect 10974 -33408 11068 -33374
rect 10924 -33424 11068 -33408
rect 11116 -33374 11260 -33358
rect 11116 -33408 11132 -33374
rect 11166 -33408 11260 -33374
rect 10399 -33449 10459 -33424
rect 10189 -33629 10363 -33491
rect 10053 -33701 10267 -33671
rect 10237 -33734 10267 -33701
rect 10333 -33734 10363 -33629
rect 10405 -33711 10459 -33449
rect 10573 -33554 10663 -33424
rect 10429 -33734 10459 -33711
rect 10525 -33584 10663 -33554
rect 10525 -33734 10555 -33584
rect 10980 -33671 11010 -33424
rect 11116 -33491 11260 -33408
rect 11308 -33374 11452 -33358
rect 11308 -33408 11324 -33374
rect 11358 -33408 11452 -33374
rect 11308 -33424 11452 -33408
rect 11500 -33374 11644 -33358
rect 11500 -33408 11516 -33374
rect 11550 -33408 11644 -33374
rect 11500 -33424 11644 -33408
rect 11326 -33449 11386 -33424
rect 11116 -33629 11290 -33491
rect 10980 -33701 11194 -33671
rect 11164 -33734 11194 -33701
rect 11260 -33734 11290 -33629
rect 11332 -33711 11386 -33449
rect 11500 -33554 11590 -33424
rect 11356 -33734 11386 -33711
rect 11452 -33584 11590 -33554
rect 11452 -33734 11482 -33584
rect -12342 -34403 -12316 -34373
rect -11766 -34403 -11276 -34373
rect -11146 -34403 -11120 -34373
rect -11735 -34436 -11301 -34403
rect -11585 -34501 -11476 -34436
rect -11565 -34533 -11498 -34501
rect -11565 -34567 -11548 -34533
rect -11514 -34567 -11498 -34533
rect 11835 -34215 11865 -34189
rect 11931 -34215 11961 -34189
rect 12027 -34215 12057 -34189
rect 12123 -34215 12153 -34189
rect 12219 -34215 12249 -34189
rect 12315 -34215 12345 -34189
rect 12411 -34215 12441 -34189
rect 12507 -34215 12537 -34189
rect 12603 -34215 12633 -34189
rect 12699 -34215 12729 -34189
rect 12826 -34379 12892 -34363
rect 11835 -34497 11865 -34471
rect 11931 -34497 11961 -34471
rect 12027 -34497 12057 -34471
rect 12123 -34497 12153 -34471
rect 12219 -34497 12249 -34471
rect 11835 -34521 12249 -34497
rect 7422 -34560 7452 -34534
rect 7518 -34560 7548 -34534
rect 7614 -34560 7644 -34534
rect 7710 -34560 7740 -34534
rect 8370 -34560 8400 -34534
rect 8466 -34560 8496 -34534
rect 8562 -34560 8592 -34534
rect 8658 -34560 8688 -34534
rect 9306 -34560 9336 -34534
rect 9402 -34560 9432 -34534
rect 9498 -34560 9528 -34534
rect 9594 -34560 9624 -34534
rect 10237 -34560 10267 -34534
rect 10333 -34560 10363 -34534
rect 10429 -34560 10459 -34534
rect 10525 -34560 10555 -34534
rect 11164 -34560 11194 -34534
rect 11260 -34560 11290 -34534
rect 11356 -34560 11386 -34534
rect 11452 -34560 11482 -34534
rect 11835 -34555 12170 -34521
rect 12204 -34555 12249 -34521
rect -11565 -34583 -11498 -34567
rect 11835 -34568 12249 -34555
rect 7422 -34662 7452 -34636
rect 7518 -34662 7548 -34636
rect 7614 -34662 7644 -34636
rect 7710 -34662 7740 -34636
rect 8370 -34662 8400 -34636
rect 8466 -34662 8496 -34636
rect 8562 -34662 8592 -34636
rect 8658 -34662 8688 -34636
rect 9306 -34662 9336 -34636
rect 9402 -34662 9432 -34636
rect 9498 -34662 9528 -34636
rect 9594 -34662 9624 -34636
rect 10237 -34661 10267 -34635
rect 10333 -34661 10363 -34635
rect 10429 -34661 10459 -34635
rect 10525 -34661 10555 -34635
rect 11164 -34662 11194 -34636
rect 11260 -34662 11290 -34636
rect 11356 -34662 11386 -34636
rect 11452 -34662 11482 -34636
rect 7422 -35495 7452 -35462
rect 7238 -35525 7452 -35495
rect 7238 -35772 7268 -35525
rect 7518 -35567 7548 -35462
rect 7614 -35485 7644 -35462
rect 7374 -35705 7548 -35567
rect 7182 -35788 7326 -35772
rect 7182 -35822 7198 -35788
rect 7232 -35822 7326 -35788
rect 7182 -35838 7326 -35822
rect 7374 -35788 7518 -35705
rect 7590 -35747 7644 -35485
rect 7710 -35612 7740 -35462
rect 8370 -35495 8400 -35462
rect 8186 -35525 8400 -35495
rect 7710 -35642 7848 -35612
rect 7584 -35772 7644 -35747
rect 7758 -35772 7848 -35642
rect 8186 -35772 8216 -35525
rect 8466 -35567 8496 -35462
rect 8562 -35485 8592 -35462
rect 8322 -35705 8496 -35567
rect 7374 -35822 7390 -35788
rect 7424 -35822 7518 -35788
rect 7374 -35838 7518 -35822
rect 7566 -35788 7710 -35772
rect 7566 -35822 7582 -35788
rect 7616 -35822 7710 -35788
rect 7566 -35838 7710 -35822
rect 7758 -35788 7902 -35772
rect 7758 -35822 7774 -35788
rect 7808 -35822 7902 -35788
rect 7758 -35838 7902 -35822
rect 8130 -35788 8274 -35772
rect 8130 -35822 8146 -35788
rect 8180 -35822 8274 -35788
rect 8130 -35838 8274 -35822
rect 8322 -35788 8466 -35705
rect 8538 -35747 8592 -35485
rect 8658 -35612 8688 -35462
rect 9306 -35495 9336 -35462
rect 9122 -35525 9336 -35495
rect 8658 -35642 8796 -35612
rect 8532 -35772 8592 -35747
rect 8706 -35772 8796 -35642
rect 9122 -35772 9152 -35525
rect 9402 -35567 9432 -35462
rect 9498 -35485 9528 -35462
rect 9258 -35705 9432 -35567
rect 8322 -35822 8338 -35788
rect 8372 -35822 8466 -35788
rect 8322 -35838 8466 -35822
rect 8514 -35788 8658 -35772
rect 8514 -35822 8530 -35788
rect 8564 -35822 8658 -35788
rect 8514 -35838 8658 -35822
rect 8706 -35788 8850 -35772
rect 8706 -35822 8722 -35788
rect 8756 -35822 8850 -35788
rect 8706 -35838 8850 -35822
rect 9066 -35788 9210 -35772
rect 9066 -35822 9082 -35788
rect 9116 -35822 9210 -35788
rect 9066 -35838 9210 -35822
rect 9258 -35788 9402 -35705
rect 9474 -35747 9528 -35485
rect 9594 -35612 9624 -35462
rect 10237 -35494 10267 -35461
rect 10053 -35524 10267 -35494
rect 9594 -35642 9732 -35612
rect 9468 -35772 9528 -35747
rect 9642 -35772 9732 -35642
rect 10053 -35771 10083 -35524
rect 10333 -35566 10363 -35461
rect 10429 -35484 10459 -35461
rect 10189 -35704 10363 -35566
rect 9258 -35822 9274 -35788
rect 9308 -35822 9402 -35788
rect 9258 -35838 9402 -35822
rect 9450 -35788 9594 -35772
rect 9450 -35822 9466 -35788
rect 9500 -35822 9594 -35788
rect 9450 -35838 9594 -35822
rect 9642 -35788 9786 -35772
rect 9642 -35822 9658 -35788
rect 9692 -35822 9786 -35788
rect 9642 -35838 9786 -35822
rect 9997 -35787 10141 -35771
rect 9997 -35821 10013 -35787
rect 10047 -35821 10141 -35787
rect 9997 -35837 10141 -35821
rect 10189 -35787 10333 -35704
rect 10405 -35746 10459 -35484
rect 10525 -35611 10555 -35461
rect 12219 -34704 12249 -34568
rect 12315 -34497 12345 -34471
rect 12411 -34497 12441 -34471
rect 12507 -34497 12537 -34471
rect 12603 -34497 12633 -34471
rect 12699 -34497 12729 -34471
rect 12315 -34568 12729 -34497
rect 12315 -34610 12345 -34568
rect 12826 -34605 12842 -34379
rect 12876 -34381 12892 -34379
rect 12876 -34411 12923 -34381
rect 13137 -34411 13163 -34381
rect 12876 -34477 12892 -34411
rect 12876 -34507 12923 -34477
rect 13137 -34507 13163 -34477
rect 12876 -34573 12892 -34507
rect 12876 -34603 12923 -34573
rect 13137 -34603 13163 -34573
rect 12876 -34605 12892 -34603
rect 12297 -34626 12363 -34610
rect 12826 -34621 12892 -34605
rect 12297 -34660 12313 -34626
rect 12347 -34660 12363 -34626
rect 12297 -34676 12363 -34660
rect 12315 -34704 12345 -34676
rect 12826 -34825 12893 -34809
rect 12826 -34859 12842 -34825
rect 12876 -34827 12893 -34825
rect 12876 -34857 12923 -34827
rect 13123 -34857 13149 -34827
rect 12876 -34859 12893 -34857
rect 12826 -34875 12893 -34859
rect 12219 -34930 12249 -34904
rect 12315 -34930 12345 -34904
rect 11164 -35495 11194 -35462
rect 10980 -35525 11194 -35495
rect 10525 -35641 10663 -35611
rect 10399 -35771 10459 -35746
rect 10573 -35771 10663 -35641
rect 10189 -35821 10205 -35787
rect 10239 -35821 10333 -35787
rect 10189 -35837 10333 -35821
rect 10381 -35787 10525 -35771
rect 10381 -35821 10397 -35787
rect 10431 -35821 10525 -35787
rect 10381 -35837 10525 -35821
rect 10573 -35787 10717 -35771
rect 10980 -35772 11010 -35525
rect 11260 -35567 11290 -35462
rect 11356 -35485 11386 -35462
rect 11116 -35705 11290 -35567
rect 10573 -35821 10589 -35787
rect 10623 -35821 10717 -35787
rect 10573 -35837 10717 -35821
rect 7200 -35869 7230 -35838
rect 7296 -35869 7326 -35838
rect 7392 -35869 7422 -35838
rect 7488 -35869 7518 -35838
rect 7584 -35869 7614 -35838
rect 7680 -35869 7710 -35838
rect 7776 -35869 7806 -35838
rect 7872 -35869 7902 -35838
rect 8148 -35869 8178 -35838
rect 8244 -35869 8274 -35838
rect 8340 -35869 8370 -35838
rect 8436 -35869 8466 -35838
rect 8532 -35869 8562 -35838
rect 8628 -35869 8658 -35838
rect 8724 -35869 8754 -35838
rect 8820 -35869 8850 -35838
rect 9084 -35869 9114 -35838
rect 9180 -35869 9210 -35838
rect 9276 -35869 9306 -35838
rect 9372 -35869 9402 -35838
rect 9468 -35869 9498 -35838
rect 9564 -35869 9594 -35838
rect 9660 -35869 9690 -35838
rect 9756 -35869 9786 -35838
rect 10015 -35868 10045 -35837
rect 10111 -35868 10141 -35837
rect 10207 -35868 10237 -35837
rect 10303 -35868 10333 -35837
rect 10399 -35868 10429 -35837
rect 10495 -35868 10525 -35837
rect 10591 -35868 10621 -35837
rect 10687 -35868 10717 -35837
rect 10924 -35788 11068 -35772
rect 10924 -35822 10940 -35788
rect 10974 -35822 11068 -35788
rect 10924 -35838 11068 -35822
rect 11116 -35788 11260 -35705
rect 11332 -35747 11386 -35485
rect 11452 -35612 11482 -35462
rect 11452 -35642 11590 -35612
rect 11326 -35772 11386 -35747
rect 11500 -35772 11590 -35642
rect 12914 -35634 12980 -35618
rect 12914 -35668 12930 -35634
rect 12964 -35668 12980 -35634
rect 12914 -35685 12980 -35668
rect 13168 -35634 13426 -35618
rect 13168 -35668 13184 -35634
rect 13410 -35668 13426 -35634
rect 13168 -35684 13426 -35668
rect 12932 -35715 12962 -35685
rect 13186 -35715 13216 -35684
rect 13282 -35715 13312 -35684
rect 13378 -35715 13408 -35684
rect 11116 -35822 11132 -35788
rect 11166 -35822 11260 -35788
rect 11116 -35838 11260 -35822
rect 11308 -35788 11452 -35772
rect 11308 -35822 11324 -35788
rect 11358 -35822 11452 -35788
rect 11308 -35838 11452 -35822
rect 11500 -35788 11644 -35772
rect 11500 -35822 11516 -35788
rect 11550 -35822 11644 -35788
rect 11500 -35838 11644 -35822
rect 10942 -35869 10972 -35838
rect 11038 -35869 11068 -35838
rect 11134 -35869 11164 -35838
rect 11230 -35869 11260 -35838
rect 11326 -35869 11356 -35838
rect 11422 -35869 11452 -35838
rect 11518 -35869 11548 -35838
rect 11614 -35869 11644 -35838
rect 7200 -36217 7230 -36191
rect 7296 -36217 7326 -36191
rect 7392 -36217 7422 -36191
rect 7488 -36217 7518 -36191
rect 7584 -36217 7614 -36191
rect 7680 -36217 7710 -36191
rect 7776 -36217 7806 -36191
rect 7872 -36217 7902 -36191
rect 8148 -36217 8178 -36191
rect 8244 -36217 8274 -36191
rect 8340 -36217 8370 -36191
rect 8436 -36217 8466 -36191
rect 8532 -36217 8562 -36191
rect 8628 -36217 8658 -36191
rect 8724 -36217 8754 -36191
rect 8820 -36217 8850 -36191
rect 9084 -36217 9114 -36191
rect 9180 -36217 9210 -36191
rect 9276 -36217 9306 -36191
rect 9372 -36217 9402 -36191
rect 9468 -36217 9498 -36191
rect 9564 -36217 9594 -36191
rect 9660 -36217 9690 -36191
rect 9756 -36217 9786 -36191
rect 10015 -36216 10045 -36190
rect 10111 -36216 10141 -36190
rect 10207 -36216 10237 -36190
rect 10303 -36216 10333 -36190
rect 10399 -36216 10429 -36190
rect 10495 -36216 10525 -36190
rect 10591 -36216 10621 -36190
rect 10687 -36216 10717 -36190
rect 12932 -35941 12962 -35915
rect 13186 -35955 13216 -35929
rect 13282 -35955 13312 -35929
rect 13378 -35955 13408 -35929
rect 12914 -36013 12980 -35997
rect 12914 -36047 12930 -36013
rect 12964 -36047 12980 -36013
rect 12914 -36064 12980 -36047
rect 13168 -36013 13426 -35997
rect 13168 -36047 13184 -36013
rect 13410 -36047 13426 -36013
rect 13168 -36063 13426 -36047
rect 12932 -36094 12962 -36064
rect 13186 -36094 13216 -36063
rect 13282 -36094 13312 -36063
rect 13378 -36094 13408 -36063
rect 10942 -36217 10972 -36191
rect 11038 -36217 11068 -36191
rect 11134 -36217 11164 -36191
rect 11230 -36217 11260 -36191
rect 11326 -36217 11356 -36191
rect 11422 -36217 11452 -36191
rect 11518 -36217 11548 -36191
rect 11614 -36217 11644 -36191
rect 12932 -36320 12962 -36294
rect 13186 -36334 13216 -36308
rect 13282 -36334 13312 -36308
rect 13378 -36334 13408 -36308
<< polycont >>
rect 2175 5430 2305 5475
rect 2506 5425 2636 5470
rect 1573 5254 1662 5343
rect 1900 5109 2030 5154
rect 2183 5101 2313 5146
rect 3781 5430 3911 5475
rect 4112 5425 4242 5470
rect 2753 5291 2818 5346
rect 3187 5254 3276 5343
rect 3506 5109 3636 5154
rect 3789 5101 3919 5146
rect 5485 5428 5615 5473
rect 5816 5423 5946 5468
rect 4359 5291 4424 5346
rect 4871 5252 4960 5341
rect 5210 5107 5340 5152
rect 5493 5099 5623 5144
rect 6063 5289 6128 5344
rect 7017 5145 7051 5180
rect 7306 5145 7340 5180
rect 7728 5185 7762 5411
rect 7101 5021 7135 5056
rect 7101 4888 7135 4923
rect 7728 4931 7762 4965
rect -23673 3701 -23543 3746
rect -23342 3706 -23212 3751
rect -23855 3567 -23790 3622
rect -22680 3547 -22488 3767
rect -20382 3701 -20252 3746
rect -20051 3706 -19921 3751
rect -20564 3567 -20499 3622
rect -23350 3377 -23220 3422
rect -23067 3385 -22937 3430
rect -19389 3547 -19197 3767
rect -17091 3701 -16961 3746
rect -16760 3706 -16630 3751
rect -17273 3567 -17208 3622
rect -20059 3377 -19929 3422
rect -19776 3385 -19646 3430
rect -16098 3547 -15906 3767
rect -13800 3701 -13670 3746
rect -13469 3706 -13339 3751
rect -13982 3567 -13917 3622
rect -16768 3377 -16638 3422
rect -16485 3385 -16355 3430
rect -12807 3547 -12615 3767
rect -10509 3701 -10379 3746
rect -10178 3706 -10048 3751
rect -10691 3567 -10626 3622
rect -13477 3377 -13347 3422
rect -13194 3385 -13064 3430
rect -9516 3547 -9324 3767
rect -7219 3701 -7089 3746
rect -6888 3706 -6758 3751
rect -7401 3567 -7336 3622
rect -10186 3377 -10056 3422
rect -9903 3385 -9773 3430
rect -6226 3547 -6034 3767
rect -3928 3701 -3798 3746
rect -3597 3706 -3467 3751
rect -4110 3567 -4045 3622
rect -6896 3377 -6766 3422
rect -6613 3385 -6483 3430
rect -2935 3547 -2743 3767
rect -637 3701 -507 3746
rect -306 3706 -176 3751
rect -819 3567 -754 3622
rect -3605 3377 -3475 3422
rect -3322 3385 -3192 3430
rect 356 3547 548 3767
rect 5577 3637 5611 3863
rect 6017 3637 6051 3863
rect 6457 3637 6491 3863
rect -314 3377 -184 3422
rect -31 3385 99 3430
rect 5577 3383 5611 3417
rect 6017 3383 6051 3417
rect 6457 3383 6491 3417
rect 7198 2816 7232 2850
rect 7390 2816 7424 2850
rect 7582 2816 7616 2850
rect 7774 2816 7808 2850
rect 8146 2816 8180 2850
rect 8338 2816 8372 2850
rect 8530 2816 8564 2850
rect 8722 2816 8756 2850
rect 9082 2816 9116 2850
rect 9274 2816 9308 2850
rect 9466 2816 9500 2850
rect 9658 2816 9692 2850
rect 10013 2816 10047 2850
rect 10205 2816 10239 2850
rect 10397 2816 10431 2850
rect 10589 2816 10623 2850
rect 10940 2816 10974 2850
rect 11132 2816 11166 2850
rect 11324 2816 11358 2850
rect 11516 2816 11550 2850
rect -24921 1828 -24874 1938
rect -24336 1922 -24206 1967
rect -24005 1917 -23875 1962
rect -24611 1601 -24481 1646
rect -24328 1593 -24198 1638
rect -23758 1783 -23693 1838
rect -22777 1922 -22647 1967
rect -22446 1917 -22316 1962
rect -23364 1753 -23291 1893
rect -23052 1601 -22922 1646
rect -22769 1593 -22639 1638
rect -22199 1783 -22134 1838
rect -21630 1828 -21583 1938
rect -21045 1922 -20915 1967
rect -20714 1917 -20584 1962
rect -21320 1601 -21190 1646
rect -21037 1593 -20907 1638
rect -20467 1783 -20402 1838
rect -19486 1922 -19356 1967
rect -19155 1917 -19025 1962
rect -20073 1753 -20000 1893
rect -19761 1601 -19631 1646
rect -19478 1593 -19348 1638
rect -18908 1783 -18843 1838
rect -18339 1828 -18292 1938
rect -17754 1922 -17624 1967
rect -17423 1917 -17293 1962
rect -18029 1601 -17899 1646
rect -17746 1593 -17616 1638
rect -17176 1783 -17111 1838
rect -16195 1922 -16065 1967
rect -15864 1917 -15734 1962
rect -16782 1753 -16709 1893
rect -16470 1601 -16340 1646
rect -16187 1593 -16057 1638
rect -15617 1783 -15552 1838
rect -15048 1828 -15001 1938
rect -14463 1922 -14333 1967
rect -14132 1917 -14002 1962
rect -14738 1601 -14608 1646
rect -14455 1593 -14325 1638
rect -13885 1783 -13820 1838
rect -12904 1922 -12774 1967
rect -12573 1917 -12443 1962
rect -13491 1753 -13418 1893
rect -13179 1601 -13049 1646
rect -12896 1593 -12766 1638
rect -12326 1783 -12261 1838
rect -11757 1828 -11710 1938
rect -11172 1922 -11042 1967
rect -10841 1917 -10711 1962
rect -11447 1601 -11317 1646
rect -11164 1593 -11034 1638
rect -10594 1783 -10529 1838
rect -9613 1922 -9483 1967
rect -9282 1917 -9152 1962
rect -10200 1753 -10127 1893
rect -9888 1601 -9758 1646
rect -9605 1593 -9475 1638
rect -9035 1783 -8970 1838
rect -8467 1828 -8420 1938
rect -7882 1922 -7752 1967
rect -7551 1917 -7421 1962
rect -8157 1601 -8027 1646
rect -7874 1593 -7744 1638
rect -7304 1783 -7239 1838
rect -6323 1922 -6193 1967
rect -5992 1917 -5862 1962
rect -6910 1753 -6837 1893
rect -6598 1601 -6468 1646
rect -6315 1593 -6185 1638
rect -5745 1783 -5680 1838
rect -5176 1828 -5129 1938
rect -4591 1922 -4461 1967
rect -4260 1917 -4130 1962
rect -4866 1601 -4736 1646
rect -4583 1593 -4453 1638
rect -4013 1783 -3948 1838
rect -3032 1922 -2902 1967
rect -2701 1917 -2571 1962
rect -3619 1753 -3546 1893
rect -3307 1601 -3177 1646
rect -3024 1593 -2894 1638
rect -2454 1783 -2389 1838
rect -1885 1828 -1838 1938
rect -1300 1922 -1170 1967
rect -969 1917 -839 1962
rect -1575 1601 -1445 1646
rect -1292 1593 -1162 1638
rect -722 1783 -657 1838
rect 259 1922 389 1967
rect 590 1917 720 1962
rect -328 1753 -255 1893
rect -16 1601 114 1646
rect 267 1593 397 1638
rect 837 1783 902 1838
rect 12170 1669 12204 1703
rect -24519 579 -24485 614
rect -24230 579 -24196 614
rect -23410 579 -23376 614
rect -23121 579 -23087 614
rect -22528 579 -22494 614
rect -22239 579 -22205 614
rect -21228 579 -21194 614
rect -20939 579 -20905 614
rect -20119 579 -20085 614
rect -19830 579 -19796 614
rect -19237 579 -19203 614
rect -18948 579 -18914 614
rect -17937 579 -17903 614
rect -17648 579 -17614 614
rect -16828 579 -16794 614
rect -16539 579 -16505 614
rect -15946 579 -15912 614
rect -15657 579 -15623 614
rect -14646 579 -14612 614
rect -14357 579 -14323 614
rect -13537 579 -13503 614
rect -13248 579 -13214 614
rect -12655 579 -12621 614
rect -12366 579 -12332 614
rect -11355 579 -11321 614
rect -11066 579 -11032 614
rect -10246 579 -10212 614
rect -9957 579 -9923 614
rect -9364 579 -9330 614
rect -9075 579 -9041 614
rect -8065 579 -8031 614
rect -7776 579 -7742 614
rect -6956 579 -6922 614
rect -6667 579 -6633 614
rect -6074 579 -6040 614
rect -5785 579 -5751 614
rect -4774 579 -4740 614
rect -4485 579 -4451 614
rect -3665 579 -3631 614
rect -3376 579 -3342 614
rect -2783 579 -2749 614
rect -2494 579 -2460 614
rect -1483 579 -1449 614
rect -1194 579 -1160 614
rect -374 579 -340 614
rect -85 579 -51 614
rect 508 579 542 614
rect 797 579 831 614
rect -24435 455 -24401 490
rect -23326 455 -23292 490
rect -22444 455 -22410 490
rect -21144 455 -21110 490
rect -20035 455 -20001 490
rect -19153 455 -19119 490
rect -17853 455 -17819 490
rect -16744 455 -16710 490
rect -15862 455 -15828 490
rect -14562 455 -14528 490
rect -13453 455 -13419 490
rect -12571 455 -12537 490
rect -11271 455 -11237 490
rect -10162 455 -10128 490
rect -9280 455 -9246 490
rect -7981 455 -7947 490
rect -6872 455 -6838 490
rect -5990 455 -5956 490
rect -4690 455 -4656 490
rect -3581 455 -3547 490
rect -2699 455 -2665 490
rect -1399 455 -1365 490
rect -290 455 -256 490
rect 592 455 626 490
rect 7198 402 7232 436
rect 7390 402 7424 436
rect 7582 402 7616 436
rect 7774 402 7808 436
rect 8146 402 8180 436
rect 8338 402 8372 436
rect 8530 402 8564 436
rect 8722 402 8756 436
rect 9082 402 9116 436
rect 9274 402 9308 436
rect 9466 402 9500 436
rect 9658 402 9692 436
rect 10013 403 10047 437
rect 12842 1619 12876 1845
rect 12313 1564 12347 1598
rect 12842 1365 12876 1399
rect 10205 403 10239 437
rect 10397 403 10431 437
rect 10589 403 10623 437
rect -24435 322 -24401 357
rect -23326 322 -23292 357
rect -22444 322 -22410 357
rect -21144 322 -21110 357
rect -20035 322 -20001 357
rect -19153 322 -19119 357
rect -17853 322 -17819 357
rect -16744 322 -16710 357
rect -15862 322 -15828 357
rect -14562 322 -14528 357
rect -13453 322 -13419 357
rect -12571 322 -12537 357
rect -11271 322 -11237 357
rect -10162 322 -10128 357
rect -9280 322 -9246 357
rect -7981 322 -7947 357
rect -6872 322 -6838 357
rect -5990 322 -5956 357
rect -4690 322 -4656 357
rect -3581 322 -3547 357
rect -2699 322 -2665 357
rect -1399 322 -1365 357
rect -290 322 -256 357
rect 592 322 626 357
rect 10940 402 10974 436
rect 11132 402 11166 436
rect 11324 402 11358 436
rect 11516 402 11550 436
rect 5577 -891 5611 -665
rect 6017 -891 6051 -665
rect 6457 -891 6491 -665
rect 5577 -1145 5611 -1111
rect 6017 -1145 6051 -1111
rect 6457 -1145 6491 -1111
rect 7198 -1712 7232 -1678
rect 7390 -1712 7424 -1678
rect 7582 -1712 7616 -1678
rect 7774 -1712 7808 -1678
rect 8146 -1712 8180 -1678
rect 8338 -1712 8372 -1678
rect 8530 -1712 8564 -1678
rect 8722 -1712 8756 -1678
rect 9082 -1712 9116 -1678
rect 9274 -1712 9308 -1678
rect 9466 -1712 9500 -1678
rect 9658 -1712 9692 -1678
rect 10013 -1712 10047 -1678
rect 10205 -1712 10239 -1678
rect 10397 -1712 10431 -1678
rect 10589 -1712 10623 -1678
rect 10940 -1712 10974 -1678
rect 11132 -1712 11166 -1678
rect 11324 -1712 11358 -1678
rect 11516 -1712 11550 -1678
rect -23709 -2593 -23675 -2367
rect -24369 -2709 -24335 -2674
rect -21689 -2593 -21655 -2367
rect -24080 -2709 -24046 -2674
rect -22332 -2709 -22298 -2674
rect -19948 -2593 -19914 -2367
rect -22043 -2709 -22009 -2674
rect -20602 -2709 -20568 -2674
rect -18169 -2593 -18135 -2367
rect -20313 -2709 -20279 -2674
rect -18842 -2709 -18808 -2674
rect -18553 -2709 -18519 -2674
rect -24285 -2833 -24251 -2798
rect -23709 -2847 -23675 -2813
rect -22248 -2833 -22214 -2798
rect -21689 -2847 -21655 -2813
rect -20518 -2833 -20484 -2798
rect -19948 -2847 -19914 -2813
rect -18758 -2833 -18724 -2798
rect -18169 -2847 -18135 -2813
rect 12170 -2859 12204 -2825
rect -24285 -2966 -24251 -2931
rect -22248 -2966 -22214 -2931
rect -20518 -2966 -20484 -2931
rect -18758 -2966 -18724 -2931
rect -23665 -4405 -23631 -4179
rect -24318 -4521 -24284 -4486
rect -21927 -4405 -21893 -4179
rect -24029 -4521 -23995 -4486
rect -22582 -4521 -22548 -4486
rect -22293 -4521 -22259 -4486
rect -24234 -4645 -24200 -4610
rect -23665 -4659 -23631 -4625
rect 7198 -4126 7232 -4092
rect 7390 -4126 7424 -4092
rect 7582 -4126 7616 -4092
rect 7774 -4126 7808 -4092
rect 8146 -4126 8180 -4092
rect 8338 -4126 8372 -4092
rect 8530 -4126 8564 -4092
rect 8722 -4126 8756 -4092
rect 9082 -4126 9116 -4092
rect 9274 -4126 9308 -4092
rect 9466 -4126 9500 -4092
rect 9658 -4126 9692 -4092
rect 10013 -4125 10047 -4091
rect 12842 -2909 12876 -2683
rect 12313 -2964 12347 -2930
rect 12842 -3163 12876 -3129
rect 10205 -4125 10239 -4091
rect 10397 -4125 10431 -4091
rect 10589 -4125 10623 -4091
rect 10940 -4126 10974 -4092
rect 11132 -4126 11166 -4092
rect 11324 -4126 11358 -4092
rect 11516 -4126 11550 -4092
rect -22498 -4645 -22464 -4610
rect -21927 -4659 -21893 -4625
rect -24234 -4778 -24200 -4743
rect -22498 -4778 -22464 -4743
rect -20854 -4732 -20807 -4622
rect -20269 -4638 -20139 -4593
rect -19938 -4643 -19808 -4598
rect -20544 -4959 -20414 -4914
rect -20261 -4967 -20131 -4922
rect -19691 -4777 -19626 -4722
rect -18710 -4638 -18580 -4593
rect -18379 -4643 -18249 -4598
rect -19297 -4807 -19224 -4667
rect -18985 -4959 -18855 -4914
rect -18702 -4967 -18572 -4922
rect -18132 -4777 -18067 -4722
rect -17563 -4732 -17516 -4622
rect -16978 -4638 -16848 -4593
rect -16647 -4643 -16517 -4598
rect -17253 -4959 -17123 -4914
rect -16970 -4967 -16840 -4922
rect -16400 -4777 -16335 -4722
rect -15419 -4638 -15289 -4593
rect -15088 -4643 -14958 -4598
rect -16006 -4807 -15933 -4667
rect -15694 -4959 -15564 -4914
rect -15411 -4967 -15281 -4922
rect -14841 -4777 -14776 -4722
rect -14272 -4732 -14225 -4622
rect -13687 -4638 -13557 -4593
rect -13356 -4643 -13226 -4598
rect -13962 -4959 -13832 -4914
rect -13679 -4967 -13549 -4922
rect -13109 -4777 -13044 -4722
rect -12128 -4638 -11998 -4593
rect -11797 -4643 -11667 -4598
rect -12715 -4807 -12642 -4667
rect -12403 -4959 -12273 -4914
rect -12120 -4967 -11990 -4922
rect -11550 -4777 -11485 -4722
rect -10981 -4732 -10934 -4622
rect -10396 -4638 -10266 -4593
rect -10065 -4643 -9935 -4598
rect -10671 -4959 -10541 -4914
rect -10388 -4967 -10258 -4922
rect -9818 -4777 -9753 -4722
rect -8837 -4638 -8707 -4593
rect -8506 -4643 -8376 -4598
rect -9424 -4807 -9351 -4667
rect -9112 -4959 -8982 -4914
rect -8829 -4967 -8699 -4922
rect -8259 -4777 -8194 -4722
rect 5577 -5319 5611 -5093
rect 6017 -5319 6051 -5093
rect 6457 -5319 6491 -5093
rect -23667 -5697 -23633 -5471
rect -24318 -5813 -24284 -5778
rect -21933 -5697 -21899 -5471
rect 5577 -5573 5611 -5539
rect 6017 -5573 6051 -5539
rect 6457 -5573 6491 -5539
rect -24029 -5813 -23995 -5778
rect -22582 -5813 -22548 -5778
rect -22293 -5813 -22259 -5778
rect -24234 -5937 -24200 -5902
rect -23667 -5951 -23633 -5917
rect -22498 -5937 -22464 -5902
rect -21933 -5951 -21899 -5917
rect -20452 -5981 -20418 -5946
rect -20163 -5981 -20129 -5946
rect -19343 -5981 -19309 -5946
rect -19054 -5981 -19020 -5946
rect -18461 -5981 -18427 -5946
rect -18172 -5981 -18138 -5946
rect -17161 -5981 -17127 -5946
rect -16872 -5981 -16838 -5946
rect -16052 -5981 -16018 -5946
rect -15763 -5981 -15729 -5946
rect -15170 -5981 -15136 -5946
rect -14881 -5981 -14847 -5946
rect -13870 -5981 -13836 -5946
rect -13581 -5981 -13547 -5946
rect -12761 -5981 -12727 -5946
rect -12472 -5981 -12438 -5946
rect -11879 -5981 -11845 -5946
rect -11590 -5981 -11556 -5946
rect -10579 -5981 -10545 -5946
rect -10290 -5981 -10256 -5946
rect -9470 -5981 -9436 -5946
rect -9181 -5981 -9147 -5946
rect -8588 -5981 -8554 -5946
rect -8299 -5981 -8265 -5946
rect -24234 -6070 -24200 -6035
rect -22498 -6070 -22464 -6035
rect -20368 -6105 -20334 -6070
rect -19259 -6105 -19225 -6070
rect -18377 -6105 -18343 -6070
rect -17077 -6105 -17043 -6070
rect -15968 -6105 -15934 -6070
rect -15086 -6105 -15052 -6070
rect -13786 -6105 -13752 -6070
rect -12677 -6105 -12643 -6070
rect -11795 -6105 -11761 -6070
rect -10495 -6105 -10461 -6070
rect -9386 -6105 -9352 -6070
rect -8504 -6105 -8470 -6070
rect 7198 -6140 7232 -6106
rect 7390 -6140 7424 -6106
rect -20368 -6238 -20334 -6203
rect -19259 -6238 -19225 -6203
rect -18377 -6238 -18343 -6203
rect -17077 -6238 -17043 -6203
rect -15968 -6238 -15934 -6203
rect -15086 -6238 -15052 -6203
rect -13786 -6238 -13752 -6203
rect -12677 -6238 -12643 -6203
rect -11795 -6238 -11761 -6203
rect -10495 -6238 -10461 -6203
rect -9386 -6238 -9352 -6203
rect -8504 -6238 -8470 -6203
rect 7582 -6140 7616 -6106
rect 7774 -6140 7808 -6106
rect 8146 -6140 8180 -6106
rect 8338 -6140 8372 -6106
rect 8530 -6140 8564 -6106
rect 8722 -6140 8756 -6106
rect 9082 -6140 9116 -6106
rect 9274 -6140 9308 -6106
rect 9466 -6140 9500 -6106
rect 9658 -6140 9692 -6106
rect 10013 -6140 10047 -6106
rect 10205 -6140 10239 -6106
rect 10397 -6140 10431 -6106
rect 10589 -6140 10623 -6106
rect 10940 -6140 10974 -6106
rect 11132 -6140 11166 -6106
rect 11324 -6140 11358 -6106
rect 11516 -6140 11550 -6106
rect -23665 -7670 -23631 -7444
rect -24318 -7786 -24284 -7751
rect -21931 -7670 -21897 -7444
rect -24029 -7786 -23995 -7751
rect -22581 -7786 -22547 -7751
rect -22292 -7786 -22258 -7751
rect -24234 -7910 -24200 -7875
rect -23665 -7924 -23631 -7890
rect 12170 -7287 12204 -7253
rect -22497 -7910 -22463 -7875
rect -21931 -7924 -21897 -7890
rect -24234 -8043 -24200 -8008
rect -22497 -8043 -22463 -8008
rect -20854 -7997 -20807 -7887
rect -20269 -7903 -20139 -7858
rect -19938 -7908 -19808 -7863
rect -20544 -8224 -20414 -8179
rect -20261 -8232 -20131 -8187
rect -19691 -8042 -19626 -7987
rect -18710 -7903 -18580 -7858
rect -18379 -7908 -18249 -7863
rect -19297 -8072 -19224 -7932
rect -18985 -8224 -18855 -8179
rect -18702 -8232 -18572 -8187
rect -18132 -8042 -18067 -7987
rect -17563 -7997 -17516 -7887
rect -16978 -7903 -16848 -7858
rect -16647 -7908 -16517 -7863
rect -17253 -8224 -17123 -8179
rect -16970 -8232 -16840 -8187
rect -16400 -8042 -16335 -7987
rect -15419 -7903 -15289 -7858
rect -15088 -7908 -14958 -7863
rect -16006 -8072 -15933 -7932
rect -15694 -8224 -15564 -8179
rect -15411 -8232 -15281 -8187
rect -14841 -8042 -14776 -7987
rect -14272 -7997 -14225 -7887
rect -13687 -7903 -13557 -7858
rect -13356 -7908 -13226 -7863
rect -13962 -8224 -13832 -8179
rect -13679 -8232 -13549 -8187
rect -13109 -8042 -13044 -7987
rect -12128 -7903 -11998 -7858
rect -11797 -7908 -11667 -7863
rect -12715 -8072 -12642 -7932
rect -12403 -8224 -12273 -8179
rect -12120 -8232 -11990 -8187
rect -11550 -8042 -11485 -7987
rect -10981 -7997 -10934 -7887
rect -10396 -7903 -10266 -7858
rect -10065 -7908 -9935 -7863
rect -10671 -8224 -10541 -8179
rect -10388 -8232 -10258 -8187
rect -9818 -8042 -9753 -7987
rect -8837 -7903 -8707 -7858
rect -8506 -7908 -8376 -7863
rect -9424 -8072 -9351 -7932
rect -9112 -8224 -8982 -8179
rect -8829 -8232 -8699 -8187
rect -8259 -8042 -8194 -7987
rect 7198 -8554 7232 -8520
rect 7390 -8554 7424 -8520
rect 7582 -8554 7616 -8520
rect 7774 -8554 7808 -8520
rect 8146 -8554 8180 -8520
rect 8338 -8554 8372 -8520
rect 8530 -8554 8564 -8520
rect 8722 -8554 8756 -8520
rect 9082 -8554 9116 -8520
rect 9274 -8554 9308 -8520
rect 9466 -8554 9500 -8520
rect 9658 -8554 9692 -8520
rect 10013 -8553 10047 -8519
rect 12842 -7337 12876 -7111
rect 12313 -7392 12347 -7358
rect 12842 -7591 12876 -7557
rect 10205 -8553 10239 -8519
rect 10397 -8553 10431 -8519
rect 10589 -8553 10623 -8519
rect 10940 -8554 10974 -8520
rect 11132 -8554 11166 -8520
rect 11324 -8554 11358 -8520
rect 11516 -8554 11550 -8520
rect -23664 -8962 -23630 -8736
rect -24318 -9078 -24284 -9043
rect -21927 -8962 -21893 -8736
rect -24029 -9078 -23995 -9043
rect -22582 -9078 -22548 -9043
rect -22293 -9078 -22259 -9043
rect -24234 -9202 -24200 -9167
rect -23664 -9216 -23630 -9182
rect -22498 -9202 -22464 -9167
rect -21927 -9216 -21893 -9182
rect -20452 -9246 -20418 -9211
rect -20163 -9246 -20129 -9211
rect -19343 -9246 -19309 -9211
rect -19054 -9246 -19020 -9211
rect -18461 -9246 -18427 -9211
rect -18172 -9246 -18138 -9211
rect -17161 -9246 -17127 -9211
rect -16872 -9246 -16838 -9211
rect -16052 -9246 -16018 -9211
rect -15763 -9246 -15729 -9211
rect -15170 -9246 -15136 -9211
rect -14881 -9246 -14847 -9211
rect -13870 -9246 -13836 -9211
rect -13581 -9246 -13547 -9211
rect -12761 -9246 -12727 -9211
rect -12472 -9246 -12438 -9211
rect -11879 -9246 -11845 -9211
rect -11590 -9246 -11556 -9211
rect -10579 -9246 -10545 -9211
rect -10290 -9246 -10256 -9211
rect -9470 -9246 -9436 -9211
rect -9181 -9246 -9147 -9211
rect -8588 -9246 -8554 -9211
rect -8299 -9246 -8265 -9211
rect -24234 -9335 -24200 -9300
rect -22498 -9335 -22464 -9300
rect -20368 -9370 -20334 -9335
rect -19259 -9370 -19225 -9335
rect -18377 -9370 -18343 -9335
rect -17077 -9370 -17043 -9335
rect -15968 -9370 -15934 -9335
rect -15086 -9370 -15052 -9335
rect -13786 -9370 -13752 -9335
rect -12677 -9370 -12643 -9335
rect -11795 -9370 -11761 -9335
rect -10495 -9370 -10461 -9335
rect -9386 -9370 -9352 -9335
rect -8504 -9370 -8470 -9335
rect -20368 -9503 -20334 -9468
rect -19259 -9503 -19225 -9468
rect -18377 -9503 -18343 -9468
rect -17077 -9503 -17043 -9468
rect -15968 -9503 -15934 -9468
rect -15086 -9503 -15052 -9468
rect -13786 -9503 -13752 -9468
rect -12677 -9503 -12643 -9468
rect -11795 -9503 -11761 -9468
rect -10495 -9503 -10461 -9468
rect -9386 -9503 -9352 -9468
rect -8504 -9503 -8470 -9468
rect 5577 -9947 5611 -9721
rect 6017 -9947 6051 -9721
rect 6457 -9947 6491 -9721
rect 5577 -10201 5611 -10167
rect 6017 -10201 6051 -10167
rect 6457 -10201 6491 -10167
rect -23664 -10934 -23630 -10708
rect -24318 -11050 -24284 -11015
rect -21931 -10934 -21897 -10708
rect -24029 -11050 -23995 -11015
rect -22581 -11050 -22547 -11015
rect -22292 -11050 -22258 -11015
rect -24234 -11174 -24200 -11139
rect -23664 -11188 -23630 -11154
rect 7198 -10768 7232 -10734
rect 7390 -10768 7424 -10734
rect 7582 -10768 7616 -10734
rect 7774 -10768 7808 -10734
rect 8146 -10768 8180 -10734
rect 8338 -10768 8372 -10734
rect -22497 -11174 -22463 -11139
rect -21931 -11188 -21897 -11154
rect -24234 -11307 -24200 -11272
rect -22497 -11307 -22463 -11272
rect -20854 -11261 -20807 -11151
rect -20269 -11167 -20139 -11122
rect -19938 -11172 -19808 -11127
rect -20544 -11488 -20414 -11443
rect -20261 -11496 -20131 -11451
rect -19691 -11306 -19626 -11251
rect -18710 -11167 -18580 -11122
rect -18379 -11172 -18249 -11127
rect -19297 -11336 -19224 -11196
rect -18985 -11488 -18855 -11443
rect -18702 -11496 -18572 -11451
rect -18132 -11306 -18067 -11251
rect -17563 -11261 -17516 -11151
rect -16978 -11167 -16848 -11122
rect -16647 -11172 -16517 -11127
rect -17253 -11488 -17123 -11443
rect -16970 -11496 -16840 -11451
rect -16400 -11306 -16335 -11251
rect -15419 -11167 -15289 -11122
rect -15088 -11172 -14958 -11127
rect -16006 -11336 -15933 -11196
rect -15694 -11488 -15564 -11443
rect -15411 -11496 -15281 -11451
rect -14841 -11306 -14776 -11251
rect -14272 -11261 -14225 -11151
rect -13687 -11167 -13557 -11122
rect -13356 -11172 -13226 -11127
rect -13962 -11488 -13832 -11443
rect -13679 -11496 -13549 -11451
rect -13109 -11306 -13044 -11251
rect -12128 -11167 -11998 -11122
rect -11797 -11172 -11667 -11127
rect -12715 -11336 -12642 -11196
rect -12403 -11488 -12273 -11443
rect -12120 -11496 -11990 -11451
rect -11550 -11306 -11485 -11251
rect -10981 -11261 -10934 -11151
rect -10396 -11167 -10266 -11122
rect -10065 -11172 -9935 -11127
rect -10671 -11488 -10541 -11443
rect -10388 -11496 -10258 -11451
rect -9818 -11306 -9753 -11251
rect -8837 -11167 -8707 -11122
rect -8506 -11172 -8376 -11127
rect 8530 -10768 8564 -10734
rect 8722 -10768 8756 -10734
rect 9082 -10768 9116 -10734
rect 9274 -10768 9308 -10734
rect 9466 -10768 9500 -10734
rect 9658 -10768 9692 -10734
rect 10013 -10768 10047 -10734
rect 10205 -10768 10239 -10734
rect 10397 -10768 10431 -10734
rect 10589 -10768 10623 -10734
rect 10940 -10768 10974 -10734
rect 11132 -10768 11166 -10734
rect 11324 -10768 11358 -10734
rect 11516 -10768 11550 -10734
rect -9424 -11336 -9351 -11196
rect -9112 -11488 -8982 -11443
rect -8829 -11496 -8699 -11451
rect -8259 -11306 -8194 -11251
rect -23664 -12226 -23630 -12000
rect 12170 -11915 12204 -11881
rect -24318 -12342 -24284 -12307
rect -21935 -12226 -21901 -12000
rect -24029 -12342 -23995 -12307
rect -22581 -12342 -22547 -12307
rect -22292 -12342 -22258 -12307
rect -24234 -12466 -24200 -12431
rect -23664 -12480 -23630 -12446
rect -22497 -12466 -22463 -12431
rect -21935 -12480 -21901 -12446
rect -20452 -12510 -20418 -12475
rect -20163 -12510 -20129 -12475
rect -19343 -12510 -19309 -12475
rect -19054 -12510 -19020 -12475
rect -18461 -12510 -18427 -12475
rect -18172 -12510 -18138 -12475
rect -17161 -12510 -17127 -12475
rect -16872 -12510 -16838 -12475
rect -16052 -12510 -16018 -12475
rect -15763 -12510 -15729 -12475
rect -15170 -12510 -15136 -12475
rect -14881 -12510 -14847 -12475
rect -13870 -12510 -13836 -12475
rect -13581 -12510 -13547 -12475
rect -12761 -12510 -12727 -12475
rect -12472 -12510 -12438 -12475
rect -11879 -12510 -11845 -12475
rect -11590 -12510 -11556 -12475
rect -10579 -12510 -10545 -12475
rect -10290 -12510 -10256 -12475
rect -9470 -12510 -9436 -12475
rect -9181 -12510 -9147 -12475
rect -8588 -12510 -8554 -12475
rect -8299 -12510 -8265 -12475
rect -24234 -12599 -24200 -12564
rect -22497 -12599 -22463 -12564
rect -20368 -12634 -20334 -12599
rect -19259 -12634 -19225 -12599
rect -18377 -12634 -18343 -12599
rect -17077 -12634 -17043 -12599
rect -15968 -12634 -15934 -12599
rect -15086 -12634 -15052 -12599
rect -13786 -12634 -13752 -12599
rect -12677 -12634 -12643 -12599
rect -11795 -12634 -11761 -12599
rect -10495 -12634 -10461 -12599
rect -9386 -12634 -9352 -12599
rect -8504 -12634 -8470 -12599
rect -20368 -12767 -20334 -12732
rect -19259 -12767 -19225 -12732
rect -18377 -12767 -18343 -12732
rect -17077 -12767 -17043 -12732
rect -15968 -12767 -15934 -12732
rect -15086 -12767 -15052 -12732
rect -13786 -12767 -13752 -12732
rect -12677 -12767 -12643 -12732
rect -11795 -12767 -11761 -12732
rect -10495 -12767 -10461 -12732
rect -9386 -12767 -9352 -12732
rect -8504 -12767 -8470 -12732
rect 7198 -13182 7232 -13148
rect 7390 -13182 7424 -13148
rect 7582 -13182 7616 -13148
rect 7774 -13182 7808 -13148
rect 8146 -13182 8180 -13148
rect 8338 -13182 8372 -13148
rect 8530 -13182 8564 -13148
rect 8722 -13182 8756 -13148
rect 9082 -13182 9116 -13148
rect 9274 -13182 9308 -13148
rect 9466 -13182 9500 -13148
rect 9658 -13182 9692 -13148
rect 10013 -13181 10047 -13147
rect 12842 -11965 12876 -11739
rect 12313 -12020 12347 -11986
rect 12842 -12219 12876 -12185
rect 10205 -13181 10239 -13147
rect 10397 -13181 10431 -13147
rect 10589 -13181 10623 -13147
rect 10940 -13182 10974 -13148
rect 11132 -13182 11166 -13148
rect 11324 -13182 11358 -13148
rect 11516 -13182 11550 -13148
rect -4768 -14156 -4542 -14122
rect -4322 -14156 -4288 -14122
rect -2052 -14113 -1826 -14079
rect -1606 -14113 -1572 -14079
rect -24188 -15183 -24153 -15149
rect -17266 -14977 -17232 -14943
rect -24064 -15388 -24029 -15354
rect -23931 -15388 -23896 -15354
rect -24188 -15472 -24153 -15438
rect -17371 -15120 -17337 -15086
rect -11578 -14433 -11523 -14368
rect -11702 -14680 -11657 -14550
rect -11707 -15011 -11662 -14881
rect -11378 -15003 -11333 -14873
rect -11386 -15286 -11341 -15156
rect -2052 -14492 -1826 -14458
rect -1606 -14492 -1572 -14458
rect 5577 -14475 5611 -14249
rect 6017 -14475 6051 -14249
rect 6457 -14475 6491 -14249
rect -4768 -14596 -4542 -14562
rect -4322 -14596 -4288 -14562
rect 5577 -14729 5611 -14695
rect 6017 -14729 6051 -14695
rect 6457 -14729 6491 -14695
rect -4768 -14975 -4542 -14941
rect -4322 -14975 -4288 -14941
rect -2052 -14932 -1826 -14898
rect -1606 -14932 -1572 -14898
rect -2052 -15311 -1826 -15277
rect -1606 -15311 -1572 -15277
rect 7198 -15296 7232 -15262
rect 7390 -15296 7424 -15262
rect -4768 -15415 -4542 -15381
rect -4322 -15415 -4288 -15381
rect -11557 -15658 -11503 -15604
rect -8119 -15641 -7893 -15607
rect -7673 -15641 -7639 -15607
rect 7582 -15296 7616 -15262
rect 7774 -15296 7808 -15262
rect 8146 -15296 8180 -15262
rect 8338 -15296 8372 -15262
rect 8530 -15296 8564 -15262
rect 8722 -15296 8756 -15262
rect 9082 -15296 9116 -15262
rect 9274 -15296 9308 -15262
rect 9466 -15296 9500 -15262
rect 9658 -15296 9692 -15262
rect 10013 -15296 10047 -15262
rect 10205 -15296 10239 -15262
rect 10397 -15296 10431 -15262
rect 10589 -15296 10623 -15262
rect 10940 -15296 10974 -15262
rect 11132 -15296 11166 -15262
rect 11324 -15296 11358 -15262
rect 11516 -15296 11550 -15262
rect -4768 -15794 -4542 -15760
rect -4322 -15794 -4288 -15760
rect -2052 -15751 -1826 -15717
rect -1606 -15751 -1572 -15717
rect -24187 -16368 -24152 -16334
rect -8118 -16141 -7892 -16107
rect -7672 -16141 -7638 -16107
rect -2052 -16130 -1826 -16096
rect -1606 -16130 -1572 -16096
rect -4768 -16234 -4542 -16200
rect -4322 -16234 -4288 -16200
rect -17266 -16377 -17232 -16343
rect -24063 -16573 -24028 -16539
rect -23930 -16573 -23895 -16539
rect -24187 -16657 -24152 -16623
rect -17371 -16520 -17337 -16486
rect 12170 -16443 12204 -16409
rect -8119 -16621 -7893 -16587
rect -7673 -16621 -7639 -16587
rect -4768 -16613 -4542 -16579
rect -4322 -16613 -4288 -16579
rect -2052 -16570 -1826 -16536
rect -1606 -16570 -1572 -16536
rect -24182 -17581 -24147 -17547
rect -24058 -17786 -24023 -17752
rect -23925 -17786 -23890 -17752
rect -24182 -17870 -24147 -17836
rect -17266 -17777 -17232 -17743
rect -21558 -18329 -21332 -18295
rect -21112 -18329 -21078 -18295
rect -17371 -17920 -17337 -17886
rect -15967 -18200 -15741 -18166
rect -15521 -18200 -15487 -18166
rect -11576 -17249 -11521 -17184
rect -11700 -17496 -11655 -17366
rect -11705 -17827 -11660 -17697
rect -11376 -17819 -11331 -17689
rect -11384 -18102 -11339 -17972
rect -2052 -16949 -1826 -16915
rect -1606 -16949 -1572 -16915
rect -4768 -17053 -4542 -17019
rect -4322 -17053 -4288 -17019
rect -8119 -17121 -7893 -17087
rect -7673 -17121 -7639 -17087
rect -4768 -17432 -4542 -17398
rect -4322 -17432 -4288 -17398
rect -2052 -17389 -1826 -17355
rect -1606 -17389 -1572 -17355
rect -8119 -17601 -7893 -17567
rect -7673 -17601 -7639 -17567
rect 7198 -17710 7232 -17676
rect -2052 -17768 -1826 -17734
rect 7390 -17710 7424 -17676
rect 7582 -17710 7616 -17676
rect 7774 -17710 7808 -17676
rect 8146 -17710 8180 -17676
rect 8338 -17710 8372 -17676
rect 8530 -17710 8564 -17676
rect 8722 -17710 8756 -17676
rect 9082 -17710 9116 -17676
rect 9274 -17710 9308 -17676
rect 9466 -17710 9500 -17676
rect 9658 -17710 9692 -17676
rect 10013 -17709 10047 -17675
rect 12842 -16493 12876 -16267
rect 12313 -16548 12347 -16514
rect 12842 -16747 12876 -16713
rect 10205 -17709 10239 -17675
rect 10397 -17709 10431 -17675
rect 10589 -17709 10623 -17675
rect -1606 -17768 -1572 -17734
rect 10940 -17710 10974 -17676
rect 15997 -17620 16031 -17586
rect 11132 -17710 11166 -17676
rect 11324 -17710 11358 -17676
rect 16285 -17620 16319 -17586
rect 16669 -17338 16703 -17304
rect 16417 -17620 16451 -17586
rect 11516 -17710 11550 -17676
rect -4768 -17872 -4542 -17838
rect -4322 -17872 -4288 -17838
rect -8119 -18061 -7893 -18027
rect -7673 -18061 -7639 -18027
rect -24167 -18700 -24132 -18666
rect -11555 -18467 -11501 -18413
rect -4768 -18251 -4542 -18217
rect -4322 -18251 -4288 -18217
rect -2052 -18208 -1826 -18174
rect -1606 -18208 -1572 -18174
rect -8133 -18521 -7907 -18487
rect -7687 -18521 -7653 -18487
rect -2052 -18587 -1826 -18553
rect -1606 -18587 -1572 -18553
rect -15966 -18700 -15740 -18666
rect -15520 -18700 -15486 -18666
rect -4768 -18691 -4542 -18657
rect -21557 -18829 -21331 -18795
rect -24043 -18905 -24008 -18871
rect -21111 -18829 -21077 -18795
rect -23910 -18905 -23875 -18871
rect -24167 -18989 -24132 -18955
rect -17266 -19177 -17232 -19143
rect 17372 -18571 17406 -18536
rect 17661 -18571 17695 -18536
rect 18015 -18533 18049 -18307
rect -4322 -18691 -4288 -18657
rect -8131 -19001 -7905 -18967
rect -7685 -19001 -7651 -18967
rect -4768 -19070 -4542 -19036
rect -4322 -19070 -4288 -19036
rect -2052 -19027 -1826 -18993
rect -1606 -19027 -1572 -18993
rect 5577 -19003 5611 -18777
rect 6017 -19003 6051 -18777
rect 6457 -19003 6491 -18777
rect -21558 -19309 -21332 -19275
rect -21112 -19309 -21078 -19275
rect -24165 -19894 -24130 -19860
rect -17371 -19320 -17337 -19286
rect -15967 -19180 -15741 -19146
rect -15521 -19180 -15487 -19146
rect 5577 -19257 5611 -19223
rect 6017 -19257 6051 -19223
rect 6457 -19257 6491 -19223
rect -2052 -19406 -1826 -19372
rect -1606 -19406 -1572 -19372
rect -4768 -19510 -4542 -19476
rect -4322 -19510 -4288 -19476
rect -15967 -19680 -15741 -19646
rect -15521 -19680 -15487 -19646
rect -21558 -19809 -21332 -19775
rect -21112 -19809 -21078 -19775
rect 17456 -18695 17490 -18660
rect 17456 -18828 17490 -18793
rect 18015 -18787 18049 -18753
rect 15997 -19586 16031 -19552
rect 16285 -19586 16319 -19552
rect -24041 -20099 -24006 -20065
rect -23908 -20099 -23873 -20065
rect -24165 -20183 -24130 -20149
rect -4768 -19889 -4542 -19855
rect -4322 -19889 -4288 -19855
rect -2052 -19846 -1826 -19812
rect -1606 -19846 -1572 -19812
rect 7198 -19824 7232 -19790
rect 7390 -19824 7424 -19790
rect -15967 -20160 -15741 -20126
rect -15521 -20160 -15487 -20126
rect -21558 -20289 -21332 -20255
rect -21112 -20289 -21078 -20255
rect -17266 -20577 -17232 -20543
rect -21558 -20749 -21332 -20715
rect -21112 -20749 -21078 -20715
rect -24134 -21094 -24099 -21060
rect -17371 -20720 -17337 -20686
rect -15967 -20620 -15741 -20586
rect -15521 -20620 -15487 -20586
rect -15981 -21080 -15755 -21046
rect -15535 -21080 -15501 -21046
rect -11576 -20206 -11521 -20141
rect -11700 -20453 -11655 -20323
rect -11705 -20784 -11660 -20654
rect -11376 -20776 -11331 -20646
rect -11384 -21059 -11339 -20929
rect -21572 -21209 -21346 -21175
rect 7582 -19824 7616 -19790
rect 7774 -19824 7808 -19790
rect 8146 -19824 8180 -19790
rect 8338 -19824 8372 -19790
rect 8530 -19824 8564 -19790
rect 8722 -19824 8756 -19790
rect 9082 -19824 9116 -19790
rect 9274 -19824 9308 -19790
rect 9466 -19824 9500 -19790
rect 9658 -19824 9692 -19790
rect 10013 -19824 10047 -19790
rect 10205 -19824 10239 -19790
rect 10397 -19824 10431 -19790
rect 10589 -19824 10623 -19790
rect 10940 -19824 10974 -19790
rect 11132 -19824 11166 -19790
rect 11324 -19824 11358 -19790
rect 11516 -19824 11550 -19790
rect 16417 -19586 16451 -19552
rect 16669 -19868 16703 -19834
rect -2052 -20225 -1826 -20191
rect -1606 -20225 -1572 -20191
rect -4768 -20329 -4542 -20295
rect -4322 -20329 -4288 -20295
rect -4768 -20708 -4542 -20674
rect -4322 -20708 -4288 -20674
rect -2052 -20665 -1826 -20631
rect -1606 -20665 -1572 -20631
rect 12170 -20971 12204 -20937
rect -21126 -21209 -21092 -21175
rect -24010 -21299 -23975 -21265
rect -23877 -21299 -23842 -21265
rect -24134 -21383 -24099 -21349
rect -11549 -21431 -11507 -21389
rect -15979 -21560 -15753 -21526
rect -15533 -21560 -15499 -21526
rect -21570 -21689 -21344 -21655
rect -21124 -21689 -21090 -21655
rect -17266 -21977 -17232 -21943
rect -24135 -22397 -24100 -22363
rect -17371 -22120 -17337 -22086
rect 7198 -22238 7232 -22204
rect 7390 -22238 7424 -22204
rect 7582 -22238 7616 -22204
rect 7774 -22238 7808 -22204
rect 8146 -22238 8180 -22204
rect 8338 -22238 8372 -22204
rect 8530 -22238 8564 -22204
rect 8722 -22238 8756 -22204
rect 9082 -22238 9116 -22204
rect 9274 -22238 9308 -22204
rect 9466 -22238 9500 -22204
rect 9658 -22238 9692 -22204
rect 10013 -22237 10047 -22203
rect 12842 -21021 12876 -20795
rect 12313 -21076 12347 -21042
rect 12842 -21275 12876 -21241
rect 10205 -22237 10239 -22203
rect 10397 -22237 10431 -22203
rect 10589 -22237 10623 -22203
rect 10940 -22238 10974 -22204
rect 11132 -22238 11166 -22204
rect 11324 -22238 11358 -22204
rect 11516 -22238 11550 -22204
rect -24011 -22602 -23976 -22568
rect -23878 -22602 -23843 -22568
rect -24135 -22686 -24100 -22652
rect -17266 -23377 -17232 -23343
rect -24135 -23706 -24100 -23672
rect -24011 -23911 -23976 -23877
rect -23878 -23911 -23843 -23877
rect -17371 -23520 -17337 -23486
rect -11576 -22785 -11521 -22720
rect -11700 -23032 -11655 -22902
rect -11705 -23363 -11660 -23233
rect -11376 -23355 -11331 -23225
rect -11384 -23638 -11339 -23508
rect 5577 -23531 5611 -23305
rect 6017 -23531 6051 -23305
rect 6457 -23531 6491 -23305
rect 5577 -23785 5611 -23751
rect 6017 -23785 6051 -23751
rect 6457 -23785 6491 -23751
rect -24135 -23995 -24100 -23961
rect -11553 -24019 -11504 -23970
rect 7198 -24352 7232 -24318
rect 7390 -24352 7424 -24318
rect 7582 -24352 7616 -24318
rect 7774 -24352 7808 -24318
rect 8146 -24352 8180 -24318
rect 8338 -24352 8372 -24318
rect 8530 -24352 8564 -24318
rect 8722 -24352 8756 -24318
rect 9082 -24352 9116 -24318
rect 9274 -24352 9308 -24318
rect 9466 -24352 9500 -24318
rect 9658 -24352 9692 -24318
rect 10013 -24352 10047 -24318
rect 10205 -24352 10239 -24318
rect 10397 -24352 10431 -24318
rect 10589 -24352 10623 -24318
rect 10940 -24352 10974 -24318
rect 11132 -24352 11166 -24318
rect 11324 -24352 11358 -24318
rect 11516 -24352 11550 -24318
rect -17266 -24777 -17232 -24743
rect -17371 -24920 -17337 -24886
rect -11576 -25553 -11521 -25488
rect -11700 -25800 -11655 -25670
rect -11705 -26131 -11660 -26001
rect -11376 -26123 -11331 -25993
rect -11384 -26406 -11339 -26276
rect 12170 -25499 12204 -25465
rect -11554 -26810 -11502 -26758
rect 7198 -26766 7232 -26732
rect 7390 -26766 7424 -26732
rect 7582 -26766 7616 -26732
rect 7774 -26766 7808 -26732
rect 8146 -26766 8180 -26732
rect 8338 -26766 8372 -26732
rect 8530 -26766 8564 -26732
rect 8722 -26766 8756 -26732
rect 9082 -26766 9116 -26732
rect 9274 -26766 9308 -26732
rect 9466 -26766 9500 -26732
rect 9658 -26766 9692 -26732
rect 10013 -26765 10047 -26731
rect 12842 -25549 12876 -25323
rect 12313 -25604 12347 -25570
rect 12842 -25803 12876 -25769
rect 10205 -26765 10239 -26731
rect 10397 -26765 10431 -26731
rect 10589 -26765 10623 -26731
rect 10940 -26766 10974 -26732
rect 11132 -26766 11166 -26732
rect 11324 -26766 11358 -26732
rect 11516 -26766 11550 -26732
rect -11576 -28186 -11521 -28121
rect -11700 -28433 -11655 -28303
rect -11705 -28764 -11660 -28634
rect -11376 -28756 -11331 -28626
rect -11384 -29039 -11339 -28909
rect 5577 -28059 5611 -27833
rect 6017 -28059 6051 -27833
rect 6457 -28059 6491 -27833
rect 5577 -28313 5611 -28279
rect 6017 -28313 6051 -28279
rect 6457 -28313 6491 -28279
rect 7198 -28880 7232 -28846
rect 7390 -28880 7424 -28846
rect 7582 -28880 7616 -28846
rect 7774 -28880 7808 -28846
rect 8146 -28880 8180 -28846
rect 8338 -28880 8372 -28846
rect 8530 -28880 8564 -28846
rect 8722 -28880 8756 -28846
rect 9082 -28880 9116 -28846
rect 9274 -28880 9308 -28846
rect 9466 -28880 9500 -28846
rect 9658 -28880 9692 -28846
rect 10013 -28880 10047 -28846
rect 10205 -28880 10239 -28846
rect 10397 -28880 10431 -28846
rect 10589 -28880 10623 -28846
rect 10940 -28880 10974 -28846
rect 11132 -28880 11166 -28846
rect 11324 -28880 11358 -28846
rect 11516 -28880 11550 -28846
rect -11552 -29443 -11504 -29395
rect 12170 -30027 12204 -29993
rect -11576 -30795 -11521 -30730
rect -11700 -31042 -11655 -30912
rect -11705 -31373 -11660 -31243
rect -11376 -31365 -11331 -31235
rect -11384 -31648 -11339 -31518
rect 7198 -31294 7232 -31260
rect 7390 -31294 7424 -31260
rect 7582 -31294 7616 -31260
rect 7774 -31294 7808 -31260
rect 8146 -31294 8180 -31260
rect 8338 -31294 8372 -31260
rect 8530 -31294 8564 -31260
rect 8722 -31294 8756 -31260
rect 9082 -31294 9116 -31260
rect 9274 -31294 9308 -31260
rect 9466 -31294 9500 -31260
rect 9658 -31294 9692 -31260
rect 10013 -31293 10047 -31259
rect 12842 -30077 12876 -29851
rect 12313 -30132 12347 -30098
rect 12842 -30331 12876 -30297
rect 10205 -31293 10239 -31259
rect 10397 -31293 10431 -31259
rect 10589 -31293 10623 -31259
rect 10940 -31294 10974 -31260
rect 11132 -31294 11166 -31260
rect 11324 -31294 11358 -31260
rect 11516 -31294 11550 -31260
rect -11554 -31988 -11503 -31937
rect 5577 -32587 5611 -32361
rect 6017 -32587 6051 -32361
rect 6457 -32587 6491 -32361
rect 5577 -32841 5611 -32807
rect 6017 -32841 6051 -32807
rect 6457 -32841 6491 -32807
rect -11578 -33415 -11523 -33350
rect -11702 -33662 -11657 -33532
rect -11707 -33993 -11662 -33863
rect -11378 -33985 -11333 -33855
rect -11386 -34268 -11341 -34138
rect 7198 -33408 7232 -33374
rect 7390 -33408 7424 -33374
rect 7582 -33408 7616 -33374
rect 7774 -33408 7808 -33374
rect 8146 -33408 8180 -33374
rect 8338 -33408 8372 -33374
rect 8530 -33408 8564 -33374
rect 8722 -33408 8756 -33374
rect 9082 -33408 9116 -33374
rect 9274 -33408 9308 -33374
rect 9466 -33408 9500 -33374
rect 9658 -33408 9692 -33374
rect 10013 -33408 10047 -33374
rect 10205 -33408 10239 -33374
rect 10397 -33408 10431 -33374
rect 10589 -33408 10623 -33374
rect 10940 -33408 10974 -33374
rect 11132 -33408 11166 -33374
rect 11324 -33408 11358 -33374
rect 11516 -33408 11550 -33374
rect -11548 -34567 -11514 -34533
rect 12170 -34555 12204 -34521
rect 7198 -35822 7232 -35788
rect 7390 -35822 7424 -35788
rect 7582 -35822 7616 -35788
rect 7774 -35822 7808 -35788
rect 8146 -35822 8180 -35788
rect 8338 -35822 8372 -35788
rect 8530 -35822 8564 -35788
rect 8722 -35822 8756 -35788
rect 9082 -35822 9116 -35788
rect 9274 -35822 9308 -35788
rect 9466 -35822 9500 -35788
rect 9658 -35822 9692 -35788
rect 10013 -35821 10047 -35787
rect 12842 -34605 12876 -34379
rect 12313 -34660 12347 -34626
rect 12842 -34859 12876 -34825
rect 10205 -35821 10239 -35787
rect 10397 -35821 10431 -35787
rect 10589 -35821 10623 -35787
rect 10940 -35822 10974 -35788
rect 12930 -35668 12964 -35634
rect 13184 -35668 13410 -35634
rect 11132 -35822 11166 -35788
rect 11324 -35822 11358 -35788
rect 11516 -35822 11550 -35788
rect 12930 -36047 12964 -36013
rect 13184 -36047 13410 -36013
<< locali >>
rect 1795 6241 3005 6269
rect 1795 6169 1841 6241
rect 2963 6169 3005 6241
rect 1795 6143 3005 6169
rect 3401 6241 4611 6269
rect 3401 6169 3447 6241
rect 4569 6169 4611 6241
rect 3401 6143 4611 6169
rect 5105 6239 6315 6267
rect 5105 6167 5151 6239
rect 6273 6167 6315 6239
rect 5105 6141 6315 6167
rect 1719 6072 1753 6088
rect 1564 5343 1673 5398
rect 1564 5254 1573 5343
rect 1662 5254 1673 5343
rect 1564 5244 1673 5254
rect 1719 5485 1753 5546
rect 1807 6072 1841 6088
rect 1807 5530 1841 5546
rect 1903 6072 1937 6088
rect 1903 5530 1937 5546
rect 1999 6072 2033 6088
rect 1999 5530 2033 5546
rect 2095 6072 2129 6088
rect 2095 5530 2129 5546
rect 2191 6072 2225 6088
rect 2191 5530 2225 5546
rect 2287 6072 2321 6088
rect 2287 5530 2321 5546
rect 2383 6072 2417 6088
rect 2383 5503 2417 5546
rect 2479 6072 2513 6088
rect 2479 5530 2513 5546
rect 2575 6072 2609 6088
rect 2575 5530 2609 5546
rect 2671 6072 2705 6088
rect 2671 5530 2705 5546
rect 2767 6072 2801 6088
rect 2767 5530 2801 5546
rect 2863 6072 2897 6088
rect 2863 5530 2897 5546
rect 2959 6072 2993 6088
rect 2959 5530 2993 5546
rect 3047 6072 3081 6088
rect 1719 5475 2321 5485
rect 1719 5430 2175 5475
rect 2305 5430 2321 5475
rect 1719 5416 2321 5430
rect 1573 5238 1662 5244
rect 1719 5032 1753 5416
rect 1855 5345 2076 5372
rect 1855 5292 1905 5345
rect 2038 5292 2076 5345
rect 1855 5154 2076 5292
rect 1855 5109 1900 5154
rect 2030 5109 2076 5154
rect 1855 5082 2076 5109
rect 2156 5146 2321 5416
rect 2156 5101 2183 5146
rect 2313 5101 2321 5146
rect 2156 5084 2321 5101
rect 2367 5203 2433 5503
rect 3047 5488 3081 5546
rect 2479 5470 3081 5488
rect 2479 5425 2506 5470
rect 2636 5425 3081 5470
rect 3325 6072 3359 6088
rect 3325 5485 3359 5546
rect 3413 6072 3447 6088
rect 3413 5530 3447 5546
rect 3509 6072 3543 6088
rect 3509 5530 3543 5546
rect 3605 6072 3639 6088
rect 3605 5530 3639 5546
rect 3701 6072 3735 6088
rect 3701 5530 3735 5546
rect 3797 6072 3831 6088
rect 3797 5530 3831 5546
rect 3893 6072 3927 6088
rect 3893 5530 3927 5546
rect 3989 6072 4023 6088
rect 3989 5503 4023 5546
rect 4085 6072 4119 6088
rect 4085 5530 4119 5546
rect 4181 6072 4215 6088
rect 4181 5530 4215 5546
rect 4277 6072 4311 6088
rect 4277 5530 4311 5546
rect 4373 6072 4407 6088
rect 4373 5530 4407 5546
rect 4469 6072 4503 6088
rect 4469 5530 4503 5546
rect 4565 6072 4599 6088
rect 4565 5530 4599 5546
rect 4653 6072 4687 6088
rect 5029 6070 5063 6086
rect 3325 5475 3927 5485
rect 2479 5411 3081 5425
rect 2479 5353 2656 5411
rect 2479 5300 2511 5353
rect 2625 5300 2656 5353
rect 2479 5271 2656 5300
rect 2728 5352 2843 5370
rect 2728 5284 2745 5352
rect 2825 5284 2843 5352
rect 2728 5264 2843 5284
rect 2367 5181 3007 5203
rect 2367 5126 2927 5181
rect 2992 5126 3007 5181
rect 2367 5107 3007 5126
rect 2367 5073 2433 5107
rect 1719 4910 1753 4926
rect 1807 5032 1841 5048
rect 1807 4910 1841 4926
rect 1903 5047 1937 5048
rect 1903 4910 1937 4926
rect 1999 5032 2033 5048
rect 1999 4910 2033 4912
rect 2095 5047 2129 5048
rect 2095 4910 2129 4926
rect 2191 5032 2225 5048
rect 2191 4910 2225 4912
rect 2287 5046 2321 5048
rect 2287 4910 2321 4926
rect 2383 5032 2417 5073
rect 2383 4910 2417 4912
rect 2479 5047 2513 5048
rect 2479 4910 2513 4926
rect 2575 5032 2609 5048
rect 2575 4910 2609 4912
rect 2671 5047 2705 5048
rect 2671 4910 2705 4926
rect 2767 5032 2801 5048
rect 2767 4910 2801 4912
rect 2863 5047 2897 5048
rect 2863 4910 2897 4926
rect 2959 5032 2993 5048
rect 2959 4910 2993 4926
rect 3047 5032 3081 5411
rect 3177 5343 3286 5371
rect 3177 5254 3187 5343
rect 3276 5254 3286 5343
rect 3177 5244 3286 5254
rect 3325 5430 3781 5475
rect 3911 5430 3927 5475
rect 3325 5416 3927 5430
rect 3187 5238 3276 5244
rect 3047 4910 3081 4926
rect 3325 5032 3359 5416
rect 3461 5345 3682 5372
rect 3461 5292 3511 5345
rect 3644 5292 3682 5345
rect 3461 5154 3682 5292
rect 3461 5109 3506 5154
rect 3636 5109 3682 5154
rect 3461 5082 3682 5109
rect 3762 5146 3927 5416
rect 3762 5101 3789 5146
rect 3919 5101 3927 5146
rect 3762 5084 3927 5101
rect 3973 5203 4039 5503
rect 4653 5488 4687 5546
rect 4085 5470 4687 5488
rect 4085 5425 4112 5470
rect 4242 5425 4687 5470
rect 4085 5411 4687 5425
rect 4085 5353 4262 5411
rect 4085 5300 4117 5353
rect 4231 5300 4262 5353
rect 4085 5271 4262 5300
rect 4334 5352 4449 5370
rect 4334 5284 4351 5352
rect 4431 5284 4449 5352
rect 4334 5264 4449 5284
rect 3973 5181 4613 5203
rect 3973 5126 4533 5181
rect 4598 5126 4613 5181
rect 3973 5107 4613 5126
rect 3973 5073 4039 5107
rect 3325 4910 3359 4926
rect 3413 5032 3447 5048
rect 3413 4910 3447 4926
rect 3509 5047 3543 5048
rect 3509 4910 3543 4926
rect 3605 5032 3639 5048
rect 3605 4910 3639 4912
rect 3701 5047 3735 5048
rect 3701 4910 3735 4926
rect 3797 5032 3831 5048
rect 3797 4910 3831 4912
rect 3893 5046 3927 5048
rect 3893 4910 3927 4926
rect 3989 5032 4023 5073
rect 3989 4910 4023 4912
rect 4085 5047 4119 5048
rect 4085 4910 4119 4926
rect 4181 5032 4215 5048
rect 4181 4910 4215 4912
rect 4277 5047 4311 5048
rect 4277 4910 4311 4926
rect 4373 5032 4407 5048
rect 4373 4910 4407 4912
rect 4469 5047 4503 5048
rect 4469 4910 4503 4926
rect 4565 5032 4599 5048
rect 4565 4910 4599 4926
rect 4653 5032 4687 5411
rect 4861 5373 4970 5516
rect 5029 5483 5063 5544
rect 5117 6070 5151 6086
rect 5117 5528 5151 5544
rect 5213 6070 5247 6086
rect 5213 5528 5247 5544
rect 5309 6070 5343 6086
rect 5309 5528 5343 5544
rect 5405 6070 5439 6086
rect 5405 5528 5439 5544
rect 5501 6070 5535 6086
rect 5501 5528 5535 5544
rect 5597 6070 5631 6086
rect 5597 5528 5631 5544
rect 5693 6070 5727 6086
rect 5693 5501 5727 5544
rect 5789 6070 5823 6086
rect 5789 5528 5823 5544
rect 5885 6070 5919 6086
rect 5885 5528 5919 5544
rect 5981 6070 6015 6086
rect 5981 5528 6015 5544
rect 6077 6070 6111 6086
rect 6077 5528 6111 5544
rect 6173 6070 6207 6086
rect 6173 5528 6207 5544
rect 6269 6070 6303 6086
rect 6269 5528 6303 5544
rect 6357 6070 6391 6086
rect 5029 5473 5631 5483
rect 5029 5428 5485 5473
rect 5615 5428 5631 5473
rect 5029 5414 5631 5428
rect 4861 5351 4977 5373
rect 4855 5341 4977 5351
rect 4855 5252 4871 5341
rect 4960 5252 4977 5341
rect 4855 5241 4977 5252
rect 4871 5238 4960 5241
rect 4653 4910 4687 4926
rect 5029 5030 5063 5414
rect 5165 5343 5386 5370
rect 5165 5290 5215 5343
rect 5348 5290 5386 5343
rect 5165 5152 5386 5290
rect 5165 5107 5210 5152
rect 5340 5107 5386 5152
rect 5165 5080 5386 5107
rect 5466 5144 5631 5414
rect 5466 5099 5493 5144
rect 5623 5099 5631 5144
rect 5466 5082 5631 5099
rect 5677 5201 5743 5501
rect 6357 5486 6391 5544
rect 6951 5507 6967 5554
rect 7536 5507 7560 5554
rect 7856 5497 7872 5531
rect 7963 5497 7979 5531
rect 5789 5468 6391 5486
rect 5789 5423 5816 5468
rect 5946 5423 6391 5468
rect 5789 5409 6391 5423
rect 5789 5351 5966 5409
rect 5789 5298 5821 5351
rect 5935 5298 5966 5351
rect 5789 5269 5966 5298
rect 6038 5350 6153 5368
rect 6038 5282 6055 5350
rect 6135 5282 6153 5350
rect 6038 5262 6153 5282
rect 5677 5179 6317 5201
rect 5677 5124 6237 5179
rect 6302 5124 6317 5179
rect 5677 5105 6317 5124
rect 5677 5071 5743 5105
rect 5029 4908 5063 4924
rect 5117 5030 5151 5046
rect 5117 4908 5151 4924
rect 5213 5045 5247 5046
rect 5213 4908 5247 4924
rect 5309 5030 5343 5046
rect 5309 4908 5343 4910
rect 5405 5045 5439 5046
rect 5405 4908 5439 4924
rect 5501 5030 5535 5046
rect 5501 4908 5535 4910
rect 5597 5044 5631 5046
rect 5597 4908 5631 4924
rect 5693 5030 5727 5071
rect 5693 4908 5727 4910
rect 5789 5045 5823 5046
rect 5789 4908 5823 4924
rect 5885 5030 5919 5046
rect 5885 4908 5919 4910
rect 5981 5045 6015 5046
rect 5981 4908 6015 4924
rect 6077 5030 6111 5046
rect 6077 4908 6111 4910
rect 6173 5045 6207 5046
rect 6173 4908 6207 4924
rect 6269 5030 6303 5046
rect 6269 4908 6303 4924
rect 6357 5030 6391 5409
rect 6951 5435 6985 5445
rect 6951 5223 6985 5239
rect 7047 5429 7081 5445
rect 7047 5223 7081 5233
rect 7143 5435 7177 5445
rect 7143 5223 7177 5239
rect 7239 5429 7273 5445
rect 7239 5223 7273 5233
rect 7335 5435 7369 5445
rect 7335 5223 7369 5239
rect 7431 5429 7465 5445
rect 7431 5223 7465 5233
rect 7527 5435 7561 5445
rect 7527 5223 7561 5239
rect 7712 5411 7762 5428
rect 7805 5425 7815 5459
rect 8011 5425 8027 5459
rect 7712 5185 7728 5411
rect 7805 5329 7821 5363
rect 8015 5329 8033 5363
rect 7805 5233 7815 5267
rect 8011 5233 8027 5267
rect 6357 4908 6391 4924
rect 7000 5145 7017 5180
rect 7051 5145 7067 5180
rect 7289 5174 7306 5180
rect 7101 5145 7306 5174
rect 7340 5145 7356 5180
rect 7000 4939 7043 5145
rect 7101 5140 7356 5145
rect 7101 5056 7135 5140
rect 7169 5051 7185 5085
rect 7561 5051 7577 5085
rect 7101 5005 7135 5021
rect 7712 4965 7762 5185
rect 7805 5137 7821 5171
rect 8015 5137 8033 5171
rect 7805 4975 7821 5009
rect 7997 4975 8013 5009
rect 7000 4923 7135 4939
rect 7000 4888 7101 4923
rect 7712 4931 7728 4965
rect 7712 4915 7762 4931
rect 7000 4872 7135 4888
rect 1800 4838 3002 4860
rect 1800 4792 1841 4838
rect 2964 4792 3002 4838
rect 1800 4769 3002 4792
rect 3406 4838 4608 4860
rect 7169 4859 7185 4893
rect 7561 4859 7577 4893
rect 7805 4887 7821 4921
rect 7997 4887 8013 4921
rect 3406 4792 3447 4838
rect 4570 4792 4608 4838
rect 3406 4769 4608 4792
rect 5110 4836 6312 4858
rect 5110 4790 5151 4836
rect 6274 4790 6312 4836
rect 5110 4767 6312 4790
rect 7173 4787 7200 4821
rect 7535 4787 7573 4821
rect 7824 4785 7840 4819
rect 7972 4785 7988 4819
rect -24042 4517 -22832 4545
rect -24042 4445 -24000 4517
rect -22878 4445 -22832 4517
rect -24042 4419 -22832 4445
rect -20751 4517 -19541 4545
rect -20751 4445 -20709 4517
rect -19587 4445 -19541 4517
rect -20751 4419 -19541 4445
rect -17460 4517 -16250 4545
rect -17460 4445 -17418 4517
rect -16296 4445 -16250 4517
rect -17460 4419 -16250 4445
rect -14169 4517 -12959 4545
rect -14169 4445 -14127 4517
rect -13005 4445 -12959 4517
rect -14169 4419 -12959 4445
rect -10878 4517 -9668 4545
rect -10878 4445 -10836 4517
rect -9714 4445 -9668 4517
rect -10878 4419 -9668 4445
rect -7588 4517 -6378 4545
rect -7588 4445 -7546 4517
rect -6424 4445 -6378 4517
rect -7588 4419 -6378 4445
rect -4297 4517 -3087 4545
rect -4297 4445 -4255 4517
rect -3133 4445 -3087 4517
rect -4297 4419 -3087 4445
rect -1006 4517 204 4545
rect -1006 4445 -964 4517
rect 158 4445 204 4517
rect -1006 4419 204 4445
rect -24118 4348 -24084 4364
rect -24118 3764 -24084 3822
rect -24030 4348 -23996 4364
rect -24030 3806 -23996 3822
rect -23934 4348 -23900 4364
rect -23934 3806 -23900 3822
rect -23838 4348 -23804 4364
rect -23838 3806 -23804 3822
rect -23742 4348 -23708 4364
rect -23742 3806 -23708 3822
rect -23646 4348 -23612 4364
rect -23646 3806 -23612 3822
rect -23550 4348 -23516 4364
rect -23550 3806 -23516 3822
rect -23454 4348 -23420 4364
rect -23454 3779 -23420 3822
rect -23358 4348 -23324 4364
rect -23358 3806 -23324 3822
rect -23262 4348 -23228 4364
rect -23262 3806 -23228 3822
rect -23166 4348 -23132 4364
rect -23166 3806 -23132 3822
rect -23070 4348 -23036 4364
rect -23070 3806 -23036 3822
rect -22974 4348 -22940 4364
rect -22974 3806 -22940 3822
rect -22878 4348 -22844 4364
rect -22878 3806 -22844 3822
rect -22790 4348 -22756 4364
rect -24118 3746 -23516 3764
rect -24118 3701 -23673 3746
rect -23543 3701 -23516 3746
rect -24118 3687 -23516 3701
rect -24118 3308 -24084 3687
rect -23880 3628 -23765 3646
rect -23880 3560 -23862 3628
rect -23782 3560 -23765 3628
rect -23880 3540 -23765 3560
rect -23693 3629 -23516 3687
rect -23693 3576 -23662 3629
rect -23548 3576 -23516 3629
rect -23693 3547 -23516 3576
rect -23470 3479 -23404 3779
rect -22790 3761 -22756 3822
rect -20827 4348 -20793 4364
rect -24044 3457 -23404 3479
rect -24044 3402 -24029 3457
rect -23964 3402 -23404 3457
rect -24044 3383 -23404 3402
rect -23470 3349 -23404 3383
rect -23358 3751 -22756 3761
rect -23358 3706 -23342 3751
rect -23212 3706 -22756 3751
rect -23358 3692 -22756 3706
rect -23358 3422 -23193 3692
rect -23358 3377 -23350 3422
rect -23220 3377 -23193 3422
rect -23358 3360 -23193 3377
rect -23113 3621 -22892 3648
rect -23113 3568 -23075 3621
rect -22942 3568 -22892 3621
rect -23113 3430 -22892 3568
rect -23113 3385 -23067 3430
rect -22937 3385 -22892 3430
rect -23113 3358 -22892 3385
rect -24118 3186 -24084 3202
rect -24030 3308 -23996 3324
rect -24030 3186 -23996 3202
rect -23934 3323 -23900 3324
rect -23934 3186 -23900 3202
rect -23838 3308 -23804 3324
rect -23838 3186 -23804 3188
rect -23742 3323 -23708 3324
rect -23742 3186 -23708 3202
rect -23646 3308 -23612 3324
rect -23646 3186 -23612 3188
rect -23550 3323 -23516 3324
rect -23550 3186 -23516 3202
rect -23454 3308 -23420 3349
rect -23454 3186 -23420 3188
rect -23358 3322 -23324 3324
rect -23358 3186 -23324 3202
rect -23262 3308 -23228 3324
rect -23262 3186 -23228 3188
rect -23166 3323 -23132 3324
rect -23166 3186 -23132 3202
rect -23070 3308 -23036 3324
rect -23070 3186 -23036 3188
rect -22974 3323 -22940 3324
rect -22974 3186 -22940 3202
rect -22878 3308 -22844 3324
rect -22878 3186 -22844 3202
rect -22790 3308 -22756 3692
rect -22712 3767 -22461 3784
rect -22712 3547 -22680 3767
rect -22488 3547 -22461 3767
rect -22712 3521 -22461 3547
rect -20827 3764 -20793 3822
rect -20739 4348 -20705 4364
rect -20739 3806 -20705 3822
rect -20643 4348 -20609 4364
rect -20643 3806 -20609 3822
rect -20547 4348 -20513 4364
rect -20547 3806 -20513 3822
rect -20451 4348 -20417 4364
rect -20451 3806 -20417 3822
rect -20355 4348 -20321 4364
rect -20355 3806 -20321 3822
rect -20259 4348 -20225 4364
rect -20259 3806 -20225 3822
rect -20163 4348 -20129 4364
rect -20163 3779 -20129 3822
rect -20067 4348 -20033 4364
rect -20067 3806 -20033 3822
rect -19971 4348 -19937 4364
rect -19971 3806 -19937 3822
rect -19875 4348 -19841 4364
rect -19875 3806 -19841 3822
rect -19779 4348 -19745 4364
rect -19779 3806 -19745 3822
rect -19683 4348 -19649 4364
rect -19683 3806 -19649 3822
rect -19587 4348 -19553 4364
rect -19587 3806 -19553 3822
rect -19499 4348 -19465 4364
rect -20827 3746 -20225 3764
rect -20827 3701 -20382 3746
rect -20252 3701 -20225 3746
rect -20827 3687 -20225 3701
rect -22790 3186 -22756 3202
rect -20827 3308 -20793 3687
rect -20589 3628 -20474 3646
rect -20589 3560 -20571 3628
rect -20491 3560 -20474 3628
rect -20589 3540 -20474 3560
rect -20402 3629 -20225 3687
rect -20402 3576 -20371 3629
rect -20257 3576 -20225 3629
rect -20402 3547 -20225 3576
rect -20179 3479 -20113 3779
rect -19499 3761 -19465 3822
rect -17536 4348 -17502 4364
rect -20753 3457 -20113 3479
rect -20753 3402 -20738 3457
rect -20673 3402 -20113 3457
rect -20753 3383 -20113 3402
rect -20179 3349 -20113 3383
rect -20067 3751 -19465 3761
rect -20067 3706 -20051 3751
rect -19921 3706 -19465 3751
rect -20067 3692 -19465 3706
rect -20067 3422 -19902 3692
rect -20067 3377 -20059 3422
rect -19929 3377 -19902 3422
rect -20067 3360 -19902 3377
rect -19822 3621 -19601 3648
rect -19822 3568 -19784 3621
rect -19651 3568 -19601 3621
rect -19822 3430 -19601 3568
rect -19822 3385 -19776 3430
rect -19646 3385 -19601 3430
rect -19822 3358 -19601 3385
rect -20827 3186 -20793 3202
rect -20739 3308 -20705 3324
rect -20739 3186 -20705 3202
rect -20643 3323 -20609 3324
rect -20643 3186 -20609 3202
rect -20547 3308 -20513 3324
rect -20547 3186 -20513 3188
rect -20451 3323 -20417 3324
rect -20451 3186 -20417 3202
rect -20355 3308 -20321 3324
rect -20355 3186 -20321 3188
rect -20259 3323 -20225 3324
rect -20259 3186 -20225 3202
rect -20163 3308 -20129 3349
rect -20163 3186 -20129 3188
rect -20067 3322 -20033 3324
rect -20067 3186 -20033 3202
rect -19971 3308 -19937 3324
rect -19971 3186 -19937 3188
rect -19875 3323 -19841 3324
rect -19875 3186 -19841 3202
rect -19779 3308 -19745 3324
rect -19779 3186 -19745 3188
rect -19683 3323 -19649 3324
rect -19683 3186 -19649 3202
rect -19587 3308 -19553 3324
rect -19587 3186 -19553 3202
rect -19499 3308 -19465 3692
rect -19421 3767 -19170 3784
rect -19421 3547 -19389 3767
rect -19197 3547 -19170 3767
rect -19421 3521 -19170 3547
rect -17536 3764 -17502 3822
rect -17448 4348 -17414 4364
rect -17448 3806 -17414 3822
rect -17352 4348 -17318 4364
rect -17352 3806 -17318 3822
rect -17256 4348 -17222 4364
rect -17256 3806 -17222 3822
rect -17160 4348 -17126 4364
rect -17160 3806 -17126 3822
rect -17064 4348 -17030 4364
rect -17064 3806 -17030 3822
rect -16968 4348 -16934 4364
rect -16968 3806 -16934 3822
rect -16872 4348 -16838 4364
rect -16872 3779 -16838 3822
rect -16776 4348 -16742 4364
rect -16776 3806 -16742 3822
rect -16680 4348 -16646 4364
rect -16680 3806 -16646 3822
rect -16584 4348 -16550 4364
rect -16584 3806 -16550 3822
rect -16488 4348 -16454 4364
rect -16488 3806 -16454 3822
rect -16392 4348 -16358 4364
rect -16392 3806 -16358 3822
rect -16296 4348 -16262 4364
rect -16296 3806 -16262 3822
rect -16208 4348 -16174 4364
rect -17536 3746 -16934 3764
rect -17536 3701 -17091 3746
rect -16961 3701 -16934 3746
rect -17536 3687 -16934 3701
rect -19499 3186 -19465 3202
rect -17536 3308 -17502 3687
rect -17298 3628 -17183 3646
rect -17298 3560 -17280 3628
rect -17200 3560 -17183 3628
rect -17298 3540 -17183 3560
rect -17111 3629 -16934 3687
rect -17111 3576 -17080 3629
rect -16966 3576 -16934 3629
rect -17111 3547 -16934 3576
rect -16888 3479 -16822 3779
rect -16208 3761 -16174 3822
rect -14245 4348 -14211 4364
rect -17462 3457 -16822 3479
rect -17462 3402 -17447 3457
rect -17382 3402 -16822 3457
rect -17462 3383 -16822 3402
rect -16888 3349 -16822 3383
rect -16776 3751 -16174 3761
rect -16776 3706 -16760 3751
rect -16630 3706 -16174 3751
rect -16776 3692 -16174 3706
rect -16776 3422 -16611 3692
rect -16776 3377 -16768 3422
rect -16638 3377 -16611 3422
rect -16776 3360 -16611 3377
rect -16531 3621 -16310 3648
rect -16531 3568 -16493 3621
rect -16360 3568 -16310 3621
rect -16531 3430 -16310 3568
rect -16531 3385 -16485 3430
rect -16355 3385 -16310 3430
rect -16531 3358 -16310 3385
rect -17536 3186 -17502 3202
rect -17448 3308 -17414 3324
rect -17448 3186 -17414 3202
rect -17352 3323 -17318 3324
rect -17352 3186 -17318 3202
rect -17256 3308 -17222 3324
rect -17256 3186 -17222 3188
rect -17160 3323 -17126 3324
rect -17160 3186 -17126 3202
rect -17064 3308 -17030 3324
rect -17064 3186 -17030 3188
rect -16968 3323 -16934 3324
rect -16968 3186 -16934 3202
rect -16872 3308 -16838 3349
rect -16872 3186 -16838 3188
rect -16776 3322 -16742 3324
rect -16776 3186 -16742 3202
rect -16680 3308 -16646 3324
rect -16680 3186 -16646 3188
rect -16584 3323 -16550 3324
rect -16584 3186 -16550 3202
rect -16488 3308 -16454 3324
rect -16488 3186 -16454 3188
rect -16392 3323 -16358 3324
rect -16392 3186 -16358 3202
rect -16296 3308 -16262 3324
rect -16296 3186 -16262 3202
rect -16208 3308 -16174 3692
rect -16130 3767 -15879 3784
rect -16130 3547 -16098 3767
rect -15906 3547 -15879 3767
rect -16130 3521 -15879 3547
rect -14245 3764 -14211 3822
rect -14157 4348 -14123 4364
rect -14157 3806 -14123 3822
rect -14061 4348 -14027 4364
rect -14061 3806 -14027 3822
rect -13965 4348 -13931 4364
rect -13965 3806 -13931 3822
rect -13869 4348 -13835 4364
rect -13869 3806 -13835 3822
rect -13773 4348 -13739 4364
rect -13773 3806 -13739 3822
rect -13677 4348 -13643 4364
rect -13677 3806 -13643 3822
rect -13581 4348 -13547 4364
rect -13581 3779 -13547 3822
rect -13485 4348 -13451 4364
rect -13485 3806 -13451 3822
rect -13389 4348 -13355 4364
rect -13389 3806 -13355 3822
rect -13293 4348 -13259 4364
rect -13293 3806 -13259 3822
rect -13197 4348 -13163 4364
rect -13197 3806 -13163 3822
rect -13101 4348 -13067 4364
rect -13101 3806 -13067 3822
rect -13005 4348 -12971 4364
rect -13005 3806 -12971 3822
rect -12917 4348 -12883 4364
rect -14245 3746 -13643 3764
rect -14245 3701 -13800 3746
rect -13670 3701 -13643 3746
rect -14245 3687 -13643 3701
rect -16208 3186 -16174 3202
rect -14245 3308 -14211 3687
rect -14007 3628 -13892 3646
rect -14007 3560 -13989 3628
rect -13909 3560 -13892 3628
rect -14007 3540 -13892 3560
rect -13820 3629 -13643 3687
rect -13820 3576 -13789 3629
rect -13675 3576 -13643 3629
rect -13820 3547 -13643 3576
rect -13597 3479 -13531 3779
rect -12917 3761 -12883 3822
rect -10954 4348 -10920 4364
rect -14171 3457 -13531 3479
rect -14171 3402 -14156 3457
rect -14091 3402 -13531 3457
rect -14171 3383 -13531 3402
rect -13597 3349 -13531 3383
rect -13485 3751 -12883 3761
rect -13485 3706 -13469 3751
rect -13339 3706 -12883 3751
rect -13485 3692 -12883 3706
rect -13485 3422 -13320 3692
rect -13485 3377 -13477 3422
rect -13347 3377 -13320 3422
rect -13485 3360 -13320 3377
rect -13240 3621 -13019 3648
rect -13240 3568 -13202 3621
rect -13069 3568 -13019 3621
rect -13240 3430 -13019 3568
rect -13240 3385 -13194 3430
rect -13064 3385 -13019 3430
rect -13240 3358 -13019 3385
rect -14245 3186 -14211 3202
rect -14157 3308 -14123 3324
rect -14157 3186 -14123 3202
rect -14061 3323 -14027 3324
rect -14061 3186 -14027 3202
rect -13965 3308 -13931 3324
rect -13965 3186 -13931 3188
rect -13869 3323 -13835 3324
rect -13869 3186 -13835 3202
rect -13773 3308 -13739 3324
rect -13773 3186 -13739 3188
rect -13677 3323 -13643 3324
rect -13677 3186 -13643 3202
rect -13581 3308 -13547 3349
rect -13581 3186 -13547 3188
rect -13485 3322 -13451 3324
rect -13485 3186 -13451 3202
rect -13389 3308 -13355 3324
rect -13389 3186 -13355 3188
rect -13293 3323 -13259 3324
rect -13293 3186 -13259 3202
rect -13197 3308 -13163 3324
rect -13197 3186 -13163 3188
rect -13101 3323 -13067 3324
rect -13101 3186 -13067 3202
rect -13005 3308 -12971 3324
rect -13005 3186 -12971 3202
rect -12917 3308 -12883 3692
rect -12839 3767 -12588 3784
rect -12839 3547 -12807 3767
rect -12615 3547 -12588 3767
rect -12839 3521 -12588 3547
rect -10954 3764 -10920 3822
rect -10866 4348 -10832 4364
rect -10866 3806 -10832 3822
rect -10770 4348 -10736 4364
rect -10770 3806 -10736 3822
rect -10674 4348 -10640 4364
rect -10674 3806 -10640 3822
rect -10578 4348 -10544 4364
rect -10578 3806 -10544 3822
rect -10482 4348 -10448 4364
rect -10482 3806 -10448 3822
rect -10386 4348 -10352 4364
rect -10386 3806 -10352 3822
rect -10290 4348 -10256 4364
rect -10290 3779 -10256 3822
rect -10194 4348 -10160 4364
rect -10194 3806 -10160 3822
rect -10098 4348 -10064 4364
rect -10098 3806 -10064 3822
rect -10002 4348 -9968 4364
rect -10002 3806 -9968 3822
rect -9906 4348 -9872 4364
rect -9906 3806 -9872 3822
rect -9810 4348 -9776 4364
rect -9810 3806 -9776 3822
rect -9714 4348 -9680 4364
rect -9714 3806 -9680 3822
rect -9626 4348 -9592 4364
rect -10954 3746 -10352 3764
rect -10954 3701 -10509 3746
rect -10379 3701 -10352 3746
rect -10954 3687 -10352 3701
rect -12917 3186 -12883 3202
rect -10954 3308 -10920 3687
rect -10716 3628 -10601 3646
rect -10716 3560 -10698 3628
rect -10618 3560 -10601 3628
rect -10716 3540 -10601 3560
rect -10529 3629 -10352 3687
rect -10529 3576 -10498 3629
rect -10384 3576 -10352 3629
rect -10529 3547 -10352 3576
rect -10306 3479 -10240 3779
rect -9626 3761 -9592 3822
rect -7664 4348 -7630 4364
rect -10880 3457 -10240 3479
rect -10880 3402 -10865 3457
rect -10800 3402 -10240 3457
rect -10880 3383 -10240 3402
rect -10306 3349 -10240 3383
rect -10194 3751 -9592 3761
rect -10194 3706 -10178 3751
rect -10048 3706 -9592 3751
rect -10194 3692 -9592 3706
rect -10194 3422 -10029 3692
rect -10194 3377 -10186 3422
rect -10056 3377 -10029 3422
rect -10194 3360 -10029 3377
rect -9949 3621 -9728 3648
rect -9949 3568 -9911 3621
rect -9778 3568 -9728 3621
rect -9949 3430 -9728 3568
rect -9949 3385 -9903 3430
rect -9773 3385 -9728 3430
rect -9949 3358 -9728 3385
rect -10954 3186 -10920 3202
rect -10866 3308 -10832 3324
rect -10866 3186 -10832 3202
rect -10770 3323 -10736 3324
rect -10770 3186 -10736 3202
rect -10674 3308 -10640 3324
rect -10674 3186 -10640 3188
rect -10578 3323 -10544 3324
rect -10578 3186 -10544 3202
rect -10482 3308 -10448 3324
rect -10482 3186 -10448 3188
rect -10386 3323 -10352 3324
rect -10386 3186 -10352 3202
rect -10290 3308 -10256 3349
rect -10290 3186 -10256 3188
rect -10194 3322 -10160 3324
rect -10194 3186 -10160 3202
rect -10098 3308 -10064 3324
rect -10098 3186 -10064 3188
rect -10002 3323 -9968 3324
rect -10002 3186 -9968 3202
rect -9906 3308 -9872 3324
rect -9906 3186 -9872 3188
rect -9810 3323 -9776 3324
rect -9810 3186 -9776 3202
rect -9714 3308 -9680 3324
rect -9714 3186 -9680 3202
rect -9626 3308 -9592 3692
rect -9548 3767 -9297 3784
rect -9548 3547 -9516 3767
rect -9324 3547 -9297 3767
rect -9548 3521 -9297 3547
rect -7664 3764 -7630 3822
rect -7576 4348 -7542 4364
rect -7576 3806 -7542 3822
rect -7480 4348 -7446 4364
rect -7480 3806 -7446 3822
rect -7384 4348 -7350 4364
rect -7384 3806 -7350 3822
rect -7288 4348 -7254 4364
rect -7288 3806 -7254 3822
rect -7192 4348 -7158 4364
rect -7192 3806 -7158 3822
rect -7096 4348 -7062 4364
rect -7096 3806 -7062 3822
rect -7000 4348 -6966 4364
rect -7000 3779 -6966 3822
rect -6904 4348 -6870 4364
rect -6904 3806 -6870 3822
rect -6808 4348 -6774 4364
rect -6808 3806 -6774 3822
rect -6712 4348 -6678 4364
rect -6712 3806 -6678 3822
rect -6616 4348 -6582 4364
rect -6616 3806 -6582 3822
rect -6520 4348 -6486 4364
rect -6520 3806 -6486 3822
rect -6424 4348 -6390 4364
rect -6424 3806 -6390 3822
rect -6336 4348 -6302 4364
rect -7664 3746 -7062 3764
rect -7664 3701 -7219 3746
rect -7089 3701 -7062 3746
rect -7664 3687 -7062 3701
rect -9626 3186 -9592 3202
rect -7664 3308 -7630 3687
rect -7426 3628 -7311 3646
rect -7426 3560 -7408 3628
rect -7328 3560 -7311 3628
rect -7426 3540 -7311 3560
rect -7239 3629 -7062 3687
rect -7239 3576 -7208 3629
rect -7094 3576 -7062 3629
rect -7239 3547 -7062 3576
rect -7016 3479 -6950 3779
rect -6336 3761 -6302 3822
rect -4373 4348 -4339 4364
rect -7590 3457 -6950 3479
rect -7590 3402 -7575 3457
rect -7510 3402 -6950 3457
rect -7590 3383 -6950 3402
rect -7016 3349 -6950 3383
rect -6904 3751 -6302 3761
rect -6904 3706 -6888 3751
rect -6758 3706 -6302 3751
rect -6904 3692 -6302 3706
rect -6904 3422 -6739 3692
rect -6904 3377 -6896 3422
rect -6766 3377 -6739 3422
rect -6904 3360 -6739 3377
rect -6659 3621 -6438 3648
rect -6659 3568 -6621 3621
rect -6488 3568 -6438 3621
rect -6659 3430 -6438 3568
rect -6659 3385 -6613 3430
rect -6483 3385 -6438 3430
rect -6659 3358 -6438 3385
rect -7664 3186 -7630 3202
rect -7576 3308 -7542 3324
rect -7576 3186 -7542 3202
rect -7480 3323 -7446 3324
rect -7480 3186 -7446 3202
rect -7384 3308 -7350 3324
rect -7384 3186 -7350 3188
rect -7288 3323 -7254 3324
rect -7288 3186 -7254 3202
rect -7192 3308 -7158 3324
rect -7192 3186 -7158 3188
rect -7096 3323 -7062 3324
rect -7096 3186 -7062 3202
rect -7000 3308 -6966 3349
rect -7000 3186 -6966 3188
rect -6904 3322 -6870 3324
rect -6904 3186 -6870 3202
rect -6808 3308 -6774 3324
rect -6808 3186 -6774 3188
rect -6712 3323 -6678 3324
rect -6712 3186 -6678 3202
rect -6616 3308 -6582 3324
rect -6616 3186 -6582 3188
rect -6520 3323 -6486 3324
rect -6520 3186 -6486 3202
rect -6424 3308 -6390 3324
rect -6424 3186 -6390 3202
rect -6336 3308 -6302 3692
rect -6258 3767 -6007 3784
rect -6258 3547 -6226 3767
rect -6034 3547 -6007 3767
rect -6258 3521 -6007 3547
rect -4373 3764 -4339 3822
rect -4285 4348 -4251 4364
rect -4285 3806 -4251 3822
rect -4189 4348 -4155 4364
rect -4189 3806 -4155 3822
rect -4093 4348 -4059 4364
rect -4093 3806 -4059 3822
rect -3997 4348 -3963 4364
rect -3997 3806 -3963 3822
rect -3901 4348 -3867 4364
rect -3901 3806 -3867 3822
rect -3805 4348 -3771 4364
rect -3805 3806 -3771 3822
rect -3709 4348 -3675 4364
rect -3709 3779 -3675 3822
rect -3613 4348 -3579 4364
rect -3613 3806 -3579 3822
rect -3517 4348 -3483 4364
rect -3517 3806 -3483 3822
rect -3421 4348 -3387 4364
rect -3421 3806 -3387 3822
rect -3325 4348 -3291 4364
rect -3325 3806 -3291 3822
rect -3229 4348 -3195 4364
rect -3229 3806 -3195 3822
rect -3133 4348 -3099 4364
rect -3133 3806 -3099 3822
rect -3045 4348 -3011 4364
rect -4373 3746 -3771 3764
rect -4373 3701 -3928 3746
rect -3798 3701 -3771 3746
rect -4373 3687 -3771 3701
rect -6336 3186 -6302 3202
rect -4373 3308 -4339 3687
rect -4135 3628 -4020 3646
rect -4135 3560 -4117 3628
rect -4037 3560 -4020 3628
rect -4135 3540 -4020 3560
rect -3948 3629 -3771 3687
rect -3948 3576 -3917 3629
rect -3803 3576 -3771 3629
rect -3948 3547 -3771 3576
rect -3725 3479 -3659 3779
rect -3045 3761 -3011 3822
rect -1082 4348 -1048 4364
rect -4299 3457 -3659 3479
rect -4299 3402 -4284 3457
rect -4219 3402 -3659 3457
rect -4299 3383 -3659 3402
rect -3725 3349 -3659 3383
rect -3613 3751 -3011 3761
rect -3613 3706 -3597 3751
rect -3467 3706 -3011 3751
rect -3613 3692 -3011 3706
rect -3613 3422 -3448 3692
rect -3613 3377 -3605 3422
rect -3475 3377 -3448 3422
rect -3613 3360 -3448 3377
rect -3368 3621 -3147 3648
rect -3368 3568 -3330 3621
rect -3197 3568 -3147 3621
rect -3368 3430 -3147 3568
rect -3368 3385 -3322 3430
rect -3192 3385 -3147 3430
rect -3368 3358 -3147 3385
rect -4373 3186 -4339 3202
rect -4285 3308 -4251 3324
rect -4285 3186 -4251 3202
rect -4189 3323 -4155 3324
rect -4189 3186 -4155 3202
rect -4093 3308 -4059 3324
rect -4093 3186 -4059 3188
rect -3997 3323 -3963 3324
rect -3997 3186 -3963 3202
rect -3901 3308 -3867 3324
rect -3901 3186 -3867 3188
rect -3805 3323 -3771 3324
rect -3805 3186 -3771 3202
rect -3709 3308 -3675 3349
rect -3709 3186 -3675 3188
rect -3613 3322 -3579 3324
rect -3613 3186 -3579 3202
rect -3517 3308 -3483 3324
rect -3517 3186 -3483 3188
rect -3421 3323 -3387 3324
rect -3421 3186 -3387 3202
rect -3325 3308 -3291 3324
rect -3325 3186 -3291 3188
rect -3229 3323 -3195 3324
rect -3229 3186 -3195 3202
rect -3133 3308 -3099 3324
rect -3133 3186 -3099 3202
rect -3045 3308 -3011 3692
rect -2967 3767 -2716 3784
rect -2967 3547 -2935 3767
rect -2743 3547 -2716 3767
rect -2967 3521 -2716 3547
rect -1082 3764 -1048 3822
rect -994 4348 -960 4364
rect -994 3806 -960 3822
rect -898 4348 -864 4364
rect -898 3806 -864 3822
rect -802 4348 -768 4364
rect -802 3806 -768 3822
rect -706 4348 -672 4364
rect -706 3806 -672 3822
rect -610 4348 -576 4364
rect -610 3806 -576 3822
rect -514 4348 -480 4364
rect -514 3806 -480 3822
rect -418 4348 -384 4364
rect -418 3779 -384 3822
rect -322 4348 -288 4364
rect -322 3806 -288 3822
rect -226 4348 -192 4364
rect -226 3806 -192 3822
rect -130 4348 -96 4364
rect -130 3806 -96 3822
rect -34 4348 0 4364
rect -34 3806 0 3822
rect 62 4348 96 4364
rect 62 3806 96 3822
rect 158 4348 192 4364
rect 158 3806 192 3822
rect 246 4348 280 4364
rect 5705 3949 5721 3983
rect 5812 3949 5828 3983
rect 6145 3949 6161 3983
rect 6252 3949 6268 3983
rect 6585 3949 6601 3983
rect 6692 3949 6708 3983
rect -1082 3746 -480 3764
rect -1082 3701 -637 3746
rect -507 3701 -480 3746
rect -1082 3687 -480 3701
rect -3045 3186 -3011 3202
rect -1082 3308 -1048 3687
rect -844 3628 -729 3646
rect -844 3560 -826 3628
rect -746 3560 -729 3628
rect -844 3540 -729 3560
rect -657 3629 -480 3687
rect -657 3576 -626 3629
rect -512 3576 -480 3629
rect -657 3547 -480 3576
rect -434 3479 -368 3779
rect 246 3761 280 3822
rect 5561 3863 5611 3880
rect 5654 3877 5664 3911
rect 5860 3877 5876 3911
rect -1008 3457 -368 3479
rect -1008 3402 -993 3457
rect -928 3402 -368 3457
rect -1008 3383 -368 3402
rect -434 3349 -368 3383
rect -322 3751 280 3761
rect -322 3706 -306 3751
rect -176 3706 280 3751
rect -322 3692 280 3706
rect -322 3422 -157 3692
rect -322 3377 -314 3422
rect -184 3377 -157 3422
rect -322 3360 -157 3377
rect -77 3621 144 3648
rect -77 3568 -39 3621
rect 94 3568 144 3621
rect -77 3430 144 3568
rect -77 3385 -31 3430
rect 99 3385 144 3430
rect -77 3358 144 3385
rect -1082 3186 -1048 3202
rect -994 3308 -960 3324
rect -994 3186 -960 3202
rect -898 3323 -864 3324
rect -898 3186 -864 3202
rect -802 3308 -768 3324
rect -802 3186 -768 3188
rect -706 3323 -672 3324
rect -706 3186 -672 3202
rect -610 3308 -576 3324
rect -610 3186 -576 3188
rect -514 3323 -480 3324
rect -514 3186 -480 3202
rect -418 3308 -384 3349
rect -418 3186 -384 3188
rect -322 3322 -288 3324
rect -322 3186 -288 3202
rect -226 3308 -192 3324
rect -226 3186 -192 3188
rect -130 3323 -96 3324
rect -130 3186 -96 3202
rect -34 3308 0 3324
rect -34 3186 0 3188
rect 62 3323 96 3324
rect 62 3186 96 3202
rect 158 3308 192 3324
rect 158 3186 192 3202
rect 246 3308 280 3692
rect 324 3767 575 3784
rect 324 3547 356 3767
rect 548 3547 575 3767
rect 324 3521 575 3547
rect 5561 3637 5577 3863
rect 6001 3863 6051 3880
rect 6094 3877 6104 3911
rect 6300 3877 6316 3911
rect 5654 3781 5670 3815
rect 5864 3781 5882 3815
rect 5654 3685 5664 3719
rect 5860 3685 5876 3719
rect 5561 3417 5611 3637
rect 6001 3637 6017 3863
rect 6441 3863 6491 3880
rect 6534 3877 6544 3911
rect 6740 3877 6756 3911
rect 6094 3781 6110 3815
rect 6304 3781 6322 3815
rect 6094 3685 6104 3719
rect 6300 3685 6316 3719
rect 5654 3589 5670 3623
rect 5864 3589 5882 3623
rect 5654 3427 5670 3461
rect 5846 3427 5862 3461
rect 5561 3383 5577 3417
rect 5561 3367 5611 3383
rect 6001 3417 6051 3637
rect 6441 3637 6457 3863
rect 6534 3781 6550 3815
rect 6744 3781 6762 3815
rect 6534 3685 6544 3719
rect 6740 3685 6756 3719
rect 6094 3589 6110 3623
rect 6304 3589 6322 3623
rect 6094 3427 6110 3461
rect 6286 3427 6302 3461
rect 6001 3383 6017 3417
rect 5654 3339 5670 3373
rect 5846 3339 5862 3373
rect 6001 3367 6051 3383
rect 6441 3417 6491 3637
rect 6534 3589 6550 3623
rect 6744 3589 6762 3623
rect 6534 3427 6550 3461
rect 6726 3427 6742 3461
rect 6441 3383 6457 3417
rect 6094 3339 6110 3373
rect 6286 3339 6302 3373
rect 6441 3367 6491 3383
rect 6534 3339 6550 3373
rect 6726 3339 6742 3373
rect 7373 3276 7389 3311
rect 7677 3276 7703 3311
rect 8321 3276 8337 3311
rect 8625 3276 8651 3311
rect 9257 3276 9273 3311
rect 9561 3276 9587 3311
rect 10188 3276 10204 3311
rect 10492 3276 10518 3311
rect 11115 3276 11131 3311
rect 11419 3276 11445 3311
rect 5673 3237 5689 3271
rect 5821 3237 5837 3271
rect 6113 3237 6129 3271
rect 6261 3237 6277 3271
rect 6553 3237 6569 3271
rect 6701 3237 6717 3271
rect 246 3186 280 3202
rect 7150 3207 7184 3223
rect -24039 3114 -22837 3136
rect -24039 3068 -24001 3114
rect -22878 3068 -22837 3114
rect -24039 3045 -22837 3068
rect -20748 3114 -19546 3136
rect -20748 3068 -20710 3114
rect -19587 3068 -19546 3114
rect -20748 3045 -19546 3068
rect -17457 3114 -16255 3136
rect -17457 3068 -17419 3114
rect -16296 3068 -16255 3114
rect -17457 3045 -16255 3068
rect -14166 3114 -12964 3136
rect -14166 3068 -14128 3114
rect -13005 3068 -12964 3114
rect -14166 3045 -12964 3068
rect -10875 3114 -9673 3136
rect -10875 3068 -10837 3114
rect -9714 3068 -9673 3114
rect -10875 3045 -9673 3068
rect -7585 3114 -6383 3136
rect -7585 3068 -7547 3114
rect -6424 3068 -6383 3114
rect -7585 3045 -6383 3068
rect -4294 3114 -3092 3136
rect -4294 3068 -4256 3114
rect -3133 3068 -3092 3114
rect -4294 3045 -3092 3068
rect -1003 3114 199 3136
rect -1003 3068 -965 3114
rect 158 3068 199 3114
rect -1003 3045 199 3068
rect 7246 3207 7280 3223
rect 7150 2893 7184 2909
rect 7246 2893 7280 2904
rect 7342 3207 7376 3223
rect 7342 2893 7376 2909
rect 7438 3207 7472 3223
rect 7534 3207 7568 3223
rect 7438 2893 7472 2904
rect 7534 2893 7568 2909
rect 7630 3207 7664 3223
rect 7726 3207 7760 3223
rect 7630 2893 7664 2904
rect 7726 2893 7760 2909
rect 7822 3207 7856 3223
rect 7918 3207 7952 3223
rect 7822 2893 7856 2904
rect 7918 2893 7952 2909
rect 8098 3207 8132 3223
rect 8194 3207 8228 3223
rect 8098 2893 8132 2909
rect 8194 2893 8228 2904
rect 8290 3207 8324 3223
rect 8290 2893 8324 2909
rect 8386 3207 8420 3223
rect 8482 3207 8516 3223
rect 8386 2893 8420 2904
rect 8482 2893 8516 2909
rect 8578 3207 8612 3223
rect 8674 3207 8708 3223
rect 8578 2893 8612 2904
rect 8674 2893 8708 2909
rect 8770 3207 8804 3223
rect 8866 3207 8900 3223
rect 8770 2893 8804 2904
rect 8866 2893 8900 2909
rect 9034 3207 9068 3223
rect 9130 3207 9164 3223
rect 9034 2893 9068 2909
rect 9130 2893 9164 2904
rect 9226 3207 9260 3223
rect 9226 2893 9260 2909
rect 9322 3207 9356 3223
rect 9418 3207 9452 3223
rect 9322 2893 9356 2904
rect 9418 2893 9452 2909
rect 9514 3207 9548 3223
rect 9610 3207 9644 3223
rect 9514 2893 9548 2904
rect 9610 2893 9644 2909
rect 9706 3207 9740 3223
rect 9802 3207 9836 3223
rect 9706 2893 9740 2904
rect 9802 2893 9836 2909
rect 9965 3207 9999 3223
rect 10061 3207 10095 3223
rect 9965 2893 9999 2909
rect 10061 2893 10095 2904
rect 10157 3207 10191 3223
rect 10157 2893 10191 2909
rect 10253 3207 10287 3223
rect 10349 3207 10383 3223
rect 10253 2893 10287 2904
rect 10349 2893 10383 2909
rect 10445 3207 10479 3223
rect 10541 3207 10575 3223
rect 10445 2893 10479 2904
rect 10541 2893 10575 2909
rect 10637 3207 10671 3223
rect 10733 3207 10767 3223
rect 10637 2893 10671 2904
rect 10733 2893 10767 2909
rect 10892 3207 10926 3223
rect 10988 3207 11022 3223
rect 10892 2893 10926 2909
rect 10988 2893 11022 2904
rect 11084 3207 11118 3223
rect 11084 2893 11118 2909
rect 11180 3207 11214 3223
rect 11276 3207 11310 3223
rect 11180 2893 11214 2904
rect 11276 2893 11310 2909
rect 11372 3207 11406 3223
rect 11468 3207 11502 3223
rect 11372 2893 11406 2904
rect 11468 2893 11502 2909
rect 11564 3207 11598 3223
rect 11660 3207 11694 3223
rect 11564 2893 11598 2904
rect 11660 2893 11694 2909
rect 7182 2816 7198 2850
rect 7232 2816 7248 2850
rect 7374 2816 7390 2850
rect 7424 2816 7440 2850
rect 7566 2816 7582 2850
rect 7616 2816 7632 2850
rect 7758 2816 7774 2850
rect 7808 2816 7824 2850
rect 8130 2816 8146 2850
rect 8180 2816 8196 2850
rect 8322 2816 8338 2850
rect 8372 2816 8388 2850
rect 8514 2816 8530 2850
rect 8564 2816 8580 2850
rect 8706 2816 8722 2850
rect 8756 2816 8772 2850
rect 9066 2816 9082 2850
rect 9116 2816 9132 2850
rect 9258 2816 9274 2850
rect 9308 2816 9324 2850
rect 9450 2816 9466 2850
rect 9500 2816 9516 2850
rect 9642 2816 9658 2850
rect 9692 2816 9708 2850
rect 9997 2816 10013 2850
rect 10047 2816 10063 2850
rect 10189 2816 10205 2850
rect 10239 2816 10255 2850
rect 10381 2816 10397 2850
rect 10431 2816 10447 2850
rect 10573 2816 10589 2850
rect 10623 2816 10639 2850
rect 10924 2816 10940 2850
rect 10974 2816 10990 2850
rect 11116 2816 11132 2850
rect 11166 2816 11182 2850
rect 11308 2816 11324 2850
rect 11358 2816 11374 2850
rect 11500 2816 11516 2850
rect 11550 2816 11566 2850
rect -24716 2733 -23506 2761
rect -24716 2661 -24670 2733
rect -23548 2661 -23506 2733
rect -24716 2635 -23506 2661
rect -23157 2733 -21947 2761
rect -23157 2661 -23111 2733
rect -21989 2661 -21947 2733
rect -23157 2635 -21947 2661
rect -21425 2733 -20215 2761
rect -21425 2661 -21379 2733
rect -20257 2661 -20215 2733
rect -21425 2635 -20215 2661
rect -19866 2733 -18656 2761
rect -19866 2661 -19820 2733
rect -18698 2661 -18656 2733
rect -19866 2635 -18656 2661
rect -18134 2733 -16924 2761
rect -18134 2661 -18088 2733
rect -16966 2661 -16924 2733
rect -18134 2635 -16924 2661
rect -16575 2733 -15365 2761
rect -16575 2661 -16529 2733
rect -15407 2661 -15365 2733
rect -16575 2635 -15365 2661
rect -14843 2733 -13633 2761
rect -14843 2661 -14797 2733
rect -13675 2661 -13633 2733
rect -14843 2635 -13633 2661
rect -13284 2733 -12074 2761
rect -13284 2661 -13238 2733
rect -12116 2661 -12074 2733
rect -13284 2635 -12074 2661
rect -11552 2733 -10342 2761
rect -11552 2661 -11506 2733
rect -10384 2661 -10342 2733
rect -11552 2635 -10342 2661
rect -9993 2733 -8783 2761
rect -9993 2661 -9947 2733
rect -8825 2661 -8783 2733
rect -9993 2635 -8783 2661
rect -8262 2733 -7052 2761
rect -8262 2661 -8216 2733
rect -7094 2661 -7052 2733
rect -8262 2635 -7052 2661
rect -6703 2733 -5493 2761
rect -6703 2661 -6657 2733
rect -5535 2661 -5493 2733
rect -6703 2635 -5493 2661
rect -4971 2733 -3761 2761
rect -4971 2661 -4925 2733
rect -3803 2661 -3761 2733
rect -4971 2635 -3761 2661
rect -3412 2733 -2202 2761
rect -3412 2661 -3366 2733
rect -2244 2661 -2202 2733
rect -3412 2635 -2202 2661
rect -1680 2733 -470 2761
rect -1680 2661 -1634 2733
rect -512 2661 -470 2733
rect -1680 2635 -470 2661
rect -121 2733 1089 2761
rect -121 2661 -75 2733
rect 1047 2661 1089 2733
rect -121 2635 1089 2661
rect -24792 2564 -24758 2580
rect -24792 1977 -24758 2038
rect -24704 2564 -24670 2580
rect -24704 2022 -24670 2038
rect -24608 2564 -24574 2580
rect -24608 2022 -24574 2038
rect -24512 2564 -24478 2580
rect -24512 2022 -24478 2038
rect -24416 2564 -24382 2580
rect -24416 2022 -24382 2038
rect -24320 2564 -24286 2580
rect -24320 2022 -24286 2038
rect -24224 2564 -24190 2580
rect -24224 2022 -24190 2038
rect -24128 2564 -24094 2580
rect -24128 1995 -24094 2038
rect -24032 2564 -23998 2580
rect -24032 2022 -23998 2038
rect -23936 2564 -23902 2580
rect -23936 2022 -23902 2038
rect -23840 2564 -23806 2580
rect -23840 2022 -23806 2038
rect -23744 2564 -23710 2580
rect -23744 2022 -23710 2038
rect -23648 2564 -23614 2580
rect -23648 2022 -23614 2038
rect -23552 2564 -23518 2580
rect -23552 2022 -23518 2038
rect -23464 2564 -23430 2580
rect -24792 1967 -24190 1977
rect -24939 1938 -24854 1961
rect -24939 1828 -24921 1938
rect -24874 1828 -24854 1938
rect -24939 1808 -24854 1828
rect -24792 1922 -24336 1967
rect -24206 1922 -24190 1967
rect -24792 1908 -24190 1922
rect -24792 1524 -24758 1908
rect -24656 1837 -24435 1864
rect -24656 1784 -24606 1837
rect -24473 1784 -24435 1837
rect -24656 1646 -24435 1784
rect -24656 1601 -24611 1646
rect -24481 1601 -24435 1646
rect -24656 1574 -24435 1601
rect -24355 1638 -24190 1908
rect -24355 1593 -24328 1638
rect -24198 1593 -24190 1638
rect -24355 1576 -24190 1593
rect -24144 1695 -24078 1995
rect -23464 1980 -23430 2038
rect -24032 1962 -23430 1980
rect -24032 1917 -24005 1962
rect -23875 1917 -23430 1962
rect -24032 1903 -23430 1917
rect -23233 2564 -23199 2580
rect -23233 1977 -23199 2038
rect -23145 2564 -23111 2580
rect -23145 2022 -23111 2038
rect -23049 2564 -23015 2580
rect -23049 2022 -23015 2038
rect -22953 2564 -22919 2580
rect -22953 2022 -22919 2038
rect -22857 2564 -22823 2580
rect -22857 2022 -22823 2038
rect -22761 2564 -22727 2580
rect -22761 2022 -22727 2038
rect -22665 2564 -22631 2580
rect -22665 2022 -22631 2038
rect -22569 2564 -22535 2580
rect -22569 1995 -22535 2038
rect -22473 2564 -22439 2580
rect -22473 2022 -22439 2038
rect -22377 2564 -22343 2580
rect -22377 2022 -22343 2038
rect -22281 2564 -22247 2580
rect -22281 2022 -22247 2038
rect -22185 2564 -22151 2580
rect -22185 2022 -22151 2038
rect -22089 2564 -22055 2580
rect -22089 2022 -22055 2038
rect -21993 2564 -21959 2580
rect -21993 2022 -21959 2038
rect -21905 2564 -21871 2580
rect -23233 1967 -22631 1977
rect -23233 1922 -22777 1967
rect -22647 1922 -22631 1967
rect -23233 1908 -22631 1922
rect -24032 1845 -23855 1903
rect -24032 1792 -24000 1845
rect -23886 1792 -23855 1845
rect -24032 1763 -23855 1792
rect -23783 1844 -23668 1862
rect -23783 1776 -23766 1844
rect -23686 1776 -23668 1844
rect -23783 1756 -23668 1776
rect -24144 1673 -23504 1695
rect -24144 1618 -23584 1673
rect -23519 1618 -23504 1673
rect -24144 1599 -23504 1618
rect -24144 1565 -24078 1599
rect -24792 1402 -24758 1418
rect -24704 1524 -24670 1540
rect -24704 1402 -24670 1418
rect -24608 1539 -24574 1540
rect -24608 1402 -24574 1418
rect -24512 1524 -24478 1540
rect -24512 1402 -24478 1404
rect -24416 1539 -24382 1540
rect -24416 1402 -24382 1418
rect -24320 1524 -24286 1540
rect -24320 1402 -24286 1404
rect -24224 1538 -24190 1540
rect -24224 1402 -24190 1418
rect -24128 1524 -24094 1565
rect -24128 1402 -24094 1404
rect -24032 1539 -23998 1540
rect -24032 1402 -23998 1418
rect -23936 1524 -23902 1540
rect -23936 1402 -23902 1404
rect -23840 1539 -23806 1540
rect -23840 1402 -23806 1418
rect -23744 1524 -23710 1540
rect -23744 1402 -23710 1404
rect -23648 1539 -23614 1540
rect -23648 1402 -23614 1418
rect -23552 1524 -23518 1540
rect -23552 1402 -23518 1418
rect -23464 1524 -23430 1903
rect -23383 1893 -23274 1908
rect -23383 1753 -23364 1893
rect -23291 1753 -23274 1893
rect -23383 1736 -23274 1753
rect -23464 1402 -23430 1418
rect -23233 1524 -23199 1908
rect -23097 1837 -22876 1864
rect -23097 1784 -23047 1837
rect -22914 1784 -22876 1837
rect -23097 1646 -22876 1784
rect -23097 1601 -23052 1646
rect -22922 1601 -22876 1646
rect -23097 1574 -22876 1601
rect -22796 1638 -22631 1908
rect -22796 1593 -22769 1638
rect -22639 1593 -22631 1638
rect -22796 1576 -22631 1593
rect -22585 1695 -22519 1995
rect -21905 1980 -21871 2038
rect -22473 1962 -21871 1980
rect -22473 1917 -22446 1962
rect -22316 1917 -21871 1962
rect -21501 2564 -21467 2580
rect -21501 1977 -21467 2038
rect -21413 2564 -21379 2580
rect -21413 2022 -21379 2038
rect -21317 2564 -21283 2580
rect -21317 2022 -21283 2038
rect -21221 2564 -21187 2580
rect -21221 2022 -21187 2038
rect -21125 2564 -21091 2580
rect -21125 2022 -21091 2038
rect -21029 2564 -20995 2580
rect -21029 2022 -20995 2038
rect -20933 2564 -20899 2580
rect -20933 2022 -20899 2038
rect -20837 2564 -20803 2580
rect -20837 1995 -20803 2038
rect -20741 2564 -20707 2580
rect -20741 2022 -20707 2038
rect -20645 2564 -20611 2580
rect -20645 2022 -20611 2038
rect -20549 2564 -20515 2580
rect -20549 2022 -20515 2038
rect -20453 2564 -20419 2580
rect -20453 2022 -20419 2038
rect -20357 2564 -20323 2580
rect -20357 2022 -20323 2038
rect -20261 2564 -20227 2580
rect -20261 2022 -20227 2038
rect -20173 2564 -20139 2580
rect -21501 1967 -20899 1977
rect -22473 1903 -21871 1917
rect -22473 1845 -22296 1903
rect -22473 1792 -22441 1845
rect -22327 1792 -22296 1845
rect -22473 1763 -22296 1792
rect -22224 1844 -22109 1862
rect -22224 1776 -22207 1844
rect -22127 1776 -22109 1844
rect -22224 1756 -22109 1776
rect -22585 1673 -21945 1695
rect -22585 1618 -22025 1673
rect -21960 1618 -21945 1673
rect -22585 1599 -21945 1618
rect -22585 1565 -22519 1599
rect -23233 1402 -23199 1418
rect -23145 1524 -23111 1540
rect -23145 1402 -23111 1418
rect -23049 1539 -23015 1540
rect -23049 1402 -23015 1418
rect -22953 1524 -22919 1540
rect -22953 1402 -22919 1404
rect -22857 1539 -22823 1540
rect -22857 1402 -22823 1418
rect -22761 1524 -22727 1540
rect -22761 1402 -22727 1404
rect -22665 1538 -22631 1540
rect -22665 1402 -22631 1418
rect -22569 1524 -22535 1565
rect -22569 1402 -22535 1404
rect -22473 1539 -22439 1540
rect -22473 1402 -22439 1418
rect -22377 1524 -22343 1540
rect -22377 1402 -22343 1404
rect -22281 1539 -22247 1540
rect -22281 1402 -22247 1418
rect -22185 1524 -22151 1540
rect -22185 1402 -22151 1404
rect -22089 1539 -22055 1540
rect -22089 1402 -22055 1418
rect -21993 1524 -21959 1540
rect -21993 1402 -21959 1418
rect -21905 1524 -21871 1903
rect -21648 1938 -21563 1961
rect -21648 1828 -21630 1938
rect -21583 1828 -21563 1938
rect -21648 1808 -21563 1828
rect -21501 1922 -21045 1967
rect -20915 1922 -20899 1967
rect -21501 1908 -20899 1922
rect -21905 1402 -21871 1418
rect -21501 1524 -21467 1908
rect -21365 1837 -21144 1864
rect -21365 1784 -21315 1837
rect -21182 1784 -21144 1837
rect -21365 1646 -21144 1784
rect -21365 1601 -21320 1646
rect -21190 1601 -21144 1646
rect -21365 1574 -21144 1601
rect -21064 1638 -20899 1908
rect -21064 1593 -21037 1638
rect -20907 1593 -20899 1638
rect -21064 1576 -20899 1593
rect -20853 1695 -20787 1995
rect -20173 1980 -20139 2038
rect -20741 1962 -20139 1980
rect -20741 1917 -20714 1962
rect -20584 1917 -20139 1962
rect -20741 1903 -20139 1917
rect -19942 2564 -19908 2580
rect -19942 1977 -19908 2038
rect -19854 2564 -19820 2580
rect -19854 2022 -19820 2038
rect -19758 2564 -19724 2580
rect -19758 2022 -19724 2038
rect -19662 2564 -19628 2580
rect -19662 2022 -19628 2038
rect -19566 2564 -19532 2580
rect -19566 2022 -19532 2038
rect -19470 2564 -19436 2580
rect -19470 2022 -19436 2038
rect -19374 2564 -19340 2580
rect -19374 2022 -19340 2038
rect -19278 2564 -19244 2580
rect -19278 1995 -19244 2038
rect -19182 2564 -19148 2580
rect -19182 2022 -19148 2038
rect -19086 2564 -19052 2580
rect -19086 2022 -19052 2038
rect -18990 2564 -18956 2580
rect -18990 2022 -18956 2038
rect -18894 2564 -18860 2580
rect -18894 2022 -18860 2038
rect -18798 2564 -18764 2580
rect -18798 2022 -18764 2038
rect -18702 2564 -18668 2580
rect -18702 2022 -18668 2038
rect -18614 2564 -18580 2580
rect -19942 1967 -19340 1977
rect -19942 1922 -19486 1967
rect -19356 1922 -19340 1967
rect -19942 1908 -19340 1922
rect -20741 1845 -20564 1903
rect -20741 1792 -20709 1845
rect -20595 1792 -20564 1845
rect -20741 1763 -20564 1792
rect -20492 1844 -20377 1862
rect -20492 1776 -20475 1844
rect -20395 1776 -20377 1844
rect -20492 1756 -20377 1776
rect -20853 1673 -20213 1695
rect -20853 1618 -20293 1673
rect -20228 1618 -20213 1673
rect -20853 1599 -20213 1618
rect -20853 1565 -20787 1599
rect -21501 1402 -21467 1418
rect -21413 1524 -21379 1540
rect -21413 1402 -21379 1418
rect -21317 1539 -21283 1540
rect -21317 1402 -21283 1418
rect -21221 1524 -21187 1540
rect -21221 1402 -21187 1404
rect -21125 1539 -21091 1540
rect -21125 1402 -21091 1418
rect -21029 1524 -20995 1540
rect -21029 1402 -20995 1404
rect -20933 1538 -20899 1540
rect -20933 1402 -20899 1418
rect -20837 1524 -20803 1565
rect -20837 1402 -20803 1404
rect -20741 1539 -20707 1540
rect -20741 1402 -20707 1418
rect -20645 1524 -20611 1540
rect -20645 1402 -20611 1404
rect -20549 1539 -20515 1540
rect -20549 1402 -20515 1418
rect -20453 1524 -20419 1540
rect -20453 1402 -20419 1404
rect -20357 1539 -20323 1540
rect -20357 1402 -20323 1418
rect -20261 1524 -20227 1540
rect -20261 1402 -20227 1418
rect -20173 1524 -20139 1903
rect -20092 1893 -19983 1908
rect -20092 1753 -20073 1893
rect -20000 1753 -19983 1893
rect -20092 1736 -19983 1753
rect -20173 1402 -20139 1418
rect -19942 1524 -19908 1908
rect -19806 1837 -19585 1864
rect -19806 1784 -19756 1837
rect -19623 1784 -19585 1837
rect -19806 1646 -19585 1784
rect -19806 1601 -19761 1646
rect -19631 1601 -19585 1646
rect -19806 1574 -19585 1601
rect -19505 1638 -19340 1908
rect -19505 1593 -19478 1638
rect -19348 1593 -19340 1638
rect -19505 1576 -19340 1593
rect -19294 1695 -19228 1995
rect -18614 1980 -18580 2038
rect -19182 1962 -18580 1980
rect -19182 1917 -19155 1962
rect -19025 1917 -18580 1962
rect -18210 2564 -18176 2580
rect -18210 1977 -18176 2038
rect -18122 2564 -18088 2580
rect -18122 2022 -18088 2038
rect -18026 2564 -17992 2580
rect -18026 2022 -17992 2038
rect -17930 2564 -17896 2580
rect -17930 2022 -17896 2038
rect -17834 2564 -17800 2580
rect -17834 2022 -17800 2038
rect -17738 2564 -17704 2580
rect -17738 2022 -17704 2038
rect -17642 2564 -17608 2580
rect -17642 2022 -17608 2038
rect -17546 2564 -17512 2580
rect -17546 1995 -17512 2038
rect -17450 2564 -17416 2580
rect -17450 2022 -17416 2038
rect -17354 2564 -17320 2580
rect -17354 2022 -17320 2038
rect -17258 2564 -17224 2580
rect -17258 2022 -17224 2038
rect -17162 2564 -17128 2580
rect -17162 2022 -17128 2038
rect -17066 2564 -17032 2580
rect -17066 2022 -17032 2038
rect -16970 2564 -16936 2580
rect -16970 2022 -16936 2038
rect -16882 2564 -16848 2580
rect -18210 1967 -17608 1977
rect -19182 1903 -18580 1917
rect -19182 1845 -19005 1903
rect -19182 1792 -19150 1845
rect -19036 1792 -19005 1845
rect -19182 1763 -19005 1792
rect -18933 1844 -18818 1862
rect -18933 1776 -18916 1844
rect -18836 1776 -18818 1844
rect -18933 1756 -18818 1776
rect -19294 1673 -18654 1695
rect -19294 1618 -18734 1673
rect -18669 1618 -18654 1673
rect -19294 1599 -18654 1618
rect -19294 1565 -19228 1599
rect -19942 1402 -19908 1418
rect -19854 1524 -19820 1540
rect -19854 1402 -19820 1418
rect -19758 1539 -19724 1540
rect -19758 1402 -19724 1418
rect -19662 1524 -19628 1540
rect -19662 1402 -19628 1404
rect -19566 1539 -19532 1540
rect -19566 1402 -19532 1418
rect -19470 1524 -19436 1540
rect -19470 1402 -19436 1404
rect -19374 1538 -19340 1540
rect -19374 1402 -19340 1418
rect -19278 1524 -19244 1565
rect -19278 1402 -19244 1404
rect -19182 1539 -19148 1540
rect -19182 1402 -19148 1418
rect -19086 1524 -19052 1540
rect -19086 1402 -19052 1404
rect -18990 1539 -18956 1540
rect -18990 1402 -18956 1418
rect -18894 1524 -18860 1540
rect -18894 1402 -18860 1404
rect -18798 1539 -18764 1540
rect -18798 1402 -18764 1418
rect -18702 1524 -18668 1540
rect -18702 1402 -18668 1418
rect -18614 1524 -18580 1903
rect -18357 1938 -18272 1961
rect -18357 1828 -18339 1938
rect -18292 1828 -18272 1938
rect -18357 1808 -18272 1828
rect -18210 1922 -17754 1967
rect -17624 1922 -17608 1967
rect -18210 1908 -17608 1922
rect -18614 1402 -18580 1418
rect -18210 1524 -18176 1908
rect -18074 1837 -17853 1864
rect -18074 1784 -18024 1837
rect -17891 1784 -17853 1837
rect -18074 1646 -17853 1784
rect -18074 1601 -18029 1646
rect -17899 1601 -17853 1646
rect -18074 1574 -17853 1601
rect -17773 1638 -17608 1908
rect -17773 1593 -17746 1638
rect -17616 1593 -17608 1638
rect -17773 1576 -17608 1593
rect -17562 1695 -17496 1995
rect -16882 1980 -16848 2038
rect -17450 1962 -16848 1980
rect -17450 1917 -17423 1962
rect -17293 1917 -16848 1962
rect -17450 1903 -16848 1917
rect -16651 2564 -16617 2580
rect -16651 1977 -16617 2038
rect -16563 2564 -16529 2580
rect -16563 2022 -16529 2038
rect -16467 2564 -16433 2580
rect -16467 2022 -16433 2038
rect -16371 2564 -16337 2580
rect -16371 2022 -16337 2038
rect -16275 2564 -16241 2580
rect -16275 2022 -16241 2038
rect -16179 2564 -16145 2580
rect -16179 2022 -16145 2038
rect -16083 2564 -16049 2580
rect -16083 2022 -16049 2038
rect -15987 2564 -15953 2580
rect -15987 1995 -15953 2038
rect -15891 2564 -15857 2580
rect -15891 2022 -15857 2038
rect -15795 2564 -15761 2580
rect -15795 2022 -15761 2038
rect -15699 2564 -15665 2580
rect -15699 2022 -15665 2038
rect -15603 2564 -15569 2580
rect -15603 2022 -15569 2038
rect -15507 2564 -15473 2580
rect -15507 2022 -15473 2038
rect -15411 2564 -15377 2580
rect -15411 2022 -15377 2038
rect -15323 2564 -15289 2580
rect -16651 1967 -16049 1977
rect -16651 1922 -16195 1967
rect -16065 1922 -16049 1967
rect -16651 1908 -16049 1922
rect -17450 1845 -17273 1903
rect -17450 1792 -17418 1845
rect -17304 1792 -17273 1845
rect -17450 1763 -17273 1792
rect -17201 1844 -17086 1862
rect -17201 1776 -17184 1844
rect -17104 1776 -17086 1844
rect -17201 1756 -17086 1776
rect -17562 1673 -16922 1695
rect -17562 1618 -17002 1673
rect -16937 1618 -16922 1673
rect -17562 1599 -16922 1618
rect -17562 1565 -17496 1599
rect -18210 1402 -18176 1418
rect -18122 1524 -18088 1540
rect -18122 1402 -18088 1418
rect -18026 1539 -17992 1540
rect -18026 1402 -17992 1418
rect -17930 1524 -17896 1540
rect -17930 1402 -17896 1404
rect -17834 1539 -17800 1540
rect -17834 1402 -17800 1418
rect -17738 1524 -17704 1540
rect -17738 1402 -17704 1404
rect -17642 1538 -17608 1540
rect -17642 1402 -17608 1418
rect -17546 1524 -17512 1565
rect -17546 1402 -17512 1404
rect -17450 1539 -17416 1540
rect -17450 1402 -17416 1418
rect -17354 1524 -17320 1540
rect -17354 1402 -17320 1404
rect -17258 1539 -17224 1540
rect -17258 1402 -17224 1418
rect -17162 1524 -17128 1540
rect -17162 1402 -17128 1404
rect -17066 1539 -17032 1540
rect -17066 1402 -17032 1418
rect -16970 1524 -16936 1540
rect -16970 1402 -16936 1418
rect -16882 1524 -16848 1903
rect -16801 1893 -16692 1908
rect -16801 1753 -16782 1893
rect -16709 1753 -16692 1893
rect -16801 1736 -16692 1753
rect -16882 1402 -16848 1418
rect -16651 1524 -16617 1908
rect -16515 1837 -16294 1864
rect -16515 1784 -16465 1837
rect -16332 1784 -16294 1837
rect -16515 1646 -16294 1784
rect -16515 1601 -16470 1646
rect -16340 1601 -16294 1646
rect -16515 1574 -16294 1601
rect -16214 1638 -16049 1908
rect -16214 1593 -16187 1638
rect -16057 1593 -16049 1638
rect -16214 1576 -16049 1593
rect -16003 1695 -15937 1995
rect -15323 1980 -15289 2038
rect -15891 1962 -15289 1980
rect -15891 1917 -15864 1962
rect -15734 1917 -15289 1962
rect -14919 2564 -14885 2580
rect -14919 1977 -14885 2038
rect -14831 2564 -14797 2580
rect -14831 2022 -14797 2038
rect -14735 2564 -14701 2580
rect -14735 2022 -14701 2038
rect -14639 2564 -14605 2580
rect -14639 2022 -14605 2038
rect -14543 2564 -14509 2580
rect -14543 2022 -14509 2038
rect -14447 2564 -14413 2580
rect -14447 2022 -14413 2038
rect -14351 2564 -14317 2580
rect -14351 2022 -14317 2038
rect -14255 2564 -14221 2580
rect -14255 1995 -14221 2038
rect -14159 2564 -14125 2580
rect -14159 2022 -14125 2038
rect -14063 2564 -14029 2580
rect -14063 2022 -14029 2038
rect -13967 2564 -13933 2580
rect -13967 2022 -13933 2038
rect -13871 2564 -13837 2580
rect -13871 2022 -13837 2038
rect -13775 2564 -13741 2580
rect -13775 2022 -13741 2038
rect -13679 2564 -13645 2580
rect -13679 2022 -13645 2038
rect -13591 2564 -13557 2580
rect -14919 1967 -14317 1977
rect -15891 1903 -15289 1917
rect -15891 1845 -15714 1903
rect -15891 1792 -15859 1845
rect -15745 1792 -15714 1845
rect -15891 1763 -15714 1792
rect -15642 1844 -15527 1862
rect -15642 1776 -15625 1844
rect -15545 1776 -15527 1844
rect -15642 1756 -15527 1776
rect -16003 1673 -15363 1695
rect -16003 1618 -15443 1673
rect -15378 1618 -15363 1673
rect -16003 1599 -15363 1618
rect -16003 1565 -15937 1599
rect -16651 1402 -16617 1418
rect -16563 1524 -16529 1540
rect -16563 1402 -16529 1418
rect -16467 1539 -16433 1540
rect -16467 1402 -16433 1418
rect -16371 1524 -16337 1540
rect -16371 1402 -16337 1404
rect -16275 1539 -16241 1540
rect -16275 1402 -16241 1418
rect -16179 1524 -16145 1540
rect -16179 1402 -16145 1404
rect -16083 1538 -16049 1540
rect -16083 1402 -16049 1418
rect -15987 1524 -15953 1565
rect -15987 1402 -15953 1404
rect -15891 1539 -15857 1540
rect -15891 1402 -15857 1418
rect -15795 1524 -15761 1540
rect -15795 1402 -15761 1404
rect -15699 1539 -15665 1540
rect -15699 1402 -15665 1418
rect -15603 1524 -15569 1540
rect -15603 1402 -15569 1404
rect -15507 1539 -15473 1540
rect -15507 1402 -15473 1418
rect -15411 1524 -15377 1540
rect -15411 1402 -15377 1418
rect -15323 1524 -15289 1903
rect -15066 1938 -14981 1961
rect -15066 1828 -15048 1938
rect -15001 1828 -14981 1938
rect -15066 1808 -14981 1828
rect -14919 1922 -14463 1967
rect -14333 1922 -14317 1967
rect -14919 1908 -14317 1922
rect -15323 1402 -15289 1418
rect -14919 1524 -14885 1908
rect -14783 1837 -14562 1864
rect -14783 1784 -14733 1837
rect -14600 1784 -14562 1837
rect -14783 1646 -14562 1784
rect -14783 1601 -14738 1646
rect -14608 1601 -14562 1646
rect -14783 1574 -14562 1601
rect -14482 1638 -14317 1908
rect -14482 1593 -14455 1638
rect -14325 1593 -14317 1638
rect -14482 1576 -14317 1593
rect -14271 1695 -14205 1995
rect -13591 1980 -13557 2038
rect -14159 1962 -13557 1980
rect -14159 1917 -14132 1962
rect -14002 1917 -13557 1962
rect -14159 1903 -13557 1917
rect -13360 2564 -13326 2580
rect -13360 1977 -13326 2038
rect -13272 2564 -13238 2580
rect -13272 2022 -13238 2038
rect -13176 2564 -13142 2580
rect -13176 2022 -13142 2038
rect -13080 2564 -13046 2580
rect -13080 2022 -13046 2038
rect -12984 2564 -12950 2580
rect -12984 2022 -12950 2038
rect -12888 2564 -12854 2580
rect -12888 2022 -12854 2038
rect -12792 2564 -12758 2580
rect -12792 2022 -12758 2038
rect -12696 2564 -12662 2580
rect -12696 1995 -12662 2038
rect -12600 2564 -12566 2580
rect -12600 2022 -12566 2038
rect -12504 2564 -12470 2580
rect -12504 2022 -12470 2038
rect -12408 2564 -12374 2580
rect -12408 2022 -12374 2038
rect -12312 2564 -12278 2580
rect -12312 2022 -12278 2038
rect -12216 2564 -12182 2580
rect -12216 2022 -12182 2038
rect -12120 2564 -12086 2580
rect -12120 2022 -12086 2038
rect -12032 2564 -11998 2580
rect -13360 1967 -12758 1977
rect -13360 1922 -12904 1967
rect -12774 1922 -12758 1967
rect -13360 1908 -12758 1922
rect -14159 1845 -13982 1903
rect -14159 1792 -14127 1845
rect -14013 1792 -13982 1845
rect -14159 1763 -13982 1792
rect -13910 1844 -13795 1862
rect -13910 1776 -13893 1844
rect -13813 1776 -13795 1844
rect -13910 1756 -13795 1776
rect -14271 1673 -13631 1695
rect -14271 1618 -13711 1673
rect -13646 1618 -13631 1673
rect -14271 1599 -13631 1618
rect -14271 1565 -14205 1599
rect -14919 1402 -14885 1418
rect -14831 1524 -14797 1540
rect -14831 1402 -14797 1418
rect -14735 1539 -14701 1540
rect -14735 1402 -14701 1418
rect -14639 1524 -14605 1540
rect -14639 1402 -14605 1404
rect -14543 1539 -14509 1540
rect -14543 1402 -14509 1418
rect -14447 1524 -14413 1540
rect -14447 1402 -14413 1404
rect -14351 1538 -14317 1540
rect -14351 1402 -14317 1418
rect -14255 1524 -14221 1565
rect -14255 1402 -14221 1404
rect -14159 1539 -14125 1540
rect -14159 1402 -14125 1418
rect -14063 1524 -14029 1540
rect -14063 1402 -14029 1404
rect -13967 1539 -13933 1540
rect -13967 1402 -13933 1418
rect -13871 1524 -13837 1540
rect -13871 1402 -13837 1404
rect -13775 1539 -13741 1540
rect -13775 1402 -13741 1418
rect -13679 1524 -13645 1540
rect -13679 1402 -13645 1418
rect -13591 1524 -13557 1903
rect -13510 1893 -13401 1908
rect -13510 1753 -13491 1893
rect -13418 1753 -13401 1893
rect -13510 1736 -13401 1753
rect -13591 1402 -13557 1418
rect -13360 1524 -13326 1908
rect -13224 1837 -13003 1864
rect -13224 1784 -13174 1837
rect -13041 1784 -13003 1837
rect -13224 1646 -13003 1784
rect -13224 1601 -13179 1646
rect -13049 1601 -13003 1646
rect -13224 1574 -13003 1601
rect -12923 1638 -12758 1908
rect -12923 1593 -12896 1638
rect -12766 1593 -12758 1638
rect -12923 1576 -12758 1593
rect -12712 1695 -12646 1995
rect -12032 1980 -11998 2038
rect -12600 1962 -11998 1980
rect -12600 1917 -12573 1962
rect -12443 1917 -11998 1962
rect -11628 2564 -11594 2580
rect -11628 1977 -11594 2038
rect -11540 2564 -11506 2580
rect -11540 2022 -11506 2038
rect -11444 2564 -11410 2580
rect -11444 2022 -11410 2038
rect -11348 2564 -11314 2580
rect -11348 2022 -11314 2038
rect -11252 2564 -11218 2580
rect -11252 2022 -11218 2038
rect -11156 2564 -11122 2580
rect -11156 2022 -11122 2038
rect -11060 2564 -11026 2580
rect -11060 2022 -11026 2038
rect -10964 2564 -10930 2580
rect -10964 1995 -10930 2038
rect -10868 2564 -10834 2580
rect -10868 2022 -10834 2038
rect -10772 2564 -10738 2580
rect -10772 2022 -10738 2038
rect -10676 2564 -10642 2580
rect -10676 2022 -10642 2038
rect -10580 2564 -10546 2580
rect -10580 2022 -10546 2038
rect -10484 2564 -10450 2580
rect -10484 2022 -10450 2038
rect -10388 2564 -10354 2580
rect -10388 2022 -10354 2038
rect -10300 2564 -10266 2580
rect -11628 1967 -11026 1977
rect -12600 1903 -11998 1917
rect -12600 1845 -12423 1903
rect -12600 1792 -12568 1845
rect -12454 1792 -12423 1845
rect -12600 1763 -12423 1792
rect -12351 1844 -12236 1862
rect -12351 1776 -12334 1844
rect -12254 1776 -12236 1844
rect -12351 1756 -12236 1776
rect -12712 1673 -12072 1695
rect -12712 1618 -12152 1673
rect -12087 1618 -12072 1673
rect -12712 1599 -12072 1618
rect -12712 1565 -12646 1599
rect -13360 1402 -13326 1418
rect -13272 1524 -13238 1540
rect -13272 1402 -13238 1418
rect -13176 1539 -13142 1540
rect -13176 1402 -13142 1418
rect -13080 1524 -13046 1540
rect -13080 1402 -13046 1404
rect -12984 1539 -12950 1540
rect -12984 1402 -12950 1418
rect -12888 1524 -12854 1540
rect -12888 1402 -12854 1404
rect -12792 1538 -12758 1540
rect -12792 1402 -12758 1418
rect -12696 1524 -12662 1565
rect -12696 1402 -12662 1404
rect -12600 1539 -12566 1540
rect -12600 1402 -12566 1418
rect -12504 1524 -12470 1540
rect -12504 1402 -12470 1404
rect -12408 1539 -12374 1540
rect -12408 1402 -12374 1418
rect -12312 1524 -12278 1540
rect -12312 1402 -12278 1404
rect -12216 1539 -12182 1540
rect -12216 1402 -12182 1418
rect -12120 1524 -12086 1540
rect -12120 1402 -12086 1418
rect -12032 1524 -11998 1903
rect -11775 1938 -11690 1961
rect -11775 1828 -11757 1938
rect -11710 1828 -11690 1938
rect -11775 1808 -11690 1828
rect -11628 1922 -11172 1967
rect -11042 1922 -11026 1967
rect -11628 1908 -11026 1922
rect -12032 1402 -11998 1418
rect -11628 1524 -11594 1908
rect -11492 1837 -11271 1864
rect -11492 1784 -11442 1837
rect -11309 1784 -11271 1837
rect -11492 1646 -11271 1784
rect -11492 1601 -11447 1646
rect -11317 1601 -11271 1646
rect -11492 1574 -11271 1601
rect -11191 1638 -11026 1908
rect -11191 1593 -11164 1638
rect -11034 1593 -11026 1638
rect -11191 1576 -11026 1593
rect -10980 1695 -10914 1995
rect -10300 1980 -10266 2038
rect -10868 1962 -10266 1980
rect -10868 1917 -10841 1962
rect -10711 1917 -10266 1962
rect -10868 1903 -10266 1917
rect -10069 2564 -10035 2580
rect -10069 1977 -10035 2038
rect -9981 2564 -9947 2580
rect -9981 2022 -9947 2038
rect -9885 2564 -9851 2580
rect -9885 2022 -9851 2038
rect -9789 2564 -9755 2580
rect -9789 2022 -9755 2038
rect -9693 2564 -9659 2580
rect -9693 2022 -9659 2038
rect -9597 2564 -9563 2580
rect -9597 2022 -9563 2038
rect -9501 2564 -9467 2580
rect -9501 2022 -9467 2038
rect -9405 2564 -9371 2580
rect -9405 1995 -9371 2038
rect -9309 2564 -9275 2580
rect -9309 2022 -9275 2038
rect -9213 2564 -9179 2580
rect -9213 2022 -9179 2038
rect -9117 2564 -9083 2580
rect -9117 2022 -9083 2038
rect -9021 2564 -8987 2580
rect -9021 2022 -8987 2038
rect -8925 2564 -8891 2580
rect -8925 2022 -8891 2038
rect -8829 2564 -8795 2580
rect -8829 2022 -8795 2038
rect -8741 2564 -8707 2580
rect -10069 1967 -9467 1977
rect -10069 1922 -9613 1967
rect -9483 1922 -9467 1967
rect -10069 1908 -9467 1922
rect -10868 1845 -10691 1903
rect -10868 1792 -10836 1845
rect -10722 1792 -10691 1845
rect -10868 1763 -10691 1792
rect -10619 1844 -10504 1862
rect -10619 1776 -10602 1844
rect -10522 1776 -10504 1844
rect -10619 1756 -10504 1776
rect -10980 1673 -10340 1695
rect -10980 1618 -10420 1673
rect -10355 1618 -10340 1673
rect -10980 1599 -10340 1618
rect -10980 1565 -10914 1599
rect -11628 1402 -11594 1418
rect -11540 1524 -11506 1540
rect -11540 1402 -11506 1418
rect -11444 1539 -11410 1540
rect -11444 1402 -11410 1418
rect -11348 1524 -11314 1540
rect -11348 1402 -11314 1404
rect -11252 1539 -11218 1540
rect -11252 1402 -11218 1418
rect -11156 1524 -11122 1540
rect -11156 1402 -11122 1404
rect -11060 1538 -11026 1540
rect -11060 1402 -11026 1418
rect -10964 1524 -10930 1565
rect -10964 1402 -10930 1404
rect -10868 1539 -10834 1540
rect -10868 1402 -10834 1418
rect -10772 1524 -10738 1540
rect -10772 1402 -10738 1404
rect -10676 1539 -10642 1540
rect -10676 1402 -10642 1418
rect -10580 1524 -10546 1540
rect -10580 1402 -10546 1404
rect -10484 1539 -10450 1540
rect -10484 1402 -10450 1418
rect -10388 1524 -10354 1540
rect -10388 1402 -10354 1418
rect -10300 1524 -10266 1903
rect -10219 1893 -10110 1908
rect -10219 1753 -10200 1893
rect -10127 1753 -10110 1893
rect -10219 1736 -10110 1753
rect -10300 1402 -10266 1418
rect -10069 1524 -10035 1908
rect -9933 1837 -9712 1864
rect -9933 1784 -9883 1837
rect -9750 1784 -9712 1837
rect -9933 1646 -9712 1784
rect -9933 1601 -9888 1646
rect -9758 1601 -9712 1646
rect -9933 1574 -9712 1601
rect -9632 1638 -9467 1908
rect -9632 1593 -9605 1638
rect -9475 1593 -9467 1638
rect -9632 1576 -9467 1593
rect -9421 1695 -9355 1995
rect -8741 1980 -8707 2038
rect -9309 1962 -8707 1980
rect -9309 1917 -9282 1962
rect -9152 1917 -8707 1962
rect -8338 2564 -8304 2580
rect -8338 1977 -8304 2038
rect -8250 2564 -8216 2580
rect -8250 2022 -8216 2038
rect -8154 2564 -8120 2580
rect -8154 2022 -8120 2038
rect -8058 2564 -8024 2580
rect -8058 2022 -8024 2038
rect -7962 2564 -7928 2580
rect -7962 2022 -7928 2038
rect -7866 2564 -7832 2580
rect -7866 2022 -7832 2038
rect -7770 2564 -7736 2580
rect -7770 2022 -7736 2038
rect -7674 2564 -7640 2580
rect -7674 1995 -7640 2038
rect -7578 2564 -7544 2580
rect -7578 2022 -7544 2038
rect -7482 2564 -7448 2580
rect -7482 2022 -7448 2038
rect -7386 2564 -7352 2580
rect -7386 2022 -7352 2038
rect -7290 2564 -7256 2580
rect -7290 2022 -7256 2038
rect -7194 2564 -7160 2580
rect -7194 2022 -7160 2038
rect -7098 2564 -7064 2580
rect -7098 2022 -7064 2038
rect -7010 2564 -6976 2580
rect -8338 1967 -7736 1977
rect -9309 1903 -8707 1917
rect -9309 1845 -9132 1903
rect -9309 1792 -9277 1845
rect -9163 1792 -9132 1845
rect -9309 1763 -9132 1792
rect -9060 1844 -8945 1862
rect -9060 1776 -9043 1844
rect -8963 1776 -8945 1844
rect -9060 1756 -8945 1776
rect -9421 1673 -8781 1695
rect -9421 1618 -8861 1673
rect -8796 1618 -8781 1673
rect -9421 1599 -8781 1618
rect -9421 1565 -9355 1599
rect -10069 1402 -10035 1418
rect -9981 1524 -9947 1540
rect -9981 1402 -9947 1418
rect -9885 1539 -9851 1540
rect -9885 1402 -9851 1418
rect -9789 1524 -9755 1540
rect -9789 1402 -9755 1404
rect -9693 1539 -9659 1540
rect -9693 1402 -9659 1418
rect -9597 1524 -9563 1540
rect -9597 1402 -9563 1404
rect -9501 1538 -9467 1540
rect -9501 1402 -9467 1418
rect -9405 1524 -9371 1565
rect -9405 1402 -9371 1404
rect -9309 1539 -9275 1540
rect -9309 1402 -9275 1418
rect -9213 1524 -9179 1540
rect -9213 1402 -9179 1404
rect -9117 1539 -9083 1540
rect -9117 1402 -9083 1418
rect -9021 1524 -8987 1540
rect -9021 1402 -8987 1404
rect -8925 1539 -8891 1540
rect -8925 1402 -8891 1418
rect -8829 1524 -8795 1540
rect -8829 1402 -8795 1418
rect -8741 1524 -8707 1903
rect -8485 1938 -8400 1961
rect -8485 1828 -8467 1938
rect -8420 1828 -8400 1938
rect -8485 1808 -8400 1828
rect -8338 1922 -7882 1967
rect -7752 1922 -7736 1967
rect -8338 1908 -7736 1922
rect -8741 1402 -8707 1418
rect -8338 1524 -8304 1908
rect -8202 1837 -7981 1864
rect -8202 1784 -8152 1837
rect -8019 1784 -7981 1837
rect -8202 1646 -7981 1784
rect -8202 1601 -8157 1646
rect -8027 1601 -7981 1646
rect -8202 1574 -7981 1601
rect -7901 1638 -7736 1908
rect -7901 1593 -7874 1638
rect -7744 1593 -7736 1638
rect -7901 1576 -7736 1593
rect -7690 1695 -7624 1995
rect -7010 1980 -6976 2038
rect -7578 1962 -6976 1980
rect -7578 1917 -7551 1962
rect -7421 1917 -6976 1962
rect -7578 1903 -6976 1917
rect -6779 2564 -6745 2580
rect -6779 1977 -6745 2038
rect -6691 2564 -6657 2580
rect -6691 2022 -6657 2038
rect -6595 2564 -6561 2580
rect -6595 2022 -6561 2038
rect -6499 2564 -6465 2580
rect -6499 2022 -6465 2038
rect -6403 2564 -6369 2580
rect -6403 2022 -6369 2038
rect -6307 2564 -6273 2580
rect -6307 2022 -6273 2038
rect -6211 2564 -6177 2580
rect -6211 2022 -6177 2038
rect -6115 2564 -6081 2580
rect -6115 1995 -6081 2038
rect -6019 2564 -5985 2580
rect -6019 2022 -5985 2038
rect -5923 2564 -5889 2580
rect -5923 2022 -5889 2038
rect -5827 2564 -5793 2580
rect -5827 2022 -5793 2038
rect -5731 2564 -5697 2580
rect -5731 2022 -5697 2038
rect -5635 2564 -5601 2580
rect -5635 2022 -5601 2038
rect -5539 2564 -5505 2580
rect -5539 2022 -5505 2038
rect -5451 2564 -5417 2580
rect -6779 1967 -6177 1977
rect -6779 1922 -6323 1967
rect -6193 1922 -6177 1967
rect -6779 1908 -6177 1922
rect -7578 1845 -7401 1903
rect -7578 1792 -7546 1845
rect -7432 1792 -7401 1845
rect -7578 1763 -7401 1792
rect -7329 1844 -7214 1862
rect -7329 1776 -7312 1844
rect -7232 1776 -7214 1844
rect -7329 1756 -7214 1776
rect -7690 1673 -7050 1695
rect -7690 1618 -7130 1673
rect -7065 1618 -7050 1673
rect -7690 1599 -7050 1618
rect -7690 1565 -7624 1599
rect -8338 1402 -8304 1418
rect -8250 1524 -8216 1540
rect -8250 1402 -8216 1418
rect -8154 1539 -8120 1540
rect -8154 1402 -8120 1418
rect -8058 1524 -8024 1540
rect -8058 1402 -8024 1404
rect -7962 1539 -7928 1540
rect -7962 1402 -7928 1418
rect -7866 1524 -7832 1540
rect -7866 1402 -7832 1404
rect -7770 1538 -7736 1540
rect -7770 1402 -7736 1418
rect -7674 1524 -7640 1565
rect -7674 1402 -7640 1404
rect -7578 1539 -7544 1540
rect -7578 1402 -7544 1418
rect -7482 1524 -7448 1540
rect -7482 1402 -7448 1404
rect -7386 1539 -7352 1540
rect -7386 1402 -7352 1418
rect -7290 1524 -7256 1540
rect -7290 1402 -7256 1404
rect -7194 1539 -7160 1540
rect -7194 1402 -7160 1418
rect -7098 1524 -7064 1540
rect -7098 1402 -7064 1418
rect -7010 1524 -6976 1903
rect -6929 1893 -6820 1908
rect -6929 1753 -6910 1893
rect -6837 1753 -6820 1893
rect -6929 1736 -6820 1753
rect -7010 1402 -6976 1418
rect -6779 1524 -6745 1908
rect -6643 1837 -6422 1864
rect -6643 1784 -6593 1837
rect -6460 1784 -6422 1837
rect -6643 1646 -6422 1784
rect -6643 1601 -6598 1646
rect -6468 1601 -6422 1646
rect -6643 1574 -6422 1601
rect -6342 1638 -6177 1908
rect -6342 1593 -6315 1638
rect -6185 1593 -6177 1638
rect -6342 1576 -6177 1593
rect -6131 1695 -6065 1995
rect -5451 1980 -5417 2038
rect -6019 1962 -5417 1980
rect -6019 1917 -5992 1962
rect -5862 1917 -5417 1962
rect -5047 2564 -5013 2580
rect -5047 1977 -5013 2038
rect -4959 2564 -4925 2580
rect -4959 2022 -4925 2038
rect -4863 2564 -4829 2580
rect -4863 2022 -4829 2038
rect -4767 2564 -4733 2580
rect -4767 2022 -4733 2038
rect -4671 2564 -4637 2580
rect -4671 2022 -4637 2038
rect -4575 2564 -4541 2580
rect -4575 2022 -4541 2038
rect -4479 2564 -4445 2580
rect -4479 2022 -4445 2038
rect -4383 2564 -4349 2580
rect -4383 1995 -4349 2038
rect -4287 2564 -4253 2580
rect -4287 2022 -4253 2038
rect -4191 2564 -4157 2580
rect -4191 2022 -4157 2038
rect -4095 2564 -4061 2580
rect -4095 2022 -4061 2038
rect -3999 2564 -3965 2580
rect -3999 2022 -3965 2038
rect -3903 2564 -3869 2580
rect -3903 2022 -3869 2038
rect -3807 2564 -3773 2580
rect -3807 2022 -3773 2038
rect -3719 2564 -3685 2580
rect -5047 1967 -4445 1977
rect -6019 1903 -5417 1917
rect -6019 1845 -5842 1903
rect -6019 1792 -5987 1845
rect -5873 1792 -5842 1845
rect -6019 1763 -5842 1792
rect -5770 1844 -5655 1862
rect -5770 1776 -5753 1844
rect -5673 1776 -5655 1844
rect -5770 1756 -5655 1776
rect -6131 1673 -5491 1695
rect -6131 1618 -5571 1673
rect -5506 1618 -5491 1673
rect -6131 1599 -5491 1618
rect -6131 1565 -6065 1599
rect -6779 1402 -6745 1418
rect -6691 1524 -6657 1540
rect -6691 1402 -6657 1418
rect -6595 1539 -6561 1540
rect -6595 1402 -6561 1418
rect -6499 1524 -6465 1540
rect -6499 1402 -6465 1404
rect -6403 1539 -6369 1540
rect -6403 1402 -6369 1418
rect -6307 1524 -6273 1540
rect -6307 1402 -6273 1404
rect -6211 1538 -6177 1540
rect -6211 1402 -6177 1418
rect -6115 1524 -6081 1565
rect -6115 1402 -6081 1404
rect -6019 1539 -5985 1540
rect -6019 1402 -5985 1418
rect -5923 1524 -5889 1540
rect -5923 1402 -5889 1404
rect -5827 1539 -5793 1540
rect -5827 1402 -5793 1418
rect -5731 1524 -5697 1540
rect -5731 1402 -5697 1404
rect -5635 1539 -5601 1540
rect -5635 1402 -5601 1418
rect -5539 1524 -5505 1540
rect -5539 1402 -5505 1418
rect -5451 1524 -5417 1903
rect -5194 1938 -5109 1961
rect -5194 1828 -5176 1938
rect -5129 1828 -5109 1938
rect -5194 1808 -5109 1828
rect -5047 1922 -4591 1967
rect -4461 1922 -4445 1967
rect -5047 1908 -4445 1922
rect -5451 1402 -5417 1418
rect -5047 1524 -5013 1908
rect -4911 1837 -4690 1864
rect -4911 1784 -4861 1837
rect -4728 1784 -4690 1837
rect -4911 1646 -4690 1784
rect -4911 1601 -4866 1646
rect -4736 1601 -4690 1646
rect -4911 1574 -4690 1601
rect -4610 1638 -4445 1908
rect -4610 1593 -4583 1638
rect -4453 1593 -4445 1638
rect -4610 1576 -4445 1593
rect -4399 1695 -4333 1995
rect -3719 1980 -3685 2038
rect -4287 1962 -3685 1980
rect -4287 1917 -4260 1962
rect -4130 1917 -3685 1962
rect -4287 1903 -3685 1917
rect -3488 2564 -3454 2580
rect -3488 1977 -3454 2038
rect -3400 2564 -3366 2580
rect -3400 2022 -3366 2038
rect -3304 2564 -3270 2580
rect -3304 2022 -3270 2038
rect -3208 2564 -3174 2580
rect -3208 2022 -3174 2038
rect -3112 2564 -3078 2580
rect -3112 2022 -3078 2038
rect -3016 2564 -2982 2580
rect -3016 2022 -2982 2038
rect -2920 2564 -2886 2580
rect -2920 2022 -2886 2038
rect -2824 2564 -2790 2580
rect -2824 1995 -2790 2038
rect -2728 2564 -2694 2580
rect -2728 2022 -2694 2038
rect -2632 2564 -2598 2580
rect -2632 2022 -2598 2038
rect -2536 2564 -2502 2580
rect -2536 2022 -2502 2038
rect -2440 2564 -2406 2580
rect -2440 2022 -2406 2038
rect -2344 2564 -2310 2580
rect -2344 2022 -2310 2038
rect -2248 2564 -2214 2580
rect -2248 2022 -2214 2038
rect -2160 2564 -2126 2580
rect -3488 1967 -2886 1977
rect -3488 1922 -3032 1967
rect -2902 1922 -2886 1967
rect -3488 1908 -2886 1922
rect -4287 1845 -4110 1903
rect -4287 1792 -4255 1845
rect -4141 1792 -4110 1845
rect -4287 1763 -4110 1792
rect -4038 1844 -3923 1862
rect -4038 1776 -4021 1844
rect -3941 1776 -3923 1844
rect -4038 1756 -3923 1776
rect -4399 1673 -3759 1695
rect -4399 1618 -3839 1673
rect -3774 1618 -3759 1673
rect -4399 1599 -3759 1618
rect -4399 1565 -4333 1599
rect -5047 1402 -5013 1418
rect -4959 1524 -4925 1540
rect -4959 1402 -4925 1418
rect -4863 1539 -4829 1540
rect -4863 1402 -4829 1418
rect -4767 1524 -4733 1540
rect -4767 1402 -4733 1404
rect -4671 1539 -4637 1540
rect -4671 1402 -4637 1418
rect -4575 1524 -4541 1540
rect -4575 1402 -4541 1404
rect -4479 1538 -4445 1540
rect -4479 1402 -4445 1418
rect -4383 1524 -4349 1565
rect -4383 1402 -4349 1404
rect -4287 1539 -4253 1540
rect -4287 1402 -4253 1418
rect -4191 1524 -4157 1540
rect -4191 1402 -4157 1404
rect -4095 1539 -4061 1540
rect -4095 1402 -4061 1418
rect -3999 1524 -3965 1540
rect -3999 1402 -3965 1404
rect -3903 1539 -3869 1540
rect -3903 1402 -3869 1418
rect -3807 1524 -3773 1540
rect -3807 1402 -3773 1418
rect -3719 1524 -3685 1903
rect -3638 1893 -3529 1908
rect -3638 1753 -3619 1893
rect -3546 1753 -3529 1893
rect -3638 1736 -3529 1753
rect -3719 1402 -3685 1418
rect -3488 1524 -3454 1908
rect -3352 1837 -3131 1864
rect -3352 1784 -3302 1837
rect -3169 1784 -3131 1837
rect -3352 1646 -3131 1784
rect -3352 1601 -3307 1646
rect -3177 1601 -3131 1646
rect -3352 1574 -3131 1601
rect -3051 1638 -2886 1908
rect -3051 1593 -3024 1638
rect -2894 1593 -2886 1638
rect -3051 1576 -2886 1593
rect -2840 1695 -2774 1995
rect -2160 1980 -2126 2038
rect -2728 1962 -2126 1980
rect -2728 1917 -2701 1962
rect -2571 1917 -2126 1962
rect -1756 2564 -1722 2580
rect -1756 1977 -1722 2038
rect -1668 2564 -1634 2580
rect -1668 2022 -1634 2038
rect -1572 2564 -1538 2580
rect -1572 2022 -1538 2038
rect -1476 2564 -1442 2580
rect -1476 2022 -1442 2038
rect -1380 2564 -1346 2580
rect -1380 2022 -1346 2038
rect -1284 2564 -1250 2580
rect -1284 2022 -1250 2038
rect -1188 2564 -1154 2580
rect -1188 2022 -1154 2038
rect -1092 2564 -1058 2580
rect -1092 1995 -1058 2038
rect -996 2564 -962 2580
rect -996 2022 -962 2038
rect -900 2564 -866 2580
rect -900 2022 -866 2038
rect -804 2564 -770 2580
rect -804 2022 -770 2038
rect -708 2564 -674 2580
rect -708 2022 -674 2038
rect -612 2564 -578 2580
rect -612 2022 -578 2038
rect -516 2564 -482 2580
rect -516 2022 -482 2038
rect -428 2564 -394 2580
rect -1756 1967 -1154 1977
rect -2728 1903 -2126 1917
rect -2728 1845 -2551 1903
rect -2728 1792 -2696 1845
rect -2582 1792 -2551 1845
rect -2728 1763 -2551 1792
rect -2479 1844 -2364 1862
rect -2479 1776 -2462 1844
rect -2382 1776 -2364 1844
rect -2479 1756 -2364 1776
rect -2840 1673 -2200 1695
rect -2840 1618 -2280 1673
rect -2215 1618 -2200 1673
rect -2840 1599 -2200 1618
rect -2840 1565 -2774 1599
rect -3488 1402 -3454 1418
rect -3400 1524 -3366 1540
rect -3400 1402 -3366 1418
rect -3304 1539 -3270 1540
rect -3304 1402 -3270 1418
rect -3208 1524 -3174 1540
rect -3208 1402 -3174 1404
rect -3112 1539 -3078 1540
rect -3112 1402 -3078 1418
rect -3016 1524 -2982 1540
rect -3016 1402 -2982 1404
rect -2920 1538 -2886 1540
rect -2920 1402 -2886 1418
rect -2824 1524 -2790 1565
rect -2824 1402 -2790 1404
rect -2728 1539 -2694 1540
rect -2728 1402 -2694 1418
rect -2632 1524 -2598 1540
rect -2632 1402 -2598 1404
rect -2536 1539 -2502 1540
rect -2536 1402 -2502 1418
rect -2440 1524 -2406 1540
rect -2440 1402 -2406 1404
rect -2344 1539 -2310 1540
rect -2344 1402 -2310 1418
rect -2248 1524 -2214 1540
rect -2248 1402 -2214 1418
rect -2160 1524 -2126 1903
rect -1903 1938 -1818 1961
rect -1903 1828 -1885 1938
rect -1838 1828 -1818 1938
rect -1903 1808 -1818 1828
rect -1756 1922 -1300 1967
rect -1170 1922 -1154 1967
rect -1756 1908 -1154 1922
rect -2160 1402 -2126 1418
rect -1756 1524 -1722 1908
rect -1620 1837 -1399 1864
rect -1620 1784 -1570 1837
rect -1437 1784 -1399 1837
rect -1620 1646 -1399 1784
rect -1620 1601 -1575 1646
rect -1445 1601 -1399 1646
rect -1620 1574 -1399 1601
rect -1319 1638 -1154 1908
rect -1319 1593 -1292 1638
rect -1162 1593 -1154 1638
rect -1319 1576 -1154 1593
rect -1108 1695 -1042 1995
rect -428 1980 -394 2038
rect -996 1962 -394 1980
rect -996 1917 -969 1962
rect -839 1917 -394 1962
rect -996 1903 -394 1917
rect -197 2564 -163 2580
rect -197 1977 -163 2038
rect -109 2564 -75 2580
rect -109 2022 -75 2038
rect -13 2564 21 2580
rect -13 2022 21 2038
rect 83 2564 117 2580
rect 83 2022 117 2038
rect 179 2564 213 2580
rect 179 2022 213 2038
rect 275 2564 309 2580
rect 275 2022 309 2038
rect 371 2564 405 2580
rect 371 2022 405 2038
rect 467 2564 501 2580
rect 467 1995 501 2038
rect 563 2564 597 2580
rect 563 2022 597 2038
rect 659 2564 693 2580
rect 659 2022 693 2038
rect 755 2564 789 2580
rect 755 2022 789 2038
rect 851 2564 885 2580
rect 851 2022 885 2038
rect 947 2564 981 2580
rect 947 2022 981 2038
rect 1043 2564 1077 2580
rect 1043 2022 1077 2038
rect 1131 2564 1165 2580
rect -197 1967 405 1977
rect -197 1922 259 1967
rect 389 1922 405 1967
rect -197 1908 405 1922
rect -996 1845 -819 1903
rect -996 1792 -964 1845
rect -850 1792 -819 1845
rect -996 1763 -819 1792
rect -747 1844 -632 1862
rect -747 1776 -730 1844
rect -650 1776 -632 1844
rect -747 1756 -632 1776
rect -1108 1673 -468 1695
rect -1108 1618 -548 1673
rect -483 1618 -468 1673
rect -1108 1599 -468 1618
rect -1108 1565 -1042 1599
rect -1756 1402 -1722 1418
rect -1668 1524 -1634 1540
rect -1668 1402 -1634 1418
rect -1572 1539 -1538 1540
rect -1572 1402 -1538 1418
rect -1476 1524 -1442 1540
rect -1476 1402 -1442 1404
rect -1380 1539 -1346 1540
rect -1380 1402 -1346 1418
rect -1284 1524 -1250 1540
rect -1284 1402 -1250 1404
rect -1188 1538 -1154 1540
rect -1188 1402 -1154 1418
rect -1092 1524 -1058 1565
rect -1092 1402 -1058 1404
rect -996 1539 -962 1540
rect -996 1402 -962 1418
rect -900 1524 -866 1540
rect -900 1402 -866 1404
rect -804 1539 -770 1540
rect -804 1402 -770 1418
rect -708 1524 -674 1540
rect -708 1402 -674 1404
rect -612 1539 -578 1540
rect -612 1402 -578 1418
rect -516 1524 -482 1540
rect -516 1402 -482 1418
rect -428 1524 -394 1903
rect -347 1893 -238 1908
rect -347 1753 -328 1893
rect -255 1753 -238 1893
rect -347 1736 -238 1753
rect -428 1402 -394 1418
rect -197 1524 -163 1908
rect -61 1837 160 1864
rect -61 1784 -11 1837
rect 122 1784 160 1837
rect -61 1646 160 1784
rect -61 1601 -16 1646
rect 114 1601 160 1646
rect -61 1574 160 1601
rect 240 1638 405 1908
rect 240 1593 267 1638
rect 397 1593 405 1638
rect 240 1576 405 1593
rect 451 1695 517 1995
rect 1131 1980 1165 2038
rect 563 1962 1165 1980
rect 563 1917 590 1962
rect 720 1917 1165 1962
rect 563 1903 1165 1917
rect 563 1845 740 1903
rect 563 1792 595 1845
rect 709 1792 740 1845
rect 563 1763 740 1792
rect 812 1844 927 1862
rect 812 1776 829 1844
rect 909 1776 927 1844
rect 812 1756 927 1776
rect 451 1673 1091 1695
rect 451 1618 1011 1673
rect 1076 1618 1091 1673
rect 451 1599 1091 1618
rect 451 1565 517 1599
rect -197 1402 -163 1418
rect -109 1524 -75 1540
rect -109 1402 -75 1418
rect -13 1539 21 1540
rect -13 1402 21 1418
rect 83 1524 117 1540
rect 83 1402 117 1404
rect 179 1539 213 1540
rect 179 1402 213 1418
rect 275 1524 309 1540
rect 275 1402 309 1404
rect 371 1538 405 1540
rect 371 1402 405 1418
rect 467 1524 501 1565
rect 467 1402 501 1404
rect 563 1539 597 1540
rect 563 1402 597 1418
rect 659 1524 693 1540
rect 659 1402 693 1404
rect 755 1539 789 1540
rect 755 1402 789 1418
rect 851 1524 885 1540
rect 851 1402 885 1404
rect 947 1539 981 1540
rect 947 1402 981 1418
rect 1043 1524 1077 1540
rect 1043 1402 1077 1418
rect 1131 1524 1165 1903
rect 7298 2494 7403 2497
rect 8246 2494 8351 2497
rect 9182 2494 9287 2497
rect 10113 2494 10218 2497
rect 11040 2494 11145 2497
rect 7298 2478 7406 2494
rect 7298 2466 7372 2478
rect 7333 1715 7372 2466
rect 7298 1702 7372 1715
rect 7298 1686 7406 1702
rect 7756 2478 7790 2494
rect 7756 1686 7790 1702
rect 8246 2478 8354 2494
rect 8246 2466 8320 2478
rect 8281 1715 8320 2466
rect 8246 1702 8320 1715
rect 8246 1686 8354 1702
rect 8704 2478 8738 2494
rect 8704 1686 8738 1702
rect 9182 2478 9290 2494
rect 9182 2466 9256 2478
rect 9217 1715 9256 2466
rect 9182 1702 9256 1715
rect 9182 1686 9290 1702
rect 9640 2478 9674 2494
rect 9640 1686 9674 1702
rect 10113 2478 10221 2494
rect 10113 2466 10187 2478
rect 10148 1715 10187 2466
rect 10113 1702 10187 1715
rect 10113 1686 10221 1702
rect 10571 2478 10605 2494
rect 10571 1686 10605 1702
rect 11040 2478 11148 2494
rect 11040 2466 11114 2478
rect 11075 1715 11114 2466
rect 11040 1702 11114 1715
rect 11040 1686 11148 1702
rect 11498 2478 11532 2494
rect 11783 2152 12203 2172
rect 11783 2101 11811 2152
rect 12168 2101 12203 2152
rect 11783 2082 12203 2101
rect 11785 1997 11819 2082
rect 11785 1749 11819 1765
rect 11881 1997 11915 2013
rect 11881 1749 11915 1765
rect 11977 1997 12011 2082
rect 11977 1749 12011 1765
rect 12073 1997 12107 2013
rect 12073 1749 12107 1765
rect 12169 1997 12203 2082
rect 12169 1749 12203 1765
rect 12265 1997 12299 2013
rect 12265 1749 12299 1765
rect 12361 1997 12395 2013
rect 12361 1749 12395 1765
rect 12457 1997 12491 2013
rect 12457 1749 12491 1765
rect 12553 1997 12587 2013
rect 12553 1749 12587 1765
rect 12649 1997 12683 2013
rect 12649 1749 12683 1765
rect 12745 1997 12779 2013
rect 12970 1931 12986 1965
rect 13077 1931 13093 1965
rect 12745 1749 12779 1765
rect 12826 1845 12876 1862
rect 12919 1859 12929 1893
rect 13125 1859 13141 1893
rect 11498 1686 11532 1702
rect 12154 1669 12170 1703
rect 12204 1669 12220 1703
rect 12826 1619 12842 1845
rect 12919 1763 12935 1797
rect 13129 1763 13147 1797
rect 12919 1667 12929 1701
rect 13125 1667 13141 1701
rect 1131 1402 1165 1418
rect 7298 1550 7406 1566
rect 7298 1537 7372 1550
rect -24711 1330 -23509 1352
rect -24711 1284 -24670 1330
rect -23547 1284 -23509 1330
rect -24711 1261 -23509 1284
rect -23152 1330 -21950 1352
rect -23152 1284 -23111 1330
rect -21988 1284 -21950 1330
rect -23152 1261 -21950 1284
rect -21420 1330 -20218 1352
rect -21420 1284 -21379 1330
rect -20256 1284 -20218 1330
rect -21420 1261 -20218 1284
rect -19861 1330 -18659 1352
rect -19861 1284 -19820 1330
rect -18697 1284 -18659 1330
rect -19861 1261 -18659 1284
rect -18129 1330 -16927 1352
rect -18129 1284 -18088 1330
rect -16965 1284 -16927 1330
rect -18129 1261 -16927 1284
rect -16570 1330 -15368 1352
rect -16570 1284 -16529 1330
rect -15406 1284 -15368 1330
rect -16570 1261 -15368 1284
rect -14838 1330 -13636 1352
rect -14838 1284 -14797 1330
rect -13674 1284 -13636 1330
rect -14838 1261 -13636 1284
rect -13279 1330 -12077 1352
rect -13279 1284 -13238 1330
rect -12115 1284 -12077 1330
rect -13279 1261 -12077 1284
rect -11547 1330 -10345 1352
rect -11547 1284 -11506 1330
rect -10383 1284 -10345 1330
rect -11547 1261 -10345 1284
rect -9988 1330 -8786 1352
rect -9988 1284 -9947 1330
rect -8824 1284 -8786 1330
rect -9988 1261 -8786 1284
rect -8257 1330 -7055 1352
rect -8257 1284 -8216 1330
rect -7093 1284 -7055 1330
rect -8257 1261 -7055 1284
rect -6698 1330 -5496 1352
rect -6698 1284 -6657 1330
rect -5534 1284 -5496 1330
rect -6698 1261 -5496 1284
rect -4966 1330 -3764 1352
rect -4966 1284 -4925 1330
rect -3802 1284 -3764 1330
rect -4966 1261 -3764 1284
rect -3407 1330 -2205 1352
rect -3407 1284 -3366 1330
rect -2243 1284 -2205 1330
rect -3407 1261 -2205 1284
rect -1675 1330 -473 1352
rect -1675 1284 -1634 1330
rect -511 1284 -473 1330
rect -1675 1261 -473 1284
rect -116 1330 1086 1352
rect -116 1284 -75 1330
rect 1048 1284 1086 1330
rect -116 1261 1086 1284
rect -24585 941 -24569 988
rect -24000 941 -23976 988
rect -23476 941 -23460 988
rect -22891 941 -22867 988
rect -22594 941 -22578 988
rect -22009 941 -21985 988
rect -21294 941 -21278 988
rect -20709 941 -20685 988
rect -20185 941 -20169 988
rect -19600 941 -19576 988
rect -19303 941 -19287 988
rect -18718 941 -18694 988
rect -18003 941 -17987 988
rect -17418 941 -17394 988
rect -16894 941 -16878 988
rect -16309 941 -16285 988
rect -16012 941 -15996 988
rect -15427 941 -15403 988
rect -14712 941 -14696 988
rect -14127 941 -14103 988
rect -13603 941 -13587 988
rect -13018 941 -12994 988
rect -12721 941 -12705 988
rect -12136 941 -12112 988
rect -11421 941 -11405 988
rect -10836 941 -10812 988
rect -10312 941 -10296 988
rect -9727 941 -9703 988
rect -9430 941 -9414 988
rect -8845 941 -8821 988
rect -8131 941 -8115 988
rect -7546 941 -7522 988
rect -7022 941 -7006 988
rect -6437 941 -6413 988
rect -6140 941 -6124 988
rect -5555 941 -5531 988
rect -4840 941 -4824 988
rect -4255 941 -4231 988
rect -3731 941 -3715 988
rect -3146 941 -3122 988
rect -2849 941 -2833 988
rect -2264 941 -2240 988
rect -1549 941 -1533 988
rect -964 941 -940 988
rect -440 941 -424 988
rect 145 941 169 988
rect 442 941 458 988
rect 1027 941 1051 988
rect -24585 869 -24551 879
rect -24585 657 -24551 673
rect -24489 863 -24455 879
rect -24489 657 -24455 667
rect -24393 869 -24359 879
rect -24393 657 -24359 673
rect -24297 863 -24263 879
rect -24297 657 -24263 667
rect -24201 869 -24167 879
rect -24201 657 -24167 673
rect -24105 863 -24071 879
rect -24105 657 -24071 667
rect -24009 869 -23975 879
rect -24009 657 -23975 673
rect -23476 869 -23442 879
rect -23476 657 -23442 673
rect -23380 863 -23346 879
rect -23380 657 -23346 667
rect -23284 869 -23250 879
rect -23284 657 -23250 673
rect -23188 863 -23154 879
rect -23188 657 -23154 667
rect -23092 869 -23058 879
rect -23092 657 -23058 673
rect -22996 863 -22962 879
rect -22996 657 -22962 667
rect -22900 869 -22866 879
rect -22900 657 -22866 673
rect -22594 869 -22560 879
rect -22594 657 -22560 673
rect -22498 863 -22464 879
rect -22498 657 -22464 667
rect -22402 869 -22368 879
rect -22402 657 -22368 673
rect -22306 863 -22272 879
rect -22306 657 -22272 667
rect -22210 869 -22176 879
rect -22210 657 -22176 673
rect -22114 863 -22080 879
rect -22114 657 -22080 667
rect -22018 869 -21984 879
rect -22018 657 -21984 673
rect -21294 869 -21260 879
rect -21294 657 -21260 673
rect -21198 863 -21164 879
rect -21198 657 -21164 667
rect -21102 869 -21068 879
rect -21102 657 -21068 673
rect -21006 863 -20972 879
rect -21006 657 -20972 667
rect -20910 869 -20876 879
rect -20910 657 -20876 673
rect -20814 863 -20780 879
rect -20814 657 -20780 667
rect -20718 869 -20684 879
rect -20718 657 -20684 673
rect -20185 869 -20151 879
rect -20185 657 -20151 673
rect -20089 863 -20055 879
rect -20089 657 -20055 667
rect -19993 869 -19959 879
rect -19993 657 -19959 673
rect -19897 863 -19863 879
rect -19897 657 -19863 667
rect -19801 869 -19767 879
rect -19801 657 -19767 673
rect -19705 863 -19671 879
rect -19705 657 -19671 667
rect -19609 869 -19575 879
rect -19609 657 -19575 673
rect -19303 869 -19269 879
rect -19303 657 -19269 673
rect -19207 863 -19173 879
rect -19207 657 -19173 667
rect -19111 869 -19077 879
rect -19111 657 -19077 673
rect -19015 863 -18981 879
rect -19015 657 -18981 667
rect -18919 869 -18885 879
rect -18919 657 -18885 673
rect -18823 863 -18789 879
rect -18823 657 -18789 667
rect -18727 869 -18693 879
rect -18727 657 -18693 673
rect -18003 869 -17969 879
rect -18003 657 -17969 673
rect -17907 863 -17873 879
rect -17907 657 -17873 667
rect -17811 869 -17777 879
rect -17811 657 -17777 673
rect -17715 863 -17681 879
rect -17715 657 -17681 667
rect -17619 869 -17585 879
rect -17619 657 -17585 673
rect -17523 863 -17489 879
rect -17523 657 -17489 667
rect -17427 869 -17393 879
rect -17427 657 -17393 673
rect -16894 869 -16860 879
rect -16894 657 -16860 673
rect -16798 863 -16764 879
rect -16798 657 -16764 667
rect -16702 869 -16668 879
rect -16702 657 -16668 673
rect -16606 863 -16572 879
rect -16606 657 -16572 667
rect -16510 869 -16476 879
rect -16510 657 -16476 673
rect -16414 863 -16380 879
rect -16414 657 -16380 667
rect -16318 869 -16284 879
rect -16318 657 -16284 673
rect -16012 869 -15978 879
rect -16012 657 -15978 673
rect -15916 863 -15882 879
rect -15916 657 -15882 667
rect -15820 869 -15786 879
rect -15820 657 -15786 673
rect -15724 863 -15690 879
rect -15724 657 -15690 667
rect -15628 869 -15594 879
rect -15628 657 -15594 673
rect -15532 863 -15498 879
rect -15532 657 -15498 667
rect -15436 869 -15402 879
rect -15436 657 -15402 673
rect -14712 869 -14678 879
rect -14712 657 -14678 673
rect -14616 863 -14582 879
rect -14616 657 -14582 667
rect -14520 869 -14486 879
rect -14520 657 -14486 673
rect -14424 863 -14390 879
rect -14424 657 -14390 667
rect -14328 869 -14294 879
rect -14328 657 -14294 673
rect -14232 863 -14198 879
rect -14232 657 -14198 667
rect -14136 869 -14102 879
rect -14136 657 -14102 673
rect -13603 869 -13569 879
rect -13603 657 -13569 673
rect -13507 863 -13473 879
rect -13507 657 -13473 667
rect -13411 869 -13377 879
rect -13411 657 -13377 673
rect -13315 863 -13281 879
rect -13315 657 -13281 667
rect -13219 869 -13185 879
rect -13219 657 -13185 673
rect -13123 863 -13089 879
rect -13123 657 -13089 667
rect -13027 869 -12993 879
rect -13027 657 -12993 673
rect -12721 869 -12687 879
rect -12721 657 -12687 673
rect -12625 863 -12591 879
rect -12625 657 -12591 667
rect -12529 869 -12495 879
rect -12529 657 -12495 673
rect -12433 863 -12399 879
rect -12433 657 -12399 667
rect -12337 869 -12303 879
rect -12337 657 -12303 673
rect -12241 863 -12207 879
rect -12241 657 -12207 667
rect -12145 869 -12111 879
rect -12145 657 -12111 673
rect -11421 869 -11387 879
rect -11421 657 -11387 673
rect -11325 863 -11291 879
rect -11325 657 -11291 667
rect -11229 869 -11195 879
rect -11229 657 -11195 673
rect -11133 863 -11099 879
rect -11133 657 -11099 667
rect -11037 869 -11003 879
rect -11037 657 -11003 673
rect -10941 863 -10907 879
rect -10941 657 -10907 667
rect -10845 869 -10811 879
rect -10845 657 -10811 673
rect -10312 869 -10278 879
rect -10312 657 -10278 673
rect -10216 863 -10182 879
rect -10216 657 -10182 667
rect -10120 869 -10086 879
rect -10120 657 -10086 673
rect -10024 863 -9990 879
rect -10024 657 -9990 667
rect -9928 869 -9894 879
rect -9928 657 -9894 673
rect -9832 863 -9798 879
rect -9832 657 -9798 667
rect -9736 869 -9702 879
rect -9736 657 -9702 673
rect -9430 869 -9396 879
rect -9430 657 -9396 673
rect -9334 863 -9300 879
rect -9334 657 -9300 667
rect -9238 869 -9204 879
rect -9238 657 -9204 673
rect -9142 863 -9108 879
rect -9142 657 -9108 667
rect -9046 869 -9012 879
rect -9046 657 -9012 673
rect -8950 863 -8916 879
rect -8950 657 -8916 667
rect -8854 869 -8820 879
rect -8854 657 -8820 673
rect -8131 869 -8097 879
rect -8131 657 -8097 673
rect -8035 863 -8001 879
rect -8035 657 -8001 667
rect -7939 869 -7905 879
rect -7939 657 -7905 673
rect -7843 863 -7809 879
rect -7843 657 -7809 667
rect -7747 869 -7713 879
rect -7747 657 -7713 673
rect -7651 863 -7617 879
rect -7651 657 -7617 667
rect -7555 869 -7521 879
rect -7555 657 -7521 673
rect -7022 869 -6988 879
rect -7022 657 -6988 673
rect -6926 863 -6892 879
rect -6926 657 -6892 667
rect -6830 869 -6796 879
rect -6830 657 -6796 673
rect -6734 863 -6700 879
rect -6734 657 -6700 667
rect -6638 869 -6604 879
rect -6638 657 -6604 673
rect -6542 863 -6508 879
rect -6542 657 -6508 667
rect -6446 869 -6412 879
rect -6446 657 -6412 673
rect -6140 869 -6106 879
rect -6140 657 -6106 673
rect -6044 863 -6010 879
rect -6044 657 -6010 667
rect -5948 869 -5914 879
rect -5948 657 -5914 673
rect -5852 863 -5818 879
rect -5852 657 -5818 667
rect -5756 869 -5722 879
rect -5756 657 -5722 673
rect -5660 863 -5626 879
rect -5660 657 -5626 667
rect -5564 869 -5530 879
rect -5564 657 -5530 673
rect -4840 869 -4806 879
rect -4840 657 -4806 673
rect -4744 863 -4710 879
rect -4744 657 -4710 667
rect -4648 869 -4614 879
rect -4648 657 -4614 673
rect -4552 863 -4518 879
rect -4552 657 -4518 667
rect -4456 869 -4422 879
rect -4456 657 -4422 673
rect -4360 863 -4326 879
rect -4360 657 -4326 667
rect -4264 869 -4230 879
rect -4264 657 -4230 673
rect -3731 869 -3697 879
rect -3731 657 -3697 673
rect -3635 863 -3601 879
rect -3635 657 -3601 667
rect -3539 869 -3505 879
rect -3539 657 -3505 673
rect -3443 863 -3409 879
rect -3443 657 -3409 667
rect -3347 869 -3313 879
rect -3347 657 -3313 673
rect -3251 863 -3217 879
rect -3251 657 -3217 667
rect -3155 869 -3121 879
rect -3155 657 -3121 673
rect -2849 869 -2815 879
rect -2849 657 -2815 673
rect -2753 863 -2719 879
rect -2753 657 -2719 667
rect -2657 869 -2623 879
rect -2657 657 -2623 673
rect -2561 863 -2527 879
rect -2561 657 -2527 667
rect -2465 869 -2431 879
rect -2465 657 -2431 673
rect -2369 863 -2335 879
rect -2369 657 -2335 667
rect -2273 869 -2239 879
rect -2273 657 -2239 673
rect -1549 869 -1515 879
rect -1549 657 -1515 673
rect -1453 863 -1419 879
rect -1453 657 -1419 667
rect -1357 869 -1323 879
rect -1357 657 -1323 673
rect -1261 863 -1227 879
rect -1261 657 -1227 667
rect -1165 869 -1131 879
rect -1165 657 -1131 673
rect -1069 863 -1035 879
rect -1069 657 -1035 667
rect -973 869 -939 879
rect -973 657 -939 673
rect -440 869 -406 879
rect -440 657 -406 673
rect -344 863 -310 879
rect -344 657 -310 667
rect -248 869 -214 879
rect -248 657 -214 673
rect -152 863 -118 879
rect -152 657 -118 667
rect -56 869 -22 879
rect -56 657 -22 673
rect 40 863 74 879
rect 40 657 74 667
rect 136 869 170 879
rect 136 657 170 673
rect 442 869 476 879
rect 442 657 476 673
rect 538 863 572 879
rect 538 657 572 667
rect 634 869 668 879
rect 634 657 668 673
rect 730 863 764 879
rect 730 657 764 667
rect 826 869 860 879
rect 826 657 860 673
rect 922 863 956 879
rect 922 657 956 667
rect 1018 869 1052 879
rect 7333 786 7372 1537
rect 7298 774 7372 786
rect 7298 758 7406 774
rect 7756 1550 7790 1566
rect 7756 758 7790 774
rect 8246 1550 8354 1566
rect 8246 1537 8320 1550
rect 8281 786 8320 1537
rect 8246 774 8320 786
rect 8246 758 8354 774
rect 8704 1550 8738 1566
rect 8704 758 8738 774
rect 9182 1550 9290 1566
rect 9182 1537 9256 1550
rect 9217 786 9256 1537
rect 9182 774 9256 786
rect 9182 758 9290 774
rect 9640 1550 9674 1566
rect 9640 758 9674 774
rect 10113 1551 10221 1567
rect 10113 1538 10187 1551
rect 10148 787 10187 1538
rect 10113 775 10187 787
rect 10113 759 10221 775
rect 10571 1551 10605 1567
rect 10571 759 10605 775
rect 11040 1550 11148 1566
rect 11040 1537 11114 1550
rect 11075 786 11114 1537
rect 11040 774 11114 786
rect 7298 755 7403 758
rect 8246 755 8351 758
rect 9182 755 9287 758
rect 10113 756 10218 759
rect 11040 758 11148 774
rect 11498 1550 11532 1566
rect 12297 1564 12313 1598
rect 12347 1564 12363 1598
rect 12169 1508 12203 1524
rect 12169 1260 12203 1332
rect 12265 1508 12299 1524
rect 12265 1316 12299 1332
rect 12361 1508 12395 1524
rect 12826 1399 12876 1619
rect 12919 1571 12935 1605
rect 13129 1571 13147 1605
rect 12919 1409 12935 1443
rect 13111 1409 13127 1443
rect 12826 1365 12842 1399
rect 12826 1349 12876 1365
rect 12361 1260 12395 1332
rect 12919 1321 12935 1355
rect 13111 1321 13127 1355
rect 12157 1249 12407 1260
rect 12157 1188 12183 1249
rect 12382 1188 12407 1249
rect 12938 1219 12954 1253
rect 13086 1219 13102 1253
rect 12157 1176 12407 1188
rect 11498 758 11532 774
rect 11040 755 11145 758
rect 1018 657 1052 673
rect -24536 579 -24519 614
rect -24485 579 -24469 614
rect -24247 608 -24230 614
rect -24435 579 -24230 608
rect -24196 579 -24180 614
rect -24536 373 -24493 579
rect -24435 574 -24180 579
rect -23427 579 -23410 614
rect -23376 579 -23360 614
rect -23138 608 -23121 614
rect -23326 579 -23121 608
rect -23087 579 -23071 614
rect -24435 490 -24401 574
rect -24367 485 -24351 519
rect -23975 485 -23959 519
rect -24435 439 -24401 455
rect -23427 373 -23384 579
rect -23326 574 -23071 579
rect -22545 579 -22528 614
rect -22494 579 -22478 614
rect -22256 608 -22239 614
rect -22444 579 -22239 608
rect -22205 579 -22189 614
rect -23326 490 -23292 574
rect -23258 485 -23242 519
rect -22866 485 -22850 519
rect -23326 439 -23292 455
rect -22545 373 -22502 579
rect -22444 574 -22189 579
rect -21245 579 -21228 614
rect -21194 579 -21178 614
rect -20956 608 -20939 614
rect -21144 579 -20939 608
rect -20905 579 -20889 614
rect -22444 490 -22410 574
rect -22376 485 -22360 519
rect -21984 485 -21968 519
rect -22444 439 -22410 455
rect -21245 373 -21202 579
rect -21144 574 -20889 579
rect -20136 579 -20119 614
rect -20085 579 -20069 614
rect -19847 608 -19830 614
rect -20035 579 -19830 608
rect -19796 579 -19780 614
rect -21144 490 -21110 574
rect -21076 485 -21060 519
rect -20684 485 -20668 519
rect -21144 439 -21110 455
rect -20136 373 -20093 579
rect -20035 574 -19780 579
rect -19254 579 -19237 614
rect -19203 579 -19187 614
rect -18965 608 -18948 614
rect -19153 579 -18948 608
rect -18914 579 -18898 614
rect -20035 490 -20001 574
rect -19967 485 -19951 519
rect -19575 485 -19559 519
rect -20035 439 -20001 455
rect -19254 373 -19211 579
rect -19153 574 -18898 579
rect -17954 579 -17937 614
rect -17903 579 -17887 614
rect -17665 608 -17648 614
rect -17853 579 -17648 608
rect -17614 579 -17598 614
rect -19153 490 -19119 574
rect -19085 485 -19069 519
rect -18693 485 -18677 519
rect -19153 439 -19119 455
rect -17954 373 -17911 579
rect -17853 574 -17598 579
rect -16845 579 -16828 614
rect -16794 579 -16778 614
rect -16556 608 -16539 614
rect -16744 579 -16539 608
rect -16505 579 -16489 614
rect -17853 490 -17819 574
rect -17785 485 -17769 519
rect -17393 485 -17377 519
rect -17853 439 -17819 455
rect -16845 373 -16802 579
rect -16744 574 -16489 579
rect -15963 579 -15946 614
rect -15912 579 -15896 614
rect -15674 608 -15657 614
rect -15862 579 -15657 608
rect -15623 579 -15607 614
rect -16744 490 -16710 574
rect -16676 485 -16660 519
rect -16284 485 -16268 519
rect -16744 439 -16710 455
rect -15963 373 -15920 579
rect -15862 574 -15607 579
rect -14663 579 -14646 614
rect -14612 579 -14596 614
rect -14374 608 -14357 614
rect -14562 579 -14357 608
rect -14323 579 -14307 614
rect -15862 490 -15828 574
rect -15794 485 -15778 519
rect -15402 485 -15386 519
rect -15862 439 -15828 455
rect -14663 373 -14620 579
rect -14562 574 -14307 579
rect -13554 579 -13537 614
rect -13503 579 -13487 614
rect -13265 608 -13248 614
rect -13453 579 -13248 608
rect -13214 579 -13198 614
rect -14562 490 -14528 574
rect -14494 485 -14478 519
rect -14102 485 -14086 519
rect -14562 439 -14528 455
rect -13554 373 -13511 579
rect -13453 574 -13198 579
rect -12672 579 -12655 614
rect -12621 579 -12605 614
rect -12383 608 -12366 614
rect -12571 579 -12366 608
rect -12332 579 -12316 614
rect -13453 490 -13419 574
rect -13385 485 -13369 519
rect -12993 485 -12977 519
rect -13453 439 -13419 455
rect -12672 373 -12629 579
rect -12571 574 -12316 579
rect -11372 579 -11355 614
rect -11321 579 -11305 614
rect -11083 608 -11066 614
rect -11271 579 -11066 608
rect -11032 579 -11016 614
rect -12571 490 -12537 574
rect -12503 485 -12487 519
rect -12111 485 -12095 519
rect -12571 439 -12537 455
rect -11372 373 -11329 579
rect -11271 574 -11016 579
rect -10263 579 -10246 614
rect -10212 579 -10196 614
rect -9974 608 -9957 614
rect -10162 579 -9957 608
rect -9923 579 -9907 614
rect -11271 490 -11237 574
rect -11203 485 -11187 519
rect -10811 485 -10795 519
rect -11271 439 -11237 455
rect -10263 373 -10220 579
rect -10162 574 -9907 579
rect -9381 579 -9364 614
rect -9330 579 -9314 614
rect -9092 608 -9075 614
rect -9280 579 -9075 608
rect -9041 579 -9025 614
rect -10162 490 -10128 574
rect -10094 485 -10078 519
rect -9702 485 -9686 519
rect -10162 439 -10128 455
rect -9381 373 -9338 579
rect -9280 574 -9025 579
rect -8082 579 -8065 614
rect -8031 579 -8015 614
rect -7793 608 -7776 614
rect -7981 579 -7776 608
rect -7742 579 -7726 614
rect -9280 490 -9246 574
rect -9212 485 -9196 519
rect -8820 485 -8804 519
rect -9280 439 -9246 455
rect -8082 373 -8039 579
rect -7981 574 -7726 579
rect -6973 579 -6956 614
rect -6922 579 -6906 614
rect -6684 608 -6667 614
rect -6872 579 -6667 608
rect -6633 579 -6617 614
rect -7981 490 -7947 574
rect -7913 485 -7897 519
rect -7521 485 -7505 519
rect -7981 439 -7947 455
rect -6973 373 -6930 579
rect -6872 574 -6617 579
rect -6091 579 -6074 614
rect -6040 579 -6024 614
rect -5802 608 -5785 614
rect -5990 579 -5785 608
rect -5751 579 -5735 614
rect -6872 490 -6838 574
rect -6804 485 -6788 519
rect -6412 485 -6396 519
rect -6872 439 -6838 455
rect -6091 373 -6048 579
rect -5990 574 -5735 579
rect -4791 579 -4774 614
rect -4740 579 -4724 614
rect -4502 608 -4485 614
rect -4690 579 -4485 608
rect -4451 579 -4435 614
rect -5990 490 -5956 574
rect -5922 485 -5906 519
rect -5530 485 -5514 519
rect -5990 439 -5956 455
rect -4791 373 -4748 579
rect -4690 574 -4435 579
rect -3682 579 -3665 614
rect -3631 579 -3615 614
rect -3393 608 -3376 614
rect -3581 579 -3376 608
rect -3342 579 -3326 614
rect -4690 490 -4656 574
rect -4622 485 -4606 519
rect -4230 485 -4214 519
rect -4690 439 -4656 455
rect -3682 373 -3639 579
rect -3581 574 -3326 579
rect -2800 579 -2783 614
rect -2749 579 -2733 614
rect -2511 608 -2494 614
rect -2699 579 -2494 608
rect -2460 579 -2444 614
rect -3581 490 -3547 574
rect -3513 485 -3497 519
rect -3121 485 -3105 519
rect -3581 439 -3547 455
rect -2800 373 -2757 579
rect -2699 574 -2444 579
rect -1500 579 -1483 614
rect -1449 579 -1433 614
rect -1211 608 -1194 614
rect -1399 579 -1194 608
rect -1160 579 -1144 614
rect -2699 490 -2665 574
rect -2631 485 -2615 519
rect -2239 485 -2223 519
rect -2699 439 -2665 455
rect -1500 373 -1457 579
rect -1399 574 -1144 579
rect -391 579 -374 614
rect -340 579 -324 614
rect -102 608 -85 614
rect -290 579 -85 608
rect -51 579 -35 614
rect -1399 490 -1365 574
rect -1331 485 -1315 519
rect -939 485 -923 519
rect -1399 439 -1365 455
rect -391 373 -348 579
rect -290 574 -35 579
rect 491 579 508 614
rect 542 579 558 614
rect 780 608 797 614
rect 592 579 797 608
rect 831 579 847 614
rect -290 490 -256 574
rect -222 485 -206 519
rect 170 485 186 519
rect -290 439 -256 455
rect 491 373 534 579
rect 592 574 847 579
rect 592 490 626 574
rect 660 485 676 519
rect 1052 485 1068 519
rect 592 439 626 455
rect 7182 402 7198 436
rect 7232 402 7248 436
rect 7374 402 7390 436
rect 7424 402 7440 436
rect 7566 402 7582 436
rect 7616 402 7632 436
rect 7758 402 7774 436
rect 7808 402 7824 436
rect 8130 402 8146 436
rect 8180 402 8196 436
rect 8322 402 8338 436
rect 8372 402 8388 436
rect 8514 402 8530 436
rect 8564 402 8580 436
rect 8706 402 8722 436
rect 8756 402 8772 436
rect 9066 402 9082 436
rect 9116 402 9132 436
rect 9258 402 9274 436
rect 9308 402 9324 436
rect 9450 402 9466 436
rect 9500 402 9516 436
rect 9642 402 9658 436
rect 9692 402 9708 436
rect 9997 403 10013 437
rect 10047 403 10063 437
rect 10189 403 10205 437
rect 10239 403 10255 437
rect 10381 403 10397 437
rect 10431 403 10447 437
rect 10573 403 10589 437
rect 10623 403 10639 437
rect 10924 402 10940 436
rect 10974 402 10990 436
rect 11116 402 11132 436
rect 11166 402 11182 436
rect 11308 402 11324 436
rect 11358 402 11374 436
rect 11500 402 11516 436
rect 11550 402 11566 436
rect -24536 357 -24401 373
rect -24536 322 -24435 357
rect -23427 357 -23292 373
rect -24536 306 -24401 322
rect -24367 293 -24351 327
rect -23975 293 -23959 327
rect -23427 322 -23326 357
rect -22545 357 -22410 373
rect -23427 306 -23292 322
rect -23258 293 -23242 327
rect -22866 293 -22850 327
rect -22545 322 -22444 357
rect -21245 357 -21110 373
rect -22545 306 -22410 322
rect -22376 293 -22360 327
rect -21984 293 -21968 327
rect -21245 322 -21144 357
rect -20136 357 -20001 373
rect -21245 306 -21110 322
rect -21076 293 -21060 327
rect -20684 293 -20668 327
rect -20136 322 -20035 357
rect -19254 357 -19119 373
rect -20136 306 -20001 322
rect -19967 293 -19951 327
rect -19575 293 -19559 327
rect -19254 322 -19153 357
rect -17954 357 -17819 373
rect -19254 306 -19119 322
rect -19085 293 -19069 327
rect -18693 293 -18677 327
rect -17954 322 -17853 357
rect -16845 357 -16710 373
rect -17954 306 -17819 322
rect -17785 293 -17769 327
rect -17393 293 -17377 327
rect -16845 322 -16744 357
rect -15963 357 -15828 373
rect -16845 306 -16710 322
rect -16676 293 -16660 327
rect -16284 293 -16268 327
rect -15963 322 -15862 357
rect -14663 357 -14528 373
rect -15963 306 -15828 322
rect -15794 293 -15778 327
rect -15402 293 -15386 327
rect -14663 322 -14562 357
rect -13554 357 -13419 373
rect -14663 306 -14528 322
rect -14494 293 -14478 327
rect -14102 293 -14086 327
rect -13554 322 -13453 357
rect -12672 357 -12537 373
rect -13554 306 -13419 322
rect -13385 293 -13369 327
rect -12993 293 -12977 327
rect -12672 322 -12571 357
rect -11372 357 -11237 373
rect -12672 306 -12537 322
rect -12503 293 -12487 327
rect -12111 293 -12095 327
rect -11372 322 -11271 357
rect -10263 357 -10128 373
rect -11372 306 -11237 322
rect -11203 293 -11187 327
rect -10811 293 -10795 327
rect -10263 322 -10162 357
rect -9381 357 -9246 373
rect -10263 306 -10128 322
rect -10094 293 -10078 327
rect -9702 293 -9686 327
rect -9381 322 -9280 357
rect -8082 357 -7947 373
rect -9381 306 -9246 322
rect -9212 293 -9196 327
rect -8820 293 -8804 327
rect -8082 322 -7981 357
rect -6973 357 -6838 373
rect -8082 306 -7947 322
rect -7913 293 -7897 327
rect -7521 293 -7505 327
rect -6973 322 -6872 357
rect -6091 357 -5956 373
rect -6973 306 -6838 322
rect -6804 293 -6788 327
rect -6412 293 -6396 327
rect -6091 322 -5990 357
rect -4791 357 -4656 373
rect -6091 306 -5956 322
rect -5922 293 -5906 327
rect -5530 293 -5514 327
rect -4791 322 -4690 357
rect -3682 357 -3547 373
rect -4791 306 -4656 322
rect -4622 293 -4606 327
rect -4230 293 -4214 327
rect -3682 322 -3581 357
rect -2800 357 -2665 373
rect -3682 306 -3547 322
rect -3513 293 -3497 327
rect -3121 293 -3105 327
rect -2800 322 -2699 357
rect -1500 357 -1365 373
rect -2800 306 -2665 322
rect -2631 293 -2615 327
rect -2239 293 -2223 327
rect -1500 322 -1399 357
rect -391 357 -256 373
rect -1500 306 -1365 322
rect -1331 293 -1315 327
rect -939 293 -923 327
rect -391 322 -290 357
rect 491 357 626 373
rect -391 306 -256 322
rect -222 293 -206 327
rect 170 293 186 327
rect 491 322 592 357
rect 7150 343 7184 359
rect 7246 348 7280 359
rect 491 306 626 322
rect 660 293 676 327
rect 1052 293 1068 327
rect -24363 221 -24336 255
rect -24001 221 -23963 255
rect -23254 221 -23227 255
rect -22892 221 -22854 255
rect -22372 221 -22345 255
rect -22010 221 -21972 255
rect -21072 221 -21045 255
rect -20710 221 -20672 255
rect -19963 221 -19936 255
rect -19601 221 -19563 255
rect -19081 221 -19054 255
rect -18719 221 -18681 255
rect -17781 221 -17754 255
rect -17419 221 -17381 255
rect -16672 221 -16645 255
rect -16310 221 -16272 255
rect -15790 221 -15763 255
rect -15428 221 -15390 255
rect -14490 221 -14463 255
rect -14128 221 -14090 255
rect -13381 221 -13354 255
rect -13019 221 -12981 255
rect -12499 221 -12472 255
rect -12137 221 -12099 255
rect -11199 221 -11172 255
rect -10837 221 -10799 255
rect -10090 221 -10063 255
rect -9728 221 -9690 255
rect -9208 221 -9181 255
rect -8846 221 -8808 255
rect -7909 221 -7882 255
rect -7547 221 -7509 255
rect -6800 221 -6773 255
rect -6438 221 -6400 255
rect -5918 221 -5891 255
rect -5556 221 -5518 255
rect -4618 221 -4591 255
rect -4256 221 -4218 255
rect -3509 221 -3482 255
rect -3147 221 -3109 255
rect -2627 221 -2600 255
rect -2265 221 -2227 255
rect -1327 221 -1300 255
rect -965 221 -927 255
rect -218 221 -191 255
rect 144 221 182 255
rect 664 221 691 255
rect 1026 221 1064 255
rect 7150 29 7184 45
rect 7246 29 7280 45
rect 7342 343 7376 359
rect 7342 29 7376 45
rect 7438 348 7472 359
rect 7534 343 7568 359
rect 7438 29 7472 45
rect 7534 29 7568 45
rect 7630 348 7664 359
rect 7726 343 7760 359
rect 7630 29 7664 45
rect 7726 29 7760 45
rect 7822 348 7856 359
rect 7918 343 7952 359
rect 7822 29 7856 45
rect 7918 29 7952 45
rect 8098 343 8132 359
rect 8194 348 8228 359
rect 8098 29 8132 45
rect 8194 29 8228 45
rect 8290 343 8324 359
rect 8290 29 8324 45
rect 8386 348 8420 359
rect 8482 343 8516 359
rect 8386 29 8420 45
rect 8482 29 8516 45
rect 8578 348 8612 359
rect 8674 343 8708 359
rect 8578 29 8612 45
rect 8674 29 8708 45
rect 8770 348 8804 359
rect 8866 343 8900 359
rect 8770 29 8804 45
rect 8866 29 8900 45
rect 9034 343 9068 359
rect 9130 348 9164 359
rect 9034 29 9068 45
rect 9130 29 9164 45
rect 9226 343 9260 359
rect 9226 29 9260 45
rect 9322 348 9356 359
rect 9418 343 9452 359
rect 9322 29 9356 45
rect 9418 29 9452 45
rect 9514 348 9548 359
rect 9610 343 9644 359
rect 9514 29 9548 45
rect 9610 29 9644 45
rect 9706 348 9740 359
rect 9802 343 9836 359
rect 9706 29 9740 45
rect 9802 29 9836 45
rect 9965 344 9999 360
rect 10061 349 10095 360
rect 9965 30 9999 46
rect 10061 30 10095 46
rect 10157 344 10191 360
rect 10157 30 10191 46
rect 10253 349 10287 360
rect 10349 344 10383 360
rect 10253 30 10287 46
rect 10349 30 10383 46
rect 10445 349 10479 360
rect 10541 344 10575 360
rect 10445 30 10479 46
rect 10541 30 10575 46
rect 10637 349 10671 360
rect 10733 344 10767 360
rect 10637 30 10671 46
rect 10733 30 10767 46
rect 10892 343 10926 359
rect 10988 348 11022 359
rect 10892 29 10926 45
rect 10988 29 11022 45
rect 11084 343 11118 359
rect 11084 29 11118 45
rect 11180 348 11214 359
rect 11276 343 11310 359
rect 11180 29 11214 45
rect 11276 29 11310 45
rect 11372 348 11406 359
rect 11468 343 11502 359
rect 11372 29 11406 45
rect 11468 29 11502 45
rect 11564 348 11598 359
rect 11660 343 11694 359
rect 11564 29 11598 45
rect 11660 29 11694 45
rect 7373 -59 7389 -24
rect 7677 -59 7703 -24
rect 8321 -59 8337 -24
rect 8625 -59 8651 -24
rect 9257 -59 9273 -24
rect 9561 -59 9587 -24
rect 10188 -58 10204 -23
rect 10492 -58 10518 -23
rect 11115 -59 11131 -24
rect 11419 -59 11445 -24
rect 5705 -579 5721 -545
rect 5812 -579 5828 -545
rect 6145 -579 6161 -545
rect 6252 -579 6268 -545
rect 6585 -579 6601 -545
rect 6692 -579 6708 -545
rect 5561 -665 5611 -648
rect 5654 -651 5664 -617
rect 5860 -651 5876 -617
rect 5561 -891 5577 -665
rect 6001 -665 6051 -648
rect 6094 -651 6104 -617
rect 6300 -651 6316 -617
rect 5654 -747 5670 -713
rect 5864 -747 5882 -713
rect 5654 -843 5664 -809
rect 5860 -843 5876 -809
rect 5561 -1111 5611 -891
rect 6001 -891 6017 -665
rect 6441 -665 6491 -648
rect 6534 -651 6544 -617
rect 6740 -651 6756 -617
rect 6094 -747 6110 -713
rect 6304 -747 6322 -713
rect 6094 -843 6104 -809
rect 6300 -843 6316 -809
rect 5654 -939 5670 -905
rect 5864 -939 5882 -905
rect 5654 -1101 5670 -1067
rect 5846 -1101 5862 -1067
rect 5561 -1145 5577 -1111
rect 5561 -1161 5611 -1145
rect 6001 -1111 6051 -891
rect 6441 -891 6457 -665
rect 6534 -747 6550 -713
rect 6744 -747 6762 -713
rect 6534 -843 6544 -809
rect 6740 -843 6756 -809
rect 6094 -939 6110 -905
rect 6304 -939 6322 -905
rect 6094 -1101 6110 -1067
rect 6286 -1101 6302 -1067
rect 6001 -1145 6017 -1111
rect 5654 -1189 5670 -1155
rect 5846 -1189 5862 -1155
rect 6001 -1161 6051 -1145
rect 6441 -1111 6491 -891
rect 6534 -939 6550 -905
rect 6744 -939 6762 -905
rect 6534 -1101 6550 -1067
rect 6726 -1101 6742 -1067
rect 6441 -1145 6457 -1111
rect 6094 -1189 6110 -1155
rect 6286 -1189 6302 -1155
rect 6441 -1161 6491 -1145
rect 6534 -1189 6550 -1155
rect 6726 -1189 6742 -1155
rect 7373 -1252 7389 -1217
rect 7677 -1252 7703 -1217
rect 8321 -1252 8337 -1217
rect 8625 -1252 8651 -1217
rect 9257 -1252 9273 -1217
rect 9561 -1252 9587 -1217
rect 10188 -1252 10204 -1217
rect 10492 -1252 10518 -1217
rect 11115 -1252 11131 -1217
rect 11419 -1252 11445 -1217
rect 5673 -1291 5689 -1257
rect 5821 -1291 5837 -1257
rect 6113 -1291 6129 -1257
rect 6261 -1291 6277 -1257
rect 6553 -1291 6569 -1257
rect 6701 -1291 6717 -1257
rect 7150 -1321 7184 -1305
rect 7246 -1321 7280 -1305
rect 7150 -1635 7184 -1619
rect 7246 -1635 7280 -1624
rect 7342 -1321 7376 -1305
rect 7342 -1635 7376 -1619
rect 7438 -1321 7472 -1305
rect 7534 -1321 7568 -1305
rect 7438 -1635 7472 -1624
rect 7534 -1635 7568 -1619
rect 7630 -1321 7664 -1305
rect 7726 -1321 7760 -1305
rect 7630 -1635 7664 -1624
rect 7726 -1635 7760 -1619
rect 7822 -1321 7856 -1305
rect 7918 -1321 7952 -1305
rect 7822 -1635 7856 -1624
rect 7918 -1635 7952 -1619
rect 8098 -1321 8132 -1305
rect 8194 -1321 8228 -1305
rect 8098 -1635 8132 -1619
rect 8194 -1635 8228 -1624
rect 8290 -1321 8324 -1305
rect 8290 -1635 8324 -1619
rect 8386 -1321 8420 -1305
rect 8482 -1321 8516 -1305
rect 8386 -1635 8420 -1624
rect 8482 -1635 8516 -1619
rect 8578 -1321 8612 -1305
rect 8674 -1321 8708 -1305
rect 8578 -1635 8612 -1624
rect 8674 -1635 8708 -1619
rect 8770 -1321 8804 -1305
rect 8866 -1321 8900 -1305
rect 8770 -1635 8804 -1624
rect 8866 -1635 8900 -1619
rect 9034 -1321 9068 -1305
rect 9130 -1321 9164 -1305
rect 9034 -1635 9068 -1619
rect 9130 -1635 9164 -1624
rect 9226 -1321 9260 -1305
rect 9226 -1635 9260 -1619
rect 9322 -1321 9356 -1305
rect 9418 -1321 9452 -1305
rect 9322 -1635 9356 -1624
rect 9418 -1635 9452 -1619
rect 9514 -1321 9548 -1305
rect 9610 -1321 9644 -1305
rect 9514 -1635 9548 -1624
rect 9610 -1635 9644 -1619
rect 9706 -1321 9740 -1305
rect 9802 -1321 9836 -1305
rect 9706 -1635 9740 -1624
rect 9802 -1635 9836 -1619
rect 9965 -1321 9999 -1305
rect 10061 -1321 10095 -1305
rect 9965 -1635 9999 -1619
rect 10061 -1635 10095 -1624
rect 10157 -1321 10191 -1305
rect 10157 -1635 10191 -1619
rect 10253 -1321 10287 -1305
rect 10349 -1321 10383 -1305
rect 10253 -1635 10287 -1624
rect 10349 -1635 10383 -1619
rect 10445 -1321 10479 -1305
rect 10541 -1321 10575 -1305
rect 10445 -1635 10479 -1624
rect 10541 -1635 10575 -1619
rect 10637 -1321 10671 -1305
rect 10733 -1321 10767 -1305
rect 10637 -1635 10671 -1624
rect 10733 -1635 10767 -1619
rect 10892 -1321 10926 -1305
rect 10988 -1321 11022 -1305
rect 10892 -1635 10926 -1619
rect 10988 -1635 11022 -1624
rect 11084 -1321 11118 -1305
rect 11084 -1635 11118 -1619
rect 11180 -1321 11214 -1305
rect 11276 -1321 11310 -1305
rect 11180 -1635 11214 -1624
rect 11276 -1635 11310 -1619
rect 11372 -1321 11406 -1305
rect 11468 -1321 11502 -1305
rect 11372 -1635 11406 -1624
rect 11468 -1635 11502 -1619
rect 11564 -1321 11598 -1305
rect 11660 -1321 11694 -1305
rect 11564 -1635 11598 -1624
rect 11660 -1635 11694 -1619
rect 7182 -1712 7198 -1678
rect 7232 -1712 7248 -1678
rect 7374 -1712 7390 -1678
rect 7424 -1712 7440 -1678
rect 7566 -1712 7582 -1678
rect 7616 -1712 7632 -1678
rect 7758 -1712 7774 -1678
rect 7808 -1712 7824 -1678
rect 8130 -1712 8146 -1678
rect 8180 -1712 8196 -1678
rect 8322 -1712 8338 -1678
rect 8372 -1712 8388 -1678
rect 8514 -1712 8530 -1678
rect 8564 -1712 8580 -1678
rect 8706 -1712 8722 -1678
rect 8756 -1712 8772 -1678
rect 9066 -1712 9082 -1678
rect 9116 -1712 9132 -1678
rect 9258 -1712 9274 -1678
rect 9308 -1712 9324 -1678
rect 9450 -1712 9466 -1678
rect 9500 -1712 9516 -1678
rect 9642 -1712 9658 -1678
rect 9692 -1712 9708 -1678
rect 9997 -1712 10013 -1678
rect 10047 -1712 10063 -1678
rect 10189 -1712 10205 -1678
rect 10239 -1712 10255 -1678
rect 10381 -1712 10397 -1678
rect 10431 -1712 10447 -1678
rect 10573 -1712 10589 -1678
rect 10623 -1712 10639 -1678
rect 10924 -1712 10940 -1678
rect 10974 -1712 10990 -1678
rect 11116 -1712 11132 -1678
rect 11166 -1712 11182 -1678
rect 11308 -1712 11324 -1678
rect 11358 -1712 11374 -1678
rect 11500 -1712 11516 -1678
rect 11550 -1712 11566 -1678
rect 7298 -2034 7403 -2031
rect 8246 -2034 8351 -2031
rect 9182 -2034 9287 -2031
rect 10113 -2034 10218 -2031
rect 11040 -2034 11145 -2031
rect 7298 -2050 7406 -2034
rect 7298 -2062 7372 -2050
rect -23581 -2281 -23565 -2247
rect -23474 -2281 -23458 -2247
rect -21561 -2281 -21545 -2247
rect -21454 -2281 -21438 -2247
rect -19820 -2281 -19804 -2247
rect -19713 -2281 -19697 -2247
rect -18041 -2281 -18025 -2247
rect -17934 -2281 -17918 -2247
rect -24435 -2347 -24419 -2300
rect -23850 -2347 -23826 -2300
rect -23725 -2367 -23675 -2350
rect -23632 -2353 -23622 -2319
rect -23426 -2353 -23410 -2319
rect -22398 -2347 -22382 -2300
rect -21813 -2347 -21789 -2300
rect -24435 -2419 -24401 -2409
rect -24435 -2631 -24401 -2615
rect -24339 -2425 -24305 -2409
rect -24339 -2631 -24305 -2621
rect -24243 -2419 -24209 -2409
rect -24243 -2631 -24209 -2615
rect -24147 -2425 -24113 -2409
rect -24147 -2631 -24113 -2621
rect -24051 -2419 -24017 -2409
rect -24051 -2631 -24017 -2615
rect -23955 -2425 -23921 -2409
rect -23955 -2631 -23921 -2621
rect -23859 -2419 -23825 -2409
rect -23859 -2631 -23825 -2615
rect -23725 -2593 -23709 -2367
rect -21705 -2367 -21655 -2350
rect -21612 -2353 -21602 -2319
rect -21406 -2353 -21390 -2319
rect -20668 -2347 -20652 -2300
rect -20083 -2347 -20059 -2300
rect -23632 -2449 -23616 -2415
rect -23422 -2449 -23404 -2415
rect -22398 -2419 -22364 -2409
rect -23632 -2545 -23622 -2511
rect -23426 -2545 -23410 -2511
rect -24386 -2709 -24369 -2674
rect -24335 -2709 -24319 -2674
rect -24097 -2680 -24080 -2674
rect -24285 -2709 -24080 -2680
rect -24046 -2709 -24030 -2674
rect -24386 -2915 -24343 -2709
rect -24285 -2714 -24030 -2709
rect -24285 -2798 -24251 -2714
rect -24217 -2803 -24201 -2769
rect -23825 -2803 -23809 -2769
rect -24285 -2849 -24251 -2833
rect -23725 -2813 -23675 -2593
rect -23632 -2641 -23616 -2607
rect -23422 -2641 -23404 -2607
rect -22398 -2631 -22364 -2615
rect -22302 -2425 -22268 -2409
rect -22302 -2631 -22268 -2621
rect -22206 -2419 -22172 -2409
rect -22206 -2631 -22172 -2615
rect -22110 -2425 -22076 -2409
rect -22110 -2631 -22076 -2621
rect -22014 -2419 -21980 -2409
rect -22014 -2631 -21980 -2615
rect -21918 -2425 -21884 -2409
rect -21918 -2631 -21884 -2621
rect -21822 -2419 -21788 -2409
rect -21822 -2631 -21788 -2615
rect -21705 -2593 -21689 -2367
rect -19964 -2367 -19914 -2350
rect -19871 -2353 -19861 -2319
rect -19665 -2353 -19649 -2319
rect -18908 -2347 -18892 -2300
rect -18323 -2347 -18299 -2300
rect -21612 -2449 -21596 -2415
rect -21402 -2449 -21384 -2415
rect -20668 -2419 -20634 -2409
rect -21612 -2545 -21602 -2511
rect -21406 -2545 -21390 -2511
rect -22349 -2709 -22332 -2674
rect -22298 -2709 -22282 -2674
rect -22060 -2680 -22043 -2674
rect -22248 -2709 -22043 -2680
rect -22009 -2709 -21993 -2674
rect -23632 -2803 -23616 -2769
rect -23440 -2803 -23424 -2769
rect -23725 -2847 -23709 -2813
rect -23725 -2863 -23675 -2847
rect -23632 -2891 -23616 -2857
rect -23440 -2891 -23424 -2857
rect -22349 -2915 -22306 -2709
rect -22248 -2714 -21993 -2709
rect -22248 -2798 -22214 -2714
rect -22180 -2803 -22164 -2769
rect -21788 -2803 -21772 -2769
rect -22248 -2849 -22214 -2833
rect -21705 -2813 -21655 -2593
rect -21612 -2641 -21596 -2607
rect -21402 -2641 -21384 -2607
rect -20668 -2631 -20634 -2615
rect -20572 -2425 -20538 -2409
rect -20572 -2631 -20538 -2621
rect -20476 -2419 -20442 -2409
rect -20476 -2631 -20442 -2615
rect -20380 -2425 -20346 -2409
rect -20380 -2631 -20346 -2621
rect -20284 -2419 -20250 -2409
rect -20284 -2631 -20250 -2615
rect -20188 -2425 -20154 -2409
rect -20188 -2631 -20154 -2621
rect -20092 -2419 -20058 -2409
rect -20092 -2631 -20058 -2615
rect -19964 -2593 -19948 -2367
rect -18185 -2367 -18135 -2350
rect -18092 -2353 -18082 -2319
rect -17886 -2353 -17870 -2319
rect -19871 -2449 -19855 -2415
rect -19661 -2449 -19643 -2415
rect -18908 -2419 -18874 -2409
rect -19871 -2545 -19861 -2511
rect -19665 -2545 -19649 -2511
rect -20619 -2709 -20602 -2674
rect -20568 -2709 -20552 -2674
rect -20330 -2680 -20313 -2674
rect -20518 -2709 -20313 -2680
rect -20279 -2709 -20263 -2674
rect -21612 -2803 -21596 -2769
rect -21420 -2803 -21404 -2769
rect -21705 -2847 -21689 -2813
rect -21705 -2863 -21655 -2847
rect -21612 -2891 -21596 -2857
rect -21420 -2891 -21404 -2857
rect -20619 -2915 -20576 -2709
rect -20518 -2714 -20263 -2709
rect -20518 -2798 -20484 -2714
rect -20450 -2803 -20434 -2769
rect -20058 -2803 -20042 -2769
rect -20518 -2849 -20484 -2833
rect -19964 -2813 -19914 -2593
rect -19871 -2641 -19855 -2607
rect -19661 -2641 -19643 -2607
rect -18908 -2631 -18874 -2615
rect -18812 -2425 -18778 -2409
rect -18812 -2631 -18778 -2621
rect -18716 -2419 -18682 -2409
rect -18716 -2631 -18682 -2615
rect -18620 -2425 -18586 -2409
rect -18620 -2631 -18586 -2621
rect -18524 -2419 -18490 -2409
rect -18524 -2631 -18490 -2615
rect -18428 -2425 -18394 -2409
rect -18428 -2631 -18394 -2621
rect -18332 -2419 -18298 -2409
rect -18332 -2631 -18298 -2615
rect -18185 -2593 -18169 -2367
rect -18092 -2449 -18076 -2415
rect -17882 -2449 -17864 -2415
rect -18092 -2545 -18082 -2511
rect -17886 -2545 -17870 -2511
rect -18859 -2709 -18842 -2674
rect -18808 -2709 -18792 -2674
rect -18570 -2680 -18553 -2674
rect -18758 -2709 -18553 -2680
rect -18519 -2709 -18503 -2674
rect -19871 -2803 -19855 -2769
rect -19679 -2803 -19663 -2769
rect -19964 -2847 -19948 -2813
rect -19964 -2863 -19914 -2847
rect -19871 -2891 -19855 -2857
rect -19679 -2891 -19663 -2857
rect -18859 -2915 -18816 -2709
rect -18758 -2714 -18503 -2709
rect -18758 -2798 -18724 -2714
rect -18690 -2803 -18674 -2769
rect -18298 -2803 -18282 -2769
rect -18758 -2849 -18724 -2833
rect -18185 -2813 -18135 -2593
rect -18092 -2641 -18076 -2607
rect -17882 -2641 -17864 -2607
rect -18092 -2803 -18076 -2769
rect -17900 -2803 -17884 -2769
rect -18185 -2847 -18169 -2813
rect 7333 -2813 7372 -2062
rect 7298 -2826 7372 -2813
rect 7298 -2842 7406 -2826
rect 7756 -2050 7790 -2034
rect 7756 -2842 7790 -2826
rect 8246 -2050 8354 -2034
rect 8246 -2062 8320 -2050
rect 8281 -2813 8320 -2062
rect 8246 -2826 8320 -2813
rect 8246 -2842 8354 -2826
rect 8704 -2050 8738 -2034
rect 8704 -2842 8738 -2826
rect 9182 -2050 9290 -2034
rect 9182 -2062 9256 -2050
rect 9217 -2813 9256 -2062
rect 9182 -2826 9256 -2813
rect 9182 -2842 9290 -2826
rect 9640 -2050 9674 -2034
rect 9640 -2842 9674 -2826
rect 10113 -2050 10221 -2034
rect 10113 -2062 10187 -2050
rect 10148 -2813 10187 -2062
rect 10113 -2826 10187 -2813
rect 10113 -2842 10221 -2826
rect 10571 -2050 10605 -2034
rect 10571 -2842 10605 -2826
rect 11040 -2050 11148 -2034
rect 11040 -2062 11114 -2050
rect 11075 -2813 11114 -2062
rect 11040 -2826 11114 -2813
rect 11040 -2842 11148 -2826
rect 11498 -2050 11532 -2034
rect 11783 -2376 12203 -2356
rect 11783 -2427 11811 -2376
rect 12168 -2427 12203 -2376
rect 11783 -2446 12203 -2427
rect 11785 -2531 11819 -2446
rect 11785 -2779 11819 -2763
rect 11881 -2531 11915 -2515
rect 11881 -2779 11915 -2763
rect 11977 -2531 12011 -2446
rect 11977 -2779 12011 -2763
rect 12073 -2531 12107 -2515
rect 12073 -2779 12107 -2763
rect 12169 -2531 12203 -2446
rect 12169 -2779 12203 -2763
rect 12265 -2531 12299 -2515
rect 12265 -2779 12299 -2763
rect 12361 -2531 12395 -2515
rect 12361 -2779 12395 -2763
rect 12457 -2531 12491 -2515
rect 12457 -2779 12491 -2763
rect 12553 -2531 12587 -2515
rect 12553 -2779 12587 -2763
rect 12649 -2531 12683 -2515
rect 12649 -2779 12683 -2763
rect 12745 -2531 12779 -2515
rect 12970 -2597 12986 -2563
rect 13077 -2597 13093 -2563
rect 12745 -2779 12779 -2763
rect 12826 -2683 12876 -2666
rect 12919 -2669 12929 -2635
rect 13125 -2669 13141 -2635
rect 11498 -2842 11532 -2826
rect -18185 -2863 -18135 -2847
rect -18092 -2891 -18076 -2857
rect -17900 -2891 -17884 -2857
rect 12154 -2859 12170 -2825
rect 12204 -2859 12220 -2825
rect 12826 -2909 12842 -2683
rect 12919 -2765 12935 -2731
rect 13129 -2765 13147 -2731
rect 12919 -2861 12929 -2827
rect 13125 -2861 13141 -2827
rect -24386 -2931 -24251 -2915
rect -24386 -2966 -24285 -2931
rect -22349 -2931 -22214 -2915
rect -24386 -2982 -24251 -2966
rect -24217 -2995 -24201 -2961
rect -23825 -2995 -23809 -2961
rect -23613 -2993 -23597 -2959
rect -23465 -2993 -23449 -2959
rect -22349 -2966 -22248 -2931
rect -20619 -2931 -20484 -2915
rect -22349 -2982 -22214 -2966
rect -22180 -2995 -22164 -2961
rect -21788 -2995 -21772 -2961
rect -21593 -2993 -21577 -2959
rect -21445 -2993 -21429 -2959
rect -20619 -2966 -20518 -2931
rect -18859 -2931 -18724 -2915
rect -20619 -2982 -20484 -2966
rect -20450 -2995 -20434 -2961
rect -20058 -2995 -20042 -2961
rect -19852 -2993 -19836 -2959
rect -19704 -2993 -19688 -2959
rect -18859 -2966 -18758 -2931
rect -18859 -2982 -18724 -2966
rect -18690 -2995 -18674 -2961
rect -18298 -2995 -18282 -2961
rect -18073 -2993 -18057 -2959
rect -17925 -2993 -17909 -2959
rect 7298 -2978 7406 -2962
rect 7298 -2991 7372 -2978
rect -24213 -3067 -24186 -3033
rect -23851 -3067 -23813 -3033
rect -22176 -3067 -22149 -3033
rect -21814 -3067 -21776 -3033
rect -20446 -3067 -20419 -3033
rect -20084 -3067 -20046 -3033
rect -18686 -3067 -18659 -3033
rect -18324 -3067 -18286 -3033
rect 7333 -3742 7372 -2991
rect 7298 -3754 7372 -3742
rect 7298 -3770 7406 -3754
rect 7756 -2978 7790 -2962
rect 7756 -3770 7790 -3754
rect 8246 -2978 8354 -2962
rect 8246 -2991 8320 -2978
rect 8281 -3742 8320 -2991
rect 8246 -3754 8320 -3742
rect 8246 -3770 8354 -3754
rect 8704 -2978 8738 -2962
rect 8704 -3770 8738 -3754
rect 9182 -2978 9290 -2962
rect 9182 -2991 9256 -2978
rect 9217 -3742 9256 -2991
rect 9182 -3754 9256 -3742
rect 9182 -3770 9290 -3754
rect 9640 -2978 9674 -2962
rect 9640 -3770 9674 -3754
rect 10113 -2977 10221 -2961
rect 10113 -2990 10187 -2977
rect 10148 -3741 10187 -2990
rect 10113 -3753 10187 -3741
rect 10113 -3769 10221 -3753
rect 10571 -2977 10605 -2961
rect 10571 -3769 10605 -3753
rect 11040 -2978 11148 -2962
rect 11040 -2991 11114 -2978
rect 11075 -3742 11114 -2991
rect 11040 -3754 11114 -3742
rect 7298 -3773 7403 -3770
rect 8246 -3773 8351 -3770
rect 9182 -3773 9287 -3770
rect 10113 -3772 10218 -3769
rect 11040 -3770 11148 -3754
rect 11498 -2978 11532 -2962
rect 12297 -2964 12313 -2930
rect 12347 -2964 12363 -2930
rect 12169 -3020 12203 -3004
rect 12169 -3268 12203 -3196
rect 12265 -3020 12299 -3004
rect 12265 -3212 12299 -3196
rect 12361 -3020 12395 -3004
rect 12826 -3129 12876 -2909
rect 12919 -2957 12935 -2923
rect 13129 -2957 13147 -2923
rect 12919 -3119 12935 -3085
rect 13111 -3119 13127 -3085
rect 12826 -3163 12842 -3129
rect 12826 -3179 12876 -3163
rect 12361 -3268 12395 -3196
rect 12919 -3207 12935 -3173
rect 13111 -3207 13127 -3173
rect 12157 -3279 12407 -3268
rect 12157 -3340 12183 -3279
rect 12382 -3340 12407 -3279
rect 12938 -3309 12954 -3275
rect 13086 -3309 13102 -3275
rect 12157 -3352 12407 -3340
rect 11498 -3770 11532 -3754
rect 11040 -3773 11145 -3770
rect -20649 -3827 -19439 -3799
rect -20649 -3899 -20603 -3827
rect -19481 -3899 -19439 -3827
rect -20649 -3925 -19439 -3899
rect -19090 -3827 -17880 -3799
rect -19090 -3899 -19044 -3827
rect -17922 -3899 -17880 -3827
rect -19090 -3925 -17880 -3899
rect -17358 -3827 -16148 -3799
rect -17358 -3899 -17312 -3827
rect -16190 -3899 -16148 -3827
rect -17358 -3925 -16148 -3899
rect -15799 -3827 -14589 -3799
rect -15799 -3899 -15753 -3827
rect -14631 -3899 -14589 -3827
rect -15799 -3925 -14589 -3899
rect -14067 -3827 -12857 -3799
rect -14067 -3899 -14021 -3827
rect -12899 -3899 -12857 -3827
rect -14067 -3925 -12857 -3899
rect -12508 -3827 -11298 -3799
rect -12508 -3899 -12462 -3827
rect -11340 -3899 -11298 -3827
rect -12508 -3925 -11298 -3899
rect -10776 -3827 -9566 -3799
rect -10776 -3899 -10730 -3827
rect -9608 -3899 -9566 -3827
rect -10776 -3925 -9566 -3899
rect -9217 -3827 -8007 -3799
rect -9217 -3899 -9171 -3827
rect -8049 -3899 -8007 -3827
rect -9217 -3925 -8007 -3899
rect -20725 -3996 -20691 -3980
rect -23537 -4093 -23521 -4059
rect -23430 -4093 -23414 -4059
rect -21799 -4093 -21783 -4059
rect -21692 -4093 -21676 -4059
rect -24384 -4159 -24368 -4112
rect -23799 -4159 -23775 -4112
rect -23681 -4179 -23631 -4162
rect -23588 -4165 -23578 -4131
rect -23382 -4165 -23366 -4131
rect -22648 -4159 -22632 -4112
rect -22063 -4159 -22039 -4112
rect -24384 -4231 -24350 -4221
rect -24384 -4443 -24350 -4427
rect -24288 -4237 -24254 -4221
rect -24288 -4443 -24254 -4433
rect -24192 -4231 -24158 -4221
rect -24192 -4443 -24158 -4427
rect -24096 -4237 -24062 -4221
rect -24096 -4443 -24062 -4433
rect -24000 -4231 -23966 -4221
rect -24000 -4443 -23966 -4427
rect -23904 -4237 -23870 -4221
rect -23904 -4443 -23870 -4433
rect -23808 -4231 -23774 -4221
rect -23808 -4443 -23774 -4427
rect -23681 -4405 -23665 -4179
rect -21943 -4179 -21893 -4162
rect -21850 -4165 -21840 -4131
rect -21644 -4165 -21628 -4131
rect -23588 -4261 -23572 -4227
rect -23378 -4261 -23360 -4227
rect -22648 -4231 -22614 -4221
rect -23588 -4357 -23578 -4323
rect -23382 -4357 -23366 -4323
rect -24335 -4521 -24318 -4486
rect -24284 -4521 -24268 -4486
rect -24046 -4492 -24029 -4486
rect -24234 -4521 -24029 -4492
rect -23995 -4521 -23979 -4486
rect -24335 -4727 -24292 -4521
rect -24234 -4526 -23979 -4521
rect -24234 -4610 -24200 -4526
rect -24166 -4615 -24150 -4581
rect -23774 -4615 -23758 -4581
rect -24234 -4661 -24200 -4645
rect -23681 -4625 -23631 -4405
rect -23588 -4453 -23572 -4419
rect -23378 -4453 -23360 -4419
rect -22648 -4443 -22614 -4427
rect -22552 -4237 -22518 -4221
rect -22552 -4443 -22518 -4433
rect -22456 -4231 -22422 -4221
rect -22456 -4443 -22422 -4427
rect -22360 -4237 -22326 -4221
rect -22360 -4443 -22326 -4433
rect -22264 -4231 -22230 -4221
rect -22264 -4443 -22230 -4427
rect -22168 -4237 -22134 -4221
rect -22168 -4443 -22134 -4433
rect -22072 -4231 -22038 -4221
rect -22072 -4443 -22038 -4427
rect -21943 -4405 -21927 -4179
rect -21850 -4261 -21834 -4227
rect -21640 -4261 -21622 -4227
rect -21850 -4357 -21840 -4323
rect -21644 -4357 -21628 -4323
rect -22599 -4521 -22582 -4486
rect -22548 -4521 -22532 -4486
rect -22310 -4492 -22293 -4486
rect -22498 -4521 -22293 -4492
rect -22259 -4521 -22243 -4486
rect -23588 -4615 -23572 -4581
rect -23396 -4615 -23380 -4581
rect -23681 -4659 -23665 -4625
rect -23681 -4675 -23631 -4659
rect -23588 -4703 -23572 -4669
rect -23396 -4703 -23380 -4669
rect -22599 -4727 -22556 -4521
rect -22498 -4526 -22243 -4521
rect -22498 -4610 -22464 -4526
rect -22430 -4615 -22414 -4581
rect -22038 -4615 -22022 -4581
rect -22498 -4661 -22464 -4645
rect -21943 -4625 -21893 -4405
rect -21850 -4453 -21834 -4419
rect -21640 -4453 -21622 -4419
rect -21850 -4615 -21834 -4581
rect -21658 -4615 -21642 -4581
rect -20725 -4583 -20691 -4522
rect -20637 -3996 -20603 -3980
rect -20637 -4538 -20603 -4522
rect -20541 -3996 -20507 -3980
rect -20541 -4538 -20507 -4522
rect -20445 -3996 -20411 -3980
rect -20445 -4538 -20411 -4522
rect -20349 -3996 -20315 -3980
rect -20349 -4538 -20315 -4522
rect -20253 -3996 -20219 -3980
rect -20253 -4538 -20219 -4522
rect -20157 -3996 -20123 -3980
rect -20157 -4538 -20123 -4522
rect -20061 -3996 -20027 -3980
rect -20061 -4565 -20027 -4522
rect -19965 -3996 -19931 -3980
rect -19965 -4538 -19931 -4522
rect -19869 -3996 -19835 -3980
rect -19869 -4538 -19835 -4522
rect -19773 -3996 -19739 -3980
rect -19773 -4538 -19739 -4522
rect -19677 -3996 -19643 -3980
rect -19677 -4538 -19643 -4522
rect -19581 -3996 -19547 -3980
rect -19581 -4538 -19547 -4522
rect -19485 -3996 -19451 -3980
rect -19485 -4538 -19451 -4522
rect -19397 -3996 -19363 -3980
rect -20725 -4593 -20123 -4583
rect -21943 -4659 -21927 -4625
rect -21943 -4675 -21893 -4659
rect -20890 -4622 -20780 -4597
rect -21850 -4703 -21834 -4669
rect -21658 -4703 -21642 -4669
rect -24335 -4743 -24200 -4727
rect -24335 -4778 -24234 -4743
rect -22599 -4743 -22464 -4727
rect -24335 -4794 -24200 -4778
rect -24166 -4807 -24150 -4773
rect -23774 -4807 -23758 -4773
rect -23569 -4805 -23553 -4771
rect -23421 -4805 -23405 -4771
rect -22599 -4778 -22498 -4743
rect -20890 -4732 -20854 -4622
rect -20807 -4732 -20780 -4622
rect -22599 -4794 -22464 -4778
rect -22430 -4807 -22414 -4773
rect -22038 -4807 -22022 -4773
rect -21831 -4805 -21815 -4771
rect -21683 -4805 -21667 -4771
rect -24162 -4879 -24135 -4845
rect -23800 -4879 -23762 -4845
rect -22426 -4879 -22399 -4845
rect -22064 -4879 -22026 -4845
rect -20890 -5225 -20780 -4732
rect -20725 -4638 -20269 -4593
rect -20139 -4638 -20123 -4593
rect -20725 -4652 -20123 -4638
rect -20725 -5036 -20691 -4652
rect -20589 -4723 -20368 -4696
rect -20589 -4776 -20539 -4723
rect -20406 -4776 -20368 -4723
rect -20589 -4914 -20368 -4776
rect -20589 -4959 -20544 -4914
rect -20414 -4959 -20368 -4914
rect -20589 -4986 -20368 -4959
rect -20288 -4922 -20123 -4652
rect -20288 -4967 -20261 -4922
rect -20131 -4967 -20123 -4922
rect -20288 -4984 -20123 -4967
rect -20077 -4865 -20011 -4565
rect -19397 -4580 -19363 -4522
rect -19965 -4598 -19363 -4580
rect -19965 -4643 -19938 -4598
rect -19808 -4643 -19363 -4598
rect -19965 -4657 -19363 -4643
rect -19166 -3996 -19132 -3980
rect -19166 -4583 -19132 -4522
rect -19078 -3996 -19044 -3980
rect -19078 -4538 -19044 -4522
rect -18982 -3996 -18948 -3980
rect -18982 -4538 -18948 -4522
rect -18886 -3996 -18852 -3980
rect -18886 -4538 -18852 -4522
rect -18790 -3996 -18756 -3980
rect -18790 -4538 -18756 -4522
rect -18694 -3996 -18660 -3980
rect -18694 -4538 -18660 -4522
rect -18598 -3996 -18564 -3980
rect -18598 -4538 -18564 -4522
rect -18502 -3996 -18468 -3980
rect -18502 -4565 -18468 -4522
rect -18406 -3996 -18372 -3980
rect -18406 -4538 -18372 -4522
rect -18310 -3996 -18276 -3980
rect -18310 -4538 -18276 -4522
rect -18214 -3996 -18180 -3980
rect -18214 -4538 -18180 -4522
rect -18118 -3996 -18084 -3980
rect -18118 -4538 -18084 -4522
rect -18022 -3996 -17988 -3980
rect -18022 -4538 -17988 -4522
rect -17926 -3996 -17892 -3980
rect -17926 -4538 -17892 -4522
rect -17838 -3996 -17804 -3980
rect -19166 -4593 -18564 -4583
rect -19166 -4638 -18710 -4593
rect -18580 -4638 -18564 -4593
rect -19166 -4652 -18564 -4638
rect -19965 -4715 -19788 -4657
rect -19965 -4768 -19933 -4715
rect -19819 -4768 -19788 -4715
rect -19965 -4797 -19788 -4768
rect -19716 -4716 -19601 -4698
rect -19716 -4784 -19699 -4716
rect -19619 -4784 -19601 -4716
rect -19716 -4804 -19601 -4784
rect -20077 -4887 -19437 -4865
rect -20077 -4942 -19517 -4887
rect -19452 -4942 -19437 -4887
rect -20077 -4961 -19437 -4942
rect -20077 -4995 -20011 -4961
rect -20725 -5158 -20691 -5142
rect -20637 -5036 -20603 -5020
rect -20637 -5158 -20603 -5142
rect -20541 -5021 -20507 -5020
rect -20541 -5158 -20507 -5142
rect -20445 -5036 -20411 -5020
rect -20445 -5158 -20411 -5156
rect -20349 -5021 -20315 -5020
rect -20349 -5158 -20315 -5142
rect -20253 -5036 -20219 -5020
rect -20253 -5158 -20219 -5156
rect -20157 -5022 -20123 -5020
rect -20157 -5158 -20123 -5142
rect -20061 -5036 -20027 -4995
rect -20061 -5158 -20027 -5156
rect -19965 -5021 -19931 -5020
rect -19965 -5158 -19931 -5142
rect -19869 -5036 -19835 -5020
rect -19869 -5158 -19835 -5156
rect -19773 -5021 -19739 -5020
rect -19773 -5158 -19739 -5142
rect -19677 -5036 -19643 -5020
rect -19677 -5158 -19643 -5156
rect -19581 -5021 -19547 -5020
rect -19581 -5158 -19547 -5142
rect -19485 -5036 -19451 -5020
rect -19485 -5158 -19451 -5142
rect -19397 -5036 -19363 -4657
rect -19316 -4667 -19207 -4652
rect -19316 -4807 -19297 -4667
rect -19224 -4807 -19207 -4667
rect -19316 -4824 -19207 -4807
rect -19397 -5158 -19363 -5142
rect -19166 -5036 -19132 -4652
rect -19030 -4723 -18809 -4696
rect -19030 -4776 -18980 -4723
rect -18847 -4776 -18809 -4723
rect -19030 -4914 -18809 -4776
rect -19030 -4959 -18985 -4914
rect -18855 -4959 -18809 -4914
rect -19030 -4986 -18809 -4959
rect -18729 -4922 -18564 -4652
rect -18729 -4967 -18702 -4922
rect -18572 -4967 -18564 -4922
rect -18729 -4984 -18564 -4967
rect -18518 -4865 -18452 -4565
rect -17838 -4580 -17804 -4522
rect -18406 -4598 -17804 -4580
rect -18406 -4643 -18379 -4598
rect -18249 -4643 -17804 -4598
rect -17434 -3996 -17400 -3980
rect -17434 -4583 -17400 -4522
rect -17346 -3996 -17312 -3980
rect -17346 -4538 -17312 -4522
rect -17250 -3996 -17216 -3980
rect -17250 -4538 -17216 -4522
rect -17154 -3996 -17120 -3980
rect -17154 -4538 -17120 -4522
rect -17058 -3996 -17024 -3980
rect -17058 -4538 -17024 -4522
rect -16962 -3996 -16928 -3980
rect -16962 -4538 -16928 -4522
rect -16866 -3996 -16832 -3980
rect -16866 -4538 -16832 -4522
rect -16770 -3996 -16736 -3980
rect -16770 -4565 -16736 -4522
rect -16674 -3996 -16640 -3980
rect -16674 -4538 -16640 -4522
rect -16578 -3996 -16544 -3980
rect -16578 -4538 -16544 -4522
rect -16482 -3996 -16448 -3980
rect -16482 -4538 -16448 -4522
rect -16386 -3996 -16352 -3980
rect -16386 -4538 -16352 -4522
rect -16290 -3996 -16256 -3980
rect -16290 -4538 -16256 -4522
rect -16194 -3996 -16160 -3980
rect -16194 -4538 -16160 -4522
rect -16106 -3996 -16072 -3980
rect -17434 -4593 -16832 -4583
rect -18406 -4657 -17804 -4643
rect -18406 -4715 -18229 -4657
rect -18406 -4768 -18374 -4715
rect -18260 -4768 -18229 -4715
rect -18406 -4797 -18229 -4768
rect -18157 -4716 -18042 -4698
rect -18157 -4784 -18140 -4716
rect -18060 -4784 -18042 -4716
rect -18157 -4804 -18042 -4784
rect -18518 -4887 -17878 -4865
rect -18518 -4942 -17958 -4887
rect -17893 -4942 -17878 -4887
rect -18518 -4961 -17878 -4942
rect -18518 -4995 -18452 -4961
rect -19166 -5158 -19132 -5142
rect -19078 -5036 -19044 -5020
rect -19078 -5158 -19044 -5142
rect -18982 -5021 -18948 -5020
rect -18982 -5158 -18948 -5142
rect -18886 -5036 -18852 -5020
rect -18886 -5158 -18852 -5156
rect -18790 -5021 -18756 -5020
rect -18790 -5158 -18756 -5142
rect -18694 -5036 -18660 -5020
rect -18694 -5158 -18660 -5156
rect -18598 -5022 -18564 -5020
rect -18598 -5158 -18564 -5142
rect -18502 -5036 -18468 -4995
rect -18502 -5158 -18468 -5156
rect -18406 -5021 -18372 -5020
rect -18406 -5158 -18372 -5142
rect -18310 -5036 -18276 -5020
rect -18310 -5158 -18276 -5156
rect -18214 -5021 -18180 -5020
rect -18214 -5158 -18180 -5142
rect -18118 -5036 -18084 -5020
rect -18118 -5158 -18084 -5156
rect -18022 -5021 -17988 -5020
rect -18022 -5158 -17988 -5142
rect -17926 -5036 -17892 -5020
rect -17926 -5158 -17892 -5142
rect -17838 -5036 -17804 -4657
rect -17581 -4622 -17496 -4599
rect -17581 -4732 -17563 -4622
rect -17516 -4732 -17496 -4622
rect -17581 -4752 -17496 -4732
rect -17434 -4638 -16978 -4593
rect -16848 -4638 -16832 -4593
rect -17434 -4652 -16832 -4638
rect -17838 -5158 -17804 -5142
rect -17434 -5036 -17400 -4652
rect -17298 -4723 -17077 -4696
rect -17298 -4776 -17248 -4723
rect -17115 -4776 -17077 -4723
rect -17298 -4914 -17077 -4776
rect -17298 -4959 -17253 -4914
rect -17123 -4959 -17077 -4914
rect -17298 -4986 -17077 -4959
rect -16997 -4922 -16832 -4652
rect -16997 -4967 -16970 -4922
rect -16840 -4967 -16832 -4922
rect -16997 -4984 -16832 -4967
rect -16786 -4865 -16720 -4565
rect -16106 -4580 -16072 -4522
rect -16674 -4598 -16072 -4580
rect -16674 -4643 -16647 -4598
rect -16517 -4643 -16072 -4598
rect -16674 -4657 -16072 -4643
rect -15875 -3996 -15841 -3980
rect -15875 -4583 -15841 -4522
rect -15787 -3996 -15753 -3980
rect -15787 -4538 -15753 -4522
rect -15691 -3996 -15657 -3980
rect -15691 -4538 -15657 -4522
rect -15595 -3996 -15561 -3980
rect -15595 -4538 -15561 -4522
rect -15499 -3996 -15465 -3980
rect -15499 -4538 -15465 -4522
rect -15403 -3996 -15369 -3980
rect -15403 -4538 -15369 -4522
rect -15307 -3996 -15273 -3980
rect -15307 -4538 -15273 -4522
rect -15211 -3996 -15177 -3980
rect -15211 -4565 -15177 -4522
rect -15115 -3996 -15081 -3980
rect -15115 -4538 -15081 -4522
rect -15019 -3996 -14985 -3980
rect -15019 -4538 -14985 -4522
rect -14923 -3996 -14889 -3980
rect -14923 -4538 -14889 -4522
rect -14827 -3996 -14793 -3980
rect -14827 -4538 -14793 -4522
rect -14731 -3996 -14697 -3980
rect -14731 -4538 -14697 -4522
rect -14635 -3996 -14601 -3980
rect -14635 -4538 -14601 -4522
rect -14547 -3996 -14513 -3980
rect -15875 -4593 -15273 -4583
rect -15875 -4638 -15419 -4593
rect -15289 -4638 -15273 -4593
rect -15875 -4652 -15273 -4638
rect -16674 -4715 -16497 -4657
rect -16674 -4768 -16642 -4715
rect -16528 -4768 -16497 -4715
rect -16674 -4797 -16497 -4768
rect -16425 -4716 -16310 -4698
rect -16425 -4784 -16408 -4716
rect -16328 -4784 -16310 -4716
rect -16425 -4804 -16310 -4784
rect -16786 -4887 -16146 -4865
rect -16786 -4942 -16226 -4887
rect -16161 -4942 -16146 -4887
rect -16786 -4961 -16146 -4942
rect -16786 -4995 -16720 -4961
rect -17434 -5158 -17400 -5142
rect -17346 -5036 -17312 -5020
rect -17346 -5158 -17312 -5142
rect -17250 -5021 -17216 -5020
rect -17250 -5158 -17216 -5142
rect -17154 -5036 -17120 -5020
rect -17154 -5158 -17120 -5156
rect -17058 -5021 -17024 -5020
rect -17058 -5158 -17024 -5142
rect -16962 -5036 -16928 -5020
rect -16962 -5158 -16928 -5156
rect -16866 -5022 -16832 -5020
rect -16866 -5158 -16832 -5142
rect -16770 -5036 -16736 -4995
rect -16770 -5158 -16736 -5156
rect -16674 -5021 -16640 -5020
rect -16674 -5158 -16640 -5142
rect -16578 -5036 -16544 -5020
rect -16578 -5158 -16544 -5156
rect -16482 -5021 -16448 -5020
rect -16482 -5158 -16448 -5142
rect -16386 -5036 -16352 -5020
rect -16386 -5158 -16352 -5156
rect -16290 -5021 -16256 -5020
rect -16290 -5158 -16256 -5142
rect -16194 -5036 -16160 -5020
rect -16194 -5158 -16160 -5142
rect -16106 -5036 -16072 -4657
rect -16025 -4667 -15916 -4652
rect -16025 -4807 -16006 -4667
rect -15933 -4807 -15916 -4667
rect -16025 -4824 -15916 -4807
rect -16106 -5158 -16072 -5142
rect -15875 -5036 -15841 -4652
rect -15739 -4723 -15518 -4696
rect -15739 -4776 -15689 -4723
rect -15556 -4776 -15518 -4723
rect -15739 -4914 -15518 -4776
rect -15739 -4959 -15694 -4914
rect -15564 -4959 -15518 -4914
rect -15739 -4986 -15518 -4959
rect -15438 -4922 -15273 -4652
rect -15438 -4967 -15411 -4922
rect -15281 -4967 -15273 -4922
rect -15438 -4984 -15273 -4967
rect -15227 -4865 -15161 -4565
rect -14547 -4580 -14513 -4522
rect -15115 -4598 -14513 -4580
rect -15115 -4643 -15088 -4598
rect -14958 -4643 -14513 -4598
rect -14143 -3996 -14109 -3980
rect -14143 -4583 -14109 -4522
rect -14055 -3996 -14021 -3980
rect -14055 -4538 -14021 -4522
rect -13959 -3996 -13925 -3980
rect -13959 -4538 -13925 -4522
rect -13863 -3996 -13829 -3980
rect -13863 -4538 -13829 -4522
rect -13767 -3996 -13733 -3980
rect -13767 -4538 -13733 -4522
rect -13671 -3996 -13637 -3980
rect -13671 -4538 -13637 -4522
rect -13575 -3996 -13541 -3980
rect -13575 -4538 -13541 -4522
rect -13479 -3996 -13445 -3980
rect -13479 -4565 -13445 -4522
rect -13383 -3996 -13349 -3980
rect -13383 -4538 -13349 -4522
rect -13287 -3996 -13253 -3980
rect -13287 -4538 -13253 -4522
rect -13191 -3996 -13157 -3980
rect -13191 -4538 -13157 -4522
rect -13095 -3996 -13061 -3980
rect -13095 -4538 -13061 -4522
rect -12999 -3996 -12965 -3980
rect -12999 -4538 -12965 -4522
rect -12903 -3996 -12869 -3980
rect -12903 -4538 -12869 -4522
rect -12815 -3996 -12781 -3980
rect -14143 -4593 -13541 -4583
rect -15115 -4657 -14513 -4643
rect -15115 -4715 -14938 -4657
rect -15115 -4768 -15083 -4715
rect -14969 -4768 -14938 -4715
rect -15115 -4797 -14938 -4768
rect -14866 -4716 -14751 -4698
rect -14866 -4784 -14849 -4716
rect -14769 -4784 -14751 -4716
rect -14866 -4804 -14751 -4784
rect -15227 -4887 -14587 -4865
rect -15227 -4942 -14667 -4887
rect -14602 -4942 -14587 -4887
rect -15227 -4961 -14587 -4942
rect -15227 -4995 -15161 -4961
rect -15875 -5158 -15841 -5142
rect -15787 -5036 -15753 -5020
rect -15787 -5158 -15753 -5142
rect -15691 -5021 -15657 -5020
rect -15691 -5158 -15657 -5142
rect -15595 -5036 -15561 -5020
rect -15595 -5158 -15561 -5156
rect -15499 -5021 -15465 -5020
rect -15499 -5158 -15465 -5142
rect -15403 -5036 -15369 -5020
rect -15403 -5158 -15369 -5156
rect -15307 -5022 -15273 -5020
rect -15307 -5158 -15273 -5142
rect -15211 -5036 -15177 -4995
rect -15211 -5158 -15177 -5156
rect -15115 -5021 -15081 -5020
rect -15115 -5158 -15081 -5142
rect -15019 -5036 -14985 -5020
rect -15019 -5158 -14985 -5156
rect -14923 -5021 -14889 -5020
rect -14923 -5158 -14889 -5142
rect -14827 -5036 -14793 -5020
rect -14827 -5158 -14793 -5156
rect -14731 -5021 -14697 -5020
rect -14731 -5158 -14697 -5142
rect -14635 -5036 -14601 -5020
rect -14635 -5158 -14601 -5142
rect -14547 -5036 -14513 -4657
rect -14290 -4622 -14205 -4599
rect -14290 -4732 -14272 -4622
rect -14225 -4732 -14205 -4622
rect -14290 -4752 -14205 -4732
rect -14143 -4638 -13687 -4593
rect -13557 -4638 -13541 -4593
rect -14143 -4652 -13541 -4638
rect -14547 -5158 -14513 -5142
rect -14143 -5036 -14109 -4652
rect -14007 -4723 -13786 -4696
rect -14007 -4776 -13957 -4723
rect -13824 -4776 -13786 -4723
rect -14007 -4914 -13786 -4776
rect -14007 -4959 -13962 -4914
rect -13832 -4959 -13786 -4914
rect -14007 -4986 -13786 -4959
rect -13706 -4922 -13541 -4652
rect -13706 -4967 -13679 -4922
rect -13549 -4967 -13541 -4922
rect -13706 -4984 -13541 -4967
rect -13495 -4865 -13429 -4565
rect -12815 -4580 -12781 -4522
rect -13383 -4598 -12781 -4580
rect -13383 -4643 -13356 -4598
rect -13226 -4643 -12781 -4598
rect -13383 -4657 -12781 -4643
rect -12584 -3996 -12550 -3980
rect -12584 -4583 -12550 -4522
rect -12496 -3996 -12462 -3980
rect -12496 -4538 -12462 -4522
rect -12400 -3996 -12366 -3980
rect -12400 -4538 -12366 -4522
rect -12304 -3996 -12270 -3980
rect -12304 -4538 -12270 -4522
rect -12208 -3996 -12174 -3980
rect -12208 -4538 -12174 -4522
rect -12112 -3996 -12078 -3980
rect -12112 -4538 -12078 -4522
rect -12016 -3996 -11982 -3980
rect -12016 -4538 -11982 -4522
rect -11920 -3996 -11886 -3980
rect -11920 -4565 -11886 -4522
rect -11824 -3996 -11790 -3980
rect -11824 -4538 -11790 -4522
rect -11728 -3996 -11694 -3980
rect -11728 -4538 -11694 -4522
rect -11632 -3996 -11598 -3980
rect -11632 -4538 -11598 -4522
rect -11536 -3996 -11502 -3980
rect -11536 -4538 -11502 -4522
rect -11440 -3996 -11406 -3980
rect -11440 -4538 -11406 -4522
rect -11344 -3996 -11310 -3980
rect -11344 -4538 -11310 -4522
rect -11256 -3996 -11222 -3980
rect -12584 -4593 -11982 -4583
rect -12584 -4638 -12128 -4593
rect -11998 -4638 -11982 -4593
rect -12584 -4652 -11982 -4638
rect -13383 -4715 -13206 -4657
rect -13383 -4768 -13351 -4715
rect -13237 -4768 -13206 -4715
rect -13383 -4797 -13206 -4768
rect -13134 -4716 -13019 -4698
rect -13134 -4784 -13117 -4716
rect -13037 -4784 -13019 -4716
rect -13134 -4804 -13019 -4784
rect -13495 -4887 -12855 -4865
rect -13495 -4942 -12935 -4887
rect -12870 -4942 -12855 -4887
rect -13495 -4961 -12855 -4942
rect -13495 -4995 -13429 -4961
rect -14143 -5158 -14109 -5142
rect -14055 -5036 -14021 -5020
rect -14055 -5158 -14021 -5142
rect -13959 -5021 -13925 -5020
rect -13959 -5158 -13925 -5142
rect -13863 -5036 -13829 -5020
rect -13863 -5158 -13829 -5156
rect -13767 -5021 -13733 -5020
rect -13767 -5158 -13733 -5142
rect -13671 -5036 -13637 -5020
rect -13671 -5158 -13637 -5156
rect -13575 -5022 -13541 -5020
rect -13575 -5158 -13541 -5142
rect -13479 -5036 -13445 -4995
rect -13479 -5158 -13445 -5156
rect -13383 -5021 -13349 -5020
rect -13383 -5158 -13349 -5142
rect -13287 -5036 -13253 -5020
rect -13287 -5158 -13253 -5156
rect -13191 -5021 -13157 -5020
rect -13191 -5158 -13157 -5142
rect -13095 -5036 -13061 -5020
rect -13095 -5158 -13061 -5156
rect -12999 -5021 -12965 -5020
rect -12999 -5158 -12965 -5142
rect -12903 -5036 -12869 -5020
rect -12903 -5158 -12869 -5142
rect -12815 -5036 -12781 -4657
rect -12734 -4667 -12625 -4652
rect -12734 -4807 -12715 -4667
rect -12642 -4807 -12625 -4667
rect -12734 -4824 -12625 -4807
rect -12815 -5158 -12781 -5142
rect -12584 -5036 -12550 -4652
rect -12448 -4723 -12227 -4696
rect -12448 -4776 -12398 -4723
rect -12265 -4776 -12227 -4723
rect -12448 -4914 -12227 -4776
rect -12448 -4959 -12403 -4914
rect -12273 -4959 -12227 -4914
rect -12448 -4986 -12227 -4959
rect -12147 -4922 -11982 -4652
rect -12147 -4967 -12120 -4922
rect -11990 -4967 -11982 -4922
rect -12147 -4984 -11982 -4967
rect -11936 -4865 -11870 -4565
rect -11256 -4580 -11222 -4522
rect -11824 -4598 -11222 -4580
rect -11824 -4643 -11797 -4598
rect -11667 -4643 -11222 -4598
rect -10852 -3996 -10818 -3980
rect -10852 -4583 -10818 -4522
rect -10764 -3996 -10730 -3980
rect -10764 -4538 -10730 -4522
rect -10668 -3996 -10634 -3980
rect -10668 -4538 -10634 -4522
rect -10572 -3996 -10538 -3980
rect -10572 -4538 -10538 -4522
rect -10476 -3996 -10442 -3980
rect -10476 -4538 -10442 -4522
rect -10380 -3996 -10346 -3980
rect -10380 -4538 -10346 -4522
rect -10284 -3996 -10250 -3980
rect -10284 -4538 -10250 -4522
rect -10188 -3996 -10154 -3980
rect -10188 -4565 -10154 -4522
rect -10092 -3996 -10058 -3980
rect -10092 -4538 -10058 -4522
rect -9996 -3996 -9962 -3980
rect -9996 -4538 -9962 -4522
rect -9900 -3996 -9866 -3980
rect -9900 -4538 -9866 -4522
rect -9804 -3996 -9770 -3980
rect -9804 -4538 -9770 -4522
rect -9708 -3996 -9674 -3980
rect -9708 -4538 -9674 -4522
rect -9612 -3996 -9578 -3980
rect -9612 -4538 -9578 -4522
rect -9524 -3996 -9490 -3980
rect -10852 -4593 -10250 -4583
rect -11824 -4657 -11222 -4643
rect -11824 -4715 -11647 -4657
rect -11824 -4768 -11792 -4715
rect -11678 -4768 -11647 -4715
rect -11824 -4797 -11647 -4768
rect -11575 -4716 -11460 -4698
rect -11575 -4784 -11558 -4716
rect -11478 -4784 -11460 -4716
rect -11575 -4804 -11460 -4784
rect -11936 -4887 -11296 -4865
rect -11936 -4942 -11376 -4887
rect -11311 -4942 -11296 -4887
rect -11936 -4961 -11296 -4942
rect -11936 -4995 -11870 -4961
rect -12584 -5158 -12550 -5142
rect -12496 -5036 -12462 -5020
rect -12496 -5158 -12462 -5142
rect -12400 -5021 -12366 -5020
rect -12400 -5158 -12366 -5142
rect -12304 -5036 -12270 -5020
rect -12304 -5158 -12270 -5156
rect -12208 -5021 -12174 -5020
rect -12208 -5158 -12174 -5142
rect -12112 -5036 -12078 -5020
rect -12112 -5158 -12078 -5156
rect -12016 -5022 -11982 -5020
rect -12016 -5158 -11982 -5142
rect -11920 -5036 -11886 -4995
rect -11920 -5158 -11886 -5156
rect -11824 -5021 -11790 -5020
rect -11824 -5158 -11790 -5142
rect -11728 -5036 -11694 -5020
rect -11728 -5158 -11694 -5156
rect -11632 -5021 -11598 -5020
rect -11632 -5158 -11598 -5142
rect -11536 -5036 -11502 -5020
rect -11536 -5158 -11502 -5156
rect -11440 -5021 -11406 -5020
rect -11440 -5158 -11406 -5142
rect -11344 -5036 -11310 -5020
rect -11344 -5158 -11310 -5142
rect -11256 -5036 -11222 -4657
rect -10999 -4622 -10914 -4599
rect -10999 -4732 -10981 -4622
rect -10934 -4732 -10914 -4622
rect -10999 -4752 -10914 -4732
rect -10852 -4638 -10396 -4593
rect -10266 -4638 -10250 -4593
rect -10852 -4652 -10250 -4638
rect -11256 -5158 -11222 -5142
rect -10852 -5036 -10818 -4652
rect -10716 -4723 -10495 -4696
rect -10716 -4776 -10666 -4723
rect -10533 -4776 -10495 -4723
rect -10716 -4914 -10495 -4776
rect -10716 -4959 -10671 -4914
rect -10541 -4959 -10495 -4914
rect -10716 -4986 -10495 -4959
rect -10415 -4922 -10250 -4652
rect -10415 -4967 -10388 -4922
rect -10258 -4967 -10250 -4922
rect -10415 -4984 -10250 -4967
rect -10204 -4865 -10138 -4565
rect -9524 -4580 -9490 -4522
rect -10092 -4598 -9490 -4580
rect -10092 -4643 -10065 -4598
rect -9935 -4643 -9490 -4598
rect -10092 -4657 -9490 -4643
rect -9293 -3996 -9259 -3980
rect -9293 -4583 -9259 -4522
rect -9205 -3996 -9171 -3980
rect -9205 -4538 -9171 -4522
rect -9109 -3996 -9075 -3980
rect -9109 -4538 -9075 -4522
rect -9013 -3996 -8979 -3980
rect -9013 -4538 -8979 -4522
rect -8917 -3996 -8883 -3980
rect -8917 -4538 -8883 -4522
rect -8821 -3996 -8787 -3980
rect -8821 -4538 -8787 -4522
rect -8725 -3996 -8691 -3980
rect -8725 -4538 -8691 -4522
rect -8629 -3996 -8595 -3980
rect -8629 -4565 -8595 -4522
rect -8533 -3996 -8499 -3980
rect -8533 -4538 -8499 -4522
rect -8437 -3996 -8403 -3980
rect -8437 -4538 -8403 -4522
rect -8341 -3996 -8307 -3980
rect -8341 -4538 -8307 -4522
rect -8245 -3996 -8211 -3980
rect -8245 -4538 -8211 -4522
rect -8149 -3996 -8115 -3980
rect -8149 -4538 -8115 -4522
rect -8053 -3996 -8019 -3980
rect -8053 -4538 -8019 -4522
rect -7965 -3996 -7931 -3980
rect 7182 -4126 7198 -4092
rect 7232 -4126 7248 -4092
rect 7374 -4126 7390 -4092
rect 7424 -4126 7440 -4092
rect 7566 -4126 7582 -4092
rect 7616 -4126 7632 -4092
rect 7758 -4126 7774 -4092
rect 7808 -4126 7824 -4092
rect 8130 -4126 8146 -4092
rect 8180 -4126 8196 -4092
rect 8322 -4126 8338 -4092
rect 8372 -4126 8388 -4092
rect 8514 -4126 8530 -4092
rect 8564 -4126 8580 -4092
rect 8706 -4126 8722 -4092
rect 8756 -4126 8772 -4092
rect 9066 -4126 9082 -4092
rect 9116 -4126 9132 -4092
rect 9258 -4126 9274 -4092
rect 9308 -4126 9324 -4092
rect 9450 -4126 9466 -4092
rect 9500 -4126 9516 -4092
rect 9642 -4126 9658 -4092
rect 9692 -4126 9708 -4092
rect 9997 -4125 10013 -4091
rect 10047 -4125 10063 -4091
rect 10189 -4125 10205 -4091
rect 10239 -4125 10255 -4091
rect 10381 -4125 10397 -4091
rect 10431 -4125 10447 -4091
rect 10573 -4125 10589 -4091
rect 10623 -4125 10639 -4091
rect 10924 -4126 10940 -4092
rect 10974 -4126 10990 -4092
rect 11116 -4126 11132 -4092
rect 11166 -4126 11182 -4092
rect 11308 -4126 11324 -4092
rect 11358 -4126 11374 -4092
rect 11500 -4126 11516 -4092
rect 11550 -4126 11566 -4092
rect 7150 -4185 7184 -4169
rect 7246 -4180 7280 -4169
rect 7150 -4499 7184 -4483
rect 7246 -4499 7280 -4483
rect 7342 -4185 7376 -4169
rect 7342 -4499 7376 -4483
rect 7438 -4180 7472 -4169
rect 7534 -4185 7568 -4169
rect 7438 -4499 7472 -4483
rect 7534 -4499 7568 -4483
rect 7630 -4180 7664 -4169
rect 7726 -4185 7760 -4169
rect 7630 -4499 7664 -4483
rect 7726 -4499 7760 -4483
rect 7822 -4180 7856 -4169
rect 7918 -4185 7952 -4169
rect 7822 -4499 7856 -4483
rect 7918 -4499 7952 -4483
rect 8098 -4185 8132 -4169
rect 8194 -4180 8228 -4169
rect 8098 -4499 8132 -4483
rect 8194 -4499 8228 -4483
rect 8290 -4185 8324 -4169
rect 8290 -4499 8324 -4483
rect 8386 -4180 8420 -4169
rect 8482 -4185 8516 -4169
rect 8386 -4499 8420 -4483
rect 8482 -4499 8516 -4483
rect 8578 -4180 8612 -4169
rect 8674 -4185 8708 -4169
rect 8578 -4499 8612 -4483
rect 8674 -4499 8708 -4483
rect 8770 -4180 8804 -4169
rect 8866 -4185 8900 -4169
rect 8770 -4499 8804 -4483
rect 8866 -4499 8900 -4483
rect 9034 -4185 9068 -4169
rect 9130 -4180 9164 -4169
rect 9034 -4499 9068 -4483
rect 9130 -4499 9164 -4483
rect 9226 -4185 9260 -4169
rect 9226 -4499 9260 -4483
rect 9322 -4180 9356 -4169
rect 9418 -4185 9452 -4169
rect 9322 -4499 9356 -4483
rect 9418 -4499 9452 -4483
rect 9514 -4180 9548 -4169
rect 9610 -4185 9644 -4169
rect 9514 -4499 9548 -4483
rect 9610 -4499 9644 -4483
rect 9706 -4180 9740 -4169
rect 9802 -4185 9836 -4169
rect 9706 -4499 9740 -4483
rect 9802 -4499 9836 -4483
rect 9965 -4184 9999 -4168
rect 10061 -4179 10095 -4168
rect 9965 -4498 9999 -4482
rect 10061 -4498 10095 -4482
rect 10157 -4184 10191 -4168
rect 10157 -4498 10191 -4482
rect 10253 -4179 10287 -4168
rect 10349 -4184 10383 -4168
rect 10253 -4498 10287 -4482
rect 10349 -4498 10383 -4482
rect 10445 -4179 10479 -4168
rect 10541 -4184 10575 -4168
rect 10445 -4498 10479 -4482
rect 10541 -4498 10575 -4482
rect 10637 -4179 10671 -4168
rect 10733 -4184 10767 -4168
rect 10637 -4498 10671 -4482
rect 10733 -4498 10767 -4482
rect 10892 -4185 10926 -4169
rect 10988 -4180 11022 -4169
rect 10892 -4499 10926 -4483
rect 10988 -4499 11022 -4483
rect 11084 -4185 11118 -4169
rect 11084 -4499 11118 -4483
rect 11180 -4180 11214 -4169
rect 11276 -4185 11310 -4169
rect 11180 -4499 11214 -4483
rect 11276 -4499 11310 -4483
rect 11372 -4180 11406 -4169
rect 11468 -4185 11502 -4169
rect 11372 -4499 11406 -4483
rect 11468 -4499 11502 -4483
rect 11564 -4180 11598 -4169
rect 11660 -4185 11694 -4169
rect 11564 -4499 11598 -4483
rect 11660 -4499 11694 -4483
rect -9293 -4593 -8691 -4583
rect -9293 -4638 -8837 -4593
rect -8707 -4638 -8691 -4593
rect -9293 -4652 -8691 -4638
rect -10092 -4715 -9915 -4657
rect -10092 -4768 -10060 -4715
rect -9946 -4768 -9915 -4715
rect -10092 -4797 -9915 -4768
rect -9843 -4716 -9728 -4698
rect -9843 -4784 -9826 -4716
rect -9746 -4784 -9728 -4716
rect -9843 -4804 -9728 -4784
rect -10204 -4887 -9564 -4865
rect -10204 -4942 -9644 -4887
rect -9579 -4942 -9564 -4887
rect -10204 -4961 -9564 -4942
rect -10204 -4995 -10138 -4961
rect -10852 -5158 -10818 -5142
rect -10764 -5036 -10730 -5020
rect -10764 -5158 -10730 -5142
rect -10668 -5021 -10634 -5020
rect -10668 -5158 -10634 -5142
rect -10572 -5036 -10538 -5020
rect -10572 -5158 -10538 -5156
rect -10476 -5021 -10442 -5020
rect -10476 -5158 -10442 -5142
rect -10380 -5036 -10346 -5020
rect -10380 -5158 -10346 -5156
rect -10284 -5022 -10250 -5020
rect -10284 -5158 -10250 -5142
rect -10188 -5036 -10154 -4995
rect -10188 -5158 -10154 -5156
rect -10092 -5021 -10058 -5020
rect -10092 -5158 -10058 -5142
rect -9996 -5036 -9962 -5020
rect -9996 -5158 -9962 -5156
rect -9900 -5021 -9866 -5020
rect -9900 -5158 -9866 -5142
rect -9804 -5036 -9770 -5020
rect -9804 -5158 -9770 -5156
rect -9708 -5021 -9674 -5020
rect -9708 -5158 -9674 -5142
rect -9612 -5036 -9578 -5020
rect -9612 -5158 -9578 -5142
rect -9524 -5036 -9490 -4657
rect -9443 -4667 -9334 -4652
rect -9443 -4807 -9424 -4667
rect -9351 -4807 -9334 -4667
rect -9443 -4824 -9334 -4807
rect -9524 -5158 -9490 -5142
rect -9293 -5036 -9259 -4652
rect -9157 -4723 -8936 -4696
rect -9157 -4776 -9107 -4723
rect -8974 -4776 -8936 -4723
rect -9157 -4914 -8936 -4776
rect -9157 -4959 -9112 -4914
rect -8982 -4959 -8936 -4914
rect -9157 -4986 -8936 -4959
rect -8856 -4922 -8691 -4652
rect -8856 -4967 -8829 -4922
rect -8699 -4967 -8691 -4922
rect -8856 -4984 -8691 -4967
rect -8645 -4865 -8579 -4565
rect -7965 -4580 -7931 -4522
rect -8533 -4598 -7931 -4580
rect 7373 -4587 7389 -4552
rect 7677 -4587 7703 -4552
rect 8321 -4587 8337 -4552
rect 8625 -4587 8651 -4552
rect 9257 -4587 9273 -4552
rect 9561 -4587 9587 -4552
rect 10188 -4586 10204 -4551
rect 10492 -4586 10518 -4551
rect 11115 -4587 11131 -4552
rect 11419 -4587 11445 -4552
rect -8533 -4643 -8506 -4598
rect -8376 -4643 -7931 -4598
rect -8533 -4657 -7931 -4643
rect -8533 -4715 -8356 -4657
rect -8533 -4768 -8501 -4715
rect -8387 -4768 -8356 -4715
rect -8533 -4797 -8356 -4768
rect -8284 -4716 -8169 -4698
rect -8284 -4784 -8267 -4716
rect -8187 -4784 -8169 -4716
rect -8284 -4804 -8169 -4784
rect -8645 -4887 -8005 -4865
rect -8645 -4942 -8085 -4887
rect -8020 -4942 -8005 -4887
rect -8645 -4961 -8005 -4942
rect -8645 -4995 -8579 -4961
rect -9293 -5158 -9259 -5142
rect -9205 -5036 -9171 -5020
rect -9205 -5158 -9171 -5142
rect -9109 -5021 -9075 -5020
rect -9109 -5158 -9075 -5142
rect -9013 -5036 -8979 -5020
rect -9013 -5158 -8979 -5156
rect -8917 -5021 -8883 -5020
rect -8917 -5158 -8883 -5142
rect -8821 -5036 -8787 -5020
rect -8821 -5158 -8787 -5156
rect -8725 -5022 -8691 -5020
rect -8725 -5158 -8691 -5142
rect -8629 -5036 -8595 -4995
rect -8629 -5158 -8595 -5156
rect -8533 -5021 -8499 -5020
rect -8533 -5158 -8499 -5142
rect -8437 -5036 -8403 -5020
rect -8437 -5158 -8403 -5156
rect -8341 -5021 -8307 -5020
rect -8341 -5158 -8307 -5142
rect -8245 -5036 -8211 -5020
rect -8245 -5158 -8211 -5156
rect -8149 -5021 -8115 -5020
rect -8149 -5158 -8115 -5142
rect -8053 -5036 -8019 -5020
rect -8053 -5158 -8019 -5142
rect -7965 -5036 -7931 -4657
rect 5705 -5007 5721 -4973
rect 5812 -5007 5828 -4973
rect 6145 -5007 6161 -4973
rect 6252 -5007 6268 -4973
rect 6585 -5007 6601 -4973
rect 6692 -5007 6708 -4973
rect -7965 -5158 -7931 -5142
rect 5561 -5093 5611 -5076
rect 5654 -5079 5664 -5045
rect 5860 -5079 5876 -5045
rect -20644 -5225 -19442 -5208
rect -20890 -5230 -19442 -5225
rect -20890 -5276 -20603 -5230
rect -19480 -5276 -19442 -5230
rect -20890 -5289 -19442 -5276
rect -20644 -5299 -19442 -5289
rect -19085 -5230 -17883 -5208
rect -19085 -5276 -19044 -5230
rect -17921 -5276 -17883 -5230
rect -19085 -5299 -17883 -5276
rect -17353 -5230 -16151 -5208
rect -17353 -5276 -17312 -5230
rect -16189 -5276 -16151 -5230
rect -17353 -5299 -16151 -5276
rect -15794 -5230 -14592 -5208
rect -15794 -5276 -15753 -5230
rect -14630 -5276 -14592 -5230
rect -15794 -5299 -14592 -5276
rect -14062 -5230 -12860 -5208
rect -14062 -5276 -14021 -5230
rect -12898 -5276 -12860 -5230
rect -14062 -5299 -12860 -5276
rect -12503 -5230 -11301 -5208
rect -12503 -5276 -12462 -5230
rect -11339 -5276 -11301 -5230
rect -12503 -5299 -11301 -5276
rect -10771 -5230 -9569 -5208
rect -10771 -5276 -10730 -5230
rect -9607 -5276 -9569 -5230
rect -10771 -5299 -9569 -5276
rect -9212 -5230 -8010 -5208
rect -9212 -5276 -9171 -5230
rect -8048 -5276 -8010 -5230
rect -9212 -5299 -8010 -5276
rect 5561 -5319 5577 -5093
rect 6001 -5093 6051 -5076
rect 6094 -5079 6104 -5045
rect 6300 -5079 6316 -5045
rect 5654 -5175 5670 -5141
rect 5864 -5175 5882 -5141
rect 5654 -5271 5664 -5237
rect 5860 -5271 5876 -5237
rect -23539 -5385 -23523 -5351
rect -23432 -5385 -23416 -5351
rect -21805 -5385 -21789 -5351
rect -21698 -5385 -21682 -5351
rect -24384 -5451 -24368 -5404
rect -23799 -5451 -23775 -5404
rect -23683 -5471 -23633 -5454
rect -23590 -5457 -23580 -5423
rect -23384 -5457 -23368 -5423
rect -22648 -5451 -22632 -5404
rect -22063 -5451 -22039 -5404
rect -24384 -5523 -24350 -5513
rect -24384 -5735 -24350 -5719
rect -24288 -5529 -24254 -5513
rect -24288 -5735 -24254 -5725
rect -24192 -5523 -24158 -5513
rect -24192 -5735 -24158 -5719
rect -24096 -5529 -24062 -5513
rect -24096 -5735 -24062 -5725
rect -24000 -5523 -23966 -5513
rect -24000 -5735 -23966 -5719
rect -23904 -5529 -23870 -5513
rect -23904 -5735 -23870 -5725
rect -23808 -5523 -23774 -5513
rect -23808 -5735 -23774 -5719
rect -23683 -5697 -23667 -5471
rect -21949 -5471 -21899 -5454
rect -21856 -5457 -21846 -5423
rect -21650 -5457 -21634 -5423
rect -23590 -5553 -23574 -5519
rect -23380 -5553 -23362 -5519
rect -22648 -5523 -22614 -5513
rect -23590 -5649 -23580 -5615
rect -23384 -5649 -23368 -5615
rect -24335 -5813 -24318 -5778
rect -24284 -5813 -24268 -5778
rect -24046 -5784 -24029 -5778
rect -24234 -5813 -24029 -5784
rect -23995 -5813 -23979 -5778
rect -24335 -6019 -24292 -5813
rect -24234 -5818 -23979 -5813
rect -24234 -5902 -24200 -5818
rect -24166 -5907 -24150 -5873
rect -23774 -5907 -23758 -5873
rect -24234 -5953 -24200 -5937
rect -23683 -5917 -23633 -5697
rect -23590 -5745 -23574 -5711
rect -23380 -5745 -23362 -5711
rect -22648 -5735 -22614 -5719
rect -22552 -5529 -22518 -5513
rect -22552 -5735 -22518 -5725
rect -22456 -5523 -22422 -5513
rect -22456 -5735 -22422 -5719
rect -22360 -5529 -22326 -5513
rect -22360 -5735 -22326 -5725
rect -22264 -5523 -22230 -5513
rect -22264 -5735 -22230 -5719
rect -22168 -5529 -22134 -5513
rect -22168 -5735 -22134 -5725
rect -22072 -5523 -22038 -5513
rect -22072 -5735 -22038 -5719
rect -21949 -5697 -21933 -5471
rect -21856 -5553 -21840 -5519
rect -21646 -5553 -21628 -5519
rect 5561 -5539 5611 -5319
rect 6001 -5319 6017 -5093
rect 6441 -5093 6491 -5076
rect 6534 -5079 6544 -5045
rect 6740 -5079 6756 -5045
rect 6094 -5175 6110 -5141
rect 6304 -5175 6322 -5141
rect 6094 -5271 6104 -5237
rect 6300 -5271 6316 -5237
rect 5654 -5367 5670 -5333
rect 5864 -5367 5882 -5333
rect 5654 -5529 5670 -5495
rect 5846 -5529 5862 -5495
rect -21856 -5649 -21846 -5615
rect -21650 -5649 -21634 -5615
rect -20518 -5619 -20502 -5572
rect -19933 -5619 -19909 -5572
rect -19409 -5619 -19393 -5572
rect -18824 -5619 -18800 -5572
rect -18527 -5619 -18511 -5572
rect -17942 -5619 -17918 -5572
rect -17227 -5619 -17211 -5572
rect -16642 -5619 -16618 -5572
rect -16118 -5619 -16102 -5572
rect -15533 -5619 -15509 -5572
rect -15236 -5619 -15220 -5572
rect -14651 -5619 -14627 -5572
rect -13936 -5619 -13920 -5572
rect -13351 -5619 -13327 -5572
rect -12827 -5619 -12811 -5572
rect -12242 -5619 -12218 -5572
rect -11945 -5619 -11929 -5572
rect -11360 -5619 -11336 -5572
rect -10645 -5619 -10629 -5572
rect -10060 -5619 -10036 -5572
rect -9536 -5619 -9520 -5572
rect -8951 -5619 -8927 -5572
rect -8654 -5619 -8638 -5572
rect -8069 -5619 -8045 -5572
rect 5561 -5573 5577 -5539
rect 5561 -5589 5611 -5573
rect 6001 -5539 6051 -5319
rect 6441 -5319 6457 -5093
rect 6534 -5175 6550 -5141
rect 6744 -5175 6762 -5141
rect 6534 -5271 6544 -5237
rect 6740 -5271 6756 -5237
rect 6094 -5367 6110 -5333
rect 6304 -5367 6322 -5333
rect 6094 -5529 6110 -5495
rect 6286 -5529 6302 -5495
rect 6001 -5573 6017 -5539
rect 5654 -5617 5670 -5583
rect 5846 -5617 5862 -5583
rect 6001 -5589 6051 -5573
rect 6441 -5539 6491 -5319
rect 6534 -5367 6550 -5333
rect 6744 -5367 6762 -5333
rect 6534 -5529 6550 -5495
rect 6726 -5529 6742 -5495
rect 6441 -5573 6457 -5539
rect 6094 -5617 6110 -5583
rect 6286 -5617 6302 -5583
rect 6441 -5589 6491 -5573
rect 6534 -5617 6550 -5583
rect 6726 -5617 6742 -5583
rect 7373 -5680 7389 -5645
rect 7677 -5680 7703 -5645
rect 8321 -5680 8337 -5645
rect 8625 -5680 8651 -5645
rect 9257 -5680 9273 -5645
rect 9561 -5680 9587 -5645
rect 10188 -5680 10204 -5645
rect 10492 -5680 10518 -5645
rect 11115 -5680 11131 -5645
rect 11419 -5680 11445 -5645
rect -22599 -5813 -22582 -5778
rect -22548 -5813 -22532 -5778
rect -22310 -5784 -22293 -5778
rect -22498 -5813 -22293 -5784
rect -22259 -5813 -22243 -5778
rect -23590 -5907 -23574 -5873
rect -23398 -5907 -23382 -5873
rect -23683 -5951 -23667 -5917
rect -23683 -5967 -23633 -5951
rect -23590 -5995 -23574 -5961
rect -23398 -5995 -23382 -5961
rect -22599 -6019 -22556 -5813
rect -22498 -5818 -22243 -5813
rect -22498 -5902 -22464 -5818
rect -22430 -5907 -22414 -5873
rect -22038 -5907 -22022 -5873
rect -22498 -5953 -22464 -5937
rect -21949 -5917 -21899 -5697
rect -20518 -5691 -20484 -5681
rect -21856 -5745 -21840 -5711
rect -21646 -5745 -21628 -5711
rect -21856 -5907 -21840 -5873
rect -21664 -5907 -21648 -5873
rect -20518 -5903 -20484 -5887
rect -20422 -5697 -20388 -5681
rect -20422 -5903 -20388 -5893
rect -20326 -5691 -20292 -5681
rect -20326 -5903 -20292 -5887
rect -20230 -5697 -20196 -5681
rect -20230 -5903 -20196 -5893
rect -20134 -5691 -20100 -5681
rect -20134 -5903 -20100 -5887
rect -20038 -5697 -20004 -5681
rect -20038 -5903 -20004 -5893
rect -19942 -5691 -19908 -5681
rect -19942 -5903 -19908 -5887
rect -19409 -5691 -19375 -5681
rect -19409 -5903 -19375 -5887
rect -19313 -5697 -19279 -5681
rect -19313 -5903 -19279 -5893
rect -19217 -5691 -19183 -5681
rect -19217 -5903 -19183 -5887
rect -19121 -5697 -19087 -5681
rect -19121 -5903 -19087 -5893
rect -19025 -5691 -18991 -5681
rect -19025 -5903 -18991 -5887
rect -18929 -5697 -18895 -5681
rect -18929 -5903 -18895 -5893
rect -18833 -5691 -18799 -5681
rect -18833 -5903 -18799 -5887
rect -18527 -5691 -18493 -5681
rect -18527 -5903 -18493 -5887
rect -18431 -5697 -18397 -5681
rect -18431 -5903 -18397 -5893
rect -18335 -5691 -18301 -5681
rect -18335 -5903 -18301 -5887
rect -18239 -5697 -18205 -5681
rect -18239 -5903 -18205 -5893
rect -18143 -5691 -18109 -5681
rect -18143 -5903 -18109 -5887
rect -18047 -5697 -18013 -5681
rect -18047 -5903 -18013 -5893
rect -17951 -5691 -17917 -5681
rect -17951 -5903 -17917 -5887
rect -17227 -5691 -17193 -5681
rect -17227 -5903 -17193 -5887
rect -17131 -5697 -17097 -5681
rect -17131 -5903 -17097 -5893
rect -17035 -5691 -17001 -5681
rect -17035 -5903 -17001 -5887
rect -16939 -5697 -16905 -5681
rect -16939 -5903 -16905 -5893
rect -16843 -5691 -16809 -5681
rect -16843 -5903 -16809 -5887
rect -16747 -5697 -16713 -5681
rect -16747 -5903 -16713 -5893
rect -16651 -5691 -16617 -5681
rect -16651 -5903 -16617 -5887
rect -16118 -5691 -16084 -5681
rect -16118 -5903 -16084 -5887
rect -16022 -5697 -15988 -5681
rect -16022 -5903 -15988 -5893
rect -15926 -5691 -15892 -5681
rect -15926 -5903 -15892 -5887
rect -15830 -5697 -15796 -5681
rect -15830 -5903 -15796 -5893
rect -15734 -5691 -15700 -5681
rect -15734 -5903 -15700 -5887
rect -15638 -5697 -15604 -5681
rect -15638 -5903 -15604 -5893
rect -15542 -5691 -15508 -5681
rect -15542 -5903 -15508 -5887
rect -15236 -5691 -15202 -5681
rect -15236 -5903 -15202 -5887
rect -15140 -5697 -15106 -5681
rect -15140 -5903 -15106 -5893
rect -15044 -5691 -15010 -5681
rect -15044 -5903 -15010 -5887
rect -14948 -5697 -14914 -5681
rect -14948 -5903 -14914 -5893
rect -14852 -5691 -14818 -5681
rect -14852 -5903 -14818 -5887
rect -14756 -5697 -14722 -5681
rect -14756 -5903 -14722 -5893
rect -14660 -5691 -14626 -5681
rect -14660 -5903 -14626 -5887
rect -13936 -5691 -13902 -5681
rect -13936 -5903 -13902 -5887
rect -13840 -5697 -13806 -5681
rect -13840 -5903 -13806 -5893
rect -13744 -5691 -13710 -5681
rect -13744 -5903 -13710 -5887
rect -13648 -5697 -13614 -5681
rect -13648 -5903 -13614 -5893
rect -13552 -5691 -13518 -5681
rect -13552 -5903 -13518 -5887
rect -13456 -5697 -13422 -5681
rect -13456 -5903 -13422 -5893
rect -13360 -5691 -13326 -5681
rect -13360 -5903 -13326 -5887
rect -12827 -5691 -12793 -5681
rect -12827 -5903 -12793 -5887
rect -12731 -5697 -12697 -5681
rect -12731 -5903 -12697 -5893
rect -12635 -5691 -12601 -5681
rect -12635 -5903 -12601 -5887
rect -12539 -5697 -12505 -5681
rect -12539 -5903 -12505 -5893
rect -12443 -5691 -12409 -5681
rect -12443 -5903 -12409 -5887
rect -12347 -5697 -12313 -5681
rect -12347 -5903 -12313 -5893
rect -12251 -5691 -12217 -5681
rect -12251 -5903 -12217 -5887
rect -11945 -5691 -11911 -5681
rect -11945 -5903 -11911 -5887
rect -11849 -5697 -11815 -5681
rect -11849 -5903 -11815 -5893
rect -11753 -5691 -11719 -5681
rect -11753 -5903 -11719 -5887
rect -11657 -5697 -11623 -5681
rect -11657 -5903 -11623 -5893
rect -11561 -5691 -11527 -5681
rect -11561 -5903 -11527 -5887
rect -11465 -5697 -11431 -5681
rect -11465 -5903 -11431 -5893
rect -11369 -5691 -11335 -5681
rect -11369 -5903 -11335 -5887
rect -10645 -5691 -10611 -5681
rect -10645 -5903 -10611 -5887
rect -10549 -5697 -10515 -5681
rect -10549 -5903 -10515 -5893
rect -10453 -5691 -10419 -5681
rect -10453 -5903 -10419 -5887
rect -10357 -5697 -10323 -5681
rect -10357 -5903 -10323 -5893
rect -10261 -5691 -10227 -5681
rect -10261 -5903 -10227 -5887
rect -10165 -5697 -10131 -5681
rect -10165 -5903 -10131 -5893
rect -10069 -5691 -10035 -5681
rect -10069 -5903 -10035 -5887
rect -9536 -5691 -9502 -5681
rect -9536 -5903 -9502 -5887
rect -9440 -5697 -9406 -5681
rect -9440 -5903 -9406 -5893
rect -9344 -5691 -9310 -5681
rect -9344 -5903 -9310 -5887
rect -9248 -5697 -9214 -5681
rect -9248 -5903 -9214 -5893
rect -9152 -5691 -9118 -5681
rect -9152 -5903 -9118 -5887
rect -9056 -5697 -9022 -5681
rect -9056 -5903 -9022 -5893
rect -8960 -5691 -8926 -5681
rect -8960 -5903 -8926 -5887
rect -8654 -5691 -8620 -5681
rect -8654 -5903 -8620 -5887
rect -8558 -5697 -8524 -5681
rect -8558 -5903 -8524 -5893
rect -8462 -5691 -8428 -5681
rect -8462 -5903 -8428 -5887
rect -8366 -5697 -8332 -5681
rect -8366 -5903 -8332 -5893
rect -8270 -5691 -8236 -5681
rect -8270 -5903 -8236 -5887
rect -8174 -5697 -8140 -5681
rect -8174 -5903 -8140 -5893
rect -8078 -5691 -8044 -5681
rect 5673 -5719 5689 -5685
rect 5821 -5719 5837 -5685
rect 6113 -5719 6129 -5685
rect 6261 -5719 6277 -5685
rect 6553 -5719 6569 -5685
rect 6701 -5719 6717 -5685
rect -8078 -5903 -8044 -5887
rect 7150 -5749 7184 -5733
rect -21949 -5951 -21933 -5917
rect -21949 -5967 -21899 -5951
rect -21856 -5995 -21840 -5961
rect -21664 -5995 -21648 -5961
rect -20469 -5981 -20452 -5946
rect -20418 -5981 -20402 -5946
rect -20180 -5952 -20163 -5946
rect -20368 -5981 -20163 -5952
rect -20129 -5981 -20113 -5946
rect -24335 -6035 -24200 -6019
rect -24335 -6070 -24234 -6035
rect -22599 -6035 -22464 -6019
rect -24335 -6086 -24200 -6070
rect -24166 -6099 -24150 -6065
rect -23774 -6099 -23758 -6065
rect -23571 -6097 -23555 -6063
rect -23423 -6097 -23407 -6063
rect -22599 -6070 -22498 -6035
rect -22599 -6086 -22464 -6070
rect -22430 -6099 -22414 -6065
rect -22038 -6099 -22022 -6065
rect -21837 -6097 -21821 -6063
rect -21689 -6097 -21673 -6063
rect -24162 -6171 -24135 -6137
rect -23800 -6171 -23762 -6137
rect -22426 -6171 -22399 -6137
rect -22064 -6171 -22026 -6137
rect -20469 -6187 -20426 -5981
rect -20368 -5986 -20113 -5981
rect -19360 -5981 -19343 -5946
rect -19309 -5981 -19293 -5946
rect -19071 -5952 -19054 -5946
rect -19259 -5981 -19054 -5952
rect -19020 -5981 -19004 -5946
rect -20368 -6070 -20334 -5986
rect -20300 -6075 -20284 -6041
rect -19908 -6075 -19892 -6041
rect -20368 -6121 -20334 -6105
rect -19360 -6187 -19317 -5981
rect -19259 -5986 -19004 -5981
rect -18478 -5981 -18461 -5946
rect -18427 -5981 -18411 -5946
rect -18189 -5952 -18172 -5946
rect -18377 -5981 -18172 -5952
rect -18138 -5981 -18122 -5946
rect -19259 -6070 -19225 -5986
rect -19191 -6075 -19175 -6041
rect -18799 -6075 -18783 -6041
rect -19259 -6121 -19225 -6105
rect -18478 -6187 -18435 -5981
rect -18377 -5986 -18122 -5981
rect -17178 -5981 -17161 -5946
rect -17127 -5981 -17111 -5946
rect -16889 -5952 -16872 -5946
rect -17077 -5981 -16872 -5952
rect -16838 -5981 -16822 -5946
rect -18377 -6070 -18343 -5986
rect -18309 -6075 -18293 -6041
rect -17917 -6075 -17901 -6041
rect -18377 -6121 -18343 -6105
rect -17178 -6187 -17135 -5981
rect -17077 -5986 -16822 -5981
rect -16069 -5981 -16052 -5946
rect -16018 -5981 -16002 -5946
rect -15780 -5952 -15763 -5946
rect -15968 -5981 -15763 -5952
rect -15729 -5981 -15713 -5946
rect -17077 -6070 -17043 -5986
rect -17009 -6075 -16993 -6041
rect -16617 -6075 -16601 -6041
rect -17077 -6121 -17043 -6105
rect -16069 -6187 -16026 -5981
rect -15968 -5986 -15713 -5981
rect -15187 -5981 -15170 -5946
rect -15136 -5981 -15120 -5946
rect -14898 -5952 -14881 -5946
rect -15086 -5981 -14881 -5952
rect -14847 -5981 -14831 -5946
rect -15968 -6070 -15934 -5986
rect -15900 -6075 -15884 -6041
rect -15508 -6075 -15492 -6041
rect -15968 -6121 -15934 -6105
rect -15187 -6187 -15144 -5981
rect -15086 -5986 -14831 -5981
rect -13887 -5981 -13870 -5946
rect -13836 -5981 -13820 -5946
rect -13598 -5952 -13581 -5946
rect -13786 -5981 -13581 -5952
rect -13547 -5981 -13531 -5946
rect -15086 -6070 -15052 -5986
rect -15018 -6075 -15002 -6041
rect -14626 -6075 -14610 -6041
rect -15086 -6121 -15052 -6105
rect -13887 -6187 -13844 -5981
rect -13786 -5986 -13531 -5981
rect -12778 -5981 -12761 -5946
rect -12727 -5981 -12711 -5946
rect -12489 -5952 -12472 -5946
rect -12677 -5981 -12472 -5952
rect -12438 -5981 -12422 -5946
rect -13786 -6070 -13752 -5986
rect -13718 -6075 -13702 -6041
rect -13326 -6075 -13310 -6041
rect -13786 -6121 -13752 -6105
rect -12778 -6187 -12735 -5981
rect -12677 -5986 -12422 -5981
rect -11896 -5981 -11879 -5946
rect -11845 -5981 -11829 -5946
rect -11607 -5952 -11590 -5946
rect -11795 -5981 -11590 -5952
rect -11556 -5981 -11540 -5946
rect -12677 -6070 -12643 -5986
rect -12609 -6075 -12593 -6041
rect -12217 -6075 -12201 -6041
rect -12677 -6121 -12643 -6105
rect -11896 -6187 -11853 -5981
rect -11795 -5986 -11540 -5981
rect -10596 -5981 -10579 -5946
rect -10545 -5981 -10529 -5946
rect -10307 -5952 -10290 -5946
rect -10495 -5981 -10290 -5952
rect -10256 -5981 -10240 -5946
rect -11795 -6070 -11761 -5986
rect -11727 -6075 -11711 -6041
rect -11335 -6075 -11319 -6041
rect -11795 -6121 -11761 -6105
rect -10596 -6187 -10553 -5981
rect -10495 -5986 -10240 -5981
rect -9487 -5981 -9470 -5946
rect -9436 -5981 -9420 -5946
rect -9198 -5952 -9181 -5946
rect -9386 -5981 -9181 -5952
rect -9147 -5981 -9131 -5946
rect -10495 -6070 -10461 -5986
rect -10427 -6075 -10411 -6041
rect -10035 -6075 -10019 -6041
rect -10495 -6121 -10461 -6105
rect -9487 -6187 -9444 -5981
rect -9386 -5986 -9131 -5981
rect -8605 -5981 -8588 -5946
rect -8554 -5981 -8538 -5946
rect -8316 -5952 -8299 -5946
rect -8504 -5981 -8299 -5952
rect -8265 -5981 -8249 -5946
rect -9386 -6070 -9352 -5986
rect -9318 -6075 -9302 -6041
rect -8926 -6075 -8910 -6041
rect -9386 -6121 -9352 -6105
rect -8605 -6187 -8562 -5981
rect -8504 -5986 -8249 -5981
rect -8504 -6070 -8470 -5986
rect -8436 -6075 -8420 -6041
rect -8044 -6075 -8028 -6041
rect 7246 -5749 7280 -5733
rect 7150 -6063 7184 -6047
rect 7246 -6063 7280 -6052
rect 7342 -5749 7376 -5733
rect 7342 -6063 7376 -6047
rect 7438 -5749 7472 -5733
rect 7534 -5749 7568 -5733
rect 7438 -6063 7472 -6052
rect 7534 -6063 7568 -6047
rect 7630 -5749 7664 -5733
rect 7726 -5749 7760 -5733
rect 7630 -6063 7664 -6052
rect 7726 -6063 7760 -6047
rect 7822 -5749 7856 -5733
rect 7918 -5749 7952 -5733
rect 7822 -6063 7856 -6052
rect 7918 -6063 7952 -6047
rect 8098 -5749 8132 -5733
rect 8194 -5749 8228 -5733
rect 8098 -6063 8132 -6047
rect 8194 -6063 8228 -6052
rect 8290 -5749 8324 -5733
rect 8290 -6063 8324 -6047
rect 8386 -5749 8420 -5733
rect 8482 -5749 8516 -5733
rect 8386 -6063 8420 -6052
rect 8482 -6063 8516 -6047
rect 8578 -5749 8612 -5733
rect 8674 -5749 8708 -5733
rect 8578 -6063 8612 -6052
rect 8674 -6063 8708 -6047
rect 8770 -5749 8804 -5733
rect 8866 -5749 8900 -5733
rect 8770 -6063 8804 -6052
rect 8866 -6063 8900 -6047
rect 9034 -5749 9068 -5733
rect 9130 -5749 9164 -5733
rect 9034 -6063 9068 -6047
rect 9130 -6063 9164 -6052
rect 9226 -5749 9260 -5733
rect 9226 -6063 9260 -6047
rect 9322 -5749 9356 -5733
rect 9418 -5749 9452 -5733
rect 9322 -6063 9356 -6052
rect 9418 -6063 9452 -6047
rect 9514 -5749 9548 -5733
rect 9610 -5749 9644 -5733
rect 9514 -6063 9548 -6052
rect 9610 -6063 9644 -6047
rect 9706 -5749 9740 -5733
rect 9802 -5749 9836 -5733
rect 9706 -6063 9740 -6052
rect 9802 -6063 9836 -6047
rect 9965 -5749 9999 -5733
rect 10061 -5749 10095 -5733
rect 9965 -6063 9999 -6047
rect 10061 -6063 10095 -6052
rect 10157 -5749 10191 -5733
rect 10157 -6063 10191 -6047
rect 10253 -5749 10287 -5733
rect 10349 -5749 10383 -5733
rect 10253 -6063 10287 -6052
rect 10349 -6063 10383 -6047
rect 10445 -5749 10479 -5733
rect 10541 -5749 10575 -5733
rect 10445 -6063 10479 -6052
rect 10541 -6063 10575 -6047
rect 10637 -5749 10671 -5733
rect 10733 -5749 10767 -5733
rect 10637 -6063 10671 -6052
rect 10733 -6063 10767 -6047
rect 10892 -5749 10926 -5733
rect 10988 -5749 11022 -5733
rect 10892 -6063 10926 -6047
rect 10988 -6063 11022 -6052
rect 11084 -5749 11118 -5733
rect 11084 -6063 11118 -6047
rect 11180 -5749 11214 -5733
rect 11276 -5749 11310 -5733
rect 11180 -6063 11214 -6052
rect 11276 -6063 11310 -6047
rect 11372 -5749 11406 -5733
rect 11468 -5749 11502 -5733
rect 11372 -6063 11406 -6052
rect 11468 -6063 11502 -6047
rect 11564 -5749 11598 -5733
rect 11660 -5749 11694 -5733
rect 11564 -6063 11598 -6052
rect 11660 -6063 11694 -6047
rect -8504 -6121 -8470 -6105
rect 7182 -6140 7198 -6106
rect 7232 -6140 7248 -6106
rect 7374 -6140 7390 -6106
rect 7424 -6140 7440 -6106
rect 7566 -6140 7582 -6106
rect 7616 -6140 7632 -6106
rect 7758 -6140 7774 -6106
rect 7808 -6140 7824 -6106
rect 8130 -6140 8146 -6106
rect 8180 -6140 8196 -6106
rect 8322 -6140 8338 -6106
rect 8372 -6140 8388 -6106
rect 8514 -6140 8530 -6106
rect 8564 -6140 8580 -6106
rect 8706 -6140 8722 -6106
rect 8756 -6140 8772 -6106
rect 9066 -6140 9082 -6106
rect 9116 -6140 9132 -6106
rect 9258 -6140 9274 -6106
rect 9308 -6140 9324 -6106
rect 9450 -6140 9466 -6106
rect 9500 -6140 9516 -6106
rect 9642 -6140 9658 -6106
rect 9692 -6140 9708 -6106
rect 9997 -6140 10013 -6106
rect 10047 -6140 10063 -6106
rect 10189 -6140 10205 -6106
rect 10239 -6140 10255 -6106
rect 10381 -6140 10397 -6106
rect 10431 -6140 10447 -6106
rect 10573 -6140 10589 -6106
rect 10623 -6140 10639 -6106
rect 10924 -6140 10940 -6106
rect 10974 -6140 10990 -6106
rect 11116 -6140 11132 -6106
rect 11166 -6140 11182 -6106
rect 11308 -6140 11324 -6106
rect 11358 -6140 11374 -6106
rect 11500 -6140 11516 -6106
rect 11550 -6140 11566 -6106
rect -20469 -6203 -20334 -6187
rect -20469 -6238 -20368 -6203
rect -19360 -6203 -19225 -6187
rect -20469 -6254 -20334 -6238
rect -20300 -6267 -20284 -6233
rect -19908 -6267 -19892 -6233
rect -19360 -6238 -19259 -6203
rect -18478 -6203 -18343 -6187
rect -19360 -6254 -19225 -6238
rect -19191 -6267 -19175 -6233
rect -18799 -6267 -18783 -6233
rect -18478 -6238 -18377 -6203
rect -17178 -6203 -17043 -6187
rect -18478 -6254 -18343 -6238
rect -18309 -6267 -18293 -6233
rect -17917 -6267 -17901 -6233
rect -17178 -6238 -17077 -6203
rect -16069 -6203 -15934 -6187
rect -17178 -6254 -17043 -6238
rect -17009 -6267 -16993 -6233
rect -16617 -6267 -16601 -6233
rect -16069 -6238 -15968 -6203
rect -15187 -6203 -15052 -6187
rect -16069 -6254 -15934 -6238
rect -15900 -6267 -15884 -6233
rect -15508 -6267 -15492 -6233
rect -15187 -6238 -15086 -6203
rect -13887 -6203 -13752 -6187
rect -15187 -6254 -15052 -6238
rect -15018 -6267 -15002 -6233
rect -14626 -6267 -14610 -6233
rect -13887 -6238 -13786 -6203
rect -12778 -6203 -12643 -6187
rect -13887 -6254 -13752 -6238
rect -13718 -6267 -13702 -6233
rect -13326 -6267 -13310 -6233
rect -12778 -6238 -12677 -6203
rect -11896 -6203 -11761 -6187
rect -12778 -6254 -12643 -6238
rect -12609 -6267 -12593 -6233
rect -12217 -6267 -12201 -6233
rect -11896 -6238 -11795 -6203
rect -10596 -6203 -10461 -6187
rect -11896 -6254 -11761 -6238
rect -11727 -6267 -11711 -6233
rect -11335 -6267 -11319 -6233
rect -10596 -6238 -10495 -6203
rect -9487 -6203 -9352 -6187
rect -10596 -6254 -10461 -6238
rect -10427 -6267 -10411 -6233
rect -10035 -6267 -10019 -6233
rect -9487 -6238 -9386 -6203
rect -8605 -6203 -8470 -6187
rect -9487 -6254 -9352 -6238
rect -9318 -6267 -9302 -6233
rect -8926 -6267 -8910 -6233
rect -8605 -6238 -8504 -6203
rect -8605 -6254 -8470 -6238
rect -8436 -6267 -8420 -6233
rect -8044 -6267 -8028 -6233
rect -20296 -6339 -20269 -6305
rect -19934 -6339 -19896 -6305
rect -19187 -6339 -19160 -6305
rect -18825 -6339 -18787 -6305
rect -18305 -6339 -18278 -6305
rect -17943 -6339 -17905 -6305
rect -17005 -6339 -16978 -6305
rect -16643 -6339 -16605 -6305
rect -15896 -6339 -15869 -6305
rect -15534 -6339 -15496 -6305
rect -15014 -6339 -14987 -6305
rect -14652 -6339 -14614 -6305
rect -13714 -6339 -13687 -6305
rect -13352 -6339 -13314 -6305
rect -12605 -6339 -12578 -6305
rect -12243 -6339 -12205 -6305
rect -11723 -6339 -11696 -6305
rect -11361 -6339 -11323 -6305
rect -10423 -6339 -10396 -6305
rect -10061 -6339 -10023 -6305
rect -9314 -6339 -9287 -6305
rect -8952 -6339 -8914 -6305
rect -8432 -6339 -8405 -6305
rect -8070 -6339 -8032 -6305
rect 7298 -6462 7403 -6459
rect 8246 -6462 8351 -6459
rect 9182 -6462 9287 -6459
rect 10113 -6462 10218 -6459
rect 11040 -6462 11145 -6459
rect 7298 -6478 7406 -6462
rect 7298 -6490 7372 -6478
rect -20649 -7092 -19439 -7064
rect -20649 -7164 -20603 -7092
rect -19481 -7164 -19439 -7092
rect -20649 -7190 -19439 -7164
rect -19090 -7092 -17880 -7064
rect -19090 -7164 -19044 -7092
rect -17922 -7164 -17880 -7092
rect -19090 -7190 -17880 -7164
rect -17358 -7092 -16148 -7064
rect -17358 -7164 -17312 -7092
rect -16190 -7164 -16148 -7092
rect -17358 -7190 -16148 -7164
rect -15799 -7092 -14589 -7064
rect -15799 -7164 -15753 -7092
rect -14631 -7164 -14589 -7092
rect -15799 -7190 -14589 -7164
rect -14067 -7092 -12857 -7064
rect -14067 -7164 -14021 -7092
rect -12899 -7164 -12857 -7092
rect -14067 -7190 -12857 -7164
rect -12508 -7092 -11298 -7064
rect -12508 -7164 -12462 -7092
rect -11340 -7164 -11298 -7092
rect -12508 -7190 -11298 -7164
rect -10776 -7092 -9566 -7064
rect -10776 -7164 -10730 -7092
rect -9608 -7164 -9566 -7092
rect -10776 -7190 -9566 -7164
rect -9217 -7092 -8007 -7064
rect -9217 -7164 -9171 -7092
rect -8049 -7164 -8007 -7092
rect -9217 -7190 -8007 -7164
rect 7333 -7241 7372 -6490
rect -20725 -7261 -20691 -7245
rect -23537 -7358 -23521 -7324
rect -23430 -7358 -23414 -7324
rect -21803 -7358 -21787 -7324
rect -21696 -7358 -21680 -7324
rect -24384 -7424 -24368 -7377
rect -23799 -7424 -23775 -7377
rect -23681 -7444 -23631 -7427
rect -23588 -7430 -23578 -7396
rect -23382 -7430 -23366 -7396
rect -22647 -7424 -22631 -7377
rect -22062 -7424 -22038 -7377
rect -24384 -7496 -24350 -7486
rect -24384 -7708 -24350 -7692
rect -24288 -7502 -24254 -7486
rect -24288 -7708 -24254 -7698
rect -24192 -7496 -24158 -7486
rect -24192 -7708 -24158 -7692
rect -24096 -7502 -24062 -7486
rect -24096 -7708 -24062 -7698
rect -24000 -7496 -23966 -7486
rect -24000 -7708 -23966 -7692
rect -23904 -7502 -23870 -7486
rect -23904 -7708 -23870 -7698
rect -23808 -7496 -23774 -7486
rect -23808 -7708 -23774 -7692
rect -23681 -7670 -23665 -7444
rect -21947 -7444 -21897 -7427
rect -21854 -7430 -21844 -7396
rect -21648 -7430 -21632 -7396
rect -23588 -7526 -23572 -7492
rect -23378 -7526 -23360 -7492
rect -22647 -7496 -22613 -7486
rect -23588 -7622 -23578 -7588
rect -23382 -7622 -23366 -7588
rect -24335 -7786 -24318 -7751
rect -24284 -7786 -24268 -7751
rect -24046 -7757 -24029 -7751
rect -24234 -7786 -24029 -7757
rect -23995 -7786 -23979 -7751
rect -24335 -7992 -24292 -7786
rect -24234 -7791 -23979 -7786
rect -24234 -7875 -24200 -7791
rect -24166 -7880 -24150 -7846
rect -23774 -7880 -23758 -7846
rect -24234 -7926 -24200 -7910
rect -23681 -7890 -23631 -7670
rect -23588 -7718 -23572 -7684
rect -23378 -7718 -23360 -7684
rect -22647 -7708 -22613 -7692
rect -22551 -7502 -22517 -7486
rect -22551 -7708 -22517 -7698
rect -22455 -7496 -22421 -7486
rect -22455 -7708 -22421 -7692
rect -22359 -7502 -22325 -7486
rect -22359 -7708 -22325 -7698
rect -22263 -7496 -22229 -7486
rect -22263 -7708 -22229 -7692
rect -22167 -7502 -22133 -7486
rect -22167 -7708 -22133 -7698
rect -22071 -7496 -22037 -7486
rect -22071 -7708 -22037 -7692
rect -21947 -7670 -21931 -7444
rect -21854 -7526 -21838 -7492
rect -21644 -7526 -21626 -7492
rect -21854 -7622 -21844 -7588
rect -21648 -7622 -21632 -7588
rect -22598 -7786 -22581 -7751
rect -22547 -7786 -22531 -7751
rect -22309 -7757 -22292 -7751
rect -22497 -7786 -22292 -7757
rect -22258 -7786 -22242 -7751
rect -23588 -7880 -23572 -7846
rect -23396 -7880 -23380 -7846
rect -23681 -7924 -23665 -7890
rect -23681 -7940 -23631 -7924
rect -23588 -7968 -23572 -7934
rect -23396 -7968 -23380 -7934
rect -22598 -7992 -22555 -7786
rect -22497 -7791 -22242 -7786
rect -22497 -7875 -22463 -7791
rect -22429 -7880 -22413 -7846
rect -22037 -7880 -22021 -7846
rect -22497 -7926 -22463 -7910
rect -21947 -7890 -21897 -7670
rect -21854 -7718 -21838 -7684
rect -21644 -7718 -21626 -7684
rect -21854 -7880 -21838 -7846
rect -21662 -7880 -21646 -7846
rect -20725 -7848 -20691 -7787
rect -20637 -7261 -20603 -7245
rect -20637 -7803 -20603 -7787
rect -20541 -7261 -20507 -7245
rect -20541 -7803 -20507 -7787
rect -20445 -7261 -20411 -7245
rect -20445 -7803 -20411 -7787
rect -20349 -7261 -20315 -7245
rect -20349 -7803 -20315 -7787
rect -20253 -7261 -20219 -7245
rect -20253 -7803 -20219 -7787
rect -20157 -7261 -20123 -7245
rect -20157 -7803 -20123 -7787
rect -20061 -7261 -20027 -7245
rect -20061 -7830 -20027 -7787
rect -19965 -7261 -19931 -7245
rect -19965 -7803 -19931 -7787
rect -19869 -7261 -19835 -7245
rect -19869 -7803 -19835 -7787
rect -19773 -7261 -19739 -7245
rect -19773 -7803 -19739 -7787
rect -19677 -7261 -19643 -7245
rect -19677 -7803 -19643 -7787
rect -19581 -7261 -19547 -7245
rect -19581 -7803 -19547 -7787
rect -19485 -7261 -19451 -7245
rect -19485 -7803 -19451 -7787
rect -19397 -7261 -19363 -7245
rect -20725 -7858 -20123 -7848
rect -21947 -7924 -21931 -7890
rect -21947 -7940 -21897 -7924
rect -20872 -7887 -20787 -7864
rect -21854 -7968 -21838 -7934
rect -21662 -7968 -21646 -7934
rect -24335 -8008 -24200 -7992
rect -24335 -8043 -24234 -8008
rect -22598 -8008 -22463 -7992
rect -24335 -8059 -24200 -8043
rect -24166 -8072 -24150 -8038
rect -23774 -8072 -23758 -8038
rect -23569 -8070 -23553 -8036
rect -23421 -8070 -23405 -8036
rect -22598 -8043 -22497 -8008
rect -20872 -7997 -20854 -7887
rect -20807 -7997 -20787 -7887
rect -20872 -8017 -20787 -7997
rect -20725 -7903 -20269 -7858
rect -20139 -7903 -20123 -7858
rect -20725 -7917 -20123 -7903
rect -22598 -8059 -22463 -8043
rect -22429 -8072 -22413 -8038
rect -22037 -8072 -22021 -8038
rect -21835 -8070 -21819 -8036
rect -21687 -8070 -21671 -8036
rect -24162 -8144 -24135 -8110
rect -23800 -8144 -23762 -8110
rect -22425 -8144 -22398 -8110
rect -22063 -8144 -22025 -8110
rect -20725 -8301 -20691 -7917
rect -20589 -7988 -20368 -7961
rect -20589 -8041 -20539 -7988
rect -20406 -8041 -20368 -7988
rect -20589 -8179 -20368 -8041
rect -20589 -8224 -20544 -8179
rect -20414 -8224 -20368 -8179
rect -20589 -8251 -20368 -8224
rect -20288 -8187 -20123 -7917
rect -20288 -8232 -20261 -8187
rect -20131 -8232 -20123 -8187
rect -20288 -8249 -20123 -8232
rect -20077 -8130 -20011 -7830
rect -19397 -7845 -19363 -7787
rect -19965 -7863 -19363 -7845
rect -19965 -7908 -19938 -7863
rect -19808 -7908 -19363 -7863
rect -19965 -7922 -19363 -7908
rect -19166 -7261 -19132 -7245
rect -19166 -7848 -19132 -7787
rect -19078 -7261 -19044 -7245
rect -19078 -7803 -19044 -7787
rect -18982 -7261 -18948 -7245
rect -18982 -7803 -18948 -7787
rect -18886 -7261 -18852 -7245
rect -18886 -7803 -18852 -7787
rect -18790 -7261 -18756 -7245
rect -18790 -7803 -18756 -7787
rect -18694 -7261 -18660 -7245
rect -18694 -7803 -18660 -7787
rect -18598 -7261 -18564 -7245
rect -18598 -7803 -18564 -7787
rect -18502 -7261 -18468 -7245
rect -18502 -7830 -18468 -7787
rect -18406 -7261 -18372 -7245
rect -18406 -7803 -18372 -7787
rect -18310 -7261 -18276 -7245
rect -18310 -7803 -18276 -7787
rect -18214 -7261 -18180 -7245
rect -18214 -7803 -18180 -7787
rect -18118 -7261 -18084 -7245
rect -18118 -7803 -18084 -7787
rect -18022 -7261 -17988 -7245
rect -18022 -7803 -17988 -7787
rect -17926 -7261 -17892 -7245
rect -17926 -7803 -17892 -7787
rect -17838 -7261 -17804 -7245
rect -19166 -7858 -18564 -7848
rect -19166 -7903 -18710 -7858
rect -18580 -7903 -18564 -7858
rect -19166 -7917 -18564 -7903
rect -19965 -7980 -19788 -7922
rect -19965 -8033 -19933 -7980
rect -19819 -8033 -19788 -7980
rect -19965 -8062 -19788 -8033
rect -19716 -7981 -19601 -7963
rect -19716 -8049 -19699 -7981
rect -19619 -8049 -19601 -7981
rect -19716 -8069 -19601 -8049
rect -20077 -8152 -19437 -8130
rect -20077 -8207 -19517 -8152
rect -19452 -8207 -19437 -8152
rect -20077 -8226 -19437 -8207
rect -20077 -8260 -20011 -8226
rect -20725 -8423 -20691 -8407
rect -20637 -8301 -20603 -8285
rect -20637 -8423 -20603 -8407
rect -20541 -8286 -20507 -8285
rect -20541 -8423 -20507 -8407
rect -20445 -8301 -20411 -8285
rect -20445 -8423 -20411 -8421
rect -20349 -8286 -20315 -8285
rect -20349 -8423 -20315 -8407
rect -20253 -8301 -20219 -8285
rect -20253 -8423 -20219 -8421
rect -20157 -8287 -20123 -8285
rect -20157 -8423 -20123 -8407
rect -20061 -8301 -20027 -8260
rect -20061 -8423 -20027 -8421
rect -19965 -8286 -19931 -8285
rect -19965 -8423 -19931 -8407
rect -19869 -8301 -19835 -8285
rect -19869 -8423 -19835 -8421
rect -19773 -8286 -19739 -8285
rect -19773 -8423 -19739 -8407
rect -19677 -8301 -19643 -8285
rect -19677 -8423 -19643 -8421
rect -19581 -8286 -19547 -8285
rect -19581 -8423 -19547 -8407
rect -19485 -8301 -19451 -8285
rect -19485 -8423 -19451 -8407
rect -19397 -8301 -19363 -7922
rect -19316 -7932 -19207 -7917
rect -19316 -8072 -19297 -7932
rect -19224 -8072 -19207 -7932
rect -19316 -8089 -19207 -8072
rect -19397 -8423 -19363 -8407
rect -19166 -8301 -19132 -7917
rect -19030 -7988 -18809 -7961
rect -19030 -8041 -18980 -7988
rect -18847 -8041 -18809 -7988
rect -19030 -8179 -18809 -8041
rect -19030 -8224 -18985 -8179
rect -18855 -8224 -18809 -8179
rect -19030 -8251 -18809 -8224
rect -18729 -8187 -18564 -7917
rect -18729 -8232 -18702 -8187
rect -18572 -8232 -18564 -8187
rect -18729 -8249 -18564 -8232
rect -18518 -8130 -18452 -7830
rect -17838 -7845 -17804 -7787
rect -18406 -7863 -17804 -7845
rect -18406 -7908 -18379 -7863
rect -18249 -7908 -17804 -7863
rect -17434 -7261 -17400 -7245
rect -17434 -7848 -17400 -7787
rect -17346 -7261 -17312 -7245
rect -17346 -7803 -17312 -7787
rect -17250 -7261 -17216 -7245
rect -17250 -7803 -17216 -7787
rect -17154 -7261 -17120 -7245
rect -17154 -7803 -17120 -7787
rect -17058 -7261 -17024 -7245
rect -17058 -7803 -17024 -7787
rect -16962 -7261 -16928 -7245
rect -16962 -7803 -16928 -7787
rect -16866 -7261 -16832 -7245
rect -16866 -7803 -16832 -7787
rect -16770 -7261 -16736 -7245
rect -16770 -7830 -16736 -7787
rect -16674 -7261 -16640 -7245
rect -16674 -7803 -16640 -7787
rect -16578 -7261 -16544 -7245
rect -16578 -7803 -16544 -7787
rect -16482 -7261 -16448 -7245
rect -16482 -7803 -16448 -7787
rect -16386 -7261 -16352 -7245
rect -16386 -7803 -16352 -7787
rect -16290 -7261 -16256 -7245
rect -16290 -7803 -16256 -7787
rect -16194 -7261 -16160 -7245
rect -16194 -7803 -16160 -7787
rect -16106 -7261 -16072 -7245
rect -17434 -7858 -16832 -7848
rect -18406 -7922 -17804 -7908
rect -18406 -7980 -18229 -7922
rect -18406 -8033 -18374 -7980
rect -18260 -8033 -18229 -7980
rect -18406 -8062 -18229 -8033
rect -18157 -7981 -18042 -7963
rect -18157 -8049 -18140 -7981
rect -18060 -8049 -18042 -7981
rect -18157 -8069 -18042 -8049
rect -18518 -8152 -17878 -8130
rect -18518 -8207 -17958 -8152
rect -17893 -8207 -17878 -8152
rect -18518 -8226 -17878 -8207
rect -18518 -8260 -18452 -8226
rect -19166 -8423 -19132 -8407
rect -19078 -8301 -19044 -8285
rect -19078 -8423 -19044 -8407
rect -18982 -8286 -18948 -8285
rect -18982 -8423 -18948 -8407
rect -18886 -8301 -18852 -8285
rect -18886 -8423 -18852 -8421
rect -18790 -8286 -18756 -8285
rect -18790 -8423 -18756 -8407
rect -18694 -8301 -18660 -8285
rect -18694 -8423 -18660 -8421
rect -18598 -8287 -18564 -8285
rect -18598 -8423 -18564 -8407
rect -18502 -8301 -18468 -8260
rect -18502 -8423 -18468 -8421
rect -18406 -8286 -18372 -8285
rect -18406 -8423 -18372 -8407
rect -18310 -8301 -18276 -8285
rect -18310 -8423 -18276 -8421
rect -18214 -8286 -18180 -8285
rect -18214 -8423 -18180 -8407
rect -18118 -8301 -18084 -8285
rect -18118 -8423 -18084 -8421
rect -18022 -8286 -17988 -8285
rect -18022 -8423 -17988 -8407
rect -17926 -8301 -17892 -8285
rect -17926 -8423 -17892 -8407
rect -17838 -8301 -17804 -7922
rect -17581 -7887 -17496 -7864
rect -17581 -7997 -17563 -7887
rect -17516 -7997 -17496 -7887
rect -17581 -8017 -17496 -7997
rect -17434 -7903 -16978 -7858
rect -16848 -7903 -16832 -7858
rect -17434 -7917 -16832 -7903
rect -17838 -8423 -17804 -8407
rect -17434 -8301 -17400 -7917
rect -17298 -7988 -17077 -7961
rect -17298 -8041 -17248 -7988
rect -17115 -8041 -17077 -7988
rect -17298 -8179 -17077 -8041
rect -17298 -8224 -17253 -8179
rect -17123 -8224 -17077 -8179
rect -17298 -8251 -17077 -8224
rect -16997 -8187 -16832 -7917
rect -16997 -8232 -16970 -8187
rect -16840 -8232 -16832 -8187
rect -16997 -8249 -16832 -8232
rect -16786 -8130 -16720 -7830
rect -16106 -7845 -16072 -7787
rect -16674 -7863 -16072 -7845
rect -16674 -7908 -16647 -7863
rect -16517 -7908 -16072 -7863
rect -16674 -7922 -16072 -7908
rect -15875 -7261 -15841 -7245
rect -15875 -7848 -15841 -7787
rect -15787 -7261 -15753 -7245
rect -15787 -7803 -15753 -7787
rect -15691 -7261 -15657 -7245
rect -15691 -7803 -15657 -7787
rect -15595 -7261 -15561 -7245
rect -15595 -7803 -15561 -7787
rect -15499 -7261 -15465 -7245
rect -15499 -7803 -15465 -7787
rect -15403 -7261 -15369 -7245
rect -15403 -7803 -15369 -7787
rect -15307 -7261 -15273 -7245
rect -15307 -7803 -15273 -7787
rect -15211 -7261 -15177 -7245
rect -15211 -7830 -15177 -7787
rect -15115 -7261 -15081 -7245
rect -15115 -7803 -15081 -7787
rect -15019 -7261 -14985 -7245
rect -15019 -7803 -14985 -7787
rect -14923 -7261 -14889 -7245
rect -14923 -7803 -14889 -7787
rect -14827 -7261 -14793 -7245
rect -14827 -7803 -14793 -7787
rect -14731 -7261 -14697 -7245
rect -14731 -7803 -14697 -7787
rect -14635 -7261 -14601 -7245
rect -14635 -7803 -14601 -7787
rect -14547 -7261 -14513 -7245
rect -15875 -7858 -15273 -7848
rect -15875 -7903 -15419 -7858
rect -15289 -7903 -15273 -7858
rect -15875 -7917 -15273 -7903
rect -16674 -7980 -16497 -7922
rect -16674 -8033 -16642 -7980
rect -16528 -8033 -16497 -7980
rect -16674 -8062 -16497 -8033
rect -16425 -7981 -16310 -7963
rect -16425 -8049 -16408 -7981
rect -16328 -8049 -16310 -7981
rect -16425 -8069 -16310 -8049
rect -16786 -8152 -16146 -8130
rect -16786 -8207 -16226 -8152
rect -16161 -8207 -16146 -8152
rect -16786 -8226 -16146 -8207
rect -16786 -8260 -16720 -8226
rect -17434 -8423 -17400 -8407
rect -17346 -8301 -17312 -8285
rect -17346 -8423 -17312 -8407
rect -17250 -8286 -17216 -8285
rect -17250 -8423 -17216 -8407
rect -17154 -8301 -17120 -8285
rect -17154 -8423 -17120 -8421
rect -17058 -8286 -17024 -8285
rect -17058 -8423 -17024 -8407
rect -16962 -8301 -16928 -8285
rect -16962 -8423 -16928 -8421
rect -16866 -8287 -16832 -8285
rect -16866 -8423 -16832 -8407
rect -16770 -8301 -16736 -8260
rect -16770 -8423 -16736 -8421
rect -16674 -8286 -16640 -8285
rect -16674 -8423 -16640 -8407
rect -16578 -8301 -16544 -8285
rect -16578 -8423 -16544 -8421
rect -16482 -8286 -16448 -8285
rect -16482 -8423 -16448 -8407
rect -16386 -8301 -16352 -8285
rect -16386 -8423 -16352 -8421
rect -16290 -8286 -16256 -8285
rect -16290 -8423 -16256 -8407
rect -16194 -8301 -16160 -8285
rect -16194 -8423 -16160 -8407
rect -16106 -8301 -16072 -7922
rect -16025 -7932 -15916 -7917
rect -16025 -8072 -16006 -7932
rect -15933 -8072 -15916 -7932
rect -16025 -8089 -15916 -8072
rect -16106 -8423 -16072 -8407
rect -15875 -8301 -15841 -7917
rect -15739 -7988 -15518 -7961
rect -15739 -8041 -15689 -7988
rect -15556 -8041 -15518 -7988
rect -15739 -8179 -15518 -8041
rect -15739 -8224 -15694 -8179
rect -15564 -8224 -15518 -8179
rect -15739 -8251 -15518 -8224
rect -15438 -8187 -15273 -7917
rect -15438 -8232 -15411 -8187
rect -15281 -8232 -15273 -8187
rect -15438 -8249 -15273 -8232
rect -15227 -8130 -15161 -7830
rect -14547 -7845 -14513 -7787
rect -15115 -7863 -14513 -7845
rect -15115 -7908 -15088 -7863
rect -14958 -7908 -14513 -7863
rect -14143 -7261 -14109 -7245
rect -14143 -7848 -14109 -7787
rect -14055 -7261 -14021 -7245
rect -14055 -7803 -14021 -7787
rect -13959 -7261 -13925 -7245
rect -13959 -7803 -13925 -7787
rect -13863 -7261 -13829 -7245
rect -13863 -7803 -13829 -7787
rect -13767 -7261 -13733 -7245
rect -13767 -7803 -13733 -7787
rect -13671 -7261 -13637 -7245
rect -13671 -7803 -13637 -7787
rect -13575 -7261 -13541 -7245
rect -13575 -7803 -13541 -7787
rect -13479 -7261 -13445 -7245
rect -13479 -7830 -13445 -7787
rect -13383 -7261 -13349 -7245
rect -13383 -7803 -13349 -7787
rect -13287 -7261 -13253 -7245
rect -13287 -7803 -13253 -7787
rect -13191 -7261 -13157 -7245
rect -13191 -7803 -13157 -7787
rect -13095 -7261 -13061 -7245
rect -13095 -7803 -13061 -7787
rect -12999 -7261 -12965 -7245
rect -12999 -7803 -12965 -7787
rect -12903 -7261 -12869 -7245
rect -12903 -7803 -12869 -7787
rect -12815 -7261 -12781 -7245
rect -14143 -7858 -13541 -7848
rect -15115 -7922 -14513 -7908
rect -15115 -7980 -14938 -7922
rect -15115 -8033 -15083 -7980
rect -14969 -8033 -14938 -7980
rect -15115 -8062 -14938 -8033
rect -14866 -7981 -14751 -7963
rect -14866 -8049 -14849 -7981
rect -14769 -8049 -14751 -7981
rect -14866 -8069 -14751 -8049
rect -15227 -8152 -14587 -8130
rect -15227 -8207 -14667 -8152
rect -14602 -8207 -14587 -8152
rect -15227 -8226 -14587 -8207
rect -15227 -8260 -15161 -8226
rect -15875 -8423 -15841 -8407
rect -15787 -8301 -15753 -8285
rect -15787 -8423 -15753 -8407
rect -15691 -8286 -15657 -8285
rect -15691 -8423 -15657 -8407
rect -15595 -8301 -15561 -8285
rect -15595 -8423 -15561 -8421
rect -15499 -8286 -15465 -8285
rect -15499 -8423 -15465 -8407
rect -15403 -8301 -15369 -8285
rect -15403 -8423 -15369 -8421
rect -15307 -8287 -15273 -8285
rect -15307 -8423 -15273 -8407
rect -15211 -8301 -15177 -8260
rect -15211 -8423 -15177 -8421
rect -15115 -8286 -15081 -8285
rect -15115 -8423 -15081 -8407
rect -15019 -8301 -14985 -8285
rect -15019 -8423 -14985 -8421
rect -14923 -8286 -14889 -8285
rect -14923 -8423 -14889 -8407
rect -14827 -8301 -14793 -8285
rect -14827 -8423 -14793 -8421
rect -14731 -8286 -14697 -8285
rect -14731 -8423 -14697 -8407
rect -14635 -8301 -14601 -8285
rect -14635 -8423 -14601 -8407
rect -14547 -8301 -14513 -7922
rect -14290 -7887 -14205 -7864
rect -14290 -7997 -14272 -7887
rect -14225 -7997 -14205 -7887
rect -14290 -8017 -14205 -7997
rect -14143 -7903 -13687 -7858
rect -13557 -7903 -13541 -7858
rect -14143 -7917 -13541 -7903
rect -14547 -8423 -14513 -8407
rect -14143 -8301 -14109 -7917
rect -14007 -7988 -13786 -7961
rect -14007 -8041 -13957 -7988
rect -13824 -8041 -13786 -7988
rect -14007 -8179 -13786 -8041
rect -14007 -8224 -13962 -8179
rect -13832 -8224 -13786 -8179
rect -14007 -8251 -13786 -8224
rect -13706 -8187 -13541 -7917
rect -13706 -8232 -13679 -8187
rect -13549 -8232 -13541 -8187
rect -13706 -8249 -13541 -8232
rect -13495 -8130 -13429 -7830
rect -12815 -7845 -12781 -7787
rect -13383 -7863 -12781 -7845
rect -13383 -7908 -13356 -7863
rect -13226 -7908 -12781 -7863
rect -13383 -7922 -12781 -7908
rect -12584 -7261 -12550 -7245
rect -12584 -7848 -12550 -7787
rect -12496 -7261 -12462 -7245
rect -12496 -7803 -12462 -7787
rect -12400 -7261 -12366 -7245
rect -12400 -7803 -12366 -7787
rect -12304 -7261 -12270 -7245
rect -12304 -7803 -12270 -7787
rect -12208 -7261 -12174 -7245
rect -12208 -7803 -12174 -7787
rect -12112 -7261 -12078 -7245
rect -12112 -7803 -12078 -7787
rect -12016 -7261 -11982 -7245
rect -12016 -7803 -11982 -7787
rect -11920 -7261 -11886 -7245
rect -11920 -7830 -11886 -7787
rect -11824 -7261 -11790 -7245
rect -11824 -7803 -11790 -7787
rect -11728 -7261 -11694 -7245
rect -11728 -7803 -11694 -7787
rect -11632 -7261 -11598 -7245
rect -11632 -7803 -11598 -7787
rect -11536 -7261 -11502 -7245
rect -11536 -7803 -11502 -7787
rect -11440 -7261 -11406 -7245
rect -11440 -7803 -11406 -7787
rect -11344 -7261 -11310 -7245
rect -11344 -7803 -11310 -7787
rect -11256 -7261 -11222 -7245
rect -12584 -7858 -11982 -7848
rect -12584 -7903 -12128 -7858
rect -11998 -7903 -11982 -7858
rect -12584 -7917 -11982 -7903
rect -13383 -7980 -13206 -7922
rect -13383 -8033 -13351 -7980
rect -13237 -8033 -13206 -7980
rect -13383 -8062 -13206 -8033
rect -13134 -7981 -13019 -7963
rect -13134 -8049 -13117 -7981
rect -13037 -8049 -13019 -7981
rect -13134 -8069 -13019 -8049
rect -13495 -8152 -12855 -8130
rect -13495 -8207 -12935 -8152
rect -12870 -8207 -12855 -8152
rect -13495 -8226 -12855 -8207
rect -13495 -8260 -13429 -8226
rect -14143 -8423 -14109 -8407
rect -14055 -8301 -14021 -8285
rect -14055 -8423 -14021 -8407
rect -13959 -8286 -13925 -8285
rect -13959 -8423 -13925 -8407
rect -13863 -8301 -13829 -8285
rect -13863 -8423 -13829 -8421
rect -13767 -8286 -13733 -8285
rect -13767 -8423 -13733 -8407
rect -13671 -8301 -13637 -8285
rect -13671 -8423 -13637 -8421
rect -13575 -8287 -13541 -8285
rect -13575 -8423 -13541 -8407
rect -13479 -8301 -13445 -8260
rect -13479 -8423 -13445 -8421
rect -13383 -8286 -13349 -8285
rect -13383 -8423 -13349 -8407
rect -13287 -8301 -13253 -8285
rect -13287 -8423 -13253 -8421
rect -13191 -8286 -13157 -8285
rect -13191 -8423 -13157 -8407
rect -13095 -8301 -13061 -8285
rect -13095 -8423 -13061 -8421
rect -12999 -8286 -12965 -8285
rect -12999 -8423 -12965 -8407
rect -12903 -8301 -12869 -8285
rect -12903 -8423 -12869 -8407
rect -12815 -8301 -12781 -7922
rect -12734 -7932 -12625 -7917
rect -12734 -8072 -12715 -7932
rect -12642 -8072 -12625 -7932
rect -12734 -8089 -12625 -8072
rect -12815 -8423 -12781 -8407
rect -12584 -8301 -12550 -7917
rect -12448 -7988 -12227 -7961
rect -12448 -8041 -12398 -7988
rect -12265 -8041 -12227 -7988
rect -12448 -8179 -12227 -8041
rect -12448 -8224 -12403 -8179
rect -12273 -8224 -12227 -8179
rect -12448 -8251 -12227 -8224
rect -12147 -8187 -11982 -7917
rect -12147 -8232 -12120 -8187
rect -11990 -8232 -11982 -8187
rect -12147 -8249 -11982 -8232
rect -11936 -8130 -11870 -7830
rect -11256 -7845 -11222 -7787
rect -11824 -7863 -11222 -7845
rect -11824 -7908 -11797 -7863
rect -11667 -7908 -11222 -7863
rect -10852 -7261 -10818 -7245
rect -10852 -7848 -10818 -7787
rect -10764 -7261 -10730 -7245
rect -10764 -7803 -10730 -7787
rect -10668 -7261 -10634 -7245
rect -10668 -7803 -10634 -7787
rect -10572 -7261 -10538 -7245
rect -10572 -7803 -10538 -7787
rect -10476 -7261 -10442 -7245
rect -10476 -7803 -10442 -7787
rect -10380 -7261 -10346 -7245
rect -10380 -7803 -10346 -7787
rect -10284 -7261 -10250 -7245
rect -10284 -7803 -10250 -7787
rect -10188 -7261 -10154 -7245
rect -10188 -7830 -10154 -7787
rect -10092 -7261 -10058 -7245
rect -10092 -7803 -10058 -7787
rect -9996 -7261 -9962 -7245
rect -9996 -7803 -9962 -7787
rect -9900 -7261 -9866 -7245
rect -9900 -7803 -9866 -7787
rect -9804 -7261 -9770 -7245
rect -9804 -7803 -9770 -7787
rect -9708 -7261 -9674 -7245
rect -9708 -7803 -9674 -7787
rect -9612 -7261 -9578 -7245
rect -9612 -7803 -9578 -7787
rect -9524 -7261 -9490 -7245
rect -10852 -7858 -10250 -7848
rect -11824 -7922 -11222 -7908
rect -11824 -7980 -11647 -7922
rect -11824 -8033 -11792 -7980
rect -11678 -8033 -11647 -7980
rect -11824 -8062 -11647 -8033
rect -11575 -7981 -11460 -7963
rect -11575 -8049 -11558 -7981
rect -11478 -8049 -11460 -7981
rect -11575 -8069 -11460 -8049
rect -11936 -8152 -11296 -8130
rect -11936 -8207 -11376 -8152
rect -11311 -8207 -11296 -8152
rect -11936 -8226 -11296 -8207
rect -11936 -8260 -11870 -8226
rect -12584 -8423 -12550 -8407
rect -12496 -8301 -12462 -8285
rect -12496 -8423 -12462 -8407
rect -12400 -8286 -12366 -8285
rect -12400 -8423 -12366 -8407
rect -12304 -8301 -12270 -8285
rect -12304 -8423 -12270 -8421
rect -12208 -8286 -12174 -8285
rect -12208 -8423 -12174 -8407
rect -12112 -8301 -12078 -8285
rect -12112 -8423 -12078 -8421
rect -12016 -8287 -11982 -8285
rect -12016 -8423 -11982 -8407
rect -11920 -8301 -11886 -8260
rect -11920 -8423 -11886 -8421
rect -11824 -8286 -11790 -8285
rect -11824 -8423 -11790 -8407
rect -11728 -8301 -11694 -8285
rect -11728 -8423 -11694 -8421
rect -11632 -8286 -11598 -8285
rect -11632 -8423 -11598 -8407
rect -11536 -8301 -11502 -8285
rect -11536 -8423 -11502 -8421
rect -11440 -8286 -11406 -8285
rect -11440 -8423 -11406 -8407
rect -11344 -8301 -11310 -8285
rect -11344 -8423 -11310 -8407
rect -11256 -8301 -11222 -7922
rect -10999 -7887 -10914 -7864
rect -10999 -7997 -10981 -7887
rect -10934 -7997 -10914 -7887
rect -10999 -8017 -10914 -7997
rect -10852 -7903 -10396 -7858
rect -10266 -7903 -10250 -7858
rect -10852 -7917 -10250 -7903
rect -11256 -8423 -11222 -8407
rect -10852 -8301 -10818 -7917
rect -10716 -7988 -10495 -7961
rect -10716 -8041 -10666 -7988
rect -10533 -8041 -10495 -7988
rect -10716 -8179 -10495 -8041
rect -10716 -8224 -10671 -8179
rect -10541 -8224 -10495 -8179
rect -10716 -8251 -10495 -8224
rect -10415 -8187 -10250 -7917
rect -10415 -8232 -10388 -8187
rect -10258 -8232 -10250 -8187
rect -10415 -8249 -10250 -8232
rect -10204 -8130 -10138 -7830
rect -9524 -7845 -9490 -7787
rect -10092 -7863 -9490 -7845
rect -10092 -7908 -10065 -7863
rect -9935 -7908 -9490 -7863
rect -10092 -7922 -9490 -7908
rect -9293 -7261 -9259 -7245
rect -9293 -7848 -9259 -7787
rect -9205 -7261 -9171 -7245
rect -9205 -7803 -9171 -7787
rect -9109 -7261 -9075 -7245
rect -9109 -7803 -9075 -7787
rect -9013 -7261 -8979 -7245
rect -9013 -7803 -8979 -7787
rect -8917 -7261 -8883 -7245
rect -8917 -7803 -8883 -7787
rect -8821 -7261 -8787 -7245
rect -8821 -7803 -8787 -7787
rect -8725 -7261 -8691 -7245
rect -8725 -7803 -8691 -7787
rect -8629 -7261 -8595 -7245
rect -8629 -7830 -8595 -7787
rect -8533 -7261 -8499 -7245
rect -8533 -7803 -8499 -7787
rect -8437 -7261 -8403 -7245
rect -8437 -7803 -8403 -7787
rect -8341 -7261 -8307 -7245
rect -8341 -7803 -8307 -7787
rect -8245 -7261 -8211 -7245
rect -8245 -7803 -8211 -7787
rect -8149 -7261 -8115 -7245
rect -8149 -7803 -8115 -7787
rect -8053 -7261 -8019 -7245
rect -8053 -7803 -8019 -7787
rect -7965 -7261 -7931 -7245
rect 7298 -7254 7372 -7241
rect 7298 -7270 7406 -7254
rect 7756 -6478 7790 -6462
rect 7756 -7270 7790 -7254
rect 8246 -6478 8354 -6462
rect 8246 -6490 8320 -6478
rect 8281 -7241 8320 -6490
rect 8246 -7254 8320 -7241
rect 8246 -7270 8354 -7254
rect 8704 -6478 8738 -6462
rect 8704 -7270 8738 -7254
rect 9182 -6478 9290 -6462
rect 9182 -6490 9256 -6478
rect 9217 -7241 9256 -6490
rect 9182 -7254 9256 -7241
rect 9182 -7270 9290 -7254
rect 9640 -6478 9674 -6462
rect 9640 -7270 9674 -7254
rect 10113 -6478 10221 -6462
rect 10113 -6490 10187 -6478
rect 10148 -7241 10187 -6490
rect 10113 -7254 10187 -7241
rect 10113 -7270 10221 -7254
rect 10571 -6478 10605 -6462
rect 10571 -7270 10605 -7254
rect 11040 -6478 11148 -6462
rect 11040 -6490 11114 -6478
rect 11075 -7241 11114 -6490
rect 11040 -7254 11114 -7241
rect 11040 -7270 11148 -7254
rect 11498 -6478 11532 -6462
rect 11783 -6804 12203 -6784
rect 11783 -6855 11811 -6804
rect 12168 -6855 12203 -6804
rect 11783 -6874 12203 -6855
rect 11785 -6959 11819 -6874
rect 11785 -7207 11819 -7191
rect 11881 -6959 11915 -6943
rect 11881 -7207 11915 -7191
rect 11977 -6959 12011 -6874
rect 11977 -7207 12011 -7191
rect 12073 -6959 12107 -6943
rect 12073 -7207 12107 -7191
rect 12169 -6959 12203 -6874
rect 12169 -7207 12203 -7191
rect 12265 -6959 12299 -6943
rect 12265 -7207 12299 -7191
rect 12361 -6959 12395 -6943
rect 12361 -7207 12395 -7191
rect 12457 -6959 12491 -6943
rect 12457 -7207 12491 -7191
rect 12553 -6959 12587 -6943
rect 12553 -7207 12587 -7191
rect 12649 -6959 12683 -6943
rect 12649 -7207 12683 -7191
rect 12745 -6959 12779 -6943
rect 12970 -7025 12986 -6991
rect 13077 -7025 13093 -6991
rect 12745 -7207 12779 -7191
rect 12826 -7111 12876 -7094
rect 12919 -7097 12929 -7063
rect 13125 -7097 13141 -7063
rect 11498 -7270 11532 -7254
rect 12154 -7287 12170 -7253
rect 12204 -7287 12220 -7253
rect 12826 -7337 12842 -7111
rect 12919 -7193 12935 -7159
rect 13129 -7193 13147 -7159
rect 12919 -7289 12929 -7255
rect 13125 -7289 13141 -7255
rect -9293 -7858 -8691 -7848
rect -9293 -7903 -8837 -7858
rect -8707 -7903 -8691 -7858
rect -9293 -7917 -8691 -7903
rect -10092 -7980 -9915 -7922
rect -10092 -8033 -10060 -7980
rect -9946 -8033 -9915 -7980
rect -10092 -8062 -9915 -8033
rect -9843 -7981 -9728 -7963
rect -9843 -8049 -9826 -7981
rect -9746 -8049 -9728 -7981
rect -9843 -8069 -9728 -8049
rect -10204 -8152 -9564 -8130
rect -10204 -8207 -9644 -8152
rect -9579 -8207 -9564 -8152
rect -10204 -8226 -9564 -8207
rect -10204 -8260 -10138 -8226
rect -10852 -8423 -10818 -8407
rect -10764 -8301 -10730 -8285
rect -10764 -8423 -10730 -8407
rect -10668 -8286 -10634 -8285
rect -10668 -8423 -10634 -8407
rect -10572 -8301 -10538 -8285
rect -10572 -8423 -10538 -8421
rect -10476 -8286 -10442 -8285
rect -10476 -8423 -10442 -8407
rect -10380 -8301 -10346 -8285
rect -10380 -8423 -10346 -8421
rect -10284 -8287 -10250 -8285
rect -10284 -8423 -10250 -8407
rect -10188 -8301 -10154 -8260
rect -10188 -8423 -10154 -8421
rect -10092 -8286 -10058 -8285
rect -10092 -8423 -10058 -8407
rect -9996 -8301 -9962 -8285
rect -9996 -8423 -9962 -8421
rect -9900 -8286 -9866 -8285
rect -9900 -8423 -9866 -8407
rect -9804 -8301 -9770 -8285
rect -9804 -8423 -9770 -8421
rect -9708 -8286 -9674 -8285
rect -9708 -8423 -9674 -8407
rect -9612 -8301 -9578 -8285
rect -9612 -8423 -9578 -8407
rect -9524 -8301 -9490 -7922
rect -9443 -7932 -9334 -7917
rect -9443 -8072 -9424 -7932
rect -9351 -8072 -9334 -7932
rect -9443 -8089 -9334 -8072
rect -9524 -8423 -9490 -8407
rect -9293 -8301 -9259 -7917
rect -9157 -7988 -8936 -7961
rect -9157 -8041 -9107 -7988
rect -8974 -8041 -8936 -7988
rect -9157 -8179 -8936 -8041
rect -9157 -8224 -9112 -8179
rect -8982 -8224 -8936 -8179
rect -9157 -8251 -8936 -8224
rect -8856 -8187 -8691 -7917
rect -8856 -8232 -8829 -8187
rect -8699 -8232 -8691 -8187
rect -8856 -8249 -8691 -8232
rect -8645 -8130 -8579 -7830
rect -7965 -7845 -7931 -7787
rect -8533 -7863 -7931 -7845
rect -8533 -7908 -8506 -7863
rect -8376 -7908 -7931 -7863
rect -8533 -7922 -7931 -7908
rect -8533 -7980 -8356 -7922
rect -8533 -8033 -8501 -7980
rect -8387 -8033 -8356 -7980
rect -8533 -8062 -8356 -8033
rect -8284 -7981 -8169 -7963
rect -8284 -8049 -8267 -7981
rect -8187 -8049 -8169 -7981
rect -8284 -8069 -8169 -8049
rect -8645 -8152 -8005 -8130
rect -8645 -8207 -8085 -8152
rect -8020 -8207 -8005 -8152
rect -8645 -8226 -8005 -8207
rect -8645 -8260 -8579 -8226
rect -9293 -8423 -9259 -8407
rect -9205 -8301 -9171 -8285
rect -9205 -8423 -9171 -8407
rect -9109 -8286 -9075 -8285
rect -9109 -8423 -9075 -8407
rect -9013 -8301 -8979 -8285
rect -9013 -8423 -8979 -8421
rect -8917 -8286 -8883 -8285
rect -8917 -8423 -8883 -8407
rect -8821 -8301 -8787 -8285
rect -8821 -8423 -8787 -8421
rect -8725 -8287 -8691 -8285
rect -8725 -8423 -8691 -8407
rect -8629 -8301 -8595 -8260
rect -8629 -8423 -8595 -8421
rect -8533 -8286 -8499 -8285
rect -8533 -8423 -8499 -8407
rect -8437 -8301 -8403 -8285
rect -8437 -8423 -8403 -8421
rect -8341 -8286 -8307 -8285
rect -8341 -8423 -8307 -8407
rect -8245 -8301 -8211 -8285
rect -8245 -8423 -8211 -8421
rect -8149 -8286 -8115 -8285
rect -8149 -8423 -8115 -8407
rect -8053 -8301 -8019 -8285
rect -8053 -8423 -8019 -8407
rect -7965 -8301 -7931 -7922
rect 7298 -7406 7406 -7390
rect 7298 -7419 7372 -7406
rect 7333 -8170 7372 -7419
rect 7298 -8182 7372 -8170
rect 7298 -8198 7406 -8182
rect 7756 -7406 7790 -7390
rect 7756 -8198 7790 -8182
rect 8246 -7406 8354 -7390
rect 8246 -7419 8320 -7406
rect 8281 -8170 8320 -7419
rect 8246 -8182 8320 -8170
rect 8246 -8198 8354 -8182
rect 8704 -7406 8738 -7390
rect 8704 -8198 8738 -8182
rect 9182 -7406 9290 -7390
rect 9182 -7419 9256 -7406
rect 9217 -8170 9256 -7419
rect 9182 -8182 9256 -8170
rect 9182 -8198 9290 -8182
rect 9640 -7406 9674 -7390
rect 9640 -8198 9674 -8182
rect 10113 -7405 10221 -7389
rect 10113 -7418 10187 -7405
rect 10148 -8169 10187 -7418
rect 10113 -8181 10187 -8169
rect 10113 -8197 10221 -8181
rect 10571 -7405 10605 -7389
rect 10571 -8197 10605 -8181
rect 11040 -7406 11148 -7390
rect 11040 -7419 11114 -7406
rect 11075 -8170 11114 -7419
rect 11040 -8182 11114 -8170
rect 7298 -8201 7403 -8198
rect 8246 -8201 8351 -8198
rect 9182 -8201 9287 -8198
rect 10113 -8200 10218 -8197
rect 11040 -8198 11148 -8182
rect 11498 -7406 11532 -7390
rect 12297 -7392 12313 -7358
rect 12347 -7392 12363 -7358
rect 12169 -7448 12203 -7432
rect 12169 -7696 12203 -7624
rect 12265 -7448 12299 -7432
rect 12265 -7640 12299 -7624
rect 12361 -7448 12395 -7432
rect 12826 -7557 12876 -7337
rect 12919 -7385 12935 -7351
rect 13129 -7385 13147 -7351
rect 12919 -7547 12935 -7513
rect 13111 -7547 13127 -7513
rect 12826 -7591 12842 -7557
rect 12826 -7607 12876 -7591
rect 12361 -7696 12395 -7624
rect 12919 -7635 12935 -7601
rect 13111 -7635 13127 -7601
rect 12157 -7707 12407 -7696
rect 12157 -7768 12183 -7707
rect 12382 -7768 12407 -7707
rect 12938 -7737 12954 -7703
rect 13086 -7737 13102 -7703
rect 12157 -7780 12407 -7768
rect 11498 -8198 11532 -8182
rect 11040 -8201 11145 -8198
rect -7965 -8423 -7931 -8407
rect -20644 -8495 -19442 -8473
rect -20644 -8541 -20603 -8495
rect -19480 -8541 -19442 -8495
rect -20644 -8564 -19442 -8541
rect -19085 -8495 -17883 -8473
rect -19085 -8541 -19044 -8495
rect -17921 -8541 -17883 -8495
rect -19085 -8564 -17883 -8541
rect -17353 -8495 -16151 -8473
rect -17353 -8541 -17312 -8495
rect -16189 -8541 -16151 -8495
rect -17353 -8564 -16151 -8541
rect -15794 -8495 -14592 -8473
rect -15794 -8541 -15753 -8495
rect -14630 -8541 -14592 -8495
rect -15794 -8564 -14592 -8541
rect -14062 -8495 -12860 -8473
rect -14062 -8541 -14021 -8495
rect -12898 -8541 -12860 -8495
rect -14062 -8564 -12860 -8541
rect -12503 -8495 -11301 -8473
rect -12503 -8541 -12462 -8495
rect -11339 -8541 -11301 -8495
rect -12503 -8564 -11301 -8541
rect -10771 -8495 -9569 -8473
rect -10771 -8541 -10730 -8495
rect -9607 -8541 -9569 -8495
rect -10771 -8564 -9569 -8541
rect -9212 -8495 -8010 -8473
rect -9212 -8541 -9171 -8495
rect -8048 -8541 -8010 -8495
rect -9212 -8564 -8010 -8541
rect 7182 -8554 7198 -8520
rect 7232 -8554 7248 -8520
rect 7374 -8554 7390 -8520
rect 7424 -8554 7440 -8520
rect 7566 -8554 7582 -8520
rect 7616 -8554 7632 -8520
rect 7758 -8554 7774 -8520
rect 7808 -8554 7824 -8520
rect 8130 -8554 8146 -8520
rect 8180 -8554 8196 -8520
rect 8322 -8554 8338 -8520
rect 8372 -8554 8388 -8520
rect 8514 -8554 8530 -8520
rect 8564 -8554 8580 -8520
rect 8706 -8554 8722 -8520
rect 8756 -8554 8772 -8520
rect 9066 -8554 9082 -8520
rect 9116 -8554 9132 -8520
rect 9258 -8554 9274 -8520
rect 9308 -8554 9324 -8520
rect 9450 -8554 9466 -8520
rect 9500 -8554 9516 -8520
rect 9642 -8554 9658 -8520
rect 9692 -8554 9708 -8520
rect 9997 -8553 10013 -8519
rect 10047 -8553 10063 -8519
rect 10189 -8553 10205 -8519
rect 10239 -8553 10255 -8519
rect 10381 -8553 10397 -8519
rect 10431 -8553 10447 -8519
rect 10573 -8553 10589 -8519
rect 10623 -8553 10639 -8519
rect 10924 -8554 10940 -8520
rect 10974 -8554 10990 -8520
rect 11116 -8554 11132 -8520
rect 11166 -8554 11182 -8520
rect 11308 -8554 11324 -8520
rect 11358 -8554 11374 -8520
rect 11500 -8554 11516 -8520
rect 11550 -8554 11566 -8520
rect 7150 -8613 7184 -8597
rect 7246 -8608 7280 -8597
rect -23536 -8650 -23520 -8616
rect -23429 -8650 -23413 -8616
rect -21799 -8650 -21783 -8616
rect -21692 -8650 -21676 -8616
rect -24384 -8716 -24368 -8669
rect -23799 -8716 -23775 -8669
rect -23680 -8736 -23630 -8719
rect -23587 -8722 -23577 -8688
rect -23381 -8722 -23365 -8688
rect -22648 -8716 -22632 -8669
rect -22063 -8716 -22039 -8669
rect -24384 -8788 -24350 -8778
rect -24384 -9000 -24350 -8984
rect -24288 -8794 -24254 -8778
rect -24288 -9000 -24254 -8990
rect -24192 -8788 -24158 -8778
rect -24192 -9000 -24158 -8984
rect -24096 -8794 -24062 -8778
rect -24096 -9000 -24062 -8990
rect -24000 -8788 -23966 -8778
rect -24000 -9000 -23966 -8984
rect -23904 -8794 -23870 -8778
rect -23904 -9000 -23870 -8990
rect -23808 -8788 -23774 -8778
rect -23808 -9000 -23774 -8984
rect -23680 -8962 -23664 -8736
rect -21943 -8736 -21893 -8719
rect -21850 -8722 -21840 -8688
rect -21644 -8722 -21628 -8688
rect -23587 -8818 -23571 -8784
rect -23377 -8818 -23359 -8784
rect -22648 -8788 -22614 -8778
rect -23587 -8914 -23577 -8880
rect -23381 -8914 -23365 -8880
rect -24335 -9078 -24318 -9043
rect -24284 -9078 -24268 -9043
rect -24046 -9049 -24029 -9043
rect -24234 -9078 -24029 -9049
rect -23995 -9078 -23979 -9043
rect -24335 -9284 -24292 -9078
rect -24234 -9083 -23979 -9078
rect -24234 -9167 -24200 -9083
rect -24166 -9172 -24150 -9138
rect -23774 -9172 -23758 -9138
rect -24234 -9218 -24200 -9202
rect -23680 -9182 -23630 -8962
rect -23587 -9010 -23571 -8976
rect -23377 -9010 -23359 -8976
rect -22648 -9000 -22614 -8984
rect -22552 -8794 -22518 -8778
rect -22552 -9000 -22518 -8990
rect -22456 -8788 -22422 -8778
rect -22456 -9000 -22422 -8984
rect -22360 -8794 -22326 -8778
rect -22360 -9000 -22326 -8990
rect -22264 -8788 -22230 -8778
rect -22264 -9000 -22230 -8984
rect -22168 -8794 -22134 -8778
rect -22168 -9000 -22134 -8990
rect -22072 -8788 -22038 -8778
rect -22072 -9000 -22038 -8984
rect -21943 -8962 -21927 -8736
rect -21850 -8818 -21834 -8784
rect -21640 -8818 -21622 -8784
rect -21850 -8914 -21840 -8880
rect -21644 -8914 -21628 -8880
rect -20518 -8884 -20502 -8837
rect -19933 -8884 -19909 -8837
rect -19409 -8884 -19393 -8837
rect -18824 -8884 -18800 -8837
rect -18527 -8884 -18511 -8837
rect -17942 -8884 -17918 -8837
rect -17227 -8884 -17211 -8837
rect -16642 -8884 -16618 -8837
rect -16118 -8884 -16102 -8837
rect -15533 -8884 -15509 -8837
rect -15236 -8884 -15220 -8837
rect -14651 -8884 -14627 -8837
rect -13936 -8884 -13920 -8837
rect -13351 -8884 -13327 -8837
rect -12827 -8884 -12811 -8837
rect -12242 -8884 -12218 -8837
rect -11945 -8884 -11929 -8837
rect -11360 -8884 -11336 -8837
rect -10645 -8884 -10629 -8837
rect -10060 -8884 -10036 -8837
rect -9536 -8884 -9520 -8837
rect -8951 -8884 -8927 -8837
rect -8654 -8884 -8638 -8837
rect -8069 -8884 -8045 -8837
rect 7150 -8927 7184 -8911
rect 7246 -8927 7280 -8911
rect 7342 -8613 7376 -8597
rect 7342 -8927 7376 -8911
rect 7438 -8608 7472 -8597
rect 7534 -8613 7568 -8597
rect 7438 -8927 7472 -8911
rect 7534 -8927 7568 -8911
rect 7630 -8608 7664 -8597
rect 7726 -8613 7760 -8597
rect 7630 -8927 7664 -8911
rect 7726 -8927 7760 -8911
rect 7822 -8608 7856 -8597
rect 7918 -8613 7952 -8597
rect 7822 -8927 7856 -8911
rect 7918 -8927 7952 -8911
rect 8098 -8613 8132 -8597
rect 8194 -8608 8228 -8597
rect 8098 -8927 8132 -8911
rect 8194 -8927 8228 -8911
rect 8290 -8613 8324 -8597
rect 8290 -8927 8324 -8911
rect 8386 -8608 8420 -8597
rect 8482 -8613 8516 -8597
rect 8386 -8927 8420 -8911
rect 8482 -8927 8516 -8911
rect 8578 -8608 8612 -8597
rect 8674 -8613 8708 -8597
rect 8578 -8927 8612 -8911
rect 8674 -8927 8708 -8911
rect 8770 -8608 8804 -8597
rect 8866 -8613 8900 -8597
rect 8770 -8927 8804 -8911
rect 8866 -8927 8900 -8911
rect 9034 -8613 9068 -8597
rect 9130 -8608 9164 -8597
rect 9034 -8927 9068 -8911
rect 9130 -8927 9164 -8911
rect 9226 -8613 9260 -8597
rect 9226 -8927 9260 -8911
rect 9322 -8608 9356 -8597
rect 9418 -8613 9452 -8597
rect 9322 -8927 9356 -8911
rect 9418 -8927 9452 -8911
rect 9514 -8608 9548 -8597
rect 9610 -8613 9644 -8597
rect 9514 -8927 9548 -8911
rect 9610 -8927 9644 -8911
rect 9706 -8608 9740 -8597
rect 9802 -8613 9836 -8597
rect 9706 -8927 9740 -8911
rect 9802 -8927 9836 -8911
rect 9965 -8612 9999 -8596
rect 10061 -8607 10095 -8596
rect 9965 -8926 9999 -8910
rect 10061 -8926 10095 -8910
rect 10157 -8612 10191 -8596
rect 10157 -8926 10191 -8910
rect 10253 -8607 10287 -8596
rect 10349 -8612 10383 -8596
rect 10253 -8926 10287 -8910
rect 10349 -8926 10383 -8910
rect 10445 -8607 10479 -8596
rect 10541 -8612 10575 -8596
rect 10445 -8926 10479 -8910
rect 10541 -8926 10575 -8910
rect 10637 -8607 10671 -8596
rect 10733 -8612 10767 -8596
rect 10637 -8926 10671 -8910
rect 10733 -8926 10767 -8910
rect 10892 -8613 10926 -8597
rect 10988 -8608 11022 -8597
rect 10892 -8927 10926 -8911
rect 10988 -8927 11022 -8911
rect 11084 -8613 11118 -8597
rect 11084 -8927 11118 -8911
rect 11180 -8608 11214 -8597
rect 11276 -8613 11310 -8597
rect 11180 -8927 11214 -8911
rect 11276 -8927 11310 -8911
rect 11372 -8608 11406 -8597
rect 11468 -8613 11502 -8597
rect 11372 -8927 11406 -8911
rect 11468 -8927 11502 -8911
rect 11564 -8608 11598 -8597
rect 11660 -8613 11694 -8597
rect 11564 -8927 11598 -8911
rect 11660 -8927 11694 -8911
rect -22599 -9078 -22582 -9043
rect -22548 -9078 -22532 -9043
rect -22310 -9049 -22293 -9043
rect -22498 -9078 -22293 -9049
rect -22259 -9078 -22243 -9043
rect -23587 -9172 -23571 -9138
rect -23395 -9172 -23379 -9138
rect -23680 -9216 -23664 -9182
rect -23680 -9232 -23630 -9216
rect -23587 -9260 -23571 -9226
rect -23395 -9260 -23379 -9226
rect -22599 -9284 -22556 -9078
rect -22498 -9083 -22243 -9078
rect -22498 -9167 -22464 -9083
rect -22430 -9172 -22414 -9138
rect -22038 -9172 -22022 -9138
rect -22498 -9218 -22464 -9202
rect -21943 -9182 -21893 -8962
rect -20518 -8956 -20484 -8946
rect -21850 -9010 -21834 -8976
rect -21640 -9010 -21622 -8976
rect -21850 -9172 -21834 -9138
rect -21658 -9172 -21642 -9138
rect -20518 -9168 -20484 -9152
rect -20422 -8962 -20388 -8946
rect -20422 -9168 -20388 -9158
rect -20326 -8956 -20292 -8946
rect -20326 -9168 -20292 -9152
rect -20230 -8962 -20196 -8946
rect -20230 -9168 -20196 -9158
rect -20134 -8956 -20100 -8946
rect -20134 -9168 -20100 -9152
rect -20038 -8962 -20004 -8946
rect -20038 -9168 -20004 -9158
rect -19942 -8956 -19908 -8946
rect -19942 -9168 -19908 -9152
rect -19409 -8956 -19375 -8946
rect -19409 -9168 -19375 -9152
rect -19313 -8962 -19279 -8946
rect -19313 -9168 -19279 -9158
rect -19217 -8956 -19183 -8946
rect -19217 -9168 -19183 -9152
rect -19121 -8962 -19087 -8946
rect -19121 -9168 -19087 -9158
rect -19025 -8956 -18991 -8946
rect -19025 -9168 -18991 -9152
rect -18929 -8962 -18895 -8946
rect -18929 -9168 -18895 -9158
rect -18833 -8956 -18799 -8946
rect -18833 -9168 -18799 -9152
rect -18527 -8956 -18493 -8946
rect -18527 -9168 -18493 -9152
rect -18431 -8962 -18397 -8946
rect -18431 -9168 -18397 -9158
rect -18335 -8956 -18301 -8946
rect -18335 -9168 -18301 -9152
rect -18239 -8962 -18205 -8946
rect -18239 -9168 -18205 -9158
rect -18143 -8956 -18109 -8946
rect -18143 -9168 -18109 -9152
rect -18047 -8962 -18013 -8946
rect -18047 -9168 -18013 -9158
rect -17951 -8956 -17917 -8946
rect -17951 -9168 -17917 -9152
rect -17227 -8956 -17193 -8946
rect -17227 -9168 -17193 -9152
rect -17131 -8962 -17097 -8946
rect -17131 -9168 -17097 -9158
rect -17035 -8956 -17001 -8946
rect -17035 -9168 -17001 -9152
rect -16939 -8962 -16905 -8946
rect -16939 -9168 -16905 -9158
rect -16843 -8956 -16809 -8946
rect -16843 -9168 -16809 -9152
rect -16747 -8962 -16713 -8946
rect -16747 -9168 -16713 -9158
rect -16651 -8956 -16617 -8946
rect -16651 -9168 -16617 -9152
rect -16118 -8956 -16084 -8946
rect -16118 -9168 -16084 -9152
rect -16022 -8962 -15988 -8946
rect -16022 -9168 -15988 -9158
rect -15926 -8956 -15892 -8946
rect -15926 -9168 -15892 -9152
rect -15830 -8962 -15796 -8946
rect -15830 -9168 -15796 -9158
rect -15734 -8956 -15700 -8946
rect -15734 -9168 -15700 -9152
rect -15638 -8962 -15604 -8946
rect -15638 -9168 -15604 -9158
rect -15542 -8956 -15508 -8946
rect -15542 -9168 -15508 -9152
rect -15236 -8956 -15202 -8946
rect -15236 -9168 -15202 -9152
rect -15140 -8962 -15106 -8946
rect -15140 -9168 -15106 -9158
rect -15044 -8956 -15010 -8946
rect -15044 -9168 -15010 -9152
rect -14948 -8962 -14914 -8946
rect -14948 -9168 -14914 -9158
rect -14852 -8956 -14818 -8946
rect -14852 -9168 -14818 -9152
rect -14756 -8962 -14722 -8946
rect -14756 -9168 -14722 -9158
rect -14660 -8956 -14626 -8946
rect -14660 -9168 -14626 -9152
rect -13936 -8956 -13902 -8946
rect -13936 -9168 -13902 -9152
rect -13840 -8962 -13806 -8946
rect -13840 -9168 -13806 -9158
rect -13744 -8956 -13710 -8946
rect -13744 -9168 -13710 -9152
rect -13648 -8962 -13614 -8946
rect -13648 -9168 -13614 -9158
rect -13552 -8956 -13518 -8946
rect -13552 -9168 -13518 -9152
rect -13456 -8962 -13422 -8946
rect -13456 -9168 -13422 -9158
rect -13360 -8956 -13326 -8946
rect -13360 -9168 -13326 -9152
rect -12827 -8956 -12793 -8946
rect -12827 -9168 -12793 -9152
rect -12731 -8962 -12697 -8946
rect -12731 -9168 -12697 -9158
rect -12635 -8956 -12601 -8946
rect -12635 -9168 -12601 -9152
rect -12539 -8962 -12505 -8946
rect -12539 -9168 -12505 -9158
rect -12443 -8956 -12409 -8946
rect -12443 -9168 -12409 -9152
rect -12347 -8962 -12313 -8946
rect -12347 -9168 -12313 -9158
rect -12251 -8956 -12217 -8946
rect -12251 -9168 -12217 -9152
rect -11945 -8956 -11911 -8946
rect -11945 -9168 -11911 -9152
rect -11849 -8962 -11815 -8946
rect -11849 -9168 -11815 -9158
rect -11753 -8956 -11719 -8946
rect -11753 -9168 -11719 -9152
rect -11657 -8962 -11623 -8946
rect -11657 -9168 -11623 -9158
rect -11561 -8956 -11527 -8946
rect -11561 -9168 -11527 -9152
rect -11465 -8962 -11431 -8946
rect -11465 -9168 -11431 -9158
rect -11369 -8956 -11335 -8946
rect -11369 -9168 -11335 -9152
rect -10645 -8956 -10611 -8946
rect -10645 -9168 -10611 -9152
rect -10549 -8962 -10515 -8946
rect -10549 -9168 -10515 -9158
rect -10453 -8956 -10419 -8946
rect -10453 -9168 -10419 -9152
rect -10357 -8962 -10323 -8946
rect -10357 -9168 -10323 -9158
rect -10261 -8956 -10227 -8946
rect -10261 -9168 -10227 -9152
rect -10165 -8962 -10131 -8946
rect -10165 -9168 -10131 -9158
rect -10069 -8956 -10035 -8946
rect -10069 -9168 -10035 -9152
rect -9536 -8956 -9502 -8946
rect -9536 -9168 -9502 -9152
rect -9440 -8962 -9406 -8946
rect -9440 -9168 -9406 -9158
rect -9344 -8956 -9310 -8946
rect -9344 -9168 -9310 -9152
rect -9248 -8962 -9214 -8946
rect -9248 -9168 -9214 -9158
rect -9152 -8956 -9118 -8946
rect -9152 -9168 -9118 -9152
rect -9056 -8962 -9022 -8946
rect -9056 -9168 -9022 -9158
rect -8960 -8956 -8926 -8946
rect -8960 -9168 -8926 -9152
rect -8654 -8956 -8620 -8946
rect -8654 -9168 -8620 -9152
rect -8558 -8962 -8524 -8946
rect -8558 -9168 -8524 -9158
rect -8462 -8956 -8428 -8946
rect -8462 -9168 -8428 -9152
rect -8366 -8962 -8332 -8946
rect -8366 -9168 -8332 -9158
rect -8270 -8956 -8236 -8946
rect -8270 -9168 -8236 -9152
rect -8174 -8962 -8140 -8946
rect -8174 -9168 -8140 -9158
rect -8078 -8956 -8044 -8946
rect 7373 -9015 7389 -8980
rect 7677 -9015 7703 -8980
rect 8321 -9015 8337 -8980
rect 8625 -9015 8651 -8980
rect 9257 -9015 9273 -8980
rect 9561 -9015 9587 -8980
rect 10188 -9014 10204 -8979
rect 10492 -9014 10518 -8979
rect 11115 -9015 11131 -8980
rect 11419 -9015 11445 -8980
rect -8078 -9168 -8044 -9152
rect -21943 -9216 -21927 -9182
rect -21943 -9232 -21893 -9216
rect -21850 -9260 -21834 -9226
rect -21658 -9260 -21642 -9226
rect -20469 -9246 -20452 -9211
rect -20418 -9246 -20402 -9211
rect -20180 -9217 -20163 -9211
rect -20368 -9246 -20163 -9217
rect -20129 -9246 -20113 -9211
rect -24335 -9300 -24200 -9284
rect -24335 -9335 -24234 -9300
rect -22599 -9300 -22464 -9284
rect -24335 -9351 -24200 -9335
rect -24166 -9364 -24150 -9330
rect -23774 -9364 -23758 -9330
rect -23568 -9362 -23552 -9328
rect -23420 -9362 -23404 -9328
rect -22599 -9335 -22498 -9300
rect -22599 -9351 -22464 -9335
rect -22430 -9364 -22414 -9330
rect -22038 -9364 -22022 -9330
rect -21831 -9362 -21815 -9328
rect -21683 -9362 -21667 -9328
rect -24162 -9436 -24135 -9402
rect -23800 -9436 -23762 -9402
rect -22426 -9436 -22399 -9402
rect -22064 -9436 -22026 -9402
rect -20469 -9452 -20426 -9246
rect -20368 -9251 -20113 -9246
rect -19360 -9246 -19343 -9211
rect -19309 -9246 -19293 -9211
rect -19071 -9217 -19054 -9211
rect -19259 -9246 -19054 -9217
rect -19020 -9246 -19004 -9211
rect -20368 -9335 -20334 -9251
rect -20300 -9340 -20284 -9306
rect -19908 -9340 -19892 -9306
rect -20368 -9386 -20334 -9370
rect -19360 -9452 -19317 -9246
rect -19259 -9251 -19004 -9246
rect -18478 -9246 -18461 -9211
rect -18427 -9246 -18411 -9211
rect -18189 -9217 -18172 -9211
rect -18377 -9246 -18172 -9217
rect -18138 -9246 -18122 -9211
rect -19259 -9335 -19225 -9251
rect -19191 -9340 -19175 -9306
rect -18799 -9340 -18783 -9306
rect -19259 -9386 -19225 -9370
rect -18478 -9452 -18435 -9246
rect -18377 -9251 -18122 -9246
rect -17178 -9246 -17161 -9211
rect -17127 -9246 -17111 -9211
rect -16889 -9217 -16872 -9211
rect -17077 -9246 -16872 -9217
rect -16838 -9246 -16822 -9211
rect -18377 -9335 -18343 -9251
rect -18309 -9340 -18293 -9306
rect -17917 -9340 -17901 -9306
rect -18377 -9386 -18343 -9370
rect -17178 -9452 -17135 -9246
rect -17077 -9251 -16822 -9246
rect -16069 -9246 -16052 -9211
rect -16018 -9246 -16002 -9211
rect -15780 -9217 -15763 -9211
rect -15968 -9246 -15763 -9217
rect -15729 -9246 -15713 -9211
rect -17077 -9335 -17043 -9251
rect -17009 -9340 -16993 -9306
rect -16617 -9340 -16601 -9306
rect -17077 -9386 -17043 -9370
rect -16069 -9452 -16026 -9246
rect -15968 -9251 -15713 -9246
rect -15187 -9246 -15170 -9211
rect -15136 -9246 -15120 -9211
rect -14898 -9217 -14881 -9211
rect -15086 -9246 -14881 -9217
rect -14847 -9246 -14831 -9211
rect -15968 -9335 -15934 -9251
rect -15900 -9340 -15884 -9306
rect -15508 -9340 -15492 -9306
rect -15968 -9386 -15934 -9370
rect -15187 -9452 -15144 -9246
rect -15086 -9251 -14831 -9246
rect -13887 -9246 -13870 -9211
rect -13836 -9246 -13820 -9211
rect -13598 -9217 -13581 -9211
rect -13786 -9246 -13581 -9217
rect -13547 -9246 -13531 -9211
rect -15086 -9335 -15052 -9251
rect -15018 -9340 -15002 -9306
rect -14626 -9340 -14610 -9306
rect -15086 -9386 -15052 -9370
rect -13887 -9452 -13844 -9246
rect -13786 -9251 -13531 -9246
rect -12778 -9246 -12761 -9211
rect -12727 -9246 -12711 -9211
rect -12489 -9217 -12472 -9211
rect -12677 -9246 -12472 -9217
rect -12438 -9246 -12422 -9211
rect -13786 -9335 -13752 -9251
rect -13718 -9340 -13702 -9306
rect -13326 -9340 -13310 -9306
rect -13786 -9386 -13752 -9370
rect -12778 -9452 -12735 -9246
rect -12677 -9251 -12422 -9246
rect -11896 -9246 -11879 -9211
rect -11845 -9246 -11829 -9211
rect -11607 -9217 -11590 -9211
rect -11795 -9246 -11590 -9217
rect -11556 -9246 -11540 -9211
rect -12677 -9335 -12643 -9251
rect -12609 -9340 -12593 -9306
rect -12217 -9340 -12201 -9306
rect -12677 -9386 -12643 -9370
rect -11896 -9452 -11853 -9246
rect -11795 -9251 -11540 -9246
rect -10596 -9246 -10579 -9211
rect -10545 -9246 -10529 -9211
rect -10307 -9217 -10290 -9211
rect -10495 -9246 -10290 -9217
rect -10256 -9246 -10240 -9211
rect -11795 -9335 -11761 -9251
rect -11727 -9340 -11711 -9306
rect -11335 -9340 -11319 -9306
rect -11795 -9386 -11761 -9370
rect -10596 -9452 -10553 -9246
rect -10495 -9251 -10240 -9246
rect -9487 -9246 -9470 -9211
rect -9436 -9246 -9420 -9211
rect -9198 -9217 -9181 -9211
rect -9386 -9246 -9181 -9217
rect -9147 -9246 -9131 -9211
rect -10495 -9335 -10461 -9251
rect -10427 -9340 -10411 -9306
rect -10035 -9340 -10019 -9306
rect -10495 -9386 -10461 -9370
rect -9487 -9452 -9444 -9246
rect -9386 -9251 -9131 -9246
rect -8605 -9246 -8588 -9211
rect -8554 -9246 -8538 -9211
rect -8316 -9217 -8299 -9211
rect -8504 -9246 -8299 -9217
rect -8265 -9246 -8249 -9211
rect -9386 -9335 -9352 -9251
rect -9318 -9340 -9302 -9306
rect -8926 -9340 -8910 -9306
rect -9386 -9386 -9352 -9370
rect -8605 -9452 -8562 -9246
rect -8504 -9251 -8249 -9246
rect -8504 -9335 -8470 -9251
rect -8436 -9340 -8420 -9306
rect -8044 -9340 -8028 -9306
rect -8504 -9386 -8470 -9370
rect -20469 -9468 -20334 -9452
rect -20469 -9503 -20368 -9468
rect -19360 -9468 -19225 -9452
rect -20469 -9519 -20334 -9503
rect -20300 -9532 -20284 -9498
rect -19908 -9532 -19892 -9498
rect -19360 -9503 -19259 -9468
rect -18478 -9468 -18343 -9452
rect -19360 -9519 -19225 -9503
rect -19191 -9532 -19175 -9498
rect -18799 -9532 -18783 -9498
rect -18478 -9503 -18377 -9468
rect -17178 -9468 -17043 -9452
rect -18478 -9519 -18343 -9503
rect -18309 -9532 -18293 -9498
rect -17917 -9532 -17901 -9498
rect -17178 -9503 -17077 -9468
rect -16069 -9468 -15934 -9452
rect -17178 -9519 -17043 -9503
rect -17009 -9532 -16993 -9498
rect -16617 -9532 -16601 -9498
rect -16069 -9503 -15968 -9468
rect -15187 -9468 -15052 -9452
rect -16069 -9519 -15934 -9503
rect -15900 -9532 -15884 -9498
rect -15508 -9532 -15492 -9498
rect -15187 -9503 -15086 -9468
rect -13887 -9468 -13752 -9452
rect -15187 -9519 -15052 -9503
rect -15018 -9532 -15002 -9498
rect -14626 -9532 -14610 -9498
rect -13887 -9503 -13786 -9468
rect -12778 -9468 -12643 -9452
rect -13887 -9519 -13752 -9503
rect -13718 -9532 -13702 -9498
rect -13326 -9532 -13310 -9498
rect -12778 -9503 -12677 -9468
rect -11896 -9468 -11761 -9452
rect -12778 -9519 -12643 -9503
rect -12609 -9532 -12593 -9498
rect -12217 -9532 -12201 -9498
rect -11896 -9503 -11795 -9468
rect -10596 -9468 -10461 -9452
rect -11896 -9519 -11761 -9503
rect -11727 -9532 -11711 -9498
rect -11335 -9532 -11319 -9498
rect -10596 -9503 -10495 -9468
rect -9487 -9468 -9352 -9452
rect -10596 -9519 -10461 -9503
rect -10427 -9532 -10411 -9498
rect -10035 -9532 -10019 -9498
rect -9487 -9503 -9386 -9468
rect -8605 -9468 -8470 -9452
rect -9487 -9519 -9352 -9503
rect -9318 -9532 -9302 -9498
rect -8926 -9532 -8910 -9498
rect -8605 -9503 -8504 -9468
rect -8605 -9519 -8470 -9503
rect -8436 -9532 -8420 -9498
rect -8044 -9532 -8028 -9498
rect -20296 -9604 -20269 -9570
rect -19934 -9604 -19896 -9570
rect -19187 -9604 -19160 -9570
rect -18825 -9604 -18787 -9570
rect -18305 -9604 -18278 -9570
rect -17943 -9604 -17905 -9570
rect -17005 -9604 -16978 -9570
rect -16643 -9604 -16605 -9570
rect -15896 -9604 -15869 -9570
rect -15534 -9604 -15496 -9570
rect -15014 -9604 -14987 -9570
rect -14652 -9604 -14614 -9570
rect -13714 -9604 -13687 -9570
rect -13352 -9604 -13314 -9570
rect -12605 -9604 -12578 -9570
rect -12243 -9604 -12205 -9570
rect -11723 -9604 -11696 -9570
rect -11361 -9604 -11323 -9570
rect -10423 -9604 -10396 -9570
rect -10061 -9604 -10023 -9570
rect -9314 -9604 -9287 -9570
rect -8952 -9604 -8914 -9570
rect -8432 -9604 -8405 -9570
rect -8070 -9604 -8032 -9570
rect 5705 -9635 5721 -9601
rect 5812 -9635 5828 -9601
rect 6145 -9635 6161 -9601
rect 6252 -9635 6268 -9601
rect 6585 -9635 6601 -9601
rect 6692 -9635 6708 -9601
rect 5561 -9721 5611 -9704
rect 5654 -9707 5664 -9673
rect 5860 -9707 5876 -9673
rect 5561 -9947 5577 -9721
rect 6001 -9721 6051 -9704
rect 6094 -9707 6104 -9673
rect 6300 -9707 6316 -9673
rect 5654 -9803 5670 -9769
rect 5864 -9803 5882 -9769
rect 5654 -9899 5664 -9865
rect 5860 -9899 5876 -9865
rect 5561 -10167 5611 -9947
rect 6001 -9947 6017 -9721
rect 6441 -9721 6491 -9704
rect 6534 -9707 6544 -9673
rect 6740 -9707 6756 -9673
rect 6094 -9803 6110 -9769
rect 6304 -9803 6322 -9769
rect 6094 -9899 6104 -9865
rect 6300 -9899 6316 -9865
rect 5654 -9995 5670 -9961
rect 5864 -9995 5882 -9961
rect 5654 -10157 5670 -10123
rect 5846 -10157 5862 -10123
rect 5561 -10201 5577 -10167
rect 5561 -10217 5611 -10201
rect 6001 -10167 6051 -9947
rect 6441 -9947 6457 -9721
rect 6534 -9803 6550 -9769
rect 6744 -9803 6762 -9769
rect 6534 -9899 6544 -9865
rect 6740 -9899 6756 -9865
rect 6094 -9995 6110 -9961
rect 6304 -9995 6322 -9961
rect 6094 -10157 6110 -10123
rect 6286 -10157 6302 -10123
rect 6001 -10201 6017 -10167
rect 5654 -10245 5670 -10211
rect 5846 -10245 5862 -10211
rect 6001 -10217 6051 -10201
rect 6441 -10167 6491 -9947
rect 6534 -9995 6550 -9961
rect 6744 -9995 6762 -9961
rect 6534 -10157 6550 -10123
rect 6726 -10157 6742 -10123
rect 6441 -10201 6457 -10167
rect 6094 -10245 6110 -10211
rect 6286 -10245 6302 -10211
rect 6441 -10217 6491 -10201
rect 6534 -10245 6550 -10211
rect 6726 -10245 6742 -10211
rect 7373 -10308 7389 -10273
rect 7677 -10308 7703 -10273
rect 8321 -10308 8337 -10273
rect 8625 -10308 8651 -10273
rect 9257 -10308 9273 -10273
rect 9561 -10308 9587 -10273
rect 10188 -10308 10204 -10273
rect 10492 -10308 10518 -10273
rect 11115 -10308 11131 -10273
rect 11419 -10308 11445 -10273
rect -20649 -10356 -19439 -10328
rect -20649 -10428 -20603 -10356
rect -19481 -10428 -19439 -10356
rect -20649 -10454 -19439 -10428
rect -19090 -10356 -17880 -10328
rect -19090 -10428 -19044 -10356
rect -17922 -10428 -17880 -10356
rect -19090 -10454 -17880 -10428
rect -17358 -10356 -16148 -10328
rect -17358 -10428 -17312 -10356
rect -16190 -10428 -16148 -10356
rect -17358 -10454 -16148 -10428
rect -15799 -10356 -14589 -10328
rect -15799 -10428 -15753 -10356
rect -14631 -10428 -14589 -10356
rect -15799 -10454 -14589 -10428
rect -14067 -10356 -12857 -10328
rect -14067 -10428 -14021 -10356
rect -12899 -10428 -12857 -10356
rect -14067 -10454 -12857 -10428
rect -12508 -10356 -11298 -10328
rect -12508 -10428 -12462 -10356
rect -11340 -10428 -11298 -10356
rect -12508 -10454 -11298 -10428
rect -10776 -10356 -9566 -10328
rect -10776 -10428 -10730 -10356
rect -9608 -10428 -9566 -10356
rect -10776 -10454 -9566 -10428
rect -9217 -10356 -8007 -10328
rect 5673 -10347 5689 -10313
rect 5821 -10347 5837 -10313
rect 6113 -10347 6129 -10313
rect 6261 -10347 6277 -10313
rect 6553 -10347 6569 -10313
rect 6701 -10347 6717 -10313
rect -9217 -10428 -9171 -10356
rect -8049 -10428 -8007 -10356
rect -9217 -10454 -8007 -10428
rect 7150 -10377 7184 -10361
rect -20725 -10525 -20691 -10509
rect -23536 -10622 -23520 -10588
rect -23429 -10622 -23413 -10588
rect -21803 -10622 -21787 -10588
rect -21696 -10622 -21680 -10588
rect -24384 -10688 -24368 -10641
rect -23799 -10688 -23775 -10641
rect -23680 -10708 -23630 -10691
rect -23587 -10694 -23577 -10660
rect -23381 -10694 -23365 -10660
rect -22647 -10688 -22631 -10641
rect -22062 -10688 -22038 -10641
rect -24384 -10760 -24350 -10750
rect -24384 -10972 -24350 -10956
rect -24288 -10766 -24254 -10750
rect -24288 -10972 -24254 -10962
rect -24192 -10760 -24158 -10750
rect -24192 -10972 -24158 -10956
rect -24096 -10766 -24062 -10750
rect -24096 -10972 -24062 -10962
rect -24000 -10760 -23966 -10750
rect -24000 -10972 -23966 -10956
rect -23904 -10766 -23870 -10750
rect -23904 -10972 -23870 -10962
rect -23808 -10760 -23774 -10750
rect -23808 -10972 -23774 -10956
rect -23680 -10934 -23664 -10708
rect -21947 -10708 -21897 -10691
rect -21854 -10694 -21844 -10660
rect -21648 -10694 -21632 -10660
rect -23587 -10790 -23571 -10756
rect -23377 -10790 -23359 -10756
rect -22647 -10760 -22613 -10750
rect -23587 -10886 -23577 -10852
rect -23381 -10886 -23365 -10852
rect -24335 -11050 -24318 -11015
rect -24284 -11050 -24268 -11015
rect -24046 -11021 -24029 -11015
rect -24234 -11050 -24029 -11021
rect -23995 -11050 -23979 -11015
rect -24335 -11256 -24292 -11050
rect -24234 -11055 -23979 -11050
rect -24234 -11139 -24200 -11055
rect -24166 -11144 -24150 -11110
rect -23774 -11144 -23758 -11110
rect -24234 -11190 -24200 -11174
rect -23680 -11154 -23630 -10934
rect -23587 -10982 -23571 -10948
rect -23377 -10982 -23359 -10948
rect -22647 -10972 -22613 -10956
rect -22551 -10766 -22517 -10750
rect -22551 -10972 -22517 -10962
rect -22455 -10760 -22421 -10750
rect -22455 -10972 -22421 -10956
rect -22359 -10766 -22325 -10750
rect -22359 -10972 -22325 -10962
rect -22263 -10760 -22229 -10750
rect -22263 -10972 -22229 -10956
rect -22167 -10766 -22133 -10750
rect -22167 -10972 -22133 -10962
rect -22071 -10760 -22037 -10750
rect -22071 -10972 -22037 -10956
rect -21947 -10934 -21931 -10708
rect -21854 -10790 -21838 -10756
rect -21644 -10790 -21626 -10756
rect -21854 -10886 -21844 -10852
rect -21648 -10886 -21632 -10852
rect -22598 -11050 -22581 -11015
rect -22547 -11050 -22531 -11015
rect -22309 -11021 -22292 -11015
rect -22497 -11050 -22292 -11021
rect -22258 -11050 -22242 -11015
rect -23587 -11144 -23571 -11110
rect -23395 -11144 -23379 -11110
rect -23680 -11188 -23664 -11154
rect -23680 -11204 -23630 -11188
rect -23587 -11232 -23571 -11198
rect -23395 -11232 -23379 -11198
rect -22598 -11256 -22555 -11050
rect -22497 -11055 -22242 -11050
rect -22497 -11139 -22463 -11055
rect -22429 -11144 -22413 -11110
rect -22037 -11144 -22021 -11110
rect -22497 -11190 -22463 -11174
rect -21947 -11154 -21897 -10934
rect -21854 -10982 -21838 -10948
rect -21644 -10982 -21626 -10948
rect -21854 -11144 -21838 -11110
rect -21662 -11144 -21646 -11110
rect -20725 -11112 -20691 -11051
rect -20637 -10525 -20603 -10509
rect -20637 -11067 -20603 -11051
rect -20541 -10525 -20507 -10509
rect -20541 -11067 -20507 -11051
rect -20445 -10525 -20411 -10509
rect -20445 -11067 -20411 -11051
rect -20349 -10525 -20315 -10509
rect -20349 -11067 -20315 -11051
rect -20253 -10525 -20219 -10509
rect -20253 -11067 -20219 -11051
rect -20157 -10525 -20123 -10509
rect -20157 -11067 -20123 -11051
rect -20061 -10525 -20027 -10509
rect -20061 -11094 -20027 -11051
rect -19965 -10525 -19931 -10509
rect -19965 -11067 -19931 -11051
rect -19869 -10525 -19835 -10509
rect -19869 -11067 -19835 -11051
rect -19773 -10525 -19739 -10509
rect -19773 -11067 -19739 -11051
rect -19677 -10525 -19643 -10509
rect -19677 -11067 -19643 -11051
rect -19581 -10525 -19547 -10509
rect -19581 -11067 -19547 -11051
rect -19485 -10525 -19451 -10509
rect -19485 -11067 -19451 -11051
rect -19397 -10525 -19363 -10509
rect -20725 -11122 -20123 -11112
rect -21947 -11188 -21931 -11154
rect -21947 -11204 -21897 -11188
rect -20872 -11151 -20787 -11128
rect -21854 -11232 -21838 -11198
rect -21662 -11232 -21646 -11198
rect -24335 -11272 -24200 -11256
rect -24335 -11307 -24234 -11272
rect -22598 -11272 -22463 -11256
rect -24335 -11323 -24200 -11307
rect -24166 -11336 -24150 -11302
rect -23774 -11336 -23758 -11302
rect -23568 -11334 -23552 -11300
rect -23420 -11334 -23404 -11300
rect -22598 -11307 -22497 -11272
rect -20872 -11261 -20854 -11151
rect -20807 -11261 -20787 -11151
rect -20872 -11281 -20787 -11261
rect -20725 -11167 -20269 -11122
rect -20139 -11167 -20123 -11122
rect -20725 -11181 -20123 -11167
rect -22598 -11323 -22463 -11307
rect -22429 -11336 -22413 -11302
rect -22037 -11336 -22021 -11302
rect -21835 -11334 -21819 -11300
rect -21687 -11334 -21671 -11300
rect -24162 -11408 -24135 -11374
rect -23800 -11408 -23762 -11374
rect -22425 -11408 -22398 -11374
rect -22063 -11408 -22025 -11374
rect -20725 -11565 -20691 -11181
rect -20589 -11252 -20368 -11225
rect -20589 -11305 -20539 -11252
rect -20406 -11305 -20368 -11252
rect -20589 -11443 -20368 -11305
rect -20589 -11488 -20544 -11443
rect -20414 -11488 -20368 -11443
rect -20589 -11515 -20368 -11488
rect -20288 -11451 -20123 -11181
rect -20288 -11496 -20261 -11451
rect -20131 -11496 -20123 -11451
rect -20288 -11513 -20123 -11496
rect -20077 -11394 -20011 -11094
rect -19397 -11109 -19363 -11051
rect -19965 -11127 -19363 -11109
rect -19965 -11172 -19938 -11127
rect -19808 -11172 -19363 -11127
rect -19965 -11186 -19363 -11172
rect -19166 -10525 -19132 -10509
rect -19166 -11112 -19132 -11051
rect -19078 -10525 -19044 -10509
rect -19078 -11067 -19044 -11051
rect -18982 -10525 -18948 -10509
rect -18982 -11067 -18948 -11051
rect -18886 -10525 -18852 -10509
rect -18886 -11067 -18852 -11051
rect -18790 -10525 -18756 -10509
rect -18790 -11067 -18756 -11051
rect -18694 -10525 -18660 -10509
rect -18694 -11067 -18660 -11051
rect -18598 -10525 -18564 -10509
rect -18598 -11067 -18564 -11051
rect -18502 -10525 -18468 -10509
rect -18502 -11094 -18468 -11051
rect -18406 -10525 -18372 -10509
rect -18406 -11067 -18372 -11051
rect -18310 -10525 -18276 -10509
rect -18310 -11067 -18276 -11051
rect -18214 -10525 -18180 -10509
rect -18214 -11067 -18180 -11051
rect -18118 -10525 -18084 -10509
rect -18118 -11067 -18084 -11051
rect -18022 -10525 -17988 -10509
rect -18022 -11067 -17988 -11051
rect -17926 -10525 -17892 -10509
rect -17926 -11067 -17892 -11051
rect -17838 -10525 -17804 -10509
rect -19166 -11122 -18564 -11112
rect -19166 -11167 -18710 -11122
rect -18580 -11167 -18564 -11122
rect -19166 -11181 -18564 -11167
rect -19965 -11244 -19788 -11186
rect -19965 -11297 -19933 -11244
rect -19819 -11297 -19788 -11244
rect -19965 -11326 -19788 -11297
rect -19716 -11245 -19601 -11227
rect -19716 -11313 -19699 -11245
rect -19619 -11313 -19601 -11245
rect -19716 -11333 -19601 -11313
rect -20077 -11416 -19437 -11394
rect -20077 -11471 -19517 -11416
rect -19452 -11471 -19437 -11416
rect -20077 -11490 -19437 -11471
rect -20077 -11524 -20011 -11490
rect -20725 -11687 -20691 -11671
rect -20637 -11565 -20603 -11549
rect -20637 -11687 -20603 -11671
rect -20541 -11550 -20507 -11549
rect -20541 -11687 -20507 -11671
rect -20445 -11565 -20411 -11549
rect -20445 -11687 -20411 -11685
rect -20349 -11550 -20315 -11549
rect -20349 -11687 -20315 -11671
rect -20253 -11565 -20219 -11549
rect -20253 -11687 -20219 -11685
rect -20157 -11551 -20123 -11549
rect -20157 -11687 -20123 -11671
rect -20061 -11565 -20027 -11524
rect -20061 -11687 -20027 -11685
rect -19965 -11550 -19931 -11549
rect -19965 -11687 -19931 -11671
rect -19869 -11565 -19835 -11549
rect -19869 -11687 -19835 -11685
rect -19773 -11550 -19739 -11549
rect -19773 -11687 -19739 -11671
rect -19677 -11565 -19643 -11549
rect -19677 -11687 -19643 -11685
rect -19581 -11550 -19547 -11549
rect -19581 -11687 -19547 -11671
rect -19485 -11565 -19451 -11549
rect -19485 -11687 -19451 -11671
rect -19397 -11565 -19363 -11186
rect -19316 -11196 -19207 -11181
rect -19316 -11336 -19297 -11196
rect -19224 -11336 -19207 -11196
rect -19316 -11353 -19207 -11336
rect -19397 -11687 -19363 -11671
rect -19166 -11565 -19132 -11181
rect -19030 -11252 -18809 -11225
rect -19030 -11305 -18980 -11252
rect -18847 -11305 -18809 -11252
rect -19030 -11443 -18809 -11305
rect -19030 -11488 -18985 -11443
rect -18855 -11488 -18809 -11443
rect -19030 -11515 -18809 -11488
rect -18729 -11451 -18564 -11181
rect -18729 -11496 -18702 -11451
rect -18572 -11496 -18564 -11451
rect -18729 -11513 -18564 -11496
rect -18518 -11394 -18452 -11094
rect -17838 -11109 -17804 -11051
rect -18406 -11127 -17804 -11109
rect -18406 -11172 -18379 -11127
rect -18249 -11172 -17804 -11127
rect -17434 -10525 -17400 -10509
rect -17434 -11112 -17400 -11051
rect -17346 -10525 -17312 -10509
rect -17346 -11067 -17312 -11051
rect -17250 -10525 -17216 -10509
rect -17250 -11067 -17216 -11051
rect -17154 -10525 -17120 -10509
rect -17154 -11067 -17120 -11051
rect -17058 -10525 -17024 -10509
rect -17058 -11067 -17024 -11051
rect -16962 -10525 -16928 -10509
rect -16962 -11067 -16928 -11051
rect -16866 -10525 -16832 -10509
rect -16866 -11067 -16832 -11051
rect -16770 -10525 -16736 -10509
rect -16770 -11094 -16736 -11051
rect -16674 -10525 -16640 -10509
rect -16674 -11067 -16640 -11051
rect -16578 -10525 -16544 -10509
rect -16578 -11067 -16544 -11051
rect -16482 -10525 -16448 -10509
rect -16482 -11067 -16448 -11051
rect -16386 -10525 -16352 -10509
rect -16386 -11067 -16352 -11051
rect -16290 -10525 -16256 -10509
rect -16290 -11067 -16256 -11051
rect -16194 -10525 -16160 -10509
rect -16194 -11067 -16160 -11051
rect -16106 -10525 -16072 -10509
rect -17434 -11122 -16832 -11112
rect -18406 -11186 -17804 -11172
rect -18406 -11244 -18229 -11186
rect -18406 -11297 -18374 -11244
rect -18260 -11297 -18229 -11244
rect -18406 -11326 -18229 -11297
rect -18157 -11245 -18042 -11227
rect -18157 -11313 -18140 -11245
rect -18060 -11313 -18042 -11245
rect -18157 -11333 -18042 -11313
rect -18518 -11416 -17878 -11394
rect -18518 -11471 -17958 -11416
rect -17893 -11471 -17878 -11416
rect -18518 -11490 -17878 -11471
rect -18518 -11524 -18452 -11490
rect -19166 -11687 -19132 -11671
rect -19078 -11565 -19044 -11549
rect -19078 -11687 -19044 -11671
rect -18982 -11550 -18948 -11549
rect -18982 -11687 -18948 -11671
rect -18886 -11565 -18852 -11549
rect -18886 -11687 -18852 -11685
rect -18790 -11550 -18756 -11549
rect -18790 -11687 -18756 -11671
rect -18694 -11565 -18660 -11549
rect -18694 -11687 -18660 -11685
rect -18598 -11551 -18564 -11549
rect -18598 -11687 -18564 -11671
rect -18502 -11565 -18468 -11524
rect -18502 -11687 -18468 -11685
rect -18406 -11550 -18372 -11549
rect -18406 -11687 -18372 -11671
rect -18310 -11565 -18276 -11549
rect -18310 -11687 -18276 -11685
rect -18214 -11550 -18180 -11549
rect -18214 -11687 -18180 -11671
rect -18118 -11565 -18084 -11549
rect -18118 -11687 -18084 -11685
rect -18022 -11550 -17988 -11549
rect -18022 -11687 -17988 -11671
rect -17926 -11565 -17892 -11549
rect -17926 -11687 -17892 -11671
rect -17838 -11565 -17804 -11186
rect -17581 -11151 -17496 -11128
rect -17581 -11261 -17563 -11151
rect -17516 -11261 -17496 -11151
rect -17581 -11281 -17496 -11261
rect -17434 -11167 -16978 -11122
rect -16848 -11167 -16832 -11122
rect -17434 -11181 -16832 -11167
rect -17838 -11687 -17804 -11671
rect -17434 -11565 -17400 -11181
rect -17298 -11252 -17077 -11225
rect -17298 -11305 -17248 -11252
rect -17115 -11305 -17077 -11252
rect -17298 -11443 -17077 -11305
rect -17298 -11488 -17253 -11443
rect -17123 -11488 -17077 -11443
rect -17298 -11515 -17077 -11488
rect -16997 -11451 -16832 -11181
rect -16997 -11496 -16970 -11451
rect -16840 -11496 -16832 -11451
rect -16997 -11513 -16832 -11496
rect -16786 -11394 -16720 -11094
rect -16106 -11109 -16072 -11051
rect -16674 -11127 -16072 -11109
rect -16674 -11172 -16647 -11127
rect -16517 -11172 -16072 -11127
rect -16674 -11186 -16072 -11172
rect -15875 -10525 -15841 -10509
rect -15875 -11112 -15841 -11051
rect -15787 -10525 -15753 -10509
rect -15787 -11067 -15753 -11051
rect -15691 -10525 -15657 -10509
rect -15691 -11067 -15657 -11051
rect -15595 -10525 -15561 -10509
rect -15595 -11067 -15561 -11051
rect -15499 -10525 -15465 -10509
rect -15499 -11067 -15465 -11051
rect -15403 -10525 -15369 -10509
rect -15403 -11067 -15369 -11051
rect -15307 -10525 -15273 -10509
rect -15307 -11067 -15273 -11051
rect -15211 -10525 -15177 -10509
rect -15211 -11094 -15177 -11051
rect -15115 -10525 -15081 -10509
rect -15115 -11067 -15081 -11051
rect -15019 -10525 -14985 -10509
rect -15019 -11067 -14985 -11051
rect -14923 -10525 -14889 -10509
rect -14923 -11067 -14889 -11051
rect -14827 -10525 -14793 -10509
rect -14827 -11067 -14793 -11051
rect -14731 -10525 -14697 -10509
rect -14731 -11067 -14697 -11051
rect -14635 -10525 -14601 -10509
rect -14635 -11067 -14601 -11051
rect -14547 -10525 -14513 -10509
rect -15875 -11122 -15273 -11112
rect -15875 -11167 -15419 -11122
rect -15289 -11167 -15273 -11122
rect -15875 -11181 -15273 -11167
rect -16674 -11244 -16497 -11186
rect -16674 -11297 -16642 -11244
rect -16528 -11297 -16497 -11244
rect -16674 -11326 -16497 -11297
rect -16425 -11245 -16310 -11227
rect -16425 -11313 -16408 -11245
rect -16328 -11313 -16310 -11245
rect -16425 -11333 -16310 -11313
rect -16786 -11416 -16146 -11394
rect -16786 -11471 -16226 -11416
rect -16161 -11471 -16146 -11416
rect -16786 -11490 -16146 -11471
rect -16786 -11524 -16720 -11490
rect -17434 -11687 -17400 -11671
rect -17346 -11565 -17312 -11549
rect -17346 -11687 -17312 -11671
rect -17250 -11550 -17216 -11549
rect -17250 -11687 -17216 -11671
rect -17154 -11565 -17120 -11549
rect -17154 -11687 -17120 -11685
rect -17058 -11550 -17024 -11549
rect -17058 -11687 -17024 -11671
rect -16962 -11565 -16928 -11549
rect -16962 -11687 -16928 -11685
rect -16866 -11551 -16832 -11549
rect -16866 -11687 -16832 -11671
rect -16770 -11565 -16736 -11524
rect -16770 -11687 -16736 -11685
rect -16674 -11550 -16640 -11549
rect -16674 -11687 -16640 -11671
rect -16578 -11565 -16544 -11549
rect -16578 -11687 -16544 -11685
rect -16482 -11550 -16448 -11549
rect -16482 -11687 -16448 -11671
rect -16386 -11565 -16352 -11549
rect -16386 -11687 -16352 -11685
rect -16290 -11550 -16256 -11549
rect -16290 -11687 -16256 -11671
rect -16194 -11565 -16160 -11549
rect -16194 -11687 -16160 -11671
rect -16106 -11565 -16072 -11186
rect -16025 -11196 -15916 -11181
rect -16025 -11336 -16006 -11196
rect -15933 -11336 -15916 -11196
rect -16025 -11353 -15916 -11336
rect -16106 -11687 -16072 -11671
rect -15875 -11565 -15841 -11181
rect -15739 -11252 -15518 -11225
rect -15739 -11305 -15689 -11252
rect -15556 -11305 -15518 -11252
rect -15739 -11443 -15518 -11305
rect -15739 -11488 -15694 -11443
rect -15564 -11488 -15518 -11443
rect -15739 -11515 -15518 -11488
rect -15438 -11451 -15273 -11181
rect -15438 -11496 -15411 -11451
rect -15281 -11496 -15273 -11451
rect -15438 -11513 -15273 -11496
rect -15227 -11394 -15161 -11094
rect -14547 -11109 -14513 -11051
rect -15115 -11127 -14513 -11109
rect -15115 -11172 -15088 -11127
rect -14958 -11172 -14513 -11127
rect -14143 -10525 -14109 -10509
rect -14143 -11112 -14109 -11051
rect -14055 -10525 -14021 -10509
rect -14055 -11067 -14021 -11051
rect -13959 -10525 -13925 -10509
rect -13959 -11067 -13925 -11051
rect -13863 -10525 -13829 -10509
rect -13863 -11067 -13829 -11051
rect -13767 -10525 -13733 -10509
rect -13767 -11067 -13733 -11051
rect -13671 -10525 -13637 -10509
rect -13671 -11067 -13637 -11051
rect -13575 -10525 -13541 -10509
rect -13575 -11067 -13541 -11051
rect -13479 -10525 -13445 -10509
rect -13479 -11094 -13445 -11051
rect -13383 -10525 -13349 -10509
rect -13383 -11067 -13349 -11051
rect -13287 -10525 -13253 -10509
rect -13287 -11067 -13253 -11051
rect -13191 -10525 -13157 -10509
rect -13191 -11067 -13157 -11051
rect -13095 -10525 -13061 -10509
rect -13095 -11067 -13061 -11051
rect -12999 -10525 -12965 -10509
rect -12999 -11067 -12965 -11051
rect -12903 -10525 -12869 -10509
rect -12903 -11067 -12869 -11051
rect -12815 -10525 -12781 -10509
rect -14143 -11122 -13541 -11112
rect -15115 -11186 -14513 -11172
rect -15115 -11244 -14938 -11186
rect -15115 -11297 -15083 -11244
rect -14969 -11297 -14938 -11244
rect -15115 -11326 -14938 -11297
rect -14866 -11245 -14751 -11227
rect -14866 -11313 -14849 -11245
rect -14769 -11313 -14751 -11245
rect -14866 -11333 -14751 -11313
rect -15227 -11416 -14587 -11394
rect -15227 -11471 -14667 -11416
rect -14602 -11471 -14587 -11416
rect -15227 -11490 -14587 -11471
rect -15227 -11524 -15161 -11490
rect -15875 -11687 -15841 -11671
rect -15787 -11565 -15753 -11549
rect -15787 -11687 -15753 -11671
rect -15691 -11550 -15657 -11549
rect -15691 -11687 -15657 -11671
rect -15595 -11565 -15561 -11549
rect -15595 -11687 -15561 -11685
rect -15499 -11550 -15465 -11549
rect -15499 -11687 -15465 -11671
rect -15403 -11565 -15369 -11549
rect -15403 -11687 -15369 -11685
rect -15307 -11551 -15273 -11549
rect -15307 -11687 -15273 -11671
rect -15211 -11565 -15177 -11524
rect -15211 -11687 -15177 -11685
rect -15115 -11550 -15081 -11549
rect -15115 -11687 -15081 -11671
rect -15019 -11565 -14985 -11549
rect -15019 -11687 -14985 -11685
rect -14923 -11550 -14889 -11549
rect -14923 -11687 -14889 -11671
rect -14827 -11565 -14793 -11549
rect -14827 -11687 -14793 -11685
rect -14731 -11550 -14697 -11549
rect -14731 -11687 -14697 -11671
rect -14635 -11565 -14601 -11549
rect -14635 -11687 -14601 -11671
rect -14547 -11565 -14513 -11186
rect -14290 -11151 -14205 -11128
rect -14290 -11261 -14272 -11151
rect -14225 -11261 -14205 -11151
rect -14290 -11281 -14205 -11261
rect -14143 -11167 -13687 -11122
rect -13557 -11167 -13541 -11122
rect -14143 -11181 -13541 -11167
rect -14547 -11687 -14513 -11671
rect -14143 -11565 -14109 -11181
rect -14007 -11252 -13786 -11225
rect -14007 -11305 -13957 -11252
rect -13824 -11305 -13786 -11252
rect -14007 -11443 -13786 -11305
rect -14007 -11488 -13962 -11443
rect -13832 -11488 -13786 -11443
rect -14007 -11515 -13786 -11488
rect -13706 -11451 -13541 -11181
rect -13706 -11496 -13679 -11451
rect -13549 -11496 -13541 -11451
rect -13706 -11513 -13541 -11496
rect -13495 -11394 -13429 -11094
rect -12815 -11109 -12781 -11051
rect -13383 -11127 -12781 -11109
rect -13383 -11172 -13356 -11127
rect -13226 -11172 -12781 -11127
rect -13383 -11186 -12781 -11172
rect -12584 -10525 -12550 -10509
rect -12584 -11112 -12550 -11051
rect -12496 -10525 -12462 -10509
rect -12496 -11067 -12462 -11051
rect -12400 -10525 -12366 -10509
rect -12400 -11067 -12366 -11051
rect -12304 -10525 -12270 -10509
rect -12304 -11067 -12270 -11051
rect -12208 -10525 -12174 -10509
rect -12208 -11067 -12174 -11051
rect -12112 -10525 -12078 -10509
rect -12112 -11067 -12078 -11051
rect -12016 -10525 -11982 -10509
rect -12016 -11067 -11982 -11051
rect -11920 -10525 -11886 -10509
rect -11920 -11094 -11886 -11051
rect -11824 -10525 -11790 -10509
rect -11824 -11067 -11790 -11051
rect -11728 -10525 -11694 -10509
rect -11728 -11067 -11694 -11051
rect -11632 -10525 -11598 -10509
rect -11632 -11067 -11598 -11051
rect -11536 -10525 -11502 -10509
rect -11536 -11067 -11502 -11051
rect -11440 -10525 -11406 -10509
rect -11440 -11067 -11406 -11051
rect -11344 -10525 -11310 -10509
rect -11344 -11067 -11310 -11051
rect -11256 -10525 -11222 -10509
rect -12584 -11122 -11982 -11112
rect -12584 -11167 -12128 -11122
rect -11998 -11167 -11982 -11122
rect -12584 -11181 -11982 -11167
rect -13383 -11244 -13206 -11186
rect -13383 -11297 -13351 -11244
rect -13237 -11297 -13206 -11244
rect -13383 -11326 -13206 -11297
rect -13134 -11245 -13019 -11227
rect -13134 -11313 -13117 -11245
rect -13037 -11313 -13019 -11245
rect -13134 -11333 -13019 -11313
rect -13495 -11416 -12855 -11394
rect -13495 -11471 -12935 -11416
rect -12870 -11471 -12855 -11416
rect -13495 -11490 -12855 -11471
rect -13495 -11524 -13429 -11490
rect -14143 -11687 -14109 -11671
rect -14055 -11565 -14021 -11549
rect -14055 -11687 -14021 -11671
rect -13959 -11550 -13925 -11549
rect -13959 -11687 -13925 -11671
rect -13863 -11565 -13829 -11549
rect -13863 -11687 -13829 -11685
rect -13767 -11550 -13733 -11549
rect -13767 -11687 -13733 -11671
rect -13671 -11565 -13637 -11549
rect -13671 -11687 -13637 -11685
rect -13575 -11551 -13541 -11549
rect -13575 -11687 -13541 -11671
rect -13479 -11565 -13445 -11524
rect -13479 -11687 -13445 -11685
rect -13383 -11550 -13349 -11549
rect -13383 -11687 -13349 -11671
rect -13287 -11565 -13253 -11549
rect -13287 -11687 -13253 -11685
rect -13191 -11550 -13157 -11549
rect -13191 -11687 -13157 -11671
rect -13095 -11565 -13061 -11549
rect -13095 -11687 -13061 -11685
rect -12999 -11550 -12965 -11549
rect -12999 -11687 -12965 -11671
rect -12903 -11565 -12869 -11549
rect -12903 -11687 -12869 -11671
rect -12815 -11565 -12781 -11186
rect -12734 -11196 -12625 -11181
rect -12734 -11336 -12715 -11196
rect -12642 -11336 -12625 -11196
rect -12734 -11353 -12625 -11336
rect -12815 -11687 -12781 -11671
rect -12584 -11565 -12550 -11181
rect -12448 -11252 -12227 -11225
rect -12448 -11305 -12398 -11252
rect -12265 -11305 -12227 -11252
rect -12448 -11443 -12227 -11305
rect -12448 -11488 -12403 -11443
rect -12273 -11488 -12227 -11443
rect -12448 -11515 -12227 -11488
rect -12147 -11451 -11982 -11181
rect -12147 -11496 -12120 -11451
rect -11990 -11496 -11982 -11451
rect -12147 -11513 -11982 -11496
rect -11936 -11394 -11870 -11094
rect -11256 -11109 -11222 -11051
rect -11824 -11127 -11222 -11109
rect -11824 -11172 -11797 -11127
rect -11667 -11172 -11222 -11127
rect -10852 -10525 -10818 -10509
rect -10852 -11112 -10818 -11051
rect -10764 -10525 -10730 -10509
rect -10764 -11067 -10730 -11051
rect -10668 -10525 -10634 -10509
rect -10668 -11067 -10634 -11051
rect -10572 -10525 -10538 -10509
rect -10572 -11067 -10538 -11051
rect -10476 -10525 -10442 -10509
rect -10476 -11067 -10442 -11051
rect -10380 -10525 -10346 -10509
rect -10380 -11067 -10346 -11051
rect -10284 -10525 -10250 -10509
rect -10284 -11067 -10250 -11051
rect -10188 -10525 -10154 -10509
rect -10188 -11094 -10154 -11051
rect -10092 -10525 -10058 -10509
rect -10092 -11067 -10058 -11051
rect -9996 -10525 -9962 -10509
rect -9996 -11067 -9962 -11051
rect -9900 -10525 -9866 -10509
rect -9900 -11067 -9866 -11051
rect -9804 -10525 -9770 -10509
rect -9804 -11067 -9770 -11051
rect -9708 -10525 -9674 -10509
rect -9708 -11067 -9674 -11051
rect -9612 -10525 -9578 -10509
rect -9612 -11067 -9578 -11051
rect -9524 -10525 -9490 -10509
rect -10852 -11122 -10250 -11112
rect -11824 -11186 -11222 -11172
rect -11824 -11244 -11647 -11186
rect -11824 -11297 -11792 -11244
rect -11678 -11297 -11647 -11244
rect -11824 -11326 -11647 -11297
rect -11575 -11245 -11460 -11227
rect -11575 -11313 -11558 -11245
rect -11478 -11313 -11460 -11245
rect -11575 -11333 -11460 -11313
rect -11936 -11416 -11296 -11394
rect -11936 -11471 -11376 -11416
rect -11311 -11471 -11296 -11416
rect -11936 -11490 -11296 -11471
rect -11936 -11524 -11870 -11490
rect -12584 -11687 -12550 -11671
rect -12496 -11565 -12462 -11549
rect -12496 -11687 -12462 -11671
rect -12400 -11550 -12366 -11549
rect -12400 -11687 -12366 -11671
rect -12304 -11565 -12270 -11549
rect -12304 -11687 -12270 -11685
rect -12208 -11550 -12174 -11549
rect -12208 -11687 -12174 -11671
rect -12112 -11565 -12078 -11549
rect -12112 -11687 -12078 -11685
rect -12016 -11551 -11982 -11549
rect -12016 -11687 -11982 -11671
rect -11920 -11565 -11886 -11524
rect -11920 -11687 -11886 -11685
rect -11824 -11550 -11790 -11549
rect -11824 -11687 -11790 -11671
rect -11728 -11565 -11694 -11549
rect -11728 -11687 -11694 -11685
rect -11632 -11550 -11598 -11549
rect -11632 -11687 -11598 -11671
rect -11536 -11565 -11502 -11549
rect -11536 -11687 -11502 -11685
rect -11440 -11550 -11406 -11549
rect -11440 -11687 -11406 -11671
rect -11344 -11565 -11310 -11549
rect -11344 -11687 -11310 -11671
rect -11256 -11565 -11222 -11186
rect -10999 -11151 -10914 -11128
rect -10999 -11261 -10981 -11151
rect -10934 -11261 -10914 -11151
rect -10999 -11281 -10914 -11261
rect -10852 -11167 -10396 -11122
rect -10266 -11167 -10250 -11122
rect -10852 -11181 -10250 -11167
rect -11256 -11687 -11222 -11671
rect -10852 -11565 -10818 -11181
rect -10716 -11252 -10495 -11225
rect -10716 -11305 -10666 -11252
rect -10533 -11305 -10495 -11252
rect -10716 -11443 -10495 -11305
rect -10716 -11488 -10671 -11443
rect -10541 -11488 -10495 -11443
rect -10716 -11515 -10495 -11488
rect -10415 -11451 -10250 -11181
rect -10415 -11496 -10388 -11451
rect -10258 -11496 -10250 -11451
rect -10415 -11513 -10250 -11496
rect -10204 -11394 -10138 -11094
rect -9524 -11109 -9490 -11051
rect -10092 -11127 -9490 -11109
rect -10092 -11172 -10065 -11127
rect -9935 -11172 -9490 -11127
rect -10092 -11186 -9490 -11172
rect -9293 -10525 -9259 -10509
rect -9293 -11112 -9259 -11051
rect -9205 -10525 -9171 -10509
rect -9205 -11067 -9171 -11051
rect -9109 -10525 -9075 -10509
rect -9109 -11067 -9075 -11051
rect -9013 -10525 -8979 -10509
rect -9013 -11067 -8979 -11051
rect -8917 -10525 -8883 -10509
rect -8917 -11067 -8883 -11051
rect -8821 -10525 -8787 -10509
rect -8821 -11067 -8787 -11051
rect -8725 -10525 -8691 -10509
rect -8725 -11067 -8691 -11051
rect -8629 -10525 -8595 -10509
rect -8629 -11094 -8595 -11051
rect -8533 -10525 -8499 -10509
rect -8533 -11067 -8499 -11051
rect -8437 -10525 -8403 -10509
rect -8437 -11067 -8403 -11051
rect -8341 -10525 -8307 -10509
rect -8341 -11067 -8307 -11051
rect -8245 -10525 -8211 -10509
rect -8245 -11067 -8211 -11051
rect -8149 -10525 -8115 -10509
rect -8149 -11067 -8115 -11051
rect -8053 -10525 -8019 -10509
rect -8053 -11067 -8019 -11051
rect -7965 -10525 -7931 -10509
rect 7246 -10377 7280 -10361
rect 7150 -10691 7184 -10675
rect 7246 -10691 7280 -10680
rect 7342 -10377 7376 -10361
rect 7342 -10691 7376 -10675
rect 7438 -10377 7472 -10361
rect 7534 -10377 7568 -10361
rect 7438 -10691 7472 -10680
rect 7534 -10691 7568 -10675
rect 7630 -10377 7664 -10361
rect 7726 -10377 7760 -10361
rect 7630 -10691 7664 -10680
rect 7726 -10691 7760 -10675
rect 7822 -10377 7856 -10361
rect 7918 -10377 7952 -10361
rect 7822 -10691 7856 -10680
rect 7918 -10691 7952 -10675
rect 8098 -10377 8132 -10361
rect 8194 -10377 8228 -10361
rect 8098 -10691 8132 -10675
rect 8194 -10691 8228 -10680
rect 8290 -10377 8324 -10361
rect 8290 -10691 8324 -10675
rect 8386 -10377 8420 -10361
rect 8482 -10377 8516 -10361
rect 8386 -10691 8420 -10680
rect 8482 -10691 8516 -10675
rect 8578 -10377 8612 -10361
rect 8674 -10377 8708 -10361
rect 8578 -10691 8612 -10680
rect 8674 -10691 8708 -10675
rect 8770 -10377 8804 -10361
rect 8866 -10377 8900 -10361
rect 8770 -10691 8804 -10680
rect 8866 -10691 8900 -10675
rect 9034 -10377 9068 -10361
rect 9130 -10377 9164 -10361
rect 9034 -10691 9068 -10675
rect 9130 -10691 9164 -10680
rect 9226 -10377 9260 -10361
rect 9226 -10691 9260 -10675
rect 9322 -10377 9356 -10361
rect 9418 -10377 9452 -10361
rect 9322 -10691 9356 -10680
rect 9418 -10691 9452 -10675
rect 9514 -10377 9548 -10361
rect 9610 -10377 9644 -10361
rect 9514 -10691 9548 -10680
rect 9610 -10691 9644 -10675
rect 9706 -10377 9740 -10361
rect 9802 -10377 9836 -10361
rect 9706 -10691 9740 -10680
rect 9802 -10691 9836 -10675
rect 9965 -10377 9999 -10361
rect 10061 -10377 10095 -10361
rect 9965 -10691 9999 -10675
rect 10061 -10691 10095 -10680
rect 10157 -10377 10191 -10361
rect 10157 -10691 10191 -10675
rect 10253 -10377 10287 -10361
rect 10349 -10377 10383 -10361
rect 10253 -10691 10287 -10680
rect 10349 -10691 10383 -10675
rect 10445 -10377 10479 -10361
rect 10541 -10377 10575 -10361
rect 10445 -10691 10479 -10680
rect 10541 -10691 10575 -10675
rect 10637 -10377 10671 -10361
rect 10733 -10377 10767 -10361
rect 10637 -10691 10671 -10680
rect 10733 -10691 10767 -10675
rect 10892 -10377 10926 -10361
rect 10988 -10377 11022 -10361
rect 10892 -10691 10926 -10675
rect 10988 -10691 11022 -10680
rect 11084 -10377 11118 -10361
rect 11084 -10691 11118 -10675
rect 11180 -10377 11214 -10361
rect 11276 -10377 11310 -10361
rect 11180 -10691 11214 -10680
rect 11276 -10691 11310 -10675
rect 11372 -10377 11406 -10361
rect 11468 -10377 11502 -10361
rect 11372 -10691 11406 -10680
rect 11468 -10691 11502 -10675
rect 11564 -10377 11598 -10361
rect 11660 -10377 11694 -10361
rect 11564 -10691 11598 -10680
rect 11660 -10691 11694 -10675
rect 7182 -10768 7198 -10734
rect 7232 -10768 7248 -10734
rect 7374 -10768 7390 -10734
rect 7424 -10768 7440 -10734
rect 7566 -10768 7582 -10734
rect 7616 -10768 7632 -10734
rect 7758 -10768 7774 -10734
rect 7808 -10768 7824 -10734
rect 8130 -10768 8146 -10734
rect 8180 -10768 8196 -10734
rect 8322 -10768 8338 -10734
rect 8372 -10768 8388 -10734
rect 8514 -10768 8530 -10734
rect 8564 -10768 8580 -10734
rect 8706 -10768 8722 -10734
rect 8756 -10768 8772 -10734
rect 9066 -10768 9082 -10734
rect 9116 -10768 9132 -10734
rect 9258 -10768 9274 -10734
rect 9308 -10768 9324 -10734
rect 9450 -10768 9466 -10734
rect 9500 -10768 9516 -10734
rect 9642 -10768 9658 -10734
rect 9692 -10768 9708 -10734
rect 9997 -10768 10013 -10734
rect 10047 -10768 10063 -10734
rect 10189 -10768 10205 -10734
rect 10239 -10768 10255 -10734
rect 10381 -10768 10397 -10734
rect 10431 -10768 10447 -10734
rect 10573 -10768 10589 -10734
rect 10623 -10768 10639 -10734
rect 10924 -10768 10940 -10734
rect 10974 -10768 10990 -10734
rect 11116 -10768 11132 -10734
rect 11166 -10768 11182 -10734
rect 11308 -10768 11324 -10734
rect 11358 -10768 11374 -10734
rect 11500 -10768 11516 -10734
rect 11550 -10768 11566 -10734
rect -9293 -11122 -8691 -11112
rect -9293 -11167 -8837 -11122
rect -8707 -11167 -8691 -11122
rect -9293 -11181 -8691 -11167
rect -10092 -11244 -9915 -11186
rect -10092 -11297 -10060 -11244
rect -9946 -11297 -9915 -11244
rect -10092 -11326 -9915 -11297
rect -9843 -11245 -9728 -11227
rect -9843 -11313 -9826 -11245
rect -9746 -11313 -9728 -11245
rect -9843 -11333 -9728 -11313
rect -10204 -11416 -9564 -11394
rect -10204 -11471 -9644 -11416
rect -9579 -11471 -9564 -11416
rect -10204 -11490 -9564 -11471
rect -10204 -11524 -10138 -11490
rect -10852 -11687 -10818 -11671
rect -10764 -11565 -10730 -11549
rect -10764 -11687 -10730 -11671
rect -10668 -11550 -10634 -11549
rect -10668 -11687 -10634 -11671
rect -10572 -11565 -10538 -11549
rect -10572 -11687 -10538 -11685
rect -10476 -11550 -10442 -11549
rect -10476 -11687 -10442 -11671
rect -10380 -11565 -10346 -11549
rect -10380 -11687 -10346 -11685
rect -10284 -11551 -10250 -11549
rect -10284 -11687 -10250 -11671
rect -10188 -11565 -10154 -11524
rect -10188 -11687 -10154 -11685
rect -10092 -11550 -10058 -11549
rect -10092 -11687 -10058 -11671
rect -9996 -11565 -9962 -11549
rect -9996 -11687 -9962 -11685
rect -9900 -11550 -9866 -11549
rect -9900 -11687 -9866 -11671
rect -9804 -11565 -9770 -11549
rect -9804 -11687 -9770 -11685
rect -9708 -11550 -9674 -11549
rect -9708 -11687 -9674 -11671
rect -9612 -11565 -9578 -11549
rect -9612 -11687 -9578 -11671
rect -9524 -11565 -9490 -11186
rect -9443 -11196 -9334 -11181
rect -9443 -11336 -9424 -11196
rect -9351 -11336 -9334 -11196
rect -9443 -11353 -9334 -11336
rect -9524 -11687 -9490 -11671
rect -9293 -11565 -9259 -11181
rect -9157 -11252 -8936 -11225
rect -9157 -11305 -9107 -11252
rect -8974 -11305 -8936 -11252
rect -9157 -11443 -8936 -11305
rect -9157 -11488 -9112 -11443
rect -8982 -11488 -8936 -11443
rect -9157 -11515 -8936 -11488
rect -8856 -11451 -8691 -11181
rect -8856 -11496 -8829 -11451
rect -8699 -11496 -8691 -11451
rect -8856 -11513 -8691 -11496
rect -8645 -11394 -8579 -11094
rect -7965 -11109 -7931 -11051
rect -8533 -11127 -7931 -11109
rect -8533 -11172 -8506 -11127
rect -8376 -11172 -7931 -11127
rect -8533 -11186 -7931 -11172
rect -8533 -11244 -8356 -11186
rect -8533 -11297 -8501 -11244
rect -8387 -11297 -8356 -11244
rect -8533 -11326 -8356 -11297
rect -8284 -11245 -8169 -11227
rect -8284 -11313 -8267 -11245
rect -8187 -11313 -8169 -11245
rect -8284 -11333 -8169 -11313
rect -8645 -11416 -8005 -11394
rect -8645 -11471 -8085 -11416
rect -8020 -11471 -8005 -11416
rect -8645 -11490 -8005 -11471
rect -8645 -11524 -8579 -11490
rect -9293 -11687 -9259 -11671
rect -9205 -11565 -9171 -11549
rect -9205 -11687 -9171 -11671
rect -9109 -11550 -9075 -11549
rect -9109 -11687 -9075 -11671
rect -9013 -11565 -8979 -11549
rect -9013 -11687 -8979 -11685
rect -8917 -11550 -8883 -11549
rect -8917 -11687 -8883 -11671
rect -8821 -11565 -8787 -11549
rect -8821 -11687 -8787 -11685
rect -8725 -11551 -8691 -11549
rect -8725 -11687 -8691 -11671
rect -8629 -11565 -8595 -11524
rect -8629 -11687 -8595 -11685
rect -8533 -11550 -8499 -11549
rect -8533 -11687 -8499 -11671
rect -8437 -11565 -8403 -11549
rect -8437 -11687 -8403 -11685
rect -8341 -11550 -8307 -11549
rect -8341 -11687 -8307 -11671
rect -8245 -11565 -8211 -11549
rect -8245 -11687 -8211 -11685
rect -8149 -11550 -8115 -11549
rect -8149 -11687 -8115 -11671
rect -8053 -11565 -8019 -11549
rect -8053 -11687 -8019 -11671
rect -7965 -11565 -7931 -11186
rect -7965 -11687 -7931 -11671
rect 7298 -11090 7403 -11087
rect 8246 -11090 8351 -11087
rect 9182 -11090 9287 -11087
rect 10113 -11090 10218 -11087
rect 11040 -11090 11145 -11087
rect 7298 -11106 7406 -11090
rect 7298 -11118 7372 -11106
rect -20644 -11759 -19442 -11737
rect -20644 -11805 -20603 -11759
rect -19480 -11805 -19442 -11759
rect -20644 -11828 -19442 -11805
rect -19085 -11759 -17883 -11737
rect -19085 -11805 -19044 -11759
rect -17921 -11805 -17883 -11759
rect -19085 -11828 -17883 -11805
rect -17353 -11759 -16151 -11737
rect -17353 -11805 -17312 -11759
rect -16189 -11805 -16151 -11759
rect -17353 -11828 -16151 -11805
rect -15794 -11759 -14592 -11737
rect -15794 -11805 -15753 -11759
rect -14630 -11805 -14592 -11759
rect -15794 -11828 -14592 -11805
rect -14062 -11759 -12860 -11737
rect -14062 -11805 -14021 -11759
rect -12898 -11805 -12860 -11759
rect -14062 -11828 -12860 -11805
rect -12503 -11759 -11301 -11737
rect -12503 -11805 -12462 -11759
rect -11339 -11805 -11301 -11759
rect -12503 -11828 -11301 -11805
rect -10771 -11759 -9569 -11737
rect -10771 -11805 -10730 -11759
rect -9607 -11805 -9569 -11759
rect -10771 -11828 -9569 -11805
rect -9212 -11759 -8010 -11737
rect -9212 -11805 -9171 -11759
rect -8048 -11805 -8010 -11759
rect -9212 -11828 -8010 -11805
rect 7333 -11869 7372 -11118
rect -23536 -11914 -23520 -11880
rect -23429 -11914 -23413 -11880
rect -21807 -11914 -21791 -11880
rect -21700 -11914 -21684 -11880
rect 7298 -11882 7372 -11869
rect 7298 -11898 7406 -11882
rect 7756 -11106 7790 -11090
rect 7756 -11898 7790 -11882
rect 8246 -11106 8354 -11090
rect 8246 -11118 8320 -11106
rect 8281 -11869 8320 -11118
rect 8246 -11882 8320 -11869
rect 8246 -11898 8354 -11882
rect 8704 -11106 8738 -11090
rect 8704 -11898 8738 -11882
rect 9182 -11106 9290 -11090
rect 9182 -11118 9256 -11106
rect 9217 -11869 9256 -11118
rect 9182 -11882 9256 -11869
rect 9182 -11898 9290 -11882
rect 9640 -11106 9674 -11090
rect 9640 -11898 9674 -11882
rect 10113 -11106 10221 -11090
rect 10113 -11118 10187 -11106
rect 10148 -11869 10187 -11118
rect 10113 -11882 10187 -11869
rect 10113 -11898 10221 -11882
rect 10571 -11106 10605 -11090
rect 10571 -11898 10605 -11882
rect 11040 -11106 11148 -11090
rect 11040 -11118 11114 -11106
rect 11075 -11869 11114 -11118
rect 11040 -11882 11114 -11869
rect 11040 -11898 11148 -11882
rect 11498 -11106 11532 -11090
rect 11783 -11432 12203 -11412
rect 11783 -11483 11811 -11432
rect 12168 -11483 12203 -11432
rect 11783 -11502 12203 -11483
rect 11785 -11587 11819 -11502
rect 11785 -11835 11819 -11819
rect 11881 -11587 11915 -11571
rect 11881 -11835 11915 -11819
rect 11977 -11587 12011 -11502
rect 11977 -11835 12011 -11819
rect 12073 -11587 12107 -11571
rect 12073 -11835 12107 -11819
rect 12169 -11587 12203 -11502
rect 12169 -11835 12203 -11819
rect 12265 -11587 12299 -11571
rect 12265 -11835 12299 -11819
rect 12361 -11587 12395 -11571
rect 12361 -11835 12395 -11819
rect 12457 -11587 12491 -11571
rect 12457 -11835 12491 -11819
rect 12553 -11587 12587 -11571
rect 12553 -11835 12587 -11819
rect 12649 -11587 12683 -11571
rect 12649 -11835 12683 -11819
rect 12745 -11587 12779 -11571
rect 12970 -11653 12986 -11619
rect 13077 -11653 13093 -11619
rect 12745 -11835 12779 -11819
rect 12826 -11739 12876 -11722
rect 12919 -11725 12929 -11691
rect 13125 -11725 13141 -11691
rect 11498 -11898 11532 -11882
rect 12154 -11915 12170 -11881
rect 12204 -11915 12220 -11881
rect -24384 -11980 -24368 -11933
rect -23799 -11980 -23775 -11933
rect -23680 -12000 -23630 -11983
rect -23587 -11986 -23577 -11952
rect -23381 -11986 -23365 -11952
rect -22647 -11980 -22631 -11933
rect -22062 -11980 -22038 -11933
rect -24384 -12052 -24350 -12042
rect -24384 -12264 -24350 -12248
rect -24288 -12058 -24254 -12042
rect -24288 -12264 -24254 -12254
rect -24192 -12052 -24158 -12042
rect -24192 -12264 -24158 -12248
rect -24096 -12058 -24062 -12042
rect -24096 -12264 -24062 -12254
rect -24000 -12052 -23966 -12042
rect -24000 -12264 -23966 -12248
rect -23904 -12058 -23870 -12042
rect -23904 -12264 -23870 -12254
rect -23808 -12052 -23774 -12042
rect -23808 -12264 -23774 -12248
rect -23680 -12226 -23664 -12000
rect -21951 -12000 -21901 -11983
rect -21858 -11986 -21848 -11952
rect -21652 -11986 -21636 -11952
rect 12826 -11965 12842 -11739
rect 12919 -11821 12935 -11787
rect 13129 -11821 13147 -11787
rect 12919 -11917 12929 -11883
rect 13125 -11917 13141 -11883
rect -23587 -12082 -23571 -12048
rect -23377 -12082 -23359 -12048
rect -22647 -12052 -22613 -12042
rect -23587 -12178 -23577 -12144
rect -23381 -12178 -23365 -12144
rect -24335 -12342 -24318 -12307
rect -24284 -12342 -24268 -12307
rect -24046 -12313 -24029 -12307
rect -24234 -12342 -24029 -12313
rect -23995 -12342 -23979 -12307
rect -24335 -12548 -24292 -12342
rect -24234 -12347 -23979 -12342
rect -24234 -12431 -24200 -12347
rect -24166 -12436 -24150 -12402
rect -23774 -12436 -23758 -12402
rect -24234 -12482 -24200 -12466
rect -23680 -12446 -23630 -12226
rect -23587 -12274 -23571 -12240
rect -23377 -12274 -23359 -12240
rect -22647 -12264 -22613 -12248
rect -22551 -12058 -22517 -12042
rect -22551 -12264 -22517 -12254
rect -22455 -12052 -22421 -12042
rect -22455 -12264 -22421 -12248
rect -22359 -12058 -22325 -12042
rect -22359 -12264 -22325 -12254
rect -22263 -12052 -22229 -12042
rect -22263 -12264 -22229 -12248
rect -22167 -12058 -22133 -12042
rect -22167 -12264 -22133 -12254
rect -22071 -12052 -22037 -12042
rect -22071 -12264 -22037 -12248
rect -21951 -12226 -21935 -12000
rect 7298 -12034 7406 -12018
rect 7298 -12047 7372 -12034
rect -21858 -12082 -21842 -12048
rect -21648 -12082 -21630 -12048
rect -21858 -12178 -21848 -12144
rect -21652 -12178 -21636 -12144
rect -20518 -12148 -20502 -12101
rect -19933 -12148 -19909 -12101
rect -19409 -12148 -19393 -12101
rect -18824 -12148 -18800 -12101
rect -18527 -12148 -18511 -12101
rect -17942 -12148 -17918 -12101
rect -17227 -12148 -17211 -12101
rect -16642 -12148 -16618 -12101
rect -16118 -12148 -16102 -12101
rect -15533 -12148 -15509 -12101
rect -15236 -12148 -15220 -12101
rect -14651 -12148 -14627 -12101
rect -13936 -12148 -13920 -12101
rect -13351 -12148 -13327 -12101
rect -12827 -12148 -12811 -12101
rect -12242 -12148 -12218 -12101
rect -11945 -12148 -11929 -12101
rect -11360 -12148 -11336 -12101
rect -10645 -12148 -10629 -12101
rect -10060 -12148 -10036 -12101
rect -9536 -12148 -9520 -12101
rect -8951 -12148 -8927 -12101
rect -8654 -12148 -8638 -12101
rect -8069 -12148 -8045 -12101
rect -22598 -12342 -22581 -12307
rect -22547 -12342 -22531 -12307
rect -22309 -12313 -22292 -12307
rect -22497 -12342 -22292 -12313
rect -22258 -12342 -22242 -12307
rect -23587 -12436 -23571 -12402
rect -23395 -12436 -23379 -12402
rect -23680 -12480 -23664 -12446
rect -23680 -12496 -23630 -12480
rect -23587 -12524 -23571 -12490
rect -23395 -12524 -23379 -12490
rect -22598 -12548 -22555 -12342
rect -22497 -12347 -22242 -12342
rect -22497 -12431 -22463 -12347
rect -22429 -12436 -22413 -12402
rect -22037 -12436 -22021 -12402
rect -22497 -12482 -22463 -12466
rect -21951 -12446 -21901 -12226
rect -20518 -12220 -20484 -12210
rect -21858 -12274 -21842 -12240
rect -21648 -12274 -21630 -12240
rect -21858 -12436 -21842 -12402
rect -21666 -12436 -21650 -12402
rect -20518 -12432 -20484 -12416
rect -20422 -12226 -20388 -12210
rect -20422 -12432 -20388 -12422
rect -20326 -12220 -20292 -12210
rect -20326 -12432 -20292 -12416
rect -20230 -12226 -20196 -12210
rect -20230 -12432 -20196 -12422
rect -20134 -12220 -20100 -12210
rect -20134 -12432 -20100 -12416
rect -20038 -12226 -20004 -12210
rect -20038 -12432 -20004 -12422
rect -19942 -12220 -19908 -12210
rect -19942 -12432 -19908 -12416
rect -19409 -12220 -19375 -12210
rect -19409 -12432 -19375 -12416
rect -19313 -12226 -19279 -12210
rect -19313 -12432 -19279 -12422
rect -19217 -12220 -19183 -12210
rect -19217 -12432 -19183 -12416
rect -19121 -12226 -19087 -12210
rect -19121 -12432 -19087 -12422
rect -19025 -12220 -18991 -12210
rect -19025 -12432 -18991 -12416
rect -18929 -12226 -18895 -12210
rect -18929 -12432 -18895 -12422
rect -18833 -12220 -18799 -12210
rect -18833 -12432 -18799 -12416
rect -18527 -12220 -18493 -12210
rect -18527 -12432 -18493 -12416
rect -18431 -12226 -18397 -12210
rect -18431 -12432 -18397 -12422
rect -18335 -12220 -18301 -12210
rect -18335 -12432 -18301 -12416
rect -18239 -12226 -18205 -12210
rect -18239 -12432 -18205 -12422
rect -18143 -12220 -18109 -12210
rect -18143 -12432 -18109 -12416
rect -18047 -12226 -18013 -12210
rect -18047 -12432 -18013 -12422
rect -17951 -12220 -17917 -12210
rect -17951 -12432 -17917 -12416
rect -17227 -12220 -17193 -12210
rect -17227 -12432 -17193 -12416
rect -17131 -12226 -17097 -12210
rect -17131 -12432 -17097 -12422
rect -17035 -12220 -17001 -12210
rect -17035 -12432 -17001 -12416
rect -16939 -12226 -16905 -12210
rect -16939 -12432 -16905 -12422
rect -16843 -12220 -16809 -12210
rect -16843 -12432 -16809 -12416
rect -16747 -12226 -16713 -12210
rect -16747 -12432 -16713 -12422
rect -16651 -12220 -16617 -12210
rect -16651 -12432 -16617 -12416
rect -16118 -12220 -16084 -12210
rect -16118 -12432 -16084 -12416
rect -16022 -12226 -15988 -12210
rect -16022 -12432 -15988 -12422
rect -15926 -12220 -15892 -12210
rect -15926 -12432 -15892 -12416
rect -15830 -12226 -15796 -12210
rect -15830 -12432 -15796 -12422
rect -15734 -12220 -15700 -12210
rect -15734 -12432 -15700 -12416
rect -15638 -12226 -15604 -12210
rect -15638 -12432 -15604 -12422
rect -15542 -12220 -15508 -12210
rect -15542 -12432 -15508 -12416
rect -15236 -12220 -15202 -12210
rect -15236 -12432 -15202 -12416
rect -15140 -12226 -15106 -12210
rect -15140 -12432 -15106 -12422
rect -15044 -12220 -15010 -12210
rect -15044 -12432 -15010 -12416
rect -14948 -12226 -14914 -12210
rect -14948 -12432 -14914 -12422
rect -14852 -12220 -14818 -12210
rect -14852 -12432 -14818 -12416
rect -14756 -12226 -14722 -12210
rect -14756 -12432 -14722 -12422
rect -14660 -12220 -14626 -12210
rect -14660 -12432 -14626 -12416
rect -13936 -12220 -13902 -12210
rect -13936 -12432 -13902 -12416
rect -13840 -12226 -13806 -12210
rect -13840 -12432 -13806 -12422
rect -13744 -12220 -13710 -12210
rect -13744 -12432 -13710 -12416
rect -13648 -12226 -13614 -12210
rect -13648 -12432 -13614 -12422
rect -13552 -12220 -13518 -12210
rect -13552 -12432 -13518 -12416
rect -13456 -12226 -13422 -12210
rect -13456 -12432 -13422 -12422
rect -13360 -12220 -13326 -12210
rect -13360 -12432 -13326 -12416
rect -12827 -12220 -12793 -12210
rect -12827 -12432 -12793 -12416
rect -12731 -12226 -12697 -12210
rect -12731 -12432 -12697 -12422
rect -12635 -12220 -12601 -12210
rect -12635 -12432 -12601 -12416
rect -12539 -12226 -12505 -12210
rect -12539 -12432 -12505 -12422
rect -12443 -12220 -12409 -12210
rect -12443 -12432 -12409 -12416
rect -12347 -12226 -12313 -12210
rect -12347 -12432 -12313 -12422
rect -12251 -12220 -12217 -12210
rect -12251 -12432 -12217 -12416
rect -11945 -12220 -11911 -12210
rect -11945 -12432 -11911 -12416
rect -11849 -12226 -11815 -12210
rect -11849 -12432 -11815 -12422
rect -11753 -12220 -11719 -12210
rect -11753 -12432 -11719 -12416
rect -11657 -12226 -11623 -12210
rect -11657 -12432 -11623 -12422
rect -11561 -12220 -11527 -12210
rect -11561 -12432 -11527 -12416
rect -11465 -12226 -11431 -12210
rect -11465 -12432 -11431 -12422
rect -11369 -12220 -11335 -12210
rect -11369 -12432 -11335 -12416
rect -10645 -12220 -10611 -12210
rect -10645 -12432 -10611 -12416
rect -10549 -12226 -10515 -12210
rect -10549 -12432 -10515 -12422
rect -10453 -12220 -10419 -12210
rect -10453 -12432 -10419 -12416
rect -10357 -12226 -10323 -12210
rect -10357 -12432 -10323 -12422
rect -10261 -12220 -10227 -12210
rect -10261 -12432 -10227 -12416
rect -10165 -12226 -10131 -12210
rect -10165 -12432 -10131 -12422
rect -10069 -12220 -10035 -12210
rect -10069 -12432 -10035 -12416
rect -9536 -12220 -9502 -12210
rect -9536 -12432 -9502 -12416
rect -9440 -12226 -9406 -12210
rect -9440 -12432 -9406 -12422
rect -9344 -12220 -9310 -12210
rect -9344 -12432 -9310 -12416
rect -9248 -12226 -9214 -12210
rect -9248 -12432 -9214 -12422
rect -9152 -12220 -9118 -12210
rect -9152 -12432 -9118 -12416
rect -9056 -12226 -9022 -12210
rect -9056 -12432 -9022 -12422
rect -8960 -12220 -8926 -12210
rect -8960 -12432 -8926 -12416
rect -8654 -12220 -8620 -12210
rect -8654 -12432 -8620 -12416
rect -8558 -12226 -8524 -12210
rect -8558 -12432 -8524 -12422
rect -8462 -12220 -8428 -12210
rect -8462 -12432 -8428 -12416
rect -8366 -12226 -8332 -12210
rect -8366 -12432 -8332 -12422
rect -8270 -12220 -8236 -12210
rect -8270 -12432 -8236 -12416
rect -8174 -12226 -8140 -12210
rect -8174 -12432 -8140 -12422
rect -8078 -12220 -8044 -12210
rect -8078 -12432 -8044 -12416
rect -21951 -12480 -21935 -12446
rect -21951 -12496 -21901 -12480
rect -21858 -12524 -21842 -12490
rect -21666 -12524 -21650 -12490
rect -20469 -12510 -20452 -12475
rect -20418 -12510 -20402 -12475
rect -20180 -12481 -20163 -12475
rect -20368 -12510 -20163 -12481
rect -20129 -12510 -20113 -12475
rect -24335 -12564 -24200 -12548
rect -24335 -12599 -24234 -12564
rect -22598 -12564 -22463 -12548
rect -24335 -12615 -24200 -12599
rect -24166 -12628 -24150 -12594
rect -23774 -12628 -23758 -12594
rect -23568 -12626 -23552 -12592
rect -23420 -12626 -23404 -12592
rect -22598 -12599 -22497 -12564
rect -22598 -12615 -22463 -12599
rect -22429 -12628 -22413 -12594
rect -22037 -12628 -22021 -12594
rect -21839 -12626 -21823 -12592
rect -21691 -12626 -21675 -12592
rect -24162 -12700 -24135 -12666
rect -23800 -12700 -23762 -12666
rect -22425 -12700 -22398 -12666
rect -22063 -12700 -22025 -12666
rect -20469 -12716 -20426 -12510
rect -20368 -12515 -20113 -12510
rect -19360 -12510 -19343 -12475
rect -19309 -12510 -19293 -12475
rect -19071 -12481 -19054 -12475
rect -19259 -12510 -19054 -12481
rect -19020 -12510 -19004 -12475
rect -20368 -12599 -20334 -12515
rect -20300 -12604 -20284 -12570
rect -19908 -12604 -19892 -12570
rect -20368 -12650 -20334 -12634
rect -19360 -12716 -19317 -12510
rect -19259 -12515 -19004 -12510
rect -18478 -12510 -18461 -12475
rect -18427 -12510 -18411 -12475
rect -18189 -12481 -18172 -12475
rect -18377 -12510 -18172 -12481
rect -18138 -12510 -18122 -12475
rect -19259 -12599 -19225 -12515
rect -19191 -12604 -19175 -12570
rect -18799 -12604 -18783 -12570
rect -19259 -12650 -19225 -12634
rect -18478 -12716 -18435 -12510
rect -18377 -12515 -18122 -12510
rect -17178 -12510 -17161 -12475
rect -17127 -12510 -17111 -12475
rect -16889 -12481 -16872 -12475
rect -17077 -12510 -16872 -12481
rect -16838 -12510 -16822 -12475
rect -18377 -12599 -18343 -12515
rect -18309 -12604 -18293 -12570
rect -17917 -12604 -17901 -12570
rect -18377 -12650 -18343 -12634
rect -17178 -12716 -17135 -12510
rect -17077 -12515 -16822 -12510
rect -16069 -12510 -16052 -12475
rect -16018 -12510 -16002 -12475
rect -15780 -12481 -15763 -12475
rect -15968 -12510 -15763 -12481
rect -15729 -12510 -15713 -12475
rect -17077 -12599 -17043 -12515
rect -17009 -12604 -16993 -12570
rect -16617 -12604 -16601 -12570
rect -17077 -12650 -17043 -12634
rect -16069 -12716 -16026 -12510
rect -15968 -12515 -15713 -12510
rect -15187 -12510 -15170 -12475
rect -15136 -12510 -15120 -12475
rect -14898 -12481 -14881 -12475
rect -15086 -12510 -14881 -12481
rect -14847 -12510 -14831 -12475
rect -15968 -12599 -15934 -12515
rect -15900 -12604 -15884 -12570
rect -15508 -12604 -15492 -12570
rect -15968 -12650 -15934 -12634
rect -15187 -12716 -15144 -12510
rect -15086 -12515 -14831 -12510
rect -13887 -12510 -13870 -12475
rect -13836 -12510 -13820 -12475
rect -13598 -12481 -13581 -12475
rect -13786 -12510 -13581 -12481
rect -13547 -12510 -13531 -12475
rect -15086 -12599 -15052 -12515
rect -15018 -12604 -15002 -12570
rect -14626 -12604 -14610 -12570
rect -15086 -12650 -15052 -12634
rect -13887 -12716 -13844 -12510
rect -13786 -12515 -13531 -12510
rect -12778 -12510 -12761 -12475
rect -12727 -12510 -12711 -12475
rect -12489 -12481 -12472 -12475
rect -12677 -12510 -12472 -12481
rect -12438 -12510 -12422 -12475
rect -13786 -12599 -13752 -12515
rect -13718 -12604 -13702 -12570
rect -13326 -12604 -13310 -12570
rect -13786 -12650 -13752 -12634
rect -12778 -12716 -12735 -12510
rect -12677 -12515 -12422 -12510
rect -11896 -12510 -11879 -12475
rect -11845 -12510 -11829 -12475
rect -11607 -12481 -11590 -12475
rect -11795 -12510 -11590 -12481
rect -11556 -12510 -11540 -12475
rect -12677 -12599 -12643 -12515
rect -12609 -12604 -12593 -12570
rect -12217 -12604 -12201 -12570
rect -12677 -12650 -12643 -12634
rect -11896 -12716 -11853 -12510
rect -11795 -12515 -11540 -12510
rect -10596 -12510 -10579 -12475
rect -10545 -12510 -10529 -12475
rect -10307 -12481 -10290 -12475
rect -10495 -12510 -10290 -12481
rect -10256 -12510 -10240 -12475
rect -11795 -12599 -11761 -12515
rect -11727 -12604 -11711 -12570
rect -11335 -12604 -11319 -12570
rect -11795 -12650 -11761 -12634
rect -10596 -12716 -10553 -12510
rect -10495 -12515 -10240 -12510
rect -9487 -12510 -9470 -12475
rect -9436 -12510 -9420 -12475
rect -9198 -12481 -9181 -12475
rect -9386 -12510 -9181 -12481
rect -9147 -12510 -9131 -12475
rect -10495 -12599 -10461 -12515
rect -10427 -12604 -10411 -12570
rect -10035 -12604 -10019 -12570
rect -10495 -12650 -10461 -12634
rect -9487 -12716 -9444 -12510
rect -9386 -12515 -9131 -12510
rect -8605 -12510 -8588 -12475
rect -8554 -12510 -8538 -12475
rect -8316 -12481 -8299 -12475
rect -8504 -12510 -8299 -12481
rect -8265 -12510 -8249 -12475
rect -9386 -12599 -9352 -12515
rect -9318 -12604 -9302 -12570
rect -8926 -12604 -8910 -12570
rect -9386 -12650 -9352 -12634
rect -8605 -12716 -8562 -12510
rect -8504 -12515 -8249 -12510
rect -8504 -12599 -8470 -12515
rect -8436 -12604 -8420 -12570
rect -8044 -12604 -8028 -12570
rect -8504 -12650 -8470 -12634
rect -20469 -12732 -20334 -12716
rect -20469 -12767 -20368 -12732
rect -19360 -12732 -19225 -12716
rect -20469 -12783 -20334 -12767
rect -20300 -12796 -20284 -12762
rect -19908 -12796 -19892 -12762
rect -19360 -12767 -19259 -12732
rect -18478 -12732 -18343 -12716
rect -19360 -12783 -19225 -12767
rect -19191 -12796 -19175 -12762
rect -18799 -12796 -18783 -12762
rect -18478 -12767 -18377 -12732
rect -17178 -12732 -17043 -12716
rect -18478 -12783 -18343 -12767
rect -18309 -12796 -18293 -12762
rect -17917 -12796 -17901 -12762
rect -17178 -12767 -17077 -12732
rect -16069 -12732 -15934 -12716
rect -17178 -12783 -17043 -12767
rect -17009 -12796 -16993 -12762
rect -16617 -12796 -16601 -12762
rect -16069 -12767 -15968 -12732
rect -15187 -12732 -15052 -12716
rect -16069 -12783 -15934 -12767
rect -15900 -12796 -15884 -12762
rect -15508 -12796 -15492 -12762
rect -15187 -12767 -15086 -12732
rect -13887 -12732 -13752 -12716
rect -15187 -12783 -15052 -12767
rect -15018 -12796 -15002 -12762
rect -14626 -12796 -14610 -12762
rect -13887 -12767 -13786 -12732
rect -12778 -12732 -12643 -12716
rect -13887 -12783 -13752 -12767
rect -13718 -12796 -13702 -12762
rect -13326 -12796 -13310 -12762
rect -12778 -12767 -12677 -12732
rect -11896 -12732 -11761 -12716
rect -12778 -12783 -12643 -12767
rect -12609 -12796 -12593 -12762
rect -12217 -12796 -12201 -12762
rect -11896 -12767 -11795 -12732
rect -10596 -12732 -10461 -12716
rect -11896 -12783 -11761 -12767
rect -11727 -12796 -11711 -12762
rect -11335 -12796 -11319 -12762
rect -10596 -12767 -10495 -12732
rect -9487 -12732 -9352 -12716
rect -10596 -12783 -10461 -12767
rect -10427 -12796 -10411 -12762
rect -10035 -12796 -10019 -12762
rect -9487 -12767 -9386 -12732
rect -8605 -12732 -8470 -12716
rect -9487 -12783 -9352 -12767
rect -9318 -12796 -9302 -12762
rect -8926 -12796 -8910 -12762
rect -8605 -12767 -8504 -12732
rect -8605 -12783 -8470 -12767
rect -8436 -12796 -8420 -12762
rect -8044 -12796 -8028 -12762
rect 7333 -12798 7372 -12047
rect 7298 -12810 7372 -12798
rect 7298 -12826 7406 -12810
rect 7756 -12034 7790 -12018
rect 7756 -12826 7790 -12810
rect 8246 -12034 8354 -12018
rect 8246 -12047 8320 -12034
rect 8281 -12798 8320 -12047
rect 8246 -12810 8320 -12798
rect 8246 -12826 8354 -12810
rect 8704 -12034 8738 -12018
rect 8704 -12826 8738 -12810
rect 9182 -12034 9290 -12018
rect 9182 -12047 9256 -12034
rect 9217 -12798 9256 -12047
rect 9182 -12810 9256 -12798
rect 9182 -12826 9290 -12810
rect 9640 -12034 9674 -12018
rect 9640 -12826 9674 -12810
rect 10113 -12033 10221 -12017
rect 10113 -12046 10187 -12033
rect 10148 -12797 10187 -12046
rect 10113 -12809 10187 -12797
rect 10113 -12825 10221 -12809
rect 10571 -12033 10605 -12017
rect 10571 -12825 10605 -12809
rect 11040 -12034 11148 -12018
rect 11040 -12047 11114 -12034
rect 11075 -12798 11114 -12047
rect 11040 -12810 11114 -12798
rect 7298 -12829 7403 -12826
rect 8246 -12829 8351 -12826
rect 9182 -12829 9287 -12826
rect 10113 -12828 10218 -12825
rect 11040 -12826 11148 -12810
rect 11498 -12034 11532 -12018
rect 12297 -12020 12313 -11986
rect 12347 -12020 12363 -11986
rect 12169 -12076 12203 -12060
rect 12169 -12324 12203 -12252
rect 12265 -12076 12299 -12060
rect 12265 -12268 12299 -12252
rect 12361 -12076 12395 -12060
rect 12826 -12185 12876 -11965
rect 12919 -12013 12935 -11979
rect 13129 -12013 13147 -11979
rect 12919 -12175 12935 -12141
rect 13111 -12175 13127 -12141
rect 12826 -12219 12842 -12185
rect 12826 -12235 12876 -12219
rect 12361 -12324 12395 -12252
rect 12919 -12263 12935 -12229
rect 13111 -12263 13127 -12229
rect 12157 -12335 12407 -12324
rect 12157 -12396 12183 -12335
rect 12382 -12396 12407 -12335
rect 12938 -12365 12954 -12331
rect 13086 -12365 13102 -12331
rect 12157 -12408 12407 -12396
rect 11498 -12826 11532 -12810
rect 11040 -12829 11145 -12826
rect -20296 -12868 -20269 -12834
rect -19934 -12868 -19896 -12834
rect -19187 -12868 -19160 -12834
rect -18825 -12868 -18787 -12834
rect -18305 -12868 -18278 -12834
rect -17943 -12868 -17905 -12834
rect -17005 -12868 -16978 -12834
rect -16643 -12868 -16605 -12834
rect -15896 -12868 -15869 -12834
rect -15534 -12868 -15496 -12834
rect -15014 -12868 -14987 -12834
rect -14652 -12868 -14614 -12834
rect -13714 -12868 -13687 -12834
rect -13352 -12868 -13314 -12834
rect -12605 -12868 -12578 -12834
rect -12243 -12868 -12205 -12834
rect -11723 -12868 -11696 -12834
rect -11361 -12868 -11323 -12834
rect -10423 -12868 -10396 -12834
rect -10061 -12868 -10023 -12834
rect -9314 -12868 -9287 -12834
rect -8952 -12868 -8914 -12834
rect -8432 -12868 -8405 -12834
rect -8070 -12868 -8032 -12834
rect 7182 -13182 7198 -13148
rect 7232 -13182 7248 -13148
rect 7374 -13182 7390 -13148
rect 7424 -13182 7440 -13148
rect 7566 -13182 7582 -13148
rect 7616 -13182 7632 -13148
rect 7758 -13182 7774 -13148
rect 7808 -13182 7824 -13148
rect 8130 -13182 8146 -13148
rect 8180 -13182 8196 -13148
rect 8322 -13182 8338 -13148
rect 8372 -13182 8388 -13148
rect 8514 -13182 8530 -13148
rect 8564 -13182 8580 -13148
rect 8706 -13182 8722 -13148
rect 8756 -13182 8772 -13148
rect 9066 -13182 9082 -13148
rect 9116 -13182 9132 -13148
rect 9258 -13182 9274 -13148
rect 9308 -13182 9324 -13148
rect 9450 -13182 9466 -13148
rect 9500 -13182 9516 -13148
rect 9642 -13182 9658 -13148
rect 9692 -13182 9708 -13148
rect 9997 -13181 10013 -13147
rect 10047 -13181 10063 -13147
rect 10189 -13181 10205 -13147
rect 10239 -13181 10255 -13147
rect 10381 -13181 10397 -13147
rect 10431 -13181 10447 -13147
rect 10573 -13181 10589 -13147
rect 10623 -13181 10639 -13147
rect 10924 -13182 10940 -13148
rect 10974 -13182 10990 -13148
rect 11116 -13182 11132 -13148
rect 11166 -13182 11182 -13148
rect 11308 -13182 11324 -13148
rect 11358 -13182 11374 -13148
rect 11500 -13182 11516 -13148
rect 11550 -13182 11566 -13148
rect 7150 -13241 7184 -13225
rect 7246 -13236 7280 -13225
rect 7150 -13555 7184 -13539
rect 7246 -13555 7280 -13539
rect 7342 -13241 7376 -13225
rect 7342 -13555 7376 -13539
rect 7438 -13236 7472 -13225
rect 7534 -13241 7568 -13225
rect 7438 -13555 7472 -13539
rect 7534 -13555 7568 -13539
rect 7630 -13236 7664 -13225
rect 7726 -13241 7760 -13225
rect 7630 -13555 7664 -13539
rect 7726 -13555 7760 -13539
rect 7822 -13236 7856 -13225
rect 7918 -13241 7952 -13225
rect 7822 -13555 7856 -13539
rect 7918 -13555 7952 -13539
rect 8098 -13241 8132 -13225
rect 8194 -13236 8228 -13225
rect 8098 -13555 8132 -13539
rect 8194 -13555 8228 -13539
rect 8290 -13241 8324 -13225
rect 8290 -13555 8324 -13539
rect 8386 -13236 8420 -13225
rect 8482 -13241 8516 -13225
rect 8386 -13555 8420 -13539
rect 8482 -13555 8516 -13539
rect 8578 -13236 8612 -13225
rect 8674 -13241 8708 -13225
rect 8578 -13555 8612 -13539
rect 8674 -13555 8708 -13539
rect 8770 -13236 8804 -13225
rect 8866 -13241 8900 -13225
rect 8770 -13555 8804 -13539
rect 8866 -13555 8900 -13539
rect 9034 -13241 9068 -13225
rect 9130 -13236 9164 -13225
rect 9034 -13555 9068 -13539
rect 9130 -13555 9164 -13539
rect 9226 -13241 9260 -13225
rect 9226 -13555 9260 -13539
rect 9322 -13236 9356 -13225
rect 9418 -13241 9452 -13225
rect 9322 -13555 9356 -13539
rect 9418 -13555 9452 -13539
rect 9514 -13236 9548 -13225
rect 9610 -13241 9644 -13225
rect 9514 -13555 9548 -13539
rect 9610 -13555 9644 -13539
rect 9706 -13236 9740 -13225
rect 9802 -13241 9836 -13225
rect 9706 -13555 9740 -13539
rect 9802 -13555 9836 -13539
rect 9965 -13240 9999 -13224
rect 10061 -13235 10095 -13224
rect 9965 -13554 9999 -13538
rect 10061 -13554 10095 -13538
rect 10157 -13240 10191 -13224
rect 10157 -13554 10191 -13538
rect 10253 -13235 10287 -13224
rect 10349 -13240 10383 -13224
rect 10253 -13554 10287 -13538
rect 10349 -13554 10383 -13538
rect 10445 -13235 10479 -13224
rect 10541 -13240 10575 -13224
rect 10445 -13554 10479 -13538
rect 10541 -13554 10575 -13538
rect 10637 -13235 10671 -13224
rect 10733 -13240 10767 -13224
rect 10637 -13554 10671 -13538
rect 10733 -13554 10767 -13538
rect 10892 -13241 10926 -13225
rect 10988 -13236 11022 -13225
rect 10892 -13555 10926 -13539
rect 10988 -13555 11022 -13539
rect 11084 -13241 11118 -13225
rect 11084 -13555 11118 -13539
rect 11180 -13236 11214 -13225
rect 11276 -13241 11310 -13225
rect 11180 -13555 11214 -13539
rect 11276 -13555 11310 -13539
rect 11372 -13236 11406 -13225
rect 11468 -13241 11502 -13225
rect 11372 -13555 11406 -13539
rect 11468 -13555 11502 -13539
rect 11564 -13236 11598 -13225
rect 11660 -13241 11694 -13225
rect 11564 -13555 11598 -13539
rect 11660 -13555 11694 -13539
rect 7373 -13643 7389 -13608
rect 7677 -13643 7703 -13608
rect 8321 -13643 8337 -13608
rect 8625 -13643 8651 -13608
rect 9257 -13643 9273 -13608
rect 9561 -13643 9587 -13608
rect 10188 -13642 10204 -13607
rect 10492 -13642 10518 -13607
rect 11115 -13643 11131 -13608
rect 11419 -13643 11445 -13608
rect -2100 -13830 -2066 -13814
rect -2172 -13878 -2138 -13862
rect -2172 -13985 -2138 -13969
rect -2100 -14036 -2066 -14026
rect -2004 -13826 -1970 -13808
rect -2004 -14036 -1970 -14020
rect -1908 -13830 -1874 -13814
rect -1908 -14036 -1874 -14026
rect -1812 -13826 -1778 -13808
rect -1812 -14036 -1778 -14020
rect -1650 -13844 -1616 -13828
rect -1650 -14036 -1616 -14020
rect -1562 -13844 -1528 -13828
rect -1460 -13869 -1426 -13853
rect -1460 -14017 -1426 -14001
rect -1562 -14036 -1528 -14020
rect -12320 -14139 -12304 -14105
rect -11778 -14139 -11264 -14105
rect -11158 -14139 -11142 -14105
rect -4785 -14122 -4272 -14106
rect -12501 -14223 -12375 -14181
rect -17681 -14545 -17665 -14511
rect -17433 -14545 -17417 -14511
rect -17681 -14641 -17665 -14607
rect -17433 -14641 -17417 -14607
rect -17681 -14737 -17665 -14703
rect -17433 -14737 -17417 -14703
rect -17681 -14833 -17665 -14799
rect -17433 -14833 -17417 -14799
rect -16928 -14895 -16844 -14883
rect -24093 -14928 -24059 -14912
rect -24562 -14953 -24515 -14929
rect -24453 -14962 -24443 -14928
rect -24247 -14962 -24231 -14928
rect -24453 -15058 -24437 -15024
rect -24241 -15058 -24231 -15024
rect -24453 -15154 -24443 -15120
rect -24247 -15154 -24231 -15120
rect -24188 -15149 -24148 -15133
rect -24153 -15183 -24148 -15149
rect -24188 -15200 -24148 -15183
rect -24453 -15250 -24437 -15216
rect -24241 -15250 -24231 -15216
rect -24453 -15346 -24443 -15312
rect -24247 -15346 -24231 -15312
rect -24182 -15354 -24148 -15200
rect -24093 -15320 -24059 -15304
rect -23901 -14928 -23867 -14912
rect -23901 -15320 -23867 -15304
rect -23829 -14954 -23795 -14916
rect -17681 -14929 -17665 -14895
rect -17433 -14929 -17417 -14895
rect -17266 -14943 -17232 -14927
rect -17192 -14929 -17176 -14895
rect -17000 -14908 -16844 -14895
rect -17000 -14929 -16917 -14908
rect -17681 -15025 -17665 -14991
rect -17433 -15025 -17417 -14991
rect -17266 -14993 -17232 -14977
rect -17192 -15025 -17176 -14991
rect -17000 -15025 -16984 -14991
rect -17371 -15086 -17337 -15070
rect -23829 -15316 -23795 -15289
rect -17840 -15121 -17665 -15087
rect -17433 -15121 -17417 -15087
rect -16928 -15087 -16917 -14929
rect -17840 -15122 -17750 -15121
rect -24182 -15388 -24064 -15354
rect -24029 -15388 -24013 -15354
rect -23947 -15388 -23931 -15354
rect -23896 -15388 -23880 -15354
rect -24453 -15442 -24437 -15408
rect -24241 -15442 -24231 -15408
rect -24188 -15438 -24153 -15422
rect -23947 -15446 -23880 -15388
rect -24153 -15472 -23880 -15446
rect -24188 -15489 -23880 -15472
rect -17840 -15479 -17820 -15122
rect -17769 -15279 -17750 -15122
rect -17371 -15136 -17337 -15120
rect -17192 -15121 -17176 -15087
rect -17000 -15107 -16917 -15087
rect -16856 -15107 -16844 -14908
rect -17000 -15121 -16844 -15107
rect -16928 -15133 -16844 -15121
rect -17681 -15217 -17665 -15183
rect -17433 -15217 -17417 -15183
rect -17769 -15313 -17665 -15279
rect -17433 -15313 -17417 -15279
rect -17769 -15471 -17750 -15313
rect -12501 -15345 -12473 -14223
rect -12401 -15345 -12375 -14223
rect -12320 -14227 -12304 -14193
rect -11778 -14227 -11762 -14193
rect -12320 -14323 -12304 -14289
rect -11778 -14323 -11762 -14289
rect -12320 -14419 -12304 -14385
rect -11778 -14419 -11762 -14385
rect -12320 -14515 -12304 -14481
rect -11778 -14515 -11762 -14481
rect -11720 -14530 -11643 -14139
rect -4785 -14156 -4768 -14122
rect -4542 -14156 -4322 -14122
rect -4288 -14156 -4272 -14122
rect -2069 -14113 -2052 -14079
rect -1826 -14113 -1606 -14079
rect -1572 -14113 -1556 -14079
rect -2069 -14129 -1556 -14113
rect 5705 -14163 5721 -14129
rect 5812 -14163 5828 -14129
rect 6145 -14163 6161 -14129
rect 6252 -14163 6268 -14129
rect 6585 -14163 6601 -14129
rect 6692 -14163 6708 -14129
rect -11435 -14194 -11339 -14179
rect -11435 -14259 -11413 -14194
rect -11358 -14259 -11339 -14194
rect -11280 -14227 -11264 -14193
rect -11158 -14227 -11142 -14193
rect -11092 -14222 -11001 -14184
rect -11602 -14361 -11496 -14343
rect -11602 -14441 -11584 -14361
rect -11516 -14441 -11496 -14361
rect -11602 -14458 -11496 -14441
rect -11720 -14550 -11503 -14530
rect -12320 -14611 -12304 -14577
rect -11778 -14611 -11762 -14577
rect -12320 -14707 -12304 -14673
rect -11778 -14707 -11762 -14673
rect -11720 -14680 -11702 -14550
rect -11657 -14561 -11503 -14550
rect -11657 -14675 -11585 -14561
rect -11532 -14675 -11503 -14561
rect -11657 -14680 -11503 -14675
rect -11720 -14707 -11503 -14680
rect -11435 -14753 -11339 -14259
rect -11280 -14323 -11279 -14289
rect -11158 -14323 -11142 -14289
rect -11280 -14419 -11264 -14385
rect -11144 -14419 -11142 -14385
rect -11280 -14515 -11279 -14481
rect -11158 -14515 -11142 -14481
rect -11280 -14611 -11264 -14577
rect -11144 -14611 -11142 -14577
rect -11280 -14707 -11279 -14673
rect -11158 -14707 -11142 -14673
rect -11735 -14769 -11305 -14753
rect -12320 -14803 -12304 -14769
rect -11778 -14803 -11264 -14769
rect -11144 -14803 -11142 -14769
rect -11735 -14819 -11305 -14803
rect -12320 -14899 -12304 -14865
rect -11778 -14899 -11762 -14865
rect -11717 -14873 -11316 -14865
rect -11717 -14881 -11378 -14873
rect -12320 -14995 -12304 -14961
rect -11778 -14995 -11762 -14961
rect -11717 -15011 -11707 -14881
rect -11662 -15003 -11378 -14881
rect -11333 -15003 -11316 -14873
rect -11280 -14899 -11278 -14865
rect -11158 -14899 -11142 -14865
rect -11280 -14995 -11264 -14961
rect -11144 -14995 -11142 -14961
rect -11662 -15011 -11316 -15003
rect -11717 -15030 -11316 -15011
rect -12320 -15091 -12304 -15057
rect -11778 -15091 -11762 -15057
rect -12320 -15187 -12304 -15153
rect -11778 -15187 -11762 -15153
rect -12320 -15283 -12304 -15249
rect -11778 -15283 -11762 -15249
rect -17681 -15409 -17665 -15375
rect -17433 -15409 -17417 -15375
rect -12501 -15391 -12375 -15345
rect -12320 -15379 -12304 -15345
rect -11778 -15379 -11762 -15345
rect -11717 -15433 -11648 -15030
rect -11280 -15091 -11279 -15057
rect -11158 -15091 -11142 -15057
rect -11604 -15148 -11314 -15110
rect -11604 -15281 -11577 -15148
rect -11524 -15156 -11314 -15148
rect -11524 -15281 -11386 -15156
rect -11604 -15286 -11386 -15281
rect -11341 -15286 -11314 -15156
rect -11280 -15187 -11264 -15153
rect -11144 -15187 -11142 -15153
rect -11280 -15283 -11279 -15249
rect -11158 -15283 -11142 -15249
rect -11604 -15331 -11314 -15286
rect -11092 -15345 -11070 -14222
rect -11024 -15345 -11001 -14222
rect -4816 -14209 -4782 -14199
rect -4888 -14266 -4854 -14250
rect -4888 -14373 -4854 -14357
rect -4816 -14421 -4782 -14405
rect -4720 -14215 -4686 -14199
rect -4720 -14427 -4686 -14409
rect -4624 -14209 -4590 -14199
rect -4624 -14421 -4590 -14405
rect -4528 -14215 -4494 -14199
rect -4366 -14215 -4332 -14199
rect -4366 -14407 -4332 -14391
rect -4278 -14215 -4244 -14199
rect -2100 -14209 -2066 -14193
rect -4176 -14234 -4142 -14218
rect -2172 -14257 -2138 -14241
rect -2172 -14364 -2138 -14348
rect -4176 -14382 -4142 -14366
rect -4278 -14407 -4244 -14391
rect -4528 -14427 -4494 -14409
rect -2100 -14415 -2066 -14405
rect -2004 -14205 -1970 -14187
rect -2004 -14415 -1970 -14399
rect -1908 -14209 -1874 -14193
rect -1908 -14415 -1874 -14405
rect -1812 -14205 -1778 -14187
rect -1812 -14415 -1778 -14399
rect -1650 -14223 -1616 -14207
rect -1650 -14415 -1616 -14399
rect -1562 -14223 -1528 -14207
rect -1460 -14248 -1426 -14232
rect -1460 -14396 -1426 -14380
rect 5561 -14249 5611 -14232
rect 5654 -14235 5664 -14201
rect 5860 -14235 5876 -14201
rect -1562 -14415 -1528 -14399
rect -2069 -14492 -2052 -14458
rect -1826 -14492 -1606 -14458
rect -1572 -14492 -1556 -14458
rect -2069 -14508 -1556 -14492
rect 5561 -14475 5577 -14249
rect 6001 -14249 6051 -14232
rect 6094 -14235 6104 -14201
rect 6300 -14235 6316 -14201
rect 5654 -14331 5670 -14297
rect 5864 -14331 5882 -14297
rect 5654 -14427 5664 -14393
rect 5860 -14427 5876 -14393
rect -4785 -14562 -4272 -14546
rect -4785 -14596 -4768 -14562
rect -4542 -14596 -4322 -14562
rect -4288 -14596 -4272 -14562
rect -4816 -14649 -4782 -14639
rect -4888 -14706 -4854 -14690
rect -4888 -14813 -4854 -14797
rect -4816 -14861 -4782 -14845
rect -4720 -14655 -4686 -14639
rect -4720 -14867 -4686 -14849
rect -4624 -14649 -4590 -14639
rect -4624 -14861 -4590 -14845
rect -4528 -14655 -4494 -14639
rect -4366 -14655 -4332 -14639
rect -4366 -14847 -4332 -14831
rect -4278 -14655 -4244 -14639
rect -2100 -14649 -2066 -14633
rect -4176 -14674 -4142 -14658
rect -2172 -14697 -2138 -14681
rect -2172 -14804 -2138 -14788
rect -4176 -14822 -4142 -14806
rect -4278 -14847 -4244 -14831
rect -4528 -14867 -4494 -14849
rect -2100 -14855 -2066 -14845
rect -2004 -14645 -1970 -14627
rect -2004 -14855 -1970 -14839
rect -1908 -14649 -1874 -14633
rect -1908 -14855 -1874 -14845
rect -1812 -14645 -1778 -14627
rect -1812 -14855 -1778 -14839
rect -1650 -14663 -1616 -14647
rect -1650 -14855 -1616 -14839
rect -1562 -14663 -1528 -14647
rect -1460 -14688 -1426 -14672
rect 5561 -14695 5611 -14475
rect 6001 -14475 6017 -14249
rect 6441 -14249 6491 -14232
rect 6534 -14235 6544 -14201
rect 6740 -14235 6756 -14201
rect 6094 -14331 6110 -14297
rect 6304 -14331 6322 -14297
rect 6094 -14427 6104 -14393
rect 6300 -14427 6316 -14393
rect 5654 -14523 5670 -14489
rect 5864 -14523 5882 -14489
rect 5654 -14685 5670 -14651
rect 5846 -14685 5862 -14651
rect 5561 -14729 5577 -14695
rect 5561 -14745 5611 -14729
rect 6001 -14695 6051 -14475
rect 6441 -14475 6457 -14249
rect 6534 -14331 6550 -14297
rect 6744 -14331 6762 -14297
rect 6534 -14427 6544 -14393
rect 6740 -14427 6756 -14393
rect 6094 -14523 6110 -14489
rect 6304 -14523 6322 -14489
rect 6094 -14685 6110 -14651
rect 6286 -14685 6302 -14651
rect 6001 -14729 6017 -14695
rect 5654 -14773 5670 -14739
rect 5846 -14773 5862 -14739
rect 6001 -14745 6051 -14729
rect 6441 -14695 6491 -14475
rect 6534 -14523 6550 -14489
rect 6744 -14523 6762 -14489
rect 6534 -14685 6550 -14651
rect 6726 -14685 6742 -14651
rect 6441 -14729 6457 -14695
rect 6094 -14773 6110 -14739
rect 6286 -14773 6302 -14739
rect 6441 -14745 6491 -14729
rect 6534 -14773 6550 -14739
rect 6726 -14773 6742 -14739
rect -1460 -14836 -1426 -14820
rect 7373 -14836 7389 -14801
rect 7677 -14836 7703 -14801
rect 8321 -14836 8337 -14801
rect 8625 -14836 8651 -14801
rect 9257 -14836 9273 -14801
rect 9561 -14836 9587 -14801
rect 10188 -14836 10204 -14801
rect 10492 -14836 10518 -14801
rect 11115 -14836 11131 -14801
rect 11419 -14836 11445 -14801
rect -1562 -14855 -1528 -14839
rect 5673 -14875 5689 -14841
rect 5821 -14875 5837 -14841
rect 6113 -14875 6129 -14841
rect 6261 -14875 6277 -14841
rect 6553 -14875 6569 -14841
rect 6701 -14875 6717 -14841
rect -4785 -14941 -4272 -14925
rect -4785 -14975 -4768 -14941
rect -4542 -14975 -4322 -14941
rect -4288 -14975 -4272 -14941
rect -2069 -14932 -2052 -14898
rect -1826 -14932 -1606 -14898
rect -1572 -14932 -1556 -14898
rect -2069 -14948 -1556 -14932
rect 7150 -14905 7184 -14889
rect -4816 -15028 -4782 -15018
rect -4888 -15085 -4854 -15069
rect -4888 -15192 -4854 -15176
rect -4816 -15240 -4782 -15224
rect -4720 -15034 -4686 -15018
rect -4720 -15246 -4686 -15228
rect -4624 -15028 -4590 -15018
rect -4624 -15240 -4590 -15224
rect -4528 -15034 -4494 -15018
rect -4366 -15034 -4332 -15018
rect -4366 -15226 -4332 -15210
rect -4278 -15034 -4244 -15018
rect -2100 -15028 -2066 -15012
rect -4176 -15053 -4142 -15037
rect -2172 -15076 -2138 -15060
rect -2172 -15183 -2138 -15167
rect -4176 -15201 -4142 -15185
rect -4278 -15226 -4244 -15210
rect -4528 -15246 -4494 -15228
rect -2100 -15234 -2066 -15224
rect -2004 -15024 -1970 -15006
rect -2004 -15234 -1970 -15218
rect -1908 -15028 -1874 -15012
rect -1908 -15234 -1874 -15224
rect -1812 -15024 -1778 -15006
rect -1812 -15234 -1778 -15218
rect -1650 -15042 -1616 -15026
rect -1650 -15234 -1616 -15218
rect -1562 -15042 -1528 -15026
rect -1460 -15067 -1426 -15051
rect -1460 -15215 -1426 -15199
rect 7246 -14905 7280 -14889
rect -1562 -15234 -1528 -15218
rect 7150 -15219 7184 -15203
rect 7246 -15219 7280 -15208
rect 7342 -14905 7376 -14889
rect 7342 -15219 7376 -15203
rect 7438 -14905 7472 -14889
rect 7534 -14905 7568 -14889
rect 7438 -15219 7472 -15208
rect 7534 -15219 7568 -15203
rect 7630 -14905 7664 -14889
rect 7726 -14905 7760 -14889
rect 7630 -15219 7664 -15208
rect 7726 -15219 7760 -15203
rect 7822 -14905 7856 -14889
rect 7918 -14905 7952 -14889
rect 7822 -15219 7856 -15208
rect 7918 -15219 7952 -15203
rect 8098 -14905 8132 -14889
rect 8194 -14905 8228 -14889
rect 8098 -15219 8132 -15203
rect 8194 -15219 8228 -15208
rect 8290 -14905 8324 -14889
rect 8290 -15219 8324 -15203
rect 8386 -14905 8420 -14889
rect 8482 -14905 8516 -14889
rect 8386 -15219 8420 -15208
rect 8482 -15219 8516 -15203
rect 8578 -14905 8612 -14889
rect 8674 -14905 8708 -14889
rect 8578 -15219 8612 -15208
rect 8674 -15219 8708 -15203
rect 8770 -14905 8804 -14889
rect 8866 -14905 8900 -14889
rect 8770 -15219 8804 -15208
rect 8866 -15219 8900 -15203
rect 9034 -14905 9068 -14889
rect 9130 -14905 9164 -14889
rect 9034 -15219 9068 -15203
rect 9130 -15219 9164 -15208
rect 9226 -14905 9260 -14889
rect 9226 -15219 9260 -15203
rect 9322 -14905 9356 -14889
rect 9418 -14905 9452 -14889
rect 9322 -15219 9356 -15208
rect 9418 -15219 9452 -15203
rect 9514 -14905 9548 -14889
rect 9610 -14905 9644 -14889
rect 9514 -15219 9548 -15208
rect 9610 -15219 9644 -15203
rect 9706 -14905 9740 -14889
rect 9802 -14905 9836 -14889
rect 9706 -15219 9740 -15208
rect 9802 -15219 9836 -15203
rect 9965 -14905 9999 -14889
rect 10061 -14905 10095 -14889
rect 9965 -15219 9999 -15203
rect 10061 -15219 10095 -15208
rect 10157 -14905 10191 -14889
rect 10157 -15219 10191 -15203
rect 10253 -14905 10287 -14889
rect 10349 -14905 10383 -14889
rect 10253 -15219 10287 -15208
rect 10349 -15219 10383 -15203
rect 10445 -14905 10479 -14889
rect 10541 -14905 10575 -14889
rect 10445 -15219 10479 -15208
rect 10541 -15219 10575 -15203
rect 10637 -14905 10671 -14889
rect 10733 -14905 10767 -14889
rect 10637 -15219 10671 -15208
rect 10733 -15219 10767 -15203
rect 10892 -14905 10926 -14889
rect 10988 -14905 11022 -14889
rect 10892 -15219 10926 -15203
rect 10988 -15219 11022 -15208
rect 11084 -14905 11118 -14889
rect 11084 -15219 11118 -15203
rect 11180 -14905 11214 -14889
rect 11276 -14905 11310 -14889
rect 11180 -15219 11214 -15208
rect 11276 -15219 11310 -15203
rect 11372 -14905 11406 -14889
rect 11468 -14905 11502 -14889
rect 11372 -15219 11406 -15208
rect 11468 -15219 11502 -15203
rect 11564 -14905 11598 -14889
rect 11660 -14905 11694 -14889
rect 11564 -15219 11598 -15208
rect 11660 -15219 11694 -15203
rect -2069 -15311 -2052 -15277
rect -1826 -15311 -1606 -15277
rect -1572 -15311 -1556 -15277
rect 7182 -15296 7198 -15262
rect 7232 -15296 7248 -15262
rect 7374 -15296 7390 -15262
rect 7424 -15296 7440 -15262
rect 7566 -15296 7582 -15262
rect 7616 -15296 7632 -15262
rect 7758 -15296 7774 -15262
rect 7808 -15296 7824 -15262
rect 8130 -15296 8146 -15262
rect 8180 -15296 8196 -15262
rect 8322 -15296 8338 -15262
rect 8372 -15296 8388 -15262
rect 8514 -15296 8530 -15262
rect 8564 -15296 8580 -15262
rect 8706 -15296 8722 -15262
rect 8756 -15296 8772 -15262
rect 9066 -15296 9082 -15262
rect 9116 -15296 9132 -15262
rect 9258 -15296 9274 -15262
rect 9308 -15296 9324 -15262
rect 9450 -15296 9466 -15262
rect 9500 -15296 9516 -15262
rect 9642 -15296 9658 -15262
rect 9692 -15296 9708 -15262
rect 9997 -15296 10013 -15262
rect 10047 -15296 10063 -15262
rect 10189 -15296 10205 -15262
rect 10239 -15296 10255 -15262
rect 10381 -15296 10397 -15262
rect 10431 -15296 10447 -15262
rect 10573 -15296 10589 -15262
rect 10623 -15296 10639 -15262
rect 10924 -15296 10940 -15262
rect 10974 -15296 10990 -15262
rect 11116 -15296 11132 -15262
rect 11166 -15296 11182 -15262
rect 11308 -15296 11324 -15262
rect 11358 -15296 11374 -15262
rect 11500 -15296 11516 -15262
rect 11550 -15296 11566 -15262
rect -2069 -15327 -1556 -15311
rect -11280 -15379 -11264 -15345
rect -11158 -15379 -11142 -15345
rect -11092 -15386 -11001 -15345
rect -8167 -15358 -8133 -15342
rect -8239 -15406 -8205 -15390
rect -12320 -15467 -12304 -15433
rect -11778 -15467 -11264 -15433
rect -11158 -15467 -11142 -15433
rect -17769 -15479 -17665 -15471
rect -24562 -15538 -24515 -15522
rect -24453 -15538 -24443 -15504
rect -24247 -15538 -24231 -15504
rect -17840 -15505 -17665 -15479
rect -17433 -15505 -17417 -15471
rect -17840 -15507 -17750 -15505
rect -8239 -15513 -8205 -15497
rect -8167 -15564 -8133 -15554
rect -8071 -15354 -8037 -15336
rect -8071 -15564 -8037 -15548
rect -7975 -15358 -7941 -15342
rect -7975 -15564 -7941 -15554
rect -7879 -15354 -7845 -15336
rect -7879 -15564 -7845 -15548
rect -7717 -15372 -7683 -15356
rect -7717 -15564 -7683 -15548
rect -7629 -15372 -7595 -15356
rect -4785 -15381 -4272 -15365
rect -7527 -15397 -7493 -15381
rect -4785 -15415 -4768 -15381
rect -4542 -15415 -4322 -15381
rect -4288 -15415 -4272 -15381
rect -4816 -15468 -4782 -15458
rect -7527 -15545 -7493 -15529
rect -4888 -15525 -4854 -15509
rect -7629 -15564 -7595 -15548
rect -11573 -15658 -11567 -15604
rect -11493 -15658 -11487 -15604
rect -8136 -15641 -8119 -15607
rect -7893 -15641 -7673 -15607
rect -7639 -15641 -7623 -15607
rect -4888 -15632 -4854 -15616
rect -8136 -15657 -7623 -15641
rect -4816 -15680 -4782 -15664
rect -4720 -15474 -4686 -15458
rect -4720 -15686 -4686 -15668
rect -4624 -15468 -4590 -15458
rect -4624 -15680 -4590 -15664
rect -4528 -15474 -4494 -15458
rect -4366 -15474 -4332 -15458
rect -4366 -15666 -4332 -15650
rect -4278 -15474 -4244 -15458
rect -2100 -15468 -2066 -15452
rect -4176 -15493 -4142 -15477
rect -2172 -15516 -2138 -15500
rect -2172 -15623 -2138 -15607
rect -4176 -15641 -4142 -15625
rect -4278 -15666 -4244 -15650
rect -4528 -15686 -4494 -15668
rect -2100 -15674 -2066 -15664
rect -2004 -15464 -1970 -15446
rect -2004 -15674 -1970 -15658
rect -1908 -15468 -1874 -15452
rect -1908 -15674 -1874 -15664
rect -1812 -15464 -1778 -15446
rect -1812 -15674 -1778 -15658
rect -1650 -15482 -1616 -15466
rect -1650 -15674 -1616 -15658
rect -1562 -15482 -1528 -15466
rect -1460 -15507 -1426 -15491
rect -1460 -15655 -1426 -15639
rect 7298 -15618 7403 -15615
rect 8246 -15618 8351 -15615
rect 9182 -15618 9287 -15615
rect 10113 -15618 10218 -15615
rect 11040 -15618 11145 -15615
rect 7298 -15634 7406 -15618
rect 7298 -15646 7372 -15634
rect -1562 -15674 -1528 -15658
rect -4785 -15760 -4272 -15744
rect -4785 -15794 -4768 -15760
rect -4542 -15794 -4322 -15760
rect -4288 -15794 -4272 -15760
rect -2069 -15751 -2052 -15717
rect -1826 -15751 -1606 -15717
rect -1572 -15751 -1556 -15717
rect -2069 -15767 -1556 -15751
rect -8166 -15858 -8132 -15842
rect -8238 -15906 -8204 -15890
rect -17681 -15945 -17665 -15911
rect -17433 -15945 -17417 -15911
rect -17681 -16041 -17665 -16007
rect -17433 -16041 -17417 -16007
rect -8238 -16013 -8204 -15997
rect -8166 -16064 -8132 -16054
rect -8070 -15854 -8036 -15836
rect -8070 -16064 -8036 -16048
rect -7974 -15858 -7940 -15842
rect -7974 -16064 -7940 -16054
rect -7878 -15854 -7844 -15836
rect -4816 -15847 -4782 -15837
rect -7878 -16064 -7844 -16048
rect -7716 -15872 -7682 -15856
rect -7716 -16064 -7682 -16048
rect -7628 -15872 -7594 -15856
rect -7526 -15897 -7492 -15881
rect -4888 -15904 -4854 -15888
rect -4888 -16011 -4854 -15995
rect -7526 -16045 -7492 -16029
rect -7628 -16064 -7594 -16048
rect -4816 -16059 -4782 -16043
rect -4720 -15853 -4686 -15837
rect -4720 -16065 -4686 -16047
rect -4624 -15847 -4590 -15837
rect -4624 -16059 -4590 -16043
rect -4528 -15853 -4494 -15837
rect -4366 -15853 -4332 -15837
rect -4366 -16045 -4332 -16029
rect -4278 -15853 -4244 -15837
rect -2100 -15847 -2066 -15831
rect -4176 -15872 -4142 -15856
rect -2172 -15895 -2138 -15879
rect -2172 -16002 -2138 -15986
rect -4176 -16020 -4142 -16004
rect -4278 -16045 -4244 -16029
rect -4528 -16065 -4494 -16047
rect -2100 -16053 -2066 -16043
rect -2004 -15843 -1970 -15825
rect -2004 -16053 -1970 -16037
rect -1908 -15847 -1874 -15831
rect -1908 -16053 -1874 -16043
rect -1812 -15843 -1778 -15825
rect -1812 -16053 -1778 -16037
rect -1650 -15861 -1616 -15845
rect -1650 -16053 -1616 -16037
rect -1562 -15861 -1528 -15845
rect -1460 -15886 -1426 -15870
rect -1460 -16034 -1426 -16018
rect -1562 -16053 -1528 -16037
rect -24092 -16113 -24058 -16097
rect -24561 -16138 -24514 -16114
rect -24452 -16147 -24442 -16113
rect -24246 -16147 -24230 -16113
rect -24452 -16243 -24436 -16209
rect -24240 -16243 -24230 -16209
rect -24452 -16339 -24442 -16305
rect -24246 -16339 -24230 -16305
rect -24187 -16334 -24147 -16318
rect -24152 -16368 -24147 -16334
rect -24187 -16385 -24147 -16368
rect -24452 -16435 -24436 -16401
rect -24240 -16435 -24230 -16401
rect -24452 -16531 -24442 -16497
rect -24246 -16531 -24230 -16497
rect -24181 -16539 -24147 -16385
rect -24092 -16505 -24058 -16489
rect -23900 -16113 -23866 -16097
rect -23900 -16505 -23866 -16489
rect -23828 -16139 -23794 -16101
rect -17681 -16137 -17665 -16103
rect -17433 -16137 -17417 -16103
rect -8135 -16141 -8118 -16107
rect -7892 -16141 -7672 -16107
rect -7638 -16141 -7622 -16107
rect -8135 -16157 -7622 -16141
rect -2069 -16130 -2052 -16096
rect -1826 -16130 -1606 -16096
rect -1572 -16130 -1556 -16096
rect -2069 -16146 -1556 -16130
rect -17681 -16233 -17665 -16199
rect -17433 -16233 -17417 -16199
rect -4785 -16200 -4272 -16184
rect -4785 -16234 -4768 -16200
rect -4542 -16234 -4322 -16200
rect -4288 -16234 -4272 -16200
rect -16928 -16295 -16844 -16283
rect -17681 -16329 -17665 -16295
rect -17433 -16329 -17417 -16295
rect -17266 -16343 -17232 -16327
rect -17192 -16329 -17176 -16295
rect -17000 -16308 -16844 -16295
rect -17000 -16329 -16917 -16308
rect -17681 -16425 -17665 -16391
rect -17433 -16425 -17417 -16391
rect -17266 -16393 -17232 -16377
rect -17192 -16425 -17176 -16391
rect -17000 -16425 -16984 -16391
rect -23828 -16501 -23794 -16474
rect -17371 -16486 -17337 -16470
rect -17840 -16521 -17665 -16487
rect -17433 -16521 -17417 -16487
rect -16928 -16487 -16917 -16329
rect -17840 -16522 -17750 -16521
rect -24181 -16573 -24063 -16539
rect -24028 -16573 -24012 -16539
rect -23946 -16573 -23930 -16539
rect -23895 -16573 -23879 -16539
rect -24452 -16627 -24436 -16593
rect -24240 -16627 -24230 -16593
rect -24187 -16623 -24152 -16607
rect -23946 -16631 -23879 -16573
rect -24152 -16657 -23879 -16631
rect -24187 -16674 -23879 -16657
rect -24561 -16723 -24514 -16707
rect -24452 -16723 -24442 -16689
rect -24246 -16723 -24230 -16689
rect -17840 -16879 -17820 -16522
rect -17769 -16679 -17750 -16522
rect -17371 -16536 -17337 -16520
rect -17192 -16521 -17176 -16487
rect -17000 -16507 -16917 -16487
rect -16856 -16507 -16844 -16308
rect -4816 -16287 -4782 -16277
rect -8167 -16338 -8133 -16322
rect -8239 -16386 -8205 -16370
rect -8239 -16493 -8205 -16477
rect -17000 -16521 -16844 -16507
rect -16928 -16533 -16844 -16521
rect -8167 -16544 -8133 -16534
rect -8071 -16334 -8037 -16316
rect -8071 -16544 -8037 -16528
rect -7975 -16338 -7941 -16322
rect -7975 -16544 -7941 -16534
rect -7879 -16334 -7845 -16316
rect -7879 -16544 -7845 -16528
rect -7717 -16352 -7683 -16336
rect -7717 -16544 -7683 -16528
rect -7629 -16352 -7595 -16336
rect -4888 -16344 -4854 -16328
rect -7527 -16377 -7493 -16361
rect -4888 -16451 -4854 -16435
rect -4816 -16499 -4782 -16483
rect -4720 -16293 -4686 -16277
rect -4720 -16505 -4686 -16487
rect -4624 -16287 -4590 -16277
rect -4624 -16499 -4590 -16483
rect -4528 -16293 -4494 -16277
rect -4366 -16293 -4332 -16277
rect -4366 -16485 -4332 -16469
rect -4278 -16293 -4244 -16277
rect -2100 -16287 -2066 -16271
rect -4176 -16312 -4142 -16296
rect -2172 -16335 -2138 -16319
rect -2172 -16442 -2138 -16426
rect -4176 -16460 -4142 -16444
rect -4278 -16485 -4244 -16469
rect -4528 -16505 -4494 -16487
rect -2100 -16493 -2066 -16483
rect -2004 -16283 -1970 -16265
rect -2004 -16493 -1970 -16477
rect -1908 -16287 -1874 -16271
rect -1908 -16493 -1874 -16483
rect -1812 -16283 -1778 -16265
rect -1812 -16493 -1778 -16477
rect -1650 -16301 -1616 -16285
rect -1650 -16493 -1616 -16477
rect -1562 -16301 -1528 -16285
rect -1460 -16326 -1426 -16310
rect 7333 -16397 7372 -15646
rect 7298 -16410 7372 -16397
rect 7298 -16426 7406 -16410
rect 7756 -15634 7790 -15618
rect 7756 -16426 7790 -16410
rect 8246 -15634 8354 -15618
rect 8246 -15646 8320 -15634
rect 8281 -16397 8320 -15646
rect 8246 -16410 8320 -16397
rect 8246 -16426 8354 -16410
rect 8704 -15634 8738 -15618
rect 8704 -16426 8738 -16410
rect 9182 -15634 9290 -15618
rect 9182 -15646 9256 -15634
rect 9217 -16397 9256 -15646
rect 9182 -16410 9256 -16397
rect 9182 -16426 9290 -16410
rect 9640 -15634 9674 -15618
rect 9640 -16426 9674 -16410
rect 10113 -15634 10221 -15618
rect 10113 -15646 10187 -15634
rect 10148 -16397 10187 -15646
rect 10113 -16410 10187 -16397
rect 10113 -16426 10221 -16410
rect 10571 -15634 10605 -15618
rect 10571 -16426 10605 -16410
rect 11040 -15634 11148 -15618
rect 11040 -15646 11114 -15634
rect 11075 -16397 11114 -15646
rect 11040 -16410 11114 -16397
rect 11040 -16426 11148 -16410
rect 11498 -15634 11532 -15618
rect 11783 -15960 12203 -15940
rect 11783 -16011 11811 -15960
rect 12168 -16011 12203 -15960
rect 11783 -16030 12203 -16011
rect 11785 -16115 11819 -16030
rect 11785 -16363 11819 -16347
rect 11881 -16115 11915 -16099
rect 11881 -16363 11915 -16347
rect 11977 -16115 12011 -16030
rect 11977 -16363 12011 -16347
rect 12073 -16115 12107 -16099
rect 12073 -16363 12107 -16347
rect 12169 -16115 12203 -16030
rect 12169 -16363 12203 -16347
rect 12265 -16115 12299 -16099
rect 12265 -16363 12299 -16347
rect 12361 -16115 12395 -16099
rect 12361 -16363 12395 -16347
rect 12457 -16115 12491 -16099
rect 12457 -16363 12491 -16347
rect 12553 -16115 12587 -16099
rect 12553 -16363 12587 -16347
rect 12649 -16115 12683 -16099
rect 12649 -16363 12683 -16347
rect 12745 -16115 12779 -16099
rect 12970 -16181 12986 -16147
rect 13077 -16181 13093 -16147
rect 12745 -16363 12779 -16347
rect 12826 -16267 12876 -16250
rect 12919 -16253 12929 -16219
rect 13125 -16253 13141 -16219
rect 11498 -16426 11532 -16410
rect 12154 -16443 12170 -16409
rect 12204 -16443 12220 -16409
rect -1460 -16474 -1426 -16458
rect -1562 -16493 -1528 -16477
rect 12826 -16493 12842 -16267
rect 12919 -16349 12935 -16315
rect 13129 -16349 13147 -16315
rect 12919 -16445 12929 -16411
rect 13125 -16445 13141 -16411
rect -7527 -16525 -7493 -16509
rect -7629 -16544 -7595 -16528
rect -4785 -16579 -4272 -16563
rect -17681 -16617 -17665 -16583
rect -17433 -16617 -17417 -16583
rect -8136 -16621 -8119 -16587
rect -7893 -16621 -7673 -16587
rect -7639 -16621 -7623 -16587
rect -4785 -16613 -4768 -16579
rect -4542 -16613 -4322 -16579
rect -4288 -16613 -4272 -16579
rect -2069 -16570 -2052 -16536
rect -1826 -16570 -1606 -16536
rect -1572 -16570 -1556 -16536
rect -2069 -16586 -1556 -16570
rect 7298 -16562 7406 -16546
rect 7298 -16575 7372 -16562
rect -8136 -16637 -7623 -16621
rect -4816 -16666 -4782 -16656
rect -17769 -16713 -17665 -16679
rect -17433 -16713 -17417 -16679
rect -17769 -16871 -17750 -16713
rect -4888 -16723 -4854 -16707
rect -17681 -16809 -17665 -16775
rect -17433 -16809 -17417 -16775
rect -8167 -16838 -8133 -16822
rect -17769 -16879 -17665 -16871
rect -17840 -16905 -17665 -16879
rect -17433 -16905 -17417 -16871
rect -8239 -16886 -8205 -16870
rect -17840 -16907 -17750 -16905
rect -12318 -16955 -12302 -16921
rect -11776 -16955 -11262 -16921
rect -11156 -16955 -11140 -16921
rect -12499 -17039 -12373 -16997
rect -24087 -17326 -24053 -17310
rect -24556 -17351 -24509 -17327
rect -24447 -17360 -24437 -17326
rect -24241 -17360 -24225 -17326
rect -24447 -17456 -24431 -17422
rect -24235 -17456 -24225 -17422
rect -24447 -17552 -24437 -17518
rect -24241 -17552 -24225 -17518
rect -24182 -17547 -24142 -17531
rect -24147 -17581 -24142 -17547
rect -24182 -17598 -24142 -17581
rect -24447 -17648 -24431 -17614
rect -24235 -17648 -24225 -17614
rect -24447 -17744 -24437 -17710
rect -24241 -17744 -24225 -17710
rect -24176 -17752 -24142 -17598
rect -24087 -17718 -24053 -17702
rect -23895 -17326 -23861 -17310
rect -23895 -17718 -23861 -17702
rect -23823 -17352 -23789 -17314
rect -17681 -17345 -17665 -17311
rect -17433 -17345 -17417 -17311
rect -17681 -17441 -17665 -17407
rect -17433 -17441 -17417 -17407
rect -17681 -17537 -17665 -17503
rect -17433 -17537 -17417 -17503
rect -17681 -17633 -17665 -17599
rect -17433 -17633 -17417 -17599
rect -23823 -17714 -23789 -17687
rect -16928 -17695 -16844 -17683
rect -17681 -17729 -17665 -17695
rect -17433 -17729 -17417 -17695
rect -17266 -17743 -17232 -17727
rect -17192 -17729 -17176 -17695
rect -17000 -17708 -16844 -17695
rect -17000 -17729 -16917 -17708
rect -24176 -17786 -24058 -17752
rect -24023 -17786 -24007 -17752
rect -23941 -17786 -23925 -17752
rect -23890 -17786 -23874 -17752
rect -24447 -17840 -24431 -17806
rect -24235 -17840 -24225 -17806
rect -24182 -17836 -24147 -17820
rect -23941 -17844 -23874 -17786
rect -17681 -17825 -17665 -17791
rect -17433 -17825 -17417 -17791
rect -17266 -17793 -17232 -17777
rect -17192 -17825 -17176 -17791
rect -17000 -17825 -16984 -17791
rect -24147 -17870 -23874 -17844
rect -24182 -17887 -23874 -17870
rect -17371 -17886 -17337 -17870
rect -24556 -17936 -24509 -17920
rect -24447 -17936 -24437 -17902
rect -24241 -17936 -24225 -17902
rect -17840 -17921 -17665 -17887
rect -17433 -17921 -17417 -17887
rect -16928 -17887 -16917 -17729
rect -17840 -17922 -17750 -17921
rect -21606 -18046 -21572 -18030
rect -21678 -18094 -21644 -18078
rect -21678 -18201 -21644 -18185
rect -21606 -18252 -21572 -18242
rect -21510 -18042 -21476 -18024
rect -21510 -18252 -21476 -18236
rect -21414 -18046 -21380 -18030
rect -21414 -18252 -21380 -18242
rect -21318 -18042 -21284 -18024
rect -21318 -18252 -21284 -18236
rect -21156 -18060 -21122 -18044
rect -21156 -18252 -21122 -18236
rect -21068 -18060 -21034 -18044
rect -20966 -18085 -20932 -18069
rect -20966 -18233 -20932 -18217
rect -21068 -18252 -21034 -18236
rect -17840 -18279 -17820 -17922
rect -17769 -18079 -17750 -17922
rect -17371 -17936 -17337 -17920
rect -17192 -17921 -17176 -17887
rect -17000 -17907 -16917 -17887
rect -16856 -17907 -16844 -17708
rect -17000 -17921 -16844 -17907
rect -16928 -17933 -16844 -17921
rect -16015 -17917 -15981 -17901
rect -16087 -17965 -16053 -17949
rect -17681 -18017 -17665 -17983
rect -17433 -18017 -17417 -17983
rect -16087 -18072 -16053 -18056
rect -17769 -18113 -17665 -18079
rect -17433 -18113 -17417 -18079
rect -17769 -18271 -17750 -18113
rect -16015 -18123 -15981 -18113
rect -15919 -17913 -15885 -17895
rect -15919 -18123 -15885 -18107
rect -15823 -17917 -15789 -17901
rect -15823 -18123 -15789 -18113
rect -15727 -17913 -15693 -17895
rect -15727 -18123 -15693 -18107
rect -15565 -17931 -15531 -17915
rect -15565 -18123 -15531 -18107
rect -15477 -17931 -15443 -17915
rect -15375 -17956 -15341 -17940
rect -15375 -18104 -15341 -18088
rect -15477 -18123 -15443 -18107
rect -12499 -18161 -12471 -17039
rect -12399 -18161 -12373 -17039
rect -12318 -17043 -12302 -17009
rect -11776 -17043 -11760 -17009
rect -12318 -17139 -12302 -17105
rect -11776 -17139 -11760 -17105
rect -12318 -17235 -12302 -17201
rect -11776 -17235 -11760 -17201
rect -12318 -17331 -12302 -17297
rect -11776 -17331 -11760 -17297
rect -11718 -17346 -11641 -16955
rect -8239 -16993 -8205 -16977
rect -11433 -17010 -11337 -16995
rect -11433 -17075 -11411 -17010
rect -11356 -17075 -11337 -17010
rect -11278 -17043 -11262 -17009
rect -11156 -17043 -11140 -17009
rect -11090 -17038 -10999 -17000
rect -11600 -17177 -11494 -17159
rect -11600 -17257 -11582 -17177
rect -11514 -17257 -11494 -17177
rect -11600 -17274 -11494 -17257
rect -11718 -17366 -11501 -17346
rect -12318 -17427 -12302 -17393
rect -11776 -17427 -11760 -17393
rect -12318 -17523 -12302 -17489
rect -11776 -17523 -11760 -17489
rect -11718 -17496 -11700 -17366
rect -11655 -17377 -11501 -17366
rect -11655 -17491 -11583 -17377
rect -11530 -17491 -11501 -17377
rect -11655 -17496 -11501 -17491
rect -11718 -17523 -11501 -17496
rect -11433 -17569 -11337 -17075
rect -11278 -17139 -11277 -17105
rect -11156 -17139 -11140 -17105
rect -11278 -17235 -11262 -17201
rect -11142 -17235 -11140 -17201
rect -11278 -17331 -11277 -17297
rect -11156 -17331 -11140 -17297
rect -11278 -17427 -11262 -17393
rect -11142 -17427 -11140 -17393
rect -11278 -17523 -11277 -17489
rect -11156 -17523 -11140 -17489
rect -11733 -17585 -11303 -17569
rect -12318 -17619 -12302 -17585
rect -11776 -17619 -11262 -17585
rect -11142 -17619 -11140 -17585
rect -11733 -17635 -11303 -17619
rect -12318 -17715 -12302 -17681
rect -11776 -17715 -11760 -17681
rect -11715 -17689 -11314 -17681
rect -11715 -17697 -11376 -17689
rect -12318 -17811 -12302 -17777
rect -11776 -17811 -11760 -17777
rect -11715 -17827 -11705 -17697
rect -11660 -17819 -11376 -17697
rect -11331 -17819 -11314 -17689
rect -11278 -17715 -11276 -17681
rect -11156 -17715 -11140 -17681
rect -11278 -17811 -11262 -17777
rect -11142 -17811 -11140 -17777
rect -11660 -17827 -11314 -17819
rect -11715 -17846 -11314 -17827
rect -12318 -17907 -12302 -17873
rect -11776 -17907 -11760 -17873
rect -12318 -18003 -12302 -17969
rect -11776 -18003 -11760 -17969
rect -12318 -18099 -12302 -18065
rect -11776 -18099 -11760 -18065
rect -17681 -18209 -17665 -18175
rect -17433 -18209 -17417 -18175
rect -15984 -18200 -15967 -18166
rect -15741 -18200 -15521 -18166
rect -15487 -18200 -15471 -18166
rect -15984 -18216 -15471 -18200
rect -12499 -18207 -12373 -18161
rect -12318 -18195 -12302 -18161
rect -11776 -18195 -11760 -18161
rect -11715 -18249 -11646 -17846
rect -11278 -17907 -11277 -17873
rect -11156 -17907 -11140 -17873
rect -11602 -17964 -11312 -17926
rect -11602 -18097 -11575 -17964
rect -11522 -17972 -11312 -17964
rect -11522 -18097 -11384 -17972
rect -11602 -18102 -11384 -18097
rect -11339 -18102 -11312 -17972
rect -11278 -18003 -11262 -17969
rect -11142 -18003 -11140 -17969
rect -11278 -18099 -11277 -18065
rect -11156 -18099 -11140 -18065
rect -11602 -18147 -11312 -18102
rect -11090 -18161 -11068 -17038
rect -11022 -18161 -10999 -17038
rect -8167 -17044 -8133 -17034
rect -8071 -16834 -8037 -16816
rect -8071 -17044 -8037 -17028
rect -7975 -16838 -7941 -16822
rect -7975 -17044 -7941 -17034
rect -7879 -16834 -7845 -16816
rect -4888 -16830 -4854 -16814
rect -7879 -17044 -7845 -17028
rect -7717 -16852 -7683 -16836
rect -7717 -17044 -7683 -17028
rect -7629 -16852 -7595 -16836
rect -7527 -16877 -7493 -16861
rect -4816 -16878 -4782 -16862
rect -4720 -16672 -4686 -16656
rect -4720 -16884 -4686 -16866
rect -4624 -16666 -4590 -16656
rect -4624 -16878 -4590 -16862
rect -4528 -16672 -4494 -16656
rect -4366 -16672 -4332 -16656
rect -4366 -16864 -4332 -16848
rect -4278 -16672 -4244 -16656
rect -2100 -16666 -2066 -16650
rect -4176 -16691 -4142 -16675
rect -2172 -16714 -2138 -16698
rect -2172 -16821 -2138 -16805
rect -4176 -16839 -4142 -16823
rect -4278 -16864 -4244 -16848
rect -4528 -16884 -4494 -16866
rect -2100 -16872 -2066 -16862
rect -2004 -16662 -1970 -16644
rect -2004 -16872 -1970 -16856
rect -1908 -16666 -1874 -16650
rect -1908 -16872 -1874 -16862
rect -1812 -16662 -1778 -16644
rect -1812 -16872 -1778 -16856
rect -1650 -16680 -1616 -16664
rect -1650 -16872 -1616 -16856
rect -1562 -16680 -1528 -16664
rect -1460 -16705 -1426 -16689
rect -1460 -16853 -1426 -16837
rect -1562 -16872 -1528 -16856
rect -2069 -16949 -2052 -16915
rect -1826 -16949 -1606 -16915
rect -1572 -16949 -1556 -16915
rect -2069 -16965 -1556 -16949
rect -7527 -17025 -7493 -17009
rect -4785 -17019 -4272 -17003
rect -7629 -17044 -7595 -17028
rect -4785 -17053 -4768 -17019
rect -4542 -17053 -4322 -17019
rect -4288 -17053 -4272 -17019
rect -8136 -17121 -8119 -17087
rect -7893 -17121 -7673 -17087
rect -7639 -17121 -7623 -17087
rect -8136 -17137 -7623 -17121
rect -4816 -17106 -4782 -17096
rect -4888 -17163 -4854 -17147
rect -4888 -17270 -4854 -17254
rect -8167 -17318 -8133 -17302
rect -8239 -17366 -8205 -17350
rect -8239 -17473 -8205 -17457
rect -8167 -17524 -8133 -17514
rect -8071 -17314 -8037 -17296
rect -8071 -17524 -8037 -17508
rect -7975 -17318 -7941 -17302
rect -7975 -17524 -7941 -17514
rect -7879 -17314 -7845 -17296
rect -7879 -17524 -7845 -17508
rect -7717 -17332 -7683 -17316
rect -7717 -17524 -7683 -17508
rect -7629 -17332 -7595 -17316
rect -4816 -17318 -4782 -17302
rect -4720 -17112 -4686 -17096
rect -4720 -17324 -4686 -17306
rect -4624 -17106 -4590 -17096
rect -4624 -17318 -4590 -17302
rect -4528 -17112 -4494 -17096
rect -4366 -17112 -4332 -17096
rect -4366 -17304 -4332 -17288
rect -4278 -17112 -4244 -17096
rect -2100 -17106 -2066 -17090
rect -4176 -17131 -4142 -17115
rect -2172 -17154 -2138 -17138
rect -2172 -17261 -2138 -17245
rect -4176 -17279 -4142 -17263
rect -4278 -17304 -4244 -17288
rect -4528 -17324 -4494 -17306
rect -2100 -17312 -2066 -17302
rect -2004 -17102 -1970 -17084
rect -2004 -17312 -1970 -17296
rect -1908 -17106 -1874 -17090
rect -1908 -17312 -1874 -17302
rect -1812 -17102 -1778 -17084
rect -1812 -17312 -1778 -17296
rect -1650 -17120 -1616 -17104
rect -1650 -17312 -1616 -17296
rect -1562 -17120 -1528 -17104
rect -1460 -17145 -1426 -17129
rect -1460 -17293 -1426 -17277
rect -1562 -17312 -1528 -17296
rect 7333 -17326 7372 -16575
rect 7298 -17338 7372 -17326
rect -7527 -17357 -7493 -17341
rect 7298 -17354 7406 -17338
rect 7756 -16562 7790 -16546
rect 7756 -17354 7790 -17338
rect 8246 -16562 8354 -16546
rect 8246 -16575 8320 -16562
rect 8281 -17326 8320 -16575
rect 8246 -17338 8320 -17326
rect 8246 -17354 8354 -17338
rect 8704 -16562 8738 -16546
rect 8704 -17354 8738 -17338
rect 9182 -16562 9290 -16546
rect 9182 -16575 9256 -16562
rect 9217 -17326 9256 -16575
rect 9182 -17338 9256 -17326
rect 9182 -17354 9290 -17338
rect 9640 -16562 9674 -16546
rect 9640 -17354 9674 -17338
rect 10113 -16561 10221 -16545
rect 10113 -16574 10187 -16561
rect 10148 -17325 10187 -16574
rect 10113 -17337 10187 -17325
rect 10113 -17353 10221 -17337
rect 10571 -16561 10605 -16545
rect 10571 -17353 10605 -17337
rect 11040 -16562 11148 -16546
rect 11040 -16575 11114 -16562
rect 11075 -17326 11114 -16575
rect 11040 -17338 11114 -17326
rect -4785 -17398 -4272 -17382
rect -4785 -17432 -4768 -17398
rect -4542 -17432 -4322 -17398
rect -4288 -17432 -4272 -17398
rect -2069 -17389 -2052 -17355
rect -1826 -17389 -1606 -17355
rect -1572 -17389 -1556 -17355
rect 7298 -17357 7403 -17354
rect 8246 -17357 8351 -17354
rect 9182 -17357 9287 -17354
rect 10113 -17356 10218 -17353
rect 11040 -17354 11148 -17338
rect 11498 -16562 11532 -16546
rect 12297 -16548 12313 -16514
rect 12347 -16548 12363 -16514
rect 12169 -16604 12203 -16588
rect 12169 -16852 12203 -16780
rect 12265 -16604 12299 -16588
rect 12265 -16796 12299 -16780
rect 12361 -16604 12395 -16588
rect 12826 -16713 12876 -16493
rect 12919 -16541 12935 -16507
rect 13129 -16541 13147 -16507
rect 12919 -16703 12935 -16669
rect 13111 -16703 13127 -16669
rect 12826 -16747 12842 -16713
rect 12826 -16763 12876 -16747
rect 12361 -16852 12395 -16780
rect 12919 -16791 12935 -16757
rect 13111 -16791 13127 -16757
rect 16159 -16814 16577 -16766
rect 12157 -16863 12407 -16852
rect 12157 -16924 12183 -16863
rect 12382 -16924 12407 -16863
rect 12938 -16893 12954 -16859
rect 13086 -16893 13102 -16859
rect 12157 -16936 12407 -16924
rect 16159 -16927 16211 -16814
rect 16541 -16927 16577 -16814
rect 16159 -16995 16577 -16927
rect 16159 -17061 16193 -16995
rect 16159 -17253 16193 -17237
rect 16255 -17061 16289 -17045
rect 16255 -17253 16289 -17237
rect 16351 -17061 16385 -16995
rect 16351 -17253 16385 -17237
rect 16447 -17061 16481 -17045
rect 16447 -17253 16481 -17237
rect 16543 -17061 16577 -16995
rect 16543 -17253 16577 -17237
rect 16653 -17338 16669 -17304
rect 16703 -17338 16719 -17304
rect 11498 -17354 11532 -17338
rect 11040 -17357 11145 -17354
rect -2069 -17405 -1556 -17389
rect -7527 -17505 -7493 -17489
rect -4816 -17485 -4782 -17475
rect -7629 -17524 -7595 -17508
rect -4888 -17542 -4854 -17526
rect -8136 -17601 -8119 -17567
rect -7893 -17601 -7673 -17567
rect -7639 -17601 -7623 -17567
rect -8136 -17617 -7623 -17601
rect -4888 -17649 -4854 -17633
rect -4816 -17697 -4782 -17681
rect -4720 -17491 -4686 -17475
rect -4720 -17703 -4686 -17685
rect -4624 -17485 -4590 -17475
rect -4624 -17697 -4590 -17681
rect -4528 -17491 -4494 -17475
rect -4366 -17491 -4332 -17475
rect -4366 -17683 -4332 -17667
rect -4278 -17491 -4244 -17475
rect -2100 -17485 -2066 -17469
rect -4176 -17510 -4142 -17494
rect -2172 -17533 -2138 -17517
rect -2172 -17640 -2138 -17624
rect -4176 -17658 -4142 -17642
rect -4278 -17683 -4244 -17667
rect -4528 -17703 -4494 -17685
rect -2100 -17691 -2066 -17681
rect -2004 -17481 -1970 -17463
rect -2004 -17691 -1970 -17675
rect -1908 -17485 -1874 -17469
rect -1908 -17691 -1874 -17681
rect -1812 -17481 -1778 -17463
rect -1812 -17691 -1778 -17675
rect -1650 -17499 -1616 -17483
rect -1650 -17691 -1616 -17675
rect -1562 -17499 -1528 -17483
rect -1460 -17524 -1426 -17508
rect 15981 -17620 15997 -17586
rect 16031 -17620 16047 -17586
rect 16269 -17620 16285 -17586
rect 16319 -17620 16335 -17586
rect 16401 -17620 16417 -17586
rect 16451 -17620 16467 -17586
rect -1460 -17672 -1426 -17656
rect -1562 -17691 -1528 -17675
rect 7182 -17710 7198 -17676
rect 7232 -17710 7248 -17676
rect 7374 -17710 7390 -17676
rect 7424 -17710 7440 -17676
rect 7566 -17710 7582 -17676
rect 7616 -17710 7632 -17676
rect 7758 -17710 7774 -17676
rect 7808 -17710 7824 -17676
rect 8130 -17710 8146 -17676
rect 8180 -17710 8196 -17676
rect 8322 -17710 8338 -17676
rect 8372 -17710 8388 -17676
rect 8514 -17710 8530 -17676
rect 8564 -17710 8580 -17676
rect 8706 -17710 8722 -17676
rect 8756 -17710 8772 -17676
rect 9066 -17710 9082 -17676
rect 9116 -17710 9132 -17676
rect 9258 -17710 9274 -17676
rect 9308 -17710 9324 -17676
rect 9450 -17710 9466 -17676
rect 9500 -17710 9516 -17676
rect 9642 -17710 9658 -17676
rect 9692 -17710 9708 -17676
rect 9997 -17709 10013 -17675
rect 10047 -17709 10063 -17675
rect 10189 -17709 10205 -17675
rect 10239 -17709 10255 -17675
rect 10381 -17709 10397 -17675
rect 10431 -17709 10447 -17675
rect 10573 -17709 10589 -17675
rect 10623 -17709 10639 -17675
rect 10924 -17710 10940 -17676
rect 10974 -17710 10990 -17676
rect 11116 -17710 11132 -17676
rect 11166 -17710 11182 -17676
rect 11308 -17710 11324 -17676
rect 11358 -17710 11374 -17676
rect 11500 -17710 11516 -17676
rect 11550 -17710 11566 -17676
rect 15703 -17679 15737 -17663
rect -8167 -17778 -8133 -17762
rect -8239 -17826 -8205 -17810
rect -8239 -17933 -8205 -17917
rect -8167 -17984 -8133 -17974
rect -8071 -17774 -8037 -17756
rect -8071 -17984 -8037 -17968
rect -7975 -17778 -7941 -17762
rect -7975 -17984 -7941 -17974
rect -7879 -17774 -7845 -17756
rect -2069 -17768 -2052 -17734
rect -1826 -17768 -1606 -17734
rect -1572 -17768 -1556 -17734
rect -7879 -17984 -7845 -17968
rect -7717 -17792 -7683 -17776
rect -7717 -17984 -7683 -17968
rect -7629 -17792 -7595 -17776
rect -2069 -17784 -1556 -17768
rect 7150 -17769 7184 -17753
rect 7246 -17764 7280 -17753
rect -7527 -17817 -7493 -17801
rect -4785 -17838 -4272 -17822
rect -4785 -17872 -4768 -17838
rect -4542 -17872 -4322 -17838
rect -4288 -17872 -4272 -17838
rect -7527 -17965 -7493 -17949
rect -4816 -17925 -4782 -17915
rect -7629 -17984 -7595 -17968
rect -4888 -17982 -4854 -17966
rect -8136 -18061 -8119 -18027
rect -7893 -18061 -7673 -18027
rect -7639 -18061 -7623 -18027
rect -8136 -18077 -7623 -18061
rect -4888 -18089 -4854 -18073
rect -4816 -18137 -4782 -18121
rect -4720 -17931 -4686 -17915
rect -4720 -18143 -4686 -18125
rect -4624 -17925 -4590 -17915
rect -4624 -18137 -4590 -18121
rect -4528 -17931 -4494 -17915
rect -4366 -17931 -4332 -17915
rect -4366 -18123 -4332 -18107
rect -4278 -17931 -4244 -17915
rect -2100 -17925 -2066 -17909
rect -4176 -17950 -4142 -17934
rect -2172 -17973 -2138 -17957
rect -2172 -18080 -2138 -18064
rect -4176 -18098 -4142 -18082
rect -4278 -18123 -4244 -18107
rect -4528 -18143 -4494 -18125
rect -2100 -18131 -2066 -18121
rect -2004 -17921 -1970 -17903
rect -2004 -18131 -1970 -18115
rect -1908 -17925 -1874 -17909
rect -1908 -18131 -1874 -18121
rect -1812 -17921 -1778 -17903
rect -1812 -18131 -1778 -18115
rect -1650 -17939 -1616 -17923
rect -1650 -18131 -1616 -18115
rect -1562 -17939 -1528 -17923
rect -1460 -17964 -1426 -17948
rect 7150 -18083 7184 -18067
rect 7246 -18083 7280 -18067
rect 7342 -17769 7376 -17753
rect 7342 -18083 7376 -18067
rect 7438 -17764 7472 -17753
rect 7534 -17769 7568 -17753
rect 7438 -18083 7472 -18067
rect 7534 -18083 7568 -18067
rect 7630 -17764 7664 -17753
rect 7726 -17769 7760 -17753
rect 7630 -18083 7664 -18067
rect 7726 -18083 7760 -18067
rect 7822 -17764 7856 -17753
rect 7918 -17769 7952 -17753
rect 7822 -18083 7856 -18067
rect 7918 -18083 7952 -18067
rect 8098 -17769 8132 -17753
rect 8194 -17764 8228 -17753
rect 8098 -18083 8132 -18067
rect 8194 -18083 8228 -18067
rect 8290 -17769 8324 -17753
rect 8290 -18083 8324 -18067
rect 8386 -17764 8420 -17753
rect 8482 -17769 8516 -17753
rect 8386 -18083 8420 -18067
rect 8482 -18083 8516 -18067
rect 8578 -17764 8612 -17753
rect 8674 -17769 8708 -17753
rect 8578 -18083 8612 -18067
rect 8674 -18083 8708 -18067
rect 8770 -17764 8804 -17753
rect 8866 -17769 8900 -17753
rect 8770 -18083 8804 -18067
rect 8866 -18083 8900 -18067
rect 9034 -17769 9068 -17753
rect 9130 -17764 9164 -17753
rect 9034 -18083 9068 -18067
rect 9130 -18083 9164 -18067
rect 9226 -17769 9260 -17753
rect 9226 -18083 9260 -18067
rect 9322 -17764 9356 -17753
rect 9418 -17769 9452 -17753
rect 9322 -18083 9356 -18067
rect 9418 -18083 9452 -18067
rect 9514 -17764 9548 -17753
rect 9610 -17769 9644 -17753
rect 9514 -18083 9548 -18067
rect 9610 -18083 9644 -18067
rect 9706 -17764 9740 -17753
rect 9802 -17769 9836 -17753
rect 9706 -18083 9740 -18067
rect 9802 -18083 9836 -18067
rect 9965 -17768 9999 -17752
rect 10061 -17763 10095 -17752
rect 9965 -18082 9999 -18066
rect 10061 -18082 10095 -18066
rect 10157 -17768 10191 -17752
rect 10157 -18082 10191 -18066
rect 10253 -17763 10287 -17752
rect 10349 -17768 10383 -17752
rect 10253 -18082 10287 -18066
rect 10349 -18082 10383 -18066
rect 10445 -17763 10479 -17752
rect 10541 -17768 10575 -17752
rect 10445 -18082 10479 -18066
rect 10541 -18082 10575 -18066
rect 10637 -17763 10671 -17752
rect 10733 -17768 10767 -17752
rect 10637 -18082 10671 -18066
rect 10733 -18082 10767 -18066
rect 10892 -17769 10926 -17753
rect 10988 -17764 11022 -17753
rect 10892 -18083 10926 -18067
rect 10988 -18083 11022 -18067
rect 11084 -17769 11118 -17753
rect 11084 -18083 11118 -18067
rect 11180 -17764 11214 -17753
rect 11276 -17769 11310 -17753
rect 11180 -18083 11214 -18067
rect 11276 -18083 11310 -18067
rect 11372 -17764 11406 -17753
rect 11468 -17769 11502 -17753
rect 11372 -18083 11406 -18067
rect 11468 -18083 11502 -18067
rect 11564 -17764 11598 -17753
rect 11660 -17769 11694 -17753
rect 11564 -18083 11598 -18067
rect 15703 -18049 15737 -18033
rect 15775 -17679 15809 -17663
rect 11660 -18083 11694 -18067
rect -1460 -18112 -1426 -18096
rect -1562 -18131 -1528 -18115
rect -11278 -18195 -11262 -18161
rect -11156 -18195 -11140 -18161
rect -11090 -18202 -10999 -18161
rect 7373 -18171 7389 -18136
rect 7677 -18171 7703 -18136
rect 8321 -18171 8337 -18136
rect 8625 -18171 8651 -18136
rect 9257 -18171 9273 -18136
rect 9561 -18171 9587 -18136
rect 10188 -18170 10204 -18135
rect 10492 -18170 10518 -18135
rect 11115 -18171 11131 -18136
rect 11419 -18171 11445 -18136
rect -8181 -18238 -8147 -18222
rect -17769 -18279 -17665 -18271
rect -21575 -18329 -21558 -18295
rect -21332 -18329 -21112 -18295
rect -21078 -18329 -21062 -18295
rect -17840 -18305 -17665 -18279
rect -17433 -18305 -17417 -18271
rect -12318 -18283 -12302 -18249
rect -11776 -18283 -11262 -18249
rect -11156 -18283 -11140 -18249
rect -8253 -18286 -8219 -18270
rect -17840 -18307 -17750 -18305
rect -21575 -18345 -21062 -18329
rect -8253 -18393 -8219 -18377
rect -16014 -18417 -15980 -18401
rect -24072 -18445 -24038 -18429
rect -24541 -18470 -24494 -18446
rect -24432 -18479 -24422 -18445
rect -24226 -18479 -24210 -18445
rect -24432 -18575 -24416 -18541
rect -24220 -18575 -24210 -18541
rect -24432 -18671 -24422 -18637
rect -24226 -18671 -24210 -18637
rect -24167 -18666 -24127 -18650
rect -24132 -18700 -24127 -18666
rect -24167 -18717 -24127 -18700
rect -24432 -18767 -24416 -18733
rect -24220 -18767 -24210 -18733
rect -24432 -18863 -24422 -18829
rect -24226 -18863 -24210 -18829
rect -24161 -18871 -24127 -18717
rect -24072 -18837 -24038 -18821
rect -23880 -18445 -23846 -18429
rect -23880 -18837 -23846 -18821
rect -23808 -18471 -23774 -18433
rect -16086 -18465 -16052 -18449
rect -21605 -18546 -21571 -18530
rect -21677 -18594 -21643 -18578
rect -21677 -18701 -21643 -18685
rect -21605 -18752 -21571 -18742
rect -21509 -18542 -21475 -18524
rect -21509 -18752 -21475 -18736
rect -21413 -18546 -21379 -18530
rect -21413 -18752 -21379 -18742
rect -21317 -18542 -21283 -18524
rect -21317 -18752 -21283 -18736
rect -21155 -18560 -21121 -18544
rect -21155 -18752 -21121 -18736
rect -21067 -18560 -21033 -18544
rect -20965 -18585 -20931 -18569
rect -16086 -18572 -16052 -18556
rect -16014 -18623 -15980 -18613
rect -15918 -18413 -15884 -18395
rect -15918 -18623 -15884 -18607
rect -15822 -18417 -15788 -18401
rect -15822 -18623 -15788 -18613
rect -15726 -18413 -15692 -18395
rect -15726 -18623 -15692 -18607
rect -15564 -18431 -15530 -18415
rect -15564 -18623 -15530 -18607
rect -15476 -18431 -15442 -18415
rect -15374 -18456 -15340 -18440
rect -11571 -18467 -11565 -18413
rect -11491 -18467 -11485 -18413
rect -8181 -18444 -8147 -18434
rect -8085 -18234 -8051 -18216
rect -8085 -18444 -8051 -18428
rect -7989 -18238 -7955 -18222
rect -7989 -18444 -7955 -18434
rect -7893 -18234 -7859 -18216
rect -4785 -18217 -4272 -18201
rect -7893 -18444 -7859 -18428
rect -7731 -18252 -7697 -18236
rect -7731 -18444 -7697 -18428
rect -7643 -18252 -7609 -18236
rect -4785 -18251 -4768 -18217
rect -4542 -18251 -4322 -18217
rect -4288 -18251 -4272 -18217
rect -2069 -18208 -2052 -18174
rect -1826 -18208 -1606 -18174
rect -1572 -18208 -1556 -18174
rect -2069 -18224 -1556 -18208
rect -7541 -18277 -7507 -18261
rect -4816 -18304 -4782 -18294
rect -7541 -18425 -7507 -18409
rect -4888 -18361 -4854 -18345
rect -7643 -18444 -7609 -18428
rect -4888 -18468 -4854 -18452
rect -8150 -18521 -8133 -18487
rect -7907 -18521 -7687 -18487
rect -7653 -18521 -7637 -18487
rect -4816 -18516 -4782 -18500
rect -4720 -18310 -4686 -18294
rect -8150 -18537 -7637 -18521
rect -4720 -18522 -4686 -18504
rect -4624 -18304 -4590 -18294
rect -4624 -18516 -4590 -18500
rect -4528 -18310 -4494 -18294
rect -4366 -18310 -4332 -18294
rect -4366 -18502 -4332 -18486
rect -4278 -18310 -4244 -18294
rect -2100 -18304 -2066 -18288
rect -4176 -18329 -4142 -18313
rect -2172 -18352 -2138 -18336
rect -2172 -18459 -2138 -18443
rect -4176 -18477 -4142 -18461
rect -4278 -18502 -4244 -18486
rect -4528 -18522 -4494 -18504
rect -2100 -18510 -2066 -18500
rect -2004 -18300 -1970 -18282
rect -2004 -18510 -1970 -18494
rect -1908 -18304 -1874 -18288
rect -1908 -18510 -1874 -18500
rect -1812 -18300 -1778 -18282
rect -1812 -18510 -1778 -18494
rect -1650 -18318 -1616 -18302
rect -1650 -18510 -1616 -18494
rect -1562 -18318 -1528 -18302
rect -1460 -18343 -1426 -18327
rect -1460 -18491 -1426 -18475
rect -1562 -18510 -1528 -18494
rect 15775 -18527 15809 -18511
rect 15871 -17679 15905 -17663
rect 15871 -18527 15905 -18511
rect 15967 -17679 16001 -17663
rect 15967 -18527 16001 -18511
rect 16063 -17679 16097 -17663
rect 16063 -18527 16097 -18511
rect 16159 -17679 16193 -17663
rect 16159 -18527 16193 -18511
rect 16255 -17679 16289 -17663
rect 16255 -18527 16289 -18511
rect 16351 -17679 16385 -17663
rect 16351 -18527 16385 -18511
rect 16447 -17679 16481 -17663
rect 16447 -18527 16481 -18511
rect 16543 -17679 16577 -17663
rect 16543 -18527 16577 -18511
rect 16639 -17679 16673 -17663
rect 16639 -18527 16673 -18511
rect 16735 -17679 16769 -17663
rect 16735 -18527 16769 -18511
rect 16831 -17679 16865 -17663
rect 16831 -18527 16865 -18511
rect 16927 -17679 16961 -17663
rect 17306 -18209 17322 -18162
rect 17891 -18209 17915 -18162
rect 18143 -18221 18159 -18187
rect 18250 -18221 18266 -18187
rect 17306 -18281 17340 -18271
rect 17306 -18493 17340 -18477
rect 17402 -18287 17436 -18271
rect 17402 -18493 17436 -18483
rect 17498 -18281 17532 -18271
rect 17498 -18493 17532 -18477
rect 17594 -18287 17628 -18271
rect 17594 -18493 17628 -18483
rect 17690 -18281 17724 -18271
rect 17690 -18493 17724 -18477
rect 17786 -18287 17820 -18271
rect 17786 -18493 17820 -18483
rect 17882 -18281 17916 -18271
rect 17882 -18493 17916 -18477
rect 17999 -18307 18049 -18290
rect 18092 -18293 18102 -18259
rect 18298 -18293 18314 -18259
rect 16927 -18527 16961 -18511
rect 17999 -18533 18015 -18307
rect 18092 -18389 18108 -18355
rect 18302 -18389 18320 -18355
rect 18092 -18485 18102 -18451
rect 18298 -18485 18314 -18451
rect -15374 -18604 -15340 -18588
rect -2069 -18587 -2052 -18553
rect -1826 -18587 -1606 -18553
rect -1572 -18587 -1556 -18553
rect -2069 -18603 -1556 -18587
rect 17355 -18571 17372 -18536
rect 17406 -18571 17422 -18536
rect 17644 -18542 17661 -18536
rect 17456 -18571 17661 -18542
rect 17695 -18571 17711 -18536
rect -15476 -18623 -15442 -18607
rect -4785 -18657 -4272 -18641
rect -15983 -18700 -15966 -18666
rect -15740 -18700 -15520 -18666
rect -15486 -18700 -15470 -18666
rect -4785 -18691 -4768 -18657
rect -4542 -18691 -4322 -18657
rect -4288 -18691 -4272 -18657
rect 5705 -18691 5721 -18657
rect 5812 -18691 5828 -18657
rect 6145 -18691 6161 -18657
rect 6252 -18691 6268 -18657
rect 6585 -18691 6601 -18657
rect 6692 -18691 6708 -18657
rect 15775 -18661 15809 -18645
rect -20965 -18733 -20931 -18717
rect -21067 -18752 -21033 -18736
rect -17681 -18745 -17665 -18711
rect -17433 -18745 -17417 -18711
rect -15983 -18716 -15470 -18700
rect -8179 -18718 -8145 -18702
rect -8251 -18766 -8217 -18750
rect -23808 -18833 -23774 -18806
rect -21574 -18829 -21557 -18795
rect -21331 -18829 -21111 -18795
rect -21077 -18829 -21061 -18795
rect -21574 -18845 -21061 -18829
rect -17681 -18841 -17665 -18807
rect -17433 -18841 -17417 -18807
rect -24161 -18905 -24043 -18871
rect -24008 -18905 -23992 -18871
rect -23926 -18905 -23910 -18871
rect -23875 -18905 -23859 -18871
rect -8251 -18873 -8217 -18857
rect -16015 -18897 -15981 -18881
rect -24432 -18959 -24416 -18925
rect -24220 -18959 -24210 -18925
rect -24167 -18955 -24132 -18939
rect -23926 -18963 -23859 -18905
rect -17681 -18937 -17665 -18903
rect -17433 -18937 -17417 -18903
rect -24132 -18989 -23859 -18963
rect -24167 -19006 -23859 -18989
rect -16087 -18945 -16053 -18929
rect -24541 -19055 -24494 -19039
rect -24432 -19055 -24422 -19021
rect -24226 -19055 -24210 -19021
rect -21606 -19026 -21572 -19010
rect -21678 -19074 -21644 -19058
rect -21678 -19181 -21644 -19165
rect -21606 -19232 -21572 -19222
rect -21510 -19022 -21476 -19004
rect -21510 -19232 -21476 -19216
rect -21414 -19026 -21380 -19010
rect -21414 -19232 -21380 -19222
rect -21318 -19022 -21284 -19004
rect -21318 -19232 -21284 -19216
rect -21156 -19040 -21122 -19024
rect -21156 -19232 -21122 -19216
rect -21068 -19040 -21034 -19024
rect -17681 -19033 -17665 -18999
rect -17433 -19033 -17417 -18999
rect -20966 -19065 -20932 -19049
rect -16087 -19052 -16053 -19036
rect -16928 -19095 -16844 -19083
rect -17681 -19129 -17665 -19095
rect -17433 -19129 -17417 -19095
rect -17266 -19143 -17232 -19127
rect -17192 -19129 -17176 -19095
rect -17000 -19108 -16844 -19095
rect -16015 -19103 -15981 -19093
rect -15919 -18893 -15885 -18875
rect -15919 -19103 -15885 -19087
rect -15823 -18897 -15789 -18881
rect -15823 -19103 -15789 -19093
rect -15727 -18893 -15693 -18875
rect -15727 -19103 -15693 -19087
rect -15565 -18911 -15531 -18895
rect -15565 -19103 -15531 -19087
rect -15477 -18911 -15443 -18895
rect -15375 -18936 -15341 -18920
rect -8179 -18924 -8145 -18914
rect -8083 -18714 -8049 -18696
rect -8083 -18924 -8049 -18908
rect -7987 -18718 -7953 -18702
rect -7987 -18924 -7953 -18914
rect -7891 -18714 -7857 -18696
rect -7891 -18924 -7857 -18908
rect -7729 -18732 -7695 -18716
rect -7729 -18924 -7695 -18908
rect -7641 -18732 -7607 -18716
rect -7539 -18757 -7505 -18741
rect -4816 -18744 -4782 -18734
rect -7539 -18905 -7505 -18889
rect -4888 -18801 -4854 -18785
rect -4888 -18908 -4854 -18892
rect -7641 -18924 -7607 -18908
rect -4816 -18956 -4782 -18940
rect -4720 -18750 -4686 -18734
rect -4720 -18962 -4686 -18944
rect -4624 -18744 -4590 -18734
rect -4624 -18956 -4590 -18940
rect -4528 -18750 -4494 -18734
rect -4366 -18750 -4332 -18734
rect -4366 -18942 -4332 -18926
rect -4278 -18750 -4244 -18734
rect -2100 -18744 -2066 -18728
rect -4176 -18769 -4142 -18753
rect -2172 -18792 -2138 -18776
rect -2172 -18899 -2138 -18883
rect -4176 -18917 -4142 -18901
rect -4278 -18942 -4244 -18926
rect -4528 -18962 -4494 -18944
rect -2100 -18950 -2066 -18940
rect -2004 -18740 -1970 -18722
rect -2004 -18950 -1970 -18934
rect -1908 -18744 -1874 -18728
rect -1908 -18950 -1874 -18940
rect -1812 -18740 -1778 -18722
rect -1812 -18950 -1778 -18934
rect -1650 -18758 -1616 -18742
rect -1650 -18950 -1616 -18934
rect -1562 -18758 -1528 -18742
rect -1460 -18783 -1426 -18767
rect -1460 -18931 -1426 -18915
rect 5561 -18777 5611 -18760
rect 5654 -18763 5664 -18729
rect 5860 -18763 5876 -18729
rect -1562 -18950 -1528 -18934
rect -8148 -19001 -8131 -18967
rect -7905 -19001 -7685 -18967
rect -7651 -19001 -7635 -18967
rect -8148 -19017 -7635 -19001
rect -15375 -19084 -15341 -19068
rect -4785 -19036 -4272 -19020
rect -4785 -19070 -4768 -19036
rect -4542 -19070 -4322 -19036
rect -4288 -19070 -4272 -19036
rect -2069 -19027 -2052 -18993
rect -1826 -19027 -1606 -18993
rect -1572 -19027 -1556 -18993
rect -2069 -19043 -1556 -19027
rect 5561 -19003 5577 -18777
rect 6001 -18777 6051 -18760
rect 6094 -18763 6104 -18729
rect 6300 -18763 6316 -18729
rect 5654 -18859 5670 -18825
rect 5864 -18859 5882 -18825
rect 5654 -18955 5664 -18921
rect 5860 -18955 5876 -18921
rect -15477 -19103 -15443 -19087
rect -17000 -19129 -16917 -19108
rect -20966 -19213 -20932 -19197
rect -21068 -19232 -21034 -19216
rect -17681 -19225 -17665 -19191
rect -17433 -19225 -17417 -19191
rect -17266 -19193 -17232 -19177
rect -17192 -19225 -17176 -19191
rect -17000 -19225 -16984 -19191
rect -21575 -19309 -21558 -19275
rect -21332 -19309 -21112 -19275
rect -21078 -19309 -21062 -19275
rect -17371 -19286 -17337 -19270
rect -21575 -19325 -21062 -19309
rect -17840 -19321 -17665 -19287
rect -17433 -19321 -17417 -19287
rect -16928 -19287 -16917 -19129
rect -17840 -19322 -17750 -19321
rect -21606 -19526 -21572 -19510
rect -21678 -19574 -21644 -19558
rect -24070 -19639 -24036 -19623
rect -24539 -19664 -24492 -19640
rect -24430 -19673 -24420 -19639
rect -24224 -19673 -24208 -19639
rect -24430 -19769 -24414 -19735
rect -24218 -19769 -24208 -19735
rect -24430 -19865 -24420 -19831
rect -24224 -19865 -24208 -19831
rect -24165 -19860 -24125 -19844
rect -24130 -19894 -24125 -19860
rect -24165 -19911 -24125 -19894
rect -24430 -19961 -24414 -19927
rect -24218 -19961 -24208 -19927
rect -24430 -20057 -24420 -20023
rect -24224 -20057 -24208 -20023
rect -24159 -20065 -24125 -19911
rect -24070 -20031 -24036 -20015
rect -23878 -19639 -23844 -19623
rect -23878 -20031 -23844 -20015
rect -23806 -19665 -23772 -19627
rect -21678 -19681 -21644 -19665
rect -21606 -19732 -21572 -19722
rect -21510 -19522 -21476 -19504
rect -21510 -19732 -21476 -19716
rect -21414 -19526 -21380 -19510
rect -21414 -19732 -21380 -19722
rect -21318 -19522 -21284 -19504
rect -21318 -19732 -21284 -19716
rect -21156 -19540 -21122 -19524
rect -21156 -19732 -21122 -19716
rect -21068 -19540 -21034 -19524
rect -20966 -19565 -20932 -19549
rect -20966 -19713 -20932 -19697
rect -17840 -19679 -17820 -19322
rect -17769 -19479 -17750 -19322
rect -17371 -19336 -17337 -19320
rect -17192 -19321 -17176 -19287
rect -17000 -19307 -16917 -19287
rect -16856 -19307 -16844 -19108
rect -4816 -19123 -4782 -19113
rect -15984 -19180 -15967 -19146
rect -15741 -19180 -15521 -19146
rect -15487 -19180 -15471 -19146
rect -15984 -19196 -15471 -19180
rect -4888 -19180 -4854 -19164
rect -4888 -19287 -4854 -19271
rect -17000 -19321 -16844 -19307
rect -16928 -19333 -16844 -19321
rect -4816 -19335 -4782 -19319
rect -4720 -19129 -4686 -19113
rect -4720 -19341 -4686 -19323
rect -4624 -19123 -4590 -19113
rect -4624 -19335 -4590 -19319
rect -4528 -19129 -4494 -19113
rect -4366 -19129 -4332 -19113
rect -4366 -19321 -4332 -19305
rect -4278 -19129 -4244 -19113
rect -2100 -19123 -2066 -19107
rect -4176 -19148 -4142 -19132
rect -2172 -19171 -2138 -19155
rect -2172 -19278 -2138 -19262
rect -4176 -19296 -4142 -19280
rect -4278 -19321 -4244 -19305
rect -4528 -19341 -4494 -19323
rect -2100 -19329 -2066 -19319
rect -2004 -19119 -1970 -19101
rect -2004 -19329 -1970 -19313
rect -1908 -19123 -1874 -19107
rect -1908 -19329 -1874 -19319
rect -1812 -19119 -1778 -19101
rect -1812 -19329 -1778 -19313
rect -1650 -19137 -1616 -19121
rect -1650 -19329 -1616 -19313
rect -1562 -19137 -1528 -19121
rect -1460 -19162 -1426 -19146
rect 5561 -19223 5611 -19003
rect 6001 -19003 6017 -18777
rect 6441 -18777 6491 -18760
rect 6534 -18763 6544 -18729
rect 6740 -18763 6756 -18729
rect 6094 -18859 6110 -18825
rect 6304 -18859 6322 -18825
rect 6094 -18955 6104 -18921
rect 6300 -18955 6316 -18921
rect 5654 -19051 5670 -19017
rect 5864 -19051 5882 -19017
rect 5654 -19213 5670 -19179
rect 5846 -19213 5862 -19179
rect 5561 -19257 5577 -19223
rect 5561 -19273 5611 -19257
rect 6001 -19223 6051 -19003
rect 6441 -19003 6457 -18777
rect 6534 -18859 6550 -18825
rect 6744 -18859 6762 -18825
rect 6534 -18955 6544 -18921
rect 6740 -18955 6756 -18921
rect 6094 -19051 6110 -19017
rect 6304 -19051 6322 -19017
rect 6094 -19213 6110 -19179
rect 6286 -19213 6302 -19179
rect 6001 -19257 6017 -19223
rect -1460 -19310 -1426 -19294
rect 5654 -19301 5670 -19267
rect 5846 -19301 5862 -19267
rect 6001 -19273 6051 -19257
rect 6441 -19223 6491 -19003
rect 6534 -19051 6550 -19017
rect 6744 -19051 6762 -19017
rect 15703 -19139 15737 -19123
rect 6534 -19213 6550 -19179
rect 6726 -19213 6742 -19179
rect 6441 -19257 6457 -19223
rect 6094 -19301 6110 -19267
rect 6286 -19301 6302 -19267
rect 6441 -19273 6491 -19257
rect 6534 -19301 6550 -19267
rect 6726 -19301 6742 -19267
rect -1562 -19329 -1528 -19313
rect 7373 -19364 7389 -19329
rect 7677 -19364 7703 -19329
rect 8321 -19364 8337 -19329
rect 8625 -19364 8651 -19329
rect 9257 -19364 9273 -19329
rect 9561 -19364 9587 -19329
rect 10188 -19364 10204 -19329
rect 10492 -19364 10518 -19329
rect 11115 -19364 11131 -19329
rect 11419 -19364 11445 -19329
rect -17681 -19417 -17665 -19383
rect -17433 -19417 -17417 -19383
rect -16015 -19397 -15981 -19381
rect -16087 -19445 -16053 -19429
rect -17769 -19513 -17665 -19479
rect -17433 -19513 -17417 -19479
rect -17769 -19671 -17750 -19513
rect -16087 -19552 -16053 -19536
rect -17681 -19609 -17665 -19575
rect -17433 -19609 -17417 -19575
rect -16015 -19603 -15981 -19593
rect -15919 -19393 -15885 -19375
rect -15919 -19603 -15885 -19587
rect -15823 -19397 -15789 -19381
rect -15823 -19603 -15789 -19593
rect -15727 -19393 -15693 -19375
rect -15727 -19603 -15693 -19587
rect -15565 -19411 -15531 -19395
rect -15565 -19603 -15531 -19587
rect -15477 -19411 -15443 -19395
rect -2069 -19406 -2052 -19372
rect -1826 -19406 -1606 -19372
rect -1572 -19406 -1556 -19372
rect 5673 -19403 5689 -19369
rect 5821 -19403 5837 -19369
rect 6113 -19403 6129 -19369
rect 6261 -19403 6277 -19369
rect 6553 -19403 6569 -19369
rect 6701 -19403 6717 -19369
rect -15375 -19436 -15341 -19420
rect -2069 -19422 -1556 -19406
rect 7150 -19433 7184 -19417
rect -4785 -19476 -4272 -19460
rect -4785 -19510 -4768 -19476
rect -4542 -19510 -4322 -19476
rect -4288 -19510 -4272 -19476
rect -15375 -19584 -15341 -19568
rect -4816 -19563 -4782 -19553
rect -15477 -19603 -15443 -19587
rect -4888 -19620 -4854 -19604
rect -17769 -19679 -17665 -19671
rect -17840 -19705 -17665 -19679
rect -17433 -19705 -17417 -19671
rect -15984 -19680 -15967 -19646
rect -15741 -19680 -15521 -19646
rect -15487 -19680 -15471 -19646
rect -15984 -19696 -15471 -19680
rect -17840 -19707 -17750 -19705
rect -21068 -19732 -21034 -19716
rect -4888 -19727 -4854 -19711
rect -4816 -19775 -4782 -19759
rect -4720 -19569 -4686 -19553
rect -21575 -19809 -21558 -19775
rect -21332 -19809 -21112 -19775
rect -21078 -19809 -21062 -19775
rect -4720 -19781 -4686 -19763
rect -4624 -19563 -4590 -19553
rect -4624 -19775 -4590 -19759
rect -4528 -19569 -4494 -19553
rect -4366 -19569 -4332 -19553
rect -4366 -19761 -4332 -19745
rect -4278 -19569 -4244 -19553
rect -2100 -19563 -2066 -19547
rect -4176 -19588 -4142 -19572
rect -2172 -19611 -2138 -19595
rect -2172 -19718 -2138 -19702
rect -4176 -19736 -4142 -19720
rect -4278 -19761 -4244 -19745
rect -4528 -19781 -4494 -19763
rect -2100 -19769 -2066 -19759
rect -2004 -19559 -1970 -19541
rect -2004 -19769 -1970 -19753
rect -1908 -19563 -1874 -19547
rect -1908 -19769 -1874 -19759
rect -1812 -19559 -1778 -19541
rect -1812 -19769 -1778 -19753
rect -1650 -19577 -1616 -19561
rect -1650 -19769 -1616 -19753
rect -1562 -19577 -1528 -19561
rect -1460 -19602 -1426 -19586
rect -1460 -19750 -1426 -19734
rect 7246 -19433 7280 -19417
rect 7150 -19747 7184 -19731
rect 7246 -19747 7280 -19736
rect 7342 -19433 7376 -19417
rect 7342 -19747 7376 -19731
rect 7438 -19433 7472 -19417
rect 7534 -19433 7568 -19417
rect 7438 -19747 7472 -19736
rect 7534 -19747 7568 -19731
rect 7630 -19433 7664 -19417
rect 7726 -19433 7760 -19417
rect 7630 -19747 7664 -19736
rect 7726 -19747 7760 -19731
rect 7822 -19433 7856 -19417
rect 7918 -19433 7952 -19417
rect 7822 -19747 7856 -19736
rect 7918 -19747 7952 -19731
rect 8098 -19433 8132 -19417
rect 8194 -19433 8228 -19417
rect 8098 -19747 8132 -19731
rect 8194 -19747 8228 -19736
rect 8290 -19433 8324 -19417
rect 8290 -19747 8324 -19731
rect 8386 -19433 8420 -19417
rect 8482 -19433 8516 -19417
rect 8386 -19747 8420 -19736
rect 8482 -19747 8516 -19731
rect 8578 -19433 8612 -19417
rect 8674 -19433 8708 -19417
rect 8578 -19747 8612 -19736
rect 8674 -19747 8708 -19731
rect 8770 -19433 8804 -19417
rect 8866 -19433 8900 -19417
rect 8770 -19747 8804 -19736
rect 8866 -19747 8900 -19731
rect 9034 -19433 9068 -19417
rect 9130 -19433 9164 -19417
rect 9034 -19747 9068 -19731
rect 9130 -19747 9164 -19736
rect 9226 -19433 9260 -19417
rect 9226 -19747 9260 -19731
rect 9322 -19433 9356 -19417
rect 9418 -19433 9452 -19417
rect 9322 -19747 9356 -19736
rect 9418 -19747 9452 -19731
rect 9514 -19433 9548 -19417
rect 9610 -19433 9644 -19417
rect 9514 -19747 9548 -19736
rect 9610 -19747 9644 -19731
rect 9706 -19433 9740 -19417
rect 9802 -19433 9836 -19417
rect 9706 -19747 9740 -19736
rect 9802 -19747 9836 -19731
rect 9965 -19433 9999 -19417
rect 10061 -19433 10095 -19417
rect 9965 -19747 9999 -19731
rect 10061 -19747 10095 -19736
rect 10157 -19433 10191 -19417
rect 10157 -19747 10191 -19731
rect 10253 -19433 10287 -19417
rect 10349 -19433 10383 -19417
rect 10253 -19747 10287 -19736
rect 10349 -19747 10383 -19731
rect 10445 -19433 10479 -19417
rect 10541 -19433 10575 -19417
rect 10445 -19747 10479 -19736
rect 10541 -19747 10575 -19731
rect 10637 -19433 10671 -19417
rect 10733 -19433 10767 -19417
rect 10637 -19747 10671 -19736
rect 10733 -19747 10767 -19731
rect 10892 -19433 10926 -19417
rect 10988 -19433 11022 -19417
rect 10892 -19747 10926 -19731
rect 10988 -19747 11022 -19736
rect 11084 -19433 11118 -19417
rect 11084 -19747 11118 -19731
rect 11180 -19433 11214 -19417
rect 11276 -19433 11310 -19417
rect 11180 -19747 11214 -19736
rect 11276 -19747 11310 -19731
rect 11372 -19433 11406 -19417
rect 11468 -19433 11502 -19417
rect 11372 -19747 11406 -19736
rect 11468 -19747 11502 -19731
rect 11564 -19433 11598 -19417
rect 11660 -19433 11694 -19417
rect 15703 -19509 15737 -19493
rect 15775 -19509 15809 -19493
rect 15871 -18661 15905 -18645
rect 15871 -19509 15905 -19493
rect 15967 -18661 16001 -18645
rect 15967 -19509 16001 -19493
rect 16063 -18661 16097 -18645
rect 16063 -19509 16097 -19493
rect 16159 -18661 16193 -18645
rect 16159 -19509 16193 -19493
rect 16255 -18661 16289 -18645
rect 16255 -19509 16289 -19493
rect 16351 -18661 16385 -18645
rect 16351 -19509 16385 -19493
rect 16447 -18661 16481 -18645
rect 16447 -19509 16481 -19493
rect 16543 -18661 16577 -18645
rect 16543 -19509 16577 -19493
rect 16639 -18661 16673 -18645
rect 16639 -19509 16673 -19493
rect 16735 -18661 16769 -18645
rect 16735 -19509 16769 -19493
rect 16831 -18661 16865 -18645
rect 16831 -19509 16865 -19493
rect 16927 -18661 16961 -18645
rect 17355 -18777 17398 -18571
rect 17456 -18576 17711 -18571
rect 17456 -18660 17490 -18576
rect 17524 -18665 17540 -18631
rect 17916 -18665 17932 -18631
rect 17456 -18711 17490 -18695
rect 17999 -18753 18049 -18533
rect 18092 -18581 18108 -18547
rect 18302 -18581 18320 -18547
rect 18092 -18743 18108 -18709
rect 18284 -18743 18300 -18709
rect 17355 -18793 17490 -18777
rect 17355 -18828 17456 -18793
rect 17999 -18787 18015 -18753
rect 17999 -18803 18049 -18787
rect 17355 -18844 17490 -18828
rect 17524 -18857 17540 -18823
rect 17916 -18857 17932 -18823
rect 18092 -18831 18108 -18797
rect 18284 -18831 18300 -18797
rect 17528 -18929 17555 -18895
rect 17890 -18929 17928 -18895
rect 18111 -18933 18127 -18899
rect 18259 -18933 18275 -18899
rect 16927 -19509 16961 -19493
rect 15981 -19586 15997 -19552
rect 16031 -19586 16047 -19552
rect 16269 -19586 16285 -19552
rect 16319 -19586 16335 -19552
rect 16401 -19586 16417 -19552
rect 16451 -19586 16467 -19552
rect 11564 -19747 11598 -19736
rect 11660 -19747 11694 -19731
rect -1562 -19769 -1528 -19753
rect -21575 -19825 -21062 -19809
rect -4785 -19855 -4272 -19839
rect -16015 -19877 -15981 -19861
rect -16087 -19925 -16053 -19909
rect -23806 -20027 -23772 -20000
rect -21606 -20006 -21572 -19990
rect -21678 -20054 -21644 -20038
rect -24159 -20099 -24041 -20065
rect -24006 -20099 -23990 -20065
rect -23924 -20099 -23908 -20065
rect -23873 -20099 -23857 -20065
rect -24430 -20153 -24414 -20119
rect -24218 -20153 -24208 -20119
rect -24165 -20149 -24130 -20133
rect -23924 -20157 -23857 -20099
rect -24130 -20183 -23857 -20157
rect -21678 -20161 -21644 -20145
rect -24165 -20200 -23857 -20183
rect -21606 -20212 -21572 -20202
rect -21510 -20002 -21476 -19984
rect -21510 -20212 -21476 -20196
rect -21414 -20006 -21380 -19990
rect -21414 -20212 -21380 -20202
rect -21318 -20002 -21284 -19984
rect -21318 -20212 -21284 -20196
rect -21156 -20020 -21122 -20004
rect -21156 -20212 -21122 -20196
rect -21068 -20020 -21034 -20004
rect -20966 -20045 -20932 -20029
rect -16087 -20032 -16053 -20016
rect -16015 -20083 -15981 -20073
rect -15919 -19873 -15885 -19855
rect -15919 -20083 -15885 -20067
rect -15823 -19877 -15789 -19861
rect -15823 -20083 -15789 -20073
rect -15727 -19873 -15693 -19855
rect -15727 -20083 -15693 -20067
rect -15565 -19891 -15531 -19875
rect -15565 -20083 -15531 -20067
rect -15477 -19891 -15443 -19875
rect -15375 -19916 -15341 -19900
rect -12318 -19912 -12302 -19878
rect -11776 -19912 -11262 -19878
rect -11156 -19912 -11140 -19878
rect -4785 -19889 -4768 -19855
rect -4542 -19889 -4322 -19855
rect -4288 -19889 -4272 -19855
rect -2069 -19846 -2052 -19812
rect -1826 -19846 -1606 -19812
rect -1572 -19846 -1556 -19812
rect 7182 -19824 7198 -19790
rect 7232 -19824 7248 -19790
rect 7374 -19824 7390 -19790
rect 7424 -19824 7440 -19790
rect 7566 -19824 7582 -19790
rect 7616 -19824 7632 -19790
rect 7758 -19824 7774 -19790
rect 7808 -19824 7824 -19790
rect 8130 -19824 8146 -19790
rect 8180 -19824 8196 -19790
rect 8322 -19824 8338 -19790
rect 8372 -19824 8388 -19790
rect 8514 -19824 8530 -19790
rect 8564 -19824 8580 -19790
rect 8706 -19824 8722 -19790
rect 8756 -19824 8772 -19790
rect 9066 -19824 9082 -19790
rect 9116 -19824 9132 -19790
rect 9258 -19824 9274 -19790
rect 9308 -19824 9324 -19790
rect 9450 -19824 9466 -19790
rect 9500 -19824 9516 -19790
rect 9642 -19824 9658 -19790
rect 9692 -19824 9708 -19790
rect 9997 -19824 10013 -19790
rect 10047 -19824 10063 -19790
rect 10189 -19824 10205 -19790
rect 10239 -19824 10255 -19790
rect 10381 -19824 10397 -19790
rect 10431 -19824 10447 -19790
rect 10573 -19824 10589 -19790
rect 10623 -19824 10639 -19790
rect 10924 -19824 10940 -19790
rect 10974 -19824 10990 -19790
rect 11116 -19824 11132 -19790
rect 11166 -19824 11182 -19790
rect 11308 -19824 11324 -19790
rect 11358 -19824 11374 -19790
rect 11500 -19824 11516 -19790
rect 11550 -19824 11566 -19790
rect -2069 -19862 -1556 -19846
rect 16653 -19868 16669 -19834
rect 16703 -19868 16719 -19834
rect -15375 -20064 -15341 -20048
rect -12499 -19996 -12373 -19954
rect -15477 -20083 -15443 -20067
rect -17681 -20145 -17665 -20111
rect -17433 -20145 -17417 -20111
rect -15984 -20160 -15967 -20126
rect -15741 -20160 -15521 -20126
rect -15487 -20160 -15471 -20126
rect -15984 -20176 -15471 -20160
rect -20966 -20193 -20932 -20177
rect -21068 -20212 -21034 -20196
rect -24539 -20249 -24492 -20233
rect -24430 -20249 -24420 -20215
rect -24224 -20249 -24208 -20215
rect -17681 -20241 -17665 -20207
rect -17433 -20241 -17417 -20207
rect -21575 -20289 -21558 -20255
rect -21332 -20289 -21112 -20255
rect -21078 -20289 -21062 -20255
rect -21575 -20305 -21062 -20289
rect -17681 -20337 -17665 -20303
rect -17433 -20337 -17417 -20303
rect -16015 -20337 -15981 -20321
rect -16087 -20385 -16053 -20369
rect -17681 -20433 -17665 -20399
rect -17433 -20433 -17417 -20399
rect -21606 -20466 -21572 -20450
rect -21678 -20514 -21644 -20498
rect -21678 -20621 -21644 -20605
rect -21606 -20672 -21572 -20662
rect -21510 -20462 -21476 -20444
rect -21510 -20672 -21476 -20656
rect -21414 -20466 -21380 -20450
rect -21414 -20672 -21380 -20662
rect -21318 -20462 -21284 -20444
rect -21318 -20672 -21284 -20656
rect -21156 -20480 -21122 -20464
rect -21156 -20672 -21122 -20656
rect -21068 -20480 -21034 -20464
rect -20966 -20505 -20932 -20489
rect -16928 -20495 -16844 -20483
rect -16087 -20492 -16053 -20476
rect -17681 -20529 -17665 -20495
rect -17433 -20529 -17417 -20495
rect -17266 -20543 -17232 -20527
rect -17192 -20529 -17176 -20495
rect -17000 -20508 -16844 -20495
rect -17000 -20529 -16917 -20508
rect -17681 -20625 -17665 -20591
rect -17433 -20625 -17417 -20591
rect -17266 -20593 -17232 -20577
rect -17192 -20625 -17176 -20591
rect -17000 -20625 -16984 -20591
rect -20966 -20653 -20932 -20637
rect -21068 -20672 -21034 -20656
rect -17371 -20686 -17337 -20670
rect -21575 -20749 -21558 -20715
rect -21332 -20749 -21112 -20715
rect -21078 -20749 -21062 -20715
rect -21575 -20765 -21062 -20749
rect -17840 -20721 -17665 -20687
rect -17433 -20721 -17417 -20687
rect -16928 -20687 -16917 -20529
rect -17840 -20722 -17750 -20721
rect -24039 -20839 -24005 -20823
rect -24508 -20864 -24461 -20840
rect -24399 -20873 -24389 -20839
rect -24193 -20873 -24177 -20839
rect -24399 -20969 -24383 -20935
rect -24187 -20969 -24177 -20935
rect -24399 -21065 -24389 -21031
rect -24193 -21065 -24177 -21031
rect -24134 -21060 -24094 -21044
rect -24099 -21094 -24094 -21060
rect -24134 -21111 -24094 -21094
rect -24399 -21161 -24383 -21127
rect -24187 -21161 -24177 -21127
rect -24399 -21257 -24389 -21223
rect -24193 -21257 -24177 -21223
rect -24128 -21265 -24094 -21111
rect -24039 -21231 -24005 -21215
rect -23847 -20839 -23813 -20823
rect -23847 -21231 -23813 -21215
rect -23775 -20865 -23741 -20827
rect -21620 -20926 -21586 -20910
rect -21692 -20974 -21658 -20958
rect -21692 -21081 -21658 -21065
rect -21620 -21132 -21586 -21122
rect -21524 -20922 -21490 -20904
rect -21524 -21132 -21490 -21116
rect -21428 -20926 -21394 -20910
rect -21428 -21132 -21394 -21122
rect -21332 -20922 -21298 -20904
rect -21332 -21132 -21298 -21116
rect -21170 -20940 -21136 -20924
rect -21170 -21132 -21136 -21116
rect -21082 -20940 -21048 -20924
rect -20980 -20965 -20946 -20949
rect -20980 -21113 -20946 -21097
rect -17840 -21079 -17820 -20722
rect -17769 -20879 -17750 -20722
rect -17371 -20736 -17337 -20720
rect -17192 -20721 -17176 -20687
rect -17000 -20707 -16917 -20687
rect -16856 -20707 -16844 -20508
rect -16015 -20543 -15981 -20533
rect -15919 -20333 -15885 -20315
rect -15919 -20543 -15885 -20527
rect -15823 -20337 -15789 -20321
rect -15823 -20543 -15789 -20533
rect -15727 -20333 -15693 -20315
rect -15727 -20543 -15693 -20527
rect -15565 -20351 -15531 -20335
rect -15565 -20543 -15531 -20527
rect -15477 -20351 -15443 -20335
rect -15375 -20376 -15341 -20360
rect -15375 -20524 -15341 -20508
rect -15477 -20543 -15443 -20527
rect -15984 -20620 -15967 -20586
rect -15741 -20620 -15521 -20586
rect -15487 -20620 -15471 -20586
rect -15984 -20636 -15471 -20620
rect -17000 -20721 -16844 -20707
rect -16928 -20733 -16844 -20721
rect -17681 -20817 -17665 -20783
rect -17433 -20817 -17417 -20783
rect -16029 -20797 -15995 -20781
rect -16101 -20845 -16067 -20829
rect -17769 -20913 -17665 -20879
rect -17433 -20913 -17417 -20879
rect -17769 -21071 -17750 -20913
rect -16101 -20952 -16067 -20936
rect -17681 -21009 -17665 -20975
rect -17433 -21009 -17417 -20975
rect -16029 -21003 -15995 -20993
rect -15933 -20793 -15899 -20775
rect -15933 -21003 -15899 -20987
rect -15837 -20797 -15803 -20781
rect -15837 -21003 -15803 -20993
rect -15741 -20793 -15707 -20775
rect -15741 -21003 -15707 -20987
rect -15579 -20811 -15545 -20795
rect -15579 -21003 -15545 -20987
rect -15491 -20811 -15457 -20795
rect -15389 -20836 -15355 -20820
rect -15389 -20984 -15355 -20968
rect -15491 -21003 -15457 -20987
rect -17769 -21079 -17665 -21071
rect -17840 -21105 -17665 -21079
rect -17433 -21105 -17417 -21071
rect -15998 -21080 -15981 -21046
rect -15755 -21080 -15535 -21046
rect -15501 -21080 -15485 -21046
rect -15998 -21096 -15485 -21080
rect -17840 -21107 -17750 -21105
rect -21082 -21132 -21048 -21116
rect -12499 -21118 -12471 -19996
rect -12399 -21118 -12373 -19996
rect -12318 -20000 -12302 -19966
rect -11776 -20000 -11760 -19966
rect -12318 -20096 -12302 -20062
rect -11776 -20096 -11760 -20062
rect -12318 -20192 -12302 -20158
rect -11776 -20192 -11760 -20158
rect -12318 -20288 -12302 -20254
rect -11776 -20288 -11760 -20254
rect -11718 -20303 -11641 -19912
rect -4816 -19942 -4782 -19932
rect -11433 -19967 -11337 -19952
rect -11433 -20032 -11411 -19967
rect -11356 -20032 -11337 -19967
rect -11278 -20000 -11262 -19966
rect -11156 -20000 -11140 -19966
rect -11090 -19995 -10999 -19957
rect -11600 -20134 -11494 -20116
rect -11600 -20214 -11582 -20134
rect -11514 -20214 -11494 -20134
rect -11600 -20231 -11494 -20214
rect -11718 -20323 -11501 -20303
rect -12318 -20384 -12302 -20350
rect -11776 -20384 -11760 -20350
rect -12318 -20480 -12302 -20446
rect -11776 -20480 -11760 -20446
rect -11718 -20453 -11700 -20323
rect -11655 -20334 -11501 -20323
rect -11655 -20448 -11583 -20334
rect -11530 -20448 -11501 -20334
rect -11655 -20453 -11501 -20448
rect -11718 -20480 -11501 -20453
rect -11433 -20526 -11337 -20032
rect -11278 -20096 -11277 -20062
rect -11156 -20096 -11140 -20062
rect -11278 -20192 -11262 -20158
rect -11142 -20192 -11140 -20158
rect -11278 -20288 -11277 -20254
rect -11156 -20288 -11140 -20254
rect -11278 -20384 -11262 -20350
rect -11142 -20384 -11140 -20350
rect -11278 -20480 -11277 -20446
rect -11156 -20480 -11140 -20446
rect -11733 -20542 -11303 -20526
rect -12318 -20576 -12302 -20542
rect -11776 -20576 -11262 -20542
rect -11142 -20576 -11140 -20542
rect -11733 -20592 -11303 -20576
rect -12318 -20672 -12302 -20638
rect -11776 -20672 -11760 -20638
rect -11715 -20646 -11314 -20638
rect -11715 -20654 -11376 -20646
rect -12318 -20768 -12302 -20734
rect -11776 -20768 -11760 -20734
rect -11715 -20784 -11705 -20654
rect -11660 -20776 -11376 -20654
rect -11331 -20776 -11314 -20646
rect -11278 -20672 -11276 -20638
rect -11156 -20672 -11140 -20638
rect -11278 -20768 -11262 -20734
rect -11142 -20768 -11140 -20734
rect -11660 -20784 -11314 -20776
rect -11715 -20803 -11314 -20784
rect -12318 -20864 -12302 -20830
rect -11776 -20864 -11760 -20830
rect -12318 -20960 -12302 -20926
rect -11776 -20960 -11760 -20926
rect -12318 -21056 -12302 -21022
rect -11776 -21056 -11760 -21022
rect -12499 -21164 -12373 -21118
rect -12318 -21152 -12302 -21118
rect -11776 -21152 -11760 -21118
rect -23775 -21227 -23741 -21200
rect -21589 -21209 -21572 -21175
rect -21346 -21209 -21126 -21175
rect -21092 -21209 -21076 -21175
rect -11715 -21206 -11646 -20803
rect -11278 -20864 -11277 -20830
rect -11156 -20864 -11140 -20830
rect -11602 -20921 -11312 -20883
rect -11602 -21054 -11575 -20921
rect -11522 -20929 -11312 -20921
rect -11522 -21054 -11384 -20929
rect -11602 -21059 -11384 -21054
rect -11339 -21059 -11312 -20929
rect -11278 -20960 -11262 -20926
rect -11142 -20960 -11140 -20926
rect -11278 -21056 -11277 -21022
rect -11156 -21056 -11140 -21022
rect -11602 -21104 -11312 -21059
rect -11090 -21118 -11068 -19995
rect -11022 -21118 -10999 -19995
rect -4888 -19999 -4854 -19983
rect -4888 -20106 -4854 -20090
rect -4816 -20154 -4782 -20138
rect -4720 -19948 -4686 -19932
rect -4720 -20160 -4686 -20142
rect -4624 -19942 -4590 -19932
rect -4624 -20154 -4590 -20138
rect -4528 -19948 -4494 -19932
rect -4366 -19948 -4332 -19932
rect -4366 -20140 -4332 -20124
rect -4278 -19948 -4244 -19932
rect -2100 -19942 -2066 -19926
rect -4176 -19967 -4142 -19951
rect -2172 -19990 -2138 -19974
rect -2172 -20097 -2138 -20081
rect -4176 -20115 -4142 -20099
rect -4278 -20140 -4244 -20124
rect -4528 -20160 -4494 -20142
rect -2100 -20148 -2066 -20138
rect -2004 -19938 -1970 -19920
rect -2004 -20148 -1970 -20132
rect -1908 -19942 -1874 -19926
rect -1908 -20148 -1874 -20138
rect -1812 -19938 -1778 -19920
rect 16159 -19935 16193 -19919
rect -1812 -20148 -1778 -20132
rect -1650 -19956 -1616 -19940
rect -1650 -20148 -1616 -20132
rect -1562 -19956 -1528 -19940
rect -1460 -19981 -1426 -19965
rect -1460 -20129 -1426 -20113
rect -1562 -20148 -1528 -20132
rect 7298 -20146 7403 -20143
rect 8246 -20146 8351 -20143
rect 9182 -20146 9287 -20143
rect 10113 -20146 10218 -20143
rect 11040 -20146 11145 -20143
rect 7298 -20162 7406 -20146
rect 7298 -20174 7372 -20162
rect -2069 -20225 -2052 -20191
rect -1826 -20225 -1606 -20191
rect -1572 -20225 -1556 -20191
rect -2069 -20241 -1556 -20225
rect -4785 -20295 -4272 -20279
rect -4785 -20329 -4768 -20295
rect -4542 -20329 -4322 -20295
rect -4288 -20329 -4272 -20295
rect -4816 -20382 -4782 -20372
rect -4888 -20439 -4854 -20423
rect -4888 -20546 -4854 -20530
rect -4816 -20594 -4782 -20578
rect -4720 -20388 -4686 -20372
rect -4720 -20600 -4686 -20582
rect -4624 -20382 -4590 -20372
rect -4624 -20594 -4590 -20578
rect -4528 -20388 -4494 -20372
rect -4366 -20388 -4332 -20372
rect -4366 -20580 -4332 -20564
rect -4278 -20388 -4244 -20372
rect -2100 -20382 -2066 -20366
rect -4176 -20407 -4142 -20391
rect -2172 -20430 -2138 -20414
rect -2172 -20537 -2138 -20521
rect -4176 -20555 -4142 -20539
rect -4278 -20580 -4244 -20564
rect -4528 -20600 -4494 -20582
rect -2100 -20588 -2066 -20578
rect -2004 -20378 -1970 -20360
rect -2004 -20588 -1970 -20572
rect -1908 -20382 -1874 -20366
rect -1908 -20588 -1874 -20578
rect -1812 -20378 -1778 -20360
rect -1812 -20588 -1778 -20572
rect -1650 -20396 -1616 -20380
rect -1650 -20588 -1616 -20572
rect -1562 -20396 -1528 -20380
rect -1460 -20421 -1426 -20405
rect -1460 -20569 -1426 -20553
rect -1562 -20588 -1528 -20572
rect -4785 -20674 -4272 -20658
rect -4785 -20708 -4768 -20674
rect -4542 -20708 -4322 -20674
rect -4288 -20708 -4272 -20674
rect -2069 -20665 -2052 -20631
rect -1826 -20665 -1606 -20631
rect -1572 -20665 -1556 -20631
rect -2069 -20681 -1556 -20665
rect -4816 -20761 -4782 -20751
rect -4888 -20818 -4854 -20802
rect -4888 -20925 -4854 -20909
rect -4816 -20973 -4782 -20957
rect -4720 -20767 -4686 -20751
rect -4720 -20979 -4686 -20961
rect -4624 -20761 -4590 -20751
rect -4624 -20973 -4590 -20957
rect -4528 -20767 -4494 -20751
rect -4366 -20767 -4332 -20751
rect -4366 -20959 -4332 -20943
rect -4278 -20767 -4244 -20751
rect -4176 -20786 -4142 -20770
rect -4176 -20934 -4142 -20918
rect 7333 -20925 7372 -20174
rect -4278 -20959 -4244 -20943
rect 7298 -20938 7372 -20925
rect 7298 -20954 7406 -20938
rect 7756 -20162 7790 -20146
rect 7756 -20954 7790 -20938
rect 8246 -20162 8354 -20146
rect 8246 -20174 8320 -20162
rect 8281 -20925 8320 -20174
rect 8246 -20938 8320 -20925
rect 8246 -20954 8354 -20938
rect 8704 -20162 8738 -20146
rect 8704 -20954 8738 -20938
rect 9182 -20162 9290 -20146
rect 9182 -20174 9256 -20162
rect 9217 -20925 9256 -20174
rect 9182 -20938 9256 -20925
rect 9182 -20954 9290 -20938
rect 9640 -20162 9674 -20146
rect 9640 -20954 9674 -20938
rect 10113 -20162 10221 -20146
rect 10113 -20174 10187 -20162
rect 10148 -20925 10187 -20174
rect 10113 -20938 10187 -20925
rect 10113 -20954 10221 -20938
rect 10571 -20162 10605 -20146
rect 10571 -20954 10605 -20938
rect 11040 -20162 11148 -20146
rect 11040 -20174 11114 -20162
rect 11075 -20925 11114 -20174
rect 11040 -20938 11114 -20925
rect 11040 -20954 11148 -20938
rect 11498 -20162 11532 -20146
rect 16159 -20177 16193 -20111
rect 16255 -19935 16289 -19919
rect 16255 -20127 16289 -20111
rect 16351 -19935 16385 -19919
rect 16351 -20177 16385 -20111
rect 16447 -19935 16481 -19919
rect 16447 -20127 16481 -20111
rect 16543 -19935 16577 -19919
rect 16543 -20177 16577 -20111
rect 16159 -20245 16577 -20177
rect 16159 -20358 16211 -20245
rect 16541 -20358 16577 -20245
rect 16159 -20406 16577 -20358
rect 11783 -20488 12203 -20468
rect 11783 -20539 11811 -20488
rect 12168 -20539 12203 -20488
rect 11783 -20558 12203 -20539
rect 11785 -20643 11819 -20558
rect 11785 -20891 11819 -20875
rect 11881 -20643 11915 -20627
rect 11881 -20891 11915 -20875
rect 11977 -20643 12011 -20558
rect 11977 -20891 12011 -20875
rect 12073 -20643 12107 -20627
rect 12073 -20891 12107 -20875
rect 12169 -20643 12203 -20558
rect 12169 -20891 12203 -20875
rect 12265 -20643 12299 -20627
rect 12265 -20891 12299 -20875
rect 12361 -20643 12395 -20627
rect 12361 -20891 12395 -20875
rect 12457 -20643 12491 -20627
rect 12457 -20891 12491 -20875
rect 12553 -20643 12587 -20627
rect 12553 -20891 12587 -20875
rect 12649 -20643 12683 -20627
rect 12649 -20891 12683 -20875
rect 12745 -20643 12779 -20627
rect 12970 -20709 12986 -20675
rect 13077 -20709 13093 -20675
rect 12745 -20891 12779 -20875
rect 12826 -20795 12876 -20778
rect 12919 -20781 12929 -20747
rect 13125 -20781 13141 -20747
rect 11498 -20954 11532 -20938
rect -4528 -20979 -4494 -20961
rect 12154 -20971 12170 -20937
rect 12204 -20971 12220 -20937
rect 12826 -21021 12842 -20795
rect 12919 -20877 12935 -20843
rect 13129 -20877 13147 -20843
rect 12919 -20973 12929 -20939
rect 13125 -20973 13141 -20939
rect -11278 -21152 -11262 -21118
rect -11156 -21152 -11140 -21118
rect -11090 -21159 -10999 -21118
rect 7298 -21090 7406 -21074
rect 7298 -21103 7372 -21090
rect -21589 -21225 -21076 -21209
rect -12318 -21240 -12302 -21206
rect -11776 -21240 -11262 -21206
rect -11156 -21240 -11140 -21206
rect -24128 -21299 -24010 -21265
rect -23975 -21299 -23959 -21265
rect -23893 -21299 -23877 -21265
rect -23842 -21299 -23826 -21265
rect -24399 -21353 -24383 -21319
rect -24187 -21353 -24177 -21319
rect -24134 -21349 -24099 -21333
rect -23893 -21357 -23826 -21299
rect -16027 -21277 -15993 -21261
rect -24099 -21383 -23826 -21357
rect -24134 -21400 -23826 -21383
rect -16099 -21325 -16065 -21309
rect -21618 -21406 -21584 -21390
rect -24508 -21449 -24461 -21433
rect -24399 -21449 -24389 -21415
rect -24193 -21449 -24177 -21415
rect -21690 -21454 -21656 -21438
rect -21690 -21561 -21656 -21545
rect -21618 -21612 -21584 -21602
rect -21522 -21402 -21488 -21384
rect -21522 -21612 -21488 -21596
rect -21426 -21406 -21392 -21390
rect -21426 -21612 -21392 -21602
rect -21330 -21402 -21296 -21384
rect -21330 -21612 -21296 -21596
rect -21168 -21420 -21134 -21404
rect -21168 -21612 -21134 -21596
rect -21080 -21420 -21046 -21404
rect -20978 -21445 -20944 -21429
rect -16099 -21432 -16065 -21416
rect -16027 -21483 -15993 -21473
rect -15931 -21273 -15897 -21255
rect -15931 -21483 -15897 -21467
rect -15835 -21277 -15801 -21261
rect -15835 -21483 -15801 -21473
rect -15739 -21273 -15705 -21255
rect -15739 -21483 -15705 -21467
rect -15577 -21291 -15543 -21275
rect -15577 -21483 -15543 -21467
rect -15489 -21291 -15455 -21275
rect -15387 -21316 -15353 -21300
rect -11565 -21431 -11559 -21389
rect -11497 -21431 -11491 -21389
rect -15387 -21464 -15353 -21448
rect -15489 -21483 -15455 -21467
rect -17681 -21545 -17665 -21511
rect -17433 -21545 -17417 -21511
rect -15996 -21560 -15979 -21526
rect -15753 -21560 -15533 -21526
rect -15499 -21560 -15483 -21526
rect -15996 -21576 -15483 -21560
rect -20978 -21593 -20944 -21577
rect -21080 -21612 -21046 -21596
rect -17681 -21641 -17665 -21607
rect -17433 -21641 -17417 -21607
rect -21587 -21689 -21570 -21655
rect -21344 -21689 -21124 -21655
rect -21090 -21689 -21074 -21655
rect -21587 -21705 -21074 -21689
rect -17681 -21737 -17665 -21703
rect -17433 -21737 -17417 -21703
rect -17681 -21833 -17665 -21799
rect -17433 -21833 -17417 -21799
rect 7333 -21854 7372 -21103
rect 7298 -21866 7372 -21854
rect 7298 -21882 7406 -21866
rect 7756 -21090 7790 -21074
rect 7756 -21882 7790 -21866
rect 8246 -21090 8354 -21074
rect 8246 -21103 8320 -21090
rect 8281 -21854 8320 -21103
rect 8246 -21866 8320 -21854
rect 8246 -21882 8354 -21866
rect 8704 -21090 8738 -21074
rect 8704 -21882 8738 -21866
rect 9182 -21090 9290 -21074
rect 9182 -21103 9256 -21090
rect 9217 -21854 9256 -21103
rect 9182 -21866 9256 -21854
rect 9182 -21882 9290 -21866
rect 9640 -21090 9674 -21074
rect 9640 -21882 9674 -21866
rect 10113 -21089 10221 -21073
rect 10113 -21102 10187 -21089
rect 10148 -21853 10187 -21102
rect 10113 -21865 10187 -21853
rect 10113 -21881 10221 -21865
rect 10571 -21089 10605 -21073
rect 10571 -21881 10605 -21865
rect 11040 -21090 11148 -21074
rect 11040 -21103 11114 -21090
rect 11075 -21854 11114 -21103
rect 11040 -21866 11114 -21854
rect -16928 -21895 -16844 -21883
rect 7298 -21885 7403 -21882
rect 8246 -21885 8351 -21882
rect 9182 -21885 9287 -21882
rect 10113 -21884 10218 -21881
rect 11040 -21882 11148 -21866
rect 11498 -21090 11532 -21074
rect 12297 -21076 12313 -21042
rect 12347 -21076 12363 -21042
rect 12169 -21132 12203 -21116
rect 12169 -21380 12203 -21308
rect 12265 -21132 12299 -21116
rect 12265 -21324 12299 -21308
rect 12361 -21132 12395 -21116
rect 12826 -21241 12876 -21021
rect 12919 -21069 12935 -21035
rect 13129 -21069 13147 -21035
rect 12919 -21231 12935 -21197
rect 13111 -21231 13127 -21197
rect 12826 -21275 12842 -21241
rect 12826 -21291 12876 -21275
rect 12361 -21380 12395 -21308
rect 12919 -21319 12935 -21285
rect 13111 -21319 13127 -21285
rect 12157 -21391 12407 -21380
rect 12157 -21452 12183 -21391
rect 12382 -21452 12407 -21391
rect 12938 -21421 12954 -21387
rect 13086 -21421 13102 -21387
rect 12157 -21464 12407 -21452
rect 11498 -21882 11532 -21866
rect 11040 -21885 11145 -21882
rect -17681 -21929 -17665 -21895
rect -17433 -21929 -17417 -21895
rect -17266 -21943 -17232 -21927
rect -17192 -21929 -17176 -21895
rect -17000 -21908 -16844 -21895
rect -17000 -21929 -16917 -21908
rect -17681 -22025 -17665 -21991
rect -17433 -22025 -17417 -21991
rect -17266 -21993 -17232 -21977
rect -17192 -22025 -17176 -21991
rect -17000 -22025 -16984 -21991
rect -17371 -22086 -17337 -22070
rect -17840 -22121 -17665 -22087
rect -17433 -22121 -17417 -22087
rect -16928 -22087 -16917 -21929
rect -17840 -22122 -17750 -22121
rect -24040 -22142 -24006 -22126
rect -24509 -22167 -24462 -22143
rect -24400 -22176 -24390 -22142
rect -24194 -22176 -24178 -22142
rect -24400 -22272 -24384 -22238
rect -24188 -22272 -24178 -22238
rect -24400 -22368 -24390 -22334
rect -24194 -22368 -24178 -22334
rect -24135 -22363 -24095 -22347
rect -24100 -22397 -24095 -22363
rect -24135 -22414 -24095 -22397
rect -24400 -22464 -24384 -22430
rect -24188 -22464 -24178 -22430
rect -24400 -22560 -24390 -22526
rect -24194 -22560 -24178 -22526
rect -24129 -22568 -24095 -22414
rect -24040 -22534 -24006 -22518
rect -23848 -22142 -23814 -22126
rect -23848 -22534 -23814 -22518
rect -23776 -22168 -23742 -22130
rect -23776 -22530 -23742 -22503
rect -17840 -22479 -17820 -22122
rect -17769 -22279 -17750 -22122
rect -17371 -22136 -17337 -22120
rect -17192 -22121 -17176 -22087
rect -17000 -22107 -16917 -22087
rect -16856 -22107 -16844 -21908
rect -17000 -22121 -16844 -22107
rect -16928 -22133 -16844 -22121
rect -17681 -22217 -17665 -22183
rect -17433 -22217 -17417 -22183
rect 7182 -22238 7198 -22204
rect 7232 -22238 7248 -22204
rect 7374 -22238 7390 -22204
rect 7424 -22238 7440 -22204
rect 7566 -22238 7582 -22204
rect 7616 -22238 7632 -22204
rect 7758 -22238 7774 -22204
rect 7808 -22238 7824 -22204
rect 8130 -22238 8146 -22204
rect 8180 -22238 8196 -22204
rect 8322 -22238 8338 -22204
rect 8372 -22238 8388 -22204
rect 8514 -22238 8530 -22204
rect 8564 -22238 8580 -22204
rect 8706 -22238 8722 -22204
rect 8756 -22238 8772 -22204
rect 9066 -22238 9082 -22204
rect 9116 -22238 9132 -22204
rect 9258 -22238 9274 -22204
rect 9308 -22238 9324 -22204
rect 9450 -22238 9466 -22204
rect 9500 -22238 9516 -22204
rect 9642 -22238 9658 -22204
rect 9692 -22238 9708 -22204
rect 9997 -22237 10013 -22203
rect 10047 -22237 10063 -22203
rect 10189 -22237 10205 -22203
rect 10239 -22237 10255 -22203
rect 10381 -22237 10397 -22203
rect 10431 -22237 10447 -22203
rect 10573 -22237 10589 -22203
rect 10623 -22237 10639 -22203
rect 10924 -22238 10940 -22204
rect 10974 -22238 10990 -22204
rect 11116 -22238 11132 -22204
rect 11166 -22238 11182 -22204
rect 11308 -22238 11324 -22204
rect 11358 -22238 11374 -22204
rect 11500 -22238 11516 -22204
rect 11550 -22238 11566 -22204
rect -17769 -22313 -17665 -22279
rect -17433 -22313 -17417 -22279
rect 7150 -22297 7184 -22281
rect 7246 -22292 7280 -22281
rect -17769 -22471 -17750 -22313
rect -17681 -22409 -17665 -22375
rect -17433 -22409 -17417 -22375
rect -17769 -22479 -17665 -22471
rect -17840 -22505 -17665 -22479
rect -17433 -22505 -17417 -22471
rect -12318 -22491 -12302 -22457
rect -11776 -22491 -11262 -22457
rect -11156 -22491 -11140 -22457
rect -17840 -22507 -17750 -22505
rect -24129 -22602 -24011 -22568
rect -23976 -22602 -23960 -22568
rect -23894 -22602 -23878 -22568
rect -23843 -22602 -23827 -22568
rect -24400 -22656 -24384 -22622
rect -24188 -22656 -24178 -22622
rect -24135 -22652 -24100 -22636
rect -23894 -22660 -23827 -22602
rect -24100 -22686 -23827 -22660
rect -24135 -22703 -23827 -22686
rect -12499 -22575 -12373 -22533
rect -24509 -22752 -24462 -22736
rect -24400 -22752 -24390 -22718
rect -24194 -22752 -24178 -22718
rect -17681 -22945 -17665 -22911
rect -17433 -22945 -17417 -22911
rect -17681 -23041 -17665 -23007
rect -17433 -23041 -17417 -23007
rect -17681 -23137 -17665 -23103
rect -17433 -23137 -17417 -23103
rect -17681 -23233 -17665 -23199
rect -17433 -23233 -17417 -23199
rect -16928 -23295 -16844 -23283
rect -17681 -23329 -17665 -23295
rect -17433 -23329 -17417 -23295
rect -17266 -23343 -17232 -23327
rect -17192 -23329 -17176 -23295
rect -17000 -23308 -16844 -23295
rect -17000 -23329 -16917 -23308
rect -17681 -23425 -17665 -23391
rect -17433 -23425 -17417 -23391
rect -17266 -23393 -17232 -23377
rect -17192 -23425 -17176 -23391
rect -17000 -23425 -16984 -23391
rect -24040 -23451 -24006 -23435
rect -24509 -23476 -24462 -23452
rect -24400 -23485 -24390 -23451
rect -24194 -23485 -24178 -23451
rect -24400 -23581 -24384 -23547
rect -24188 -23581 -24178 -23547
rect -24400 -23677 -24390 -23643
rect -24194 -23677 -24178 -23643
rect -24135 -23672 -24095 -23656
rect -24100 -23706 -24095 -23672
rect -24135 -23723 -24095 -23706
rect -24400 -23773 -24384 -23739
rect -24188 -23773 -24178 -23739
rect -24400 -23869 -24390 -23835
rect -24194 -23869 -24178 -23835
rect -24129 -23877 -24095 -23723
rect -24040 -23843 -24006 -23827
rect -23848 -23451 -23814 -23435
rect -23848 -23843 -23814 -23827
rect -23776 -23477 -23742 -23439
rect -17371 -23486 -17337 -23470
rect -23776 -23839 -23742 -23812
rect -17840 -23521 -17665 -23487
rect -17433 -23521 -17417 -23487
rect -16928 -23487 -16917 -23329
rect -17840 -23522 -17750 -23521
rect -24129 -23911 -24011 -23877
rect -23976 -23911 -23960 -23877
rect -23894 -23911 -23878 -23877
rect -23843 -23911 -23827 -23877
rect -17840 -23879 -17820 -23522
rect -17769 -23679 -17750 -23522
rect -17371 -23536 -17337 -23520
rect -17192 -23521 -17176 -23487
rect -17000 -23507 -16917 -23487
rect -16856 -23507 -16844 -23308
rect -17000 -23521 -16844 -23507
rect -16928 -23533 -16844 -23521
rect -17681 -23617 -17665 -23583
rect -17433 -23617 -17417 -23583
rect -17769 -23713 -17665 -23679
rect -17433 -23713 -17417 -23679
rect -12499 -23697 -12471 -22575
rect -12399 -23697 -12373 -22575
rect -12318 -22579 -12302 -22545
rect -11776 -22579 -11760 -22545
rect -12318 -22675 -12302 -22641
rect -11776 -22675 -11760 -22641
rect -12318 -22771 -12302 -22737
rect -11776 -22771 -11760 -22737
rect -12318 -22867 -12302 -22833
rect -11776 -22867 -11760 -22833
rect -11718 -22882 -11641 -22491
rect -11433 -22546 -11337 -22531
rect -11433 -22611 -11411 -22546
rect -11356 -22611 -11337 -22546
rect -11278 -22579 -11262 -22545
rect -11156 -22579 -11140 -22545
rect -11090 -22574 -10999 -22536
rect -11600 -22713 -11494 -22695
rect -11600 -22793 -11582 -22713
rect -11514 -22793 -11494 -22713
rect -11600 -22810 -11494 -22793
rect -11718 -22902 -11501 -22882
rect -12318 -22963 -12302 -22929
rect -11776 -22963 -11760 -22929
rect -12318 -23059 -12302 -23025
rect -11776 -23059 -11760 -23025
rect -11718 -23032 -11700 -22902
rect -11655 -22913 -11501 -22902
rect -11655 -23027 -11583 -22913
rect -11530 -23027 -11501 -22913
rect -11655 -23032 -11501 -23027
rect -11718 -23059 -11501 -23032
rect -11433 -23105 -11337 -22611
rect -11278 -22675 -11277 -22641
rect -11156 -22675 -11140 -22641
rect -11278 -22771 -11262 -22737
rect -11142 -22771 -11140 -22737
rect -11278 -22867 -11277 -22833
rect -11156 -22867 -11140 -22833
rect -11278 -22963 -11262 -22929
rect -11142 -22963 -11140 -22929
rect -11278 -23059 -11277 -23025
rect -11156 -23059 -11140 -23025
rect -11733 -23121 -11303 -23105
rect -12318 -23155 -12302 -23121
rect -11776 -23155 -11262 -23121
rect -11142 -23155 -11140 -23121
rect -11733 -23171 -11303 -23155
rect -12318 -23251 -12302 -23217
rect -11776 -23251 -11760 -23217
rect -11715 -23225 -11314 -23217
rect -11715 -23233 -11376 -23225
rect -12318 -23347 -12302 -23313
rect -11776 -23347 -11760 -23313
rect -11715 -23363 -11705 -23233
rect -11660 -23355 -11376 -23233
rect -11331 -23355 -11314 -23225
rect -11278 -23251 -11276 -23217
rect -11156 -23251 -11140 -23217
rect -11278 -23347 -11262 -23313
rect -11142 -23347 -11140 -23313
rect -11660 -23363 -11314 -23355
rect -11715 -23382 -11314 -23363
rect -12318 -23443 -12302 -23409
rect -11776 -23443 -11760 -23409
rect -12318 -23539 -12302 -23505
rect -11776 -23539 -11760 -23505
rect -12318 -23635 -12302 -23601
rect -11776 -23635 -11760 -23601
rect -17769 -23871 -17750 -23713
rect -12499 -23743 -12373 -23697
rect -12318 -23731 -12302 -23697
rect -11776 -23731 -11760 -23697
rect -17681 -23809 -17665 -23775
rect -17433 -23809 -17417 -23775
rect -11715 -23785 -11646 -23382
rect -11278 -23443 -11277 -23409
rect -11156 -23443 -11140 -23409
rect -11602 -23500 -11312 -23462
rect -11602 -23633 -11575 -23500
rect -11522 -23508 -11312 -23500
rect -11522 -23633 -11384 -23508
rect -11602 -23638 -11384 -23633
rect -11339 -23638 -11312 -23508
rect -11278 -23539 -11262 -23505
rect -11142 -23539 -11140 -23505
rect -11278 -23635 -11277 -23601
rect -11156 -23635 -11140 -23601
rect -11602 -23683 -11312 -23638
rect -11090 -23697 -11068 -22574
rect -11022 -23697 -10999 -22574
rect 7150 -22611 7184 -22595
rect 7246 -22611 7280 -22595
rect 7342 -22297 7376 -22281
rect 7342 -22611 7376 -22595
rect 7438 -22292 7472 -22281
rect 7534 -22297 7568 -22281
rect 7438 -22611 7472 -22595
rect 7534 -22611 7568 -22595
rect 7630 -22292 7664 -22281
rect 7726 -22297 7760 -22281
rect 7630 -22611 7664 -22595
rect 7726 -22611 7760 -22595
rect 7822 -22292 7856 -22281
rect 7918 -22297 7952 -22281
rect 7822 -22611 7856 -22595
rect 7918 -22611 7952 -22595
rect 8098 -22297 8132 -22281
rect 8194 -22292 8228 -22281
rect 8098 -22611 8132 -22595
rect 8194 -22611 8228 -22595
rect 8290 -22297 8324 -22281
rect 8290 -22611 8324 -22595
rect 8386 -22292 8420 -22281
rect 8482 -22297 8516 -22281
rect 8386 -22611 8420 -22595
rect 8482 -22611 8516 -22595
rect 8578 -22292 8612 -22281
rect 8674 -22297 8708 -22281
rect 8578 -22611 8612 -22595
rect 8674 -22611 8708 -22595
rect 8770 -22292 8804 -22281
rect 8866 -22297 8900 -22281
rect 8770 -22611 8804 -22595
rect 8866 -22611 8900 -22595
rect 9034 -22297 9068 -22281
rect 9130 -22292 9164 -22281
rect 9034 -22611 9068 -22595
rect 9130 -22611 9164 -22595
rect 9226 -22297 9260 -22281
rect 9226 -22611 9260 -22595
rect 9322 -22292 9356 -22281
rect 9418 -22297 9452 -22281
rect 9322 -22611 9356 -22595
rect 9418 -22611 9452 -22595
rect 9514 -22292 9548 -22281
rect 9610 -22297 9644 -22281
rect 9514 -22611 9548 -22595
rect 9610 -22611 9644 -22595
rect 9706 -22292 9740 -22281
rect 9802 -22297 9836 -22281
rect 9706 -22611 9740 -22595
rect 9802 -22611 9836 -22595
rect 9965 -22296 9999 -22280
rect 10061 -22291 10095 -22280
rect 9965 -22610 9999 -22594
rect 10061 -22610 10095 -22594
rect 10157 -22296 10191 -22280
rect 10157 -22610 10191 -22594
rect 10253 -22291 10287 -22280
rect 10349 -22296 10383 -22280
rect 10253 -22610 10287 -22594
rect 10349 -22610 10383 -22594
rect 10445 -22291 10479 -22280
rect 10541 -22296 10575 -22280
rect 10445 -22610 10479 -22594
rect 10541 -22610 10575 -22594
rect 10637 -22291 10671 -22280
rect 10733 -22296 10767 -22280
rect 10637 -22610 10671 -22594
rect 10733 -22610 10767 -22594
rect 10892 -22297 10926 -22281
rect 10988 -22292 11022 -22281
rect 10892 -22611 10926 -22595
rect 10988 -22611 11022 -22595
rect 11084 -22297 11118 -22281
rect 11084 -22611 11118 -22595
rect 11180 -22292 11214 -22281
rect 11276 -22297 11310 -22281
rect 11180 -22611 11214 -22595
rect 11276 -22611 11310 -22595
rect 11372 -22292 11406 -22281
rect 11468 -22297 11502 -22281
rect 11372 -22611 11406 -22595
rect 11468 -22611 11502 -22595
rect 11564 -22292 11598 -22281
rect 11660 -22297 11694 -22281
rect 11564 -22611 11598 -22595
rect 11660 -22611 11694 -22595
rect 7373 -22699 7389 -22664
rect 7677 -22699 7703 -22664
rect 8321 -22699 8337 -22664
rect 8625 -22699 8651 -22664
rect 9257 -22699 9273 -22664
rect 9561 -22699 9587 -22664
rect 10188 -22698 10204 -22663
rect 10492 -22698 10518 -22663
rect 11115 -22699 11131 -22664
rect 11419 -22699 11445 -22664
rect 5705 -23219 5721 -23185
rect 5812 -23219 5828 -23185
rect 6145 -23219 6161 -23185
rect 6252 -23219 6268 -23185
rect 6585 -23219 6601 -23185
rect 6692 -23219 6708 -23185
rect -11278 -23731 -11262 -23697
rect -11156 -23731 -11140 -23697
rect -11090 -23738 -10999 -23697
rect 5561 -23305 5611 -23288
rect 5654 -23291 5664 -23257
rect 5860 -23291 5876 -23257
rect 5561 -23531 5577 -23305
rect 6001 -23305 6051 -23288
rect 6094 -23291 6104 -23257
rect 6300 -23291 6316 -23257
rect 5654 -23387 5670 -23353
rect 5864 -23387 5882 -23353
rect 5654 -23483 5664 -23449
rect 5860 -23483 5876 -23449
rect 5561 -23751 5611 -23531
rect 6001 -23531 6017 -23305
rect 6441 -23305 6491 -23288
rect 6534 -23291 6544 -23257
rect 6740 -23291 6756 -23257
rect 6094 -23387 6110 -23353
rect 6304 -23387 6322 -23353
rect 6094 -23483 6104 -23449
rect 6300 -23483 6316 -23449
rect 5654 -23579 5670 -23545
rect 5864 -23579 5882 -23545
rect 5654 -23741 5670 -23707
rect 5846 -23741 5862 -23707
rect 5561 -23785 5577 -23751
rect -12318 -23819 -12302 -23785
rect -11776 -23819 -11262 -23785
rect -11156 -23819 -11140 -23785
rect 5561 -23801 5611 -23785
rect 6001 -23751 6051 -23531
rect 6441 -23531 6457 -23305
rect 6534 -23387 6550 -23353
rect 6744 -23387 6762 -23353
rect 6534 -23483 6544 -23449
rect 6740 -23483 6756 -23449
rect 6094 -23579 6110 -23545
rect 6304 -23579 6322 -23545
rect 6094 -23741 6110 -23707
rect 6286 -23741 6302 -23707
rect 6001 -23785 6017 -23751
rect 5654 -23829 5670 -23795
rect 5846 -23829 5862 -23795
rect 6001 -23801 6051 -23785
rect 6441 -23751 6491 -23531
rect 6534 -23579 6550 -23545
rect 6744 -23579 6762 -23545
rect 6534 -23741 6550 -23707
rect 6726 -23741 6742 -23707
rect 6441 -23785 6457 -23751
rect 6094 -23829 6110 -23795
rect 6286 -23829 6302 -23795
rect 6441 -23801 6491 -23785
rect 6534 -23829 6550 -23795
rect 6726 -23829 6742 -23795
rect -17769 -23879 -17665 -23871
rect -17840 -23905 -17665 -23879
rect -17433 -23905 -17417 -23871
rect 7373 -23892 7389 -23857
rect 7677 -23892 7703 -23857
rect 8321 -23892 8337 -23857
rect 8625 -23892 8651 -23857
rect 9257 -23892 9273 -23857
rect 9561 -23892 9587 -23857
rect 10188 -23892 10204 -23857
rect 10492 -23892 10518 -23857
rect 11115 -23892 11131 -23857
rect 11419 -23892 11445 -23857
rect -17840 -23907 -17750 -23905
rect -24400 -23965 -24384 -23931
rect -24188 -23965 -24178 -23931
rect -24135 -23961 -24100 -23945
rect -23894 -23969 -23827 -23911
rect 5673 -23931 5689 -23897
rect 5821 -23931 5837 -23897
rect 6113 -23931 6129 -23897
rect 6261 -23931 6277 -23897
rect 6553 -23931 6569 -23897
rect 6701 -23931 6717 -23897
rect -24100 -23995 -23827 -23969
rect 7150 -23961 7184 -23945
rect -24135 -24012 -23827 -23995
rect -11569 -24019 -11563 -23970
rect -11494 -24019 -11488 -23970
rect -24509 -24061 -24462 -24045
rect -24400 -24061 -24390 -24027
rect -24194 -24061 -24178 -24027
rect 7246 -23961 7280 -23945
rect 7150 -24275 7184 -24259
rect 7246 -24275 7280 -24264
rect 7342 -23961 7376 -23945
rect 7342 -24275 7376 -24259
rect 7438 -23961 7472 -23945
rect 7534 -23961 7568 -23945
rect 7438 -24275 7472 -24264
rect 7534 -24275 7568 -24259
rect 7630 -23961 7664 -23945
rect 7726 -23961 7760 -23945
rect 7630 -24275 7664 -24264
rect 7726 -24275 7760 -24259
rect 7822 -23961 7856 -23945
rect 7918 -23961 7952 -23945
rect 7822 -24275 7856 -24264
rect 7918 -24275 7952 -24259
rect 8098 -23961 8132 -23945
rect 8194 -23961 8228 -23945
rect 8098 -24275 8132 -24259
rect 8194 -24275 8228 -24264
rect 8290 -23961 8324 -23945
rect 8290 -24275 8324 -24259
rect 8386 -23961 8420 -23945
rect 8482 -23961 8516 -23945
rect 8386 -24275 8420 -24264
rect 8482 -24275 8516 -24259
rect 8578 -23961 8612 -23945
rect 8674 -23961 8708 -23945
rect 8578 -24275 8612 -24264
rect 8674 -24275 8708 -24259
rect 8770 -23961 8804 -23945
rect 8866 -23961 8900 -23945
rect 8770 -24275 8804 -24264
rect 8866 -24275 8900 -24259
rect 9034 -23961 9068 -23945
rect 9130 -23961 9164 -23945
rect 9034 -24275 9068 -24259
rect 9130 -24275 9164 -24264
rect 9226 -23961 9260 -23945
rect 9226 -24275 9260 -24259
rect 9322 -23961 9356 -23945
rect 9418 -23961 9452 -23945
rect 9322 -24275 9356 -24264
rect 9418 -24275 9452 -24259
rect 9514 -23961 9548 -23945
rect 9610 -23961 9644 -23945
rect 9514 -24275 9548 -24264
rect 9610 -24275 9644 -24259
rect 9706 -23961 9740 -23945
rect 9802 -23961 9836 -23945
rect 9706 -24275 9740 -24264
rect 9802 -24275 9836 -24259
rect 9965 -23961 9999 -23945
rect 10061 -23961 10095 -23945
rect 9965 -24275 9999 -24259
rect 10061 -24275 10095 -24264
rect 10157 -23961 10191 -23945
rect 10157 -24275 10191 -24259
rect 10253 -23961 10287 -23945
rect 10349 -23961 10383 -23945
rect 10253 -24275 10287 -24264
rect 10349 -24275 10383 -24259
rect 10445 -23961 10479 -23945
rect 10541 -23961 10575 -23945
rect 10445 -24275 10479 -24264
rect 10541 -24275 10575 -24259
rect 10637 -23961 10671 -23945
rect 10733 -23961 10767 -23945
rect 10637 -24275 10671 -24264
rect 10733 -24275 10767 -24259
rect 10892 -23961 10926 -23945
rect 10988 -23961 11022 -23945
rect 10892 -24275 10926 -24259
rect 10988 -24275 11022 -24264
rect 11084 -23961 11118 -23945
rect 11084 -24275 11118 -24259
rect 11180 -23961 11214 -23945
rect 11276 -23961 11310 -23945
rect 11180 -24275 11214 -24264
rect 11276 -24275 11310 -24259
rect 11372 -23961 11406 -23945
rect 11468 -23961 11502 -23945
rect 11372 -24275 11406 -24264
rect 11468 -24275 11502 -24259
rect 11564 -23961 11598 -23945
rect 11660 -23961 11694 -23945
rect 11564 -24275 11598 -24264
rect 11660 -24275 11694 -24259
rect -17681 -24345 -17665 -24311
rect -17433 -24345 -17417 -24311
rect 7182 -24352 7198 -24318
rect 7232 -24352 7248 -24318
rect 7374 -24352 7390 -24318
rect 7424 -24352 7440 -24318
rect 7566 -24352 7582 -24318
rect 7616 -24352 7632 -24318
rect 7758 -24352 7774 -24318
rect 7808 -24352 7824 -24318
rect 8130 -24352 8146 -24318
rect 8180 -24352 8196 -24318
rect 8322 -24352 8338 -24318
rect 8372 -24352 8388 -24318
rect 8514 -24352 8530 -24318
rect 8564 -24352 8580 -24318
rect 8706 -24352 8722 -24318
rect 8756 -24352 8772 -24318
rect 9066 -24352 9082 -24318
rect 9116 -24352 9132 -24318
rect 9258 -24352 9274 -24318
rect 9308 -24352 9324 -24318
rect 9450 -24352 9466 -24318
rect 9500 -24352 9516 -24318
rect 9642 -24352 9658 -24318
rect 9692 -24352 9708 -24318
rect 9997 -24352 10013 -24318
rect 10047 -24352 10063 -24318
rect 10189 -24352 10205 -24318
rect 10239 -24352 10255 -24318
rect 10381 -24352 10397 -24318
rect 10431 -24352 10447 -24318
rect 10573 -24352 10589 -24318
rect 10623 -24352 10639 -24318
rect 10924 -24352 10940 -24318
rect 10974 -24352 10990 -24318
rect 11116 -24352 11132 -24318
rect 11166 -24352 11182 -24318
rect 11308 -24352 11324 -24318
rect 11358 -24352 11374 -24318
rect 11500 -24352 11516 -24318
rect 11550 -24352 11566 -24318
rect -17681 -24441 -17665 -24407
rect -17433 -24441 -17417 -24407
rect -17681 -24537 -17665 -24503
rect -17433 -24537 -17417 -24503
rect -17681 -24633 -17665 -24599
rect -17433 -24633 -17417 -24599
rect 7298 -24674 7403 -24671
rect 8246 -24674 8351 -24671
rect 9182 -24674 9287 -24671
rect 10113 -24674 10218 -24671
rect 11040 -24674 11145 -24671
rect -16928 -24695 -16844 -24683
rect -17681 -24729 -17665 -24695
rect -17433 -24729 -17417 -24695
rect -17266 -24743 -17232 -24727
rect -17192 -24729 -17176 -24695
rect -17000 -24708 -16844 -24695
rect -17000 -24729 -16917 -24708
rect -17681 -24825 -17665 -24791
rect -17433 -24825 -17417 -24791
rect -17266 -24793 -17232 -24777
rect -17192 -24825 -17176 -24791
rect -17000 -24825 -16984 -24791
rect -17371 -24886 -17337 -24870
rect -17840 -24921 -17665 -24887
rect -17433 -24921 -17417 -24887
rect -16928 -24887 -16917 -24729
rect -17840 -24922 -17750 -24921
rect -17840 -25279 -17820 -24922
rect -17769 -25079 -17750 -24922
rect -17371 -24936 -17337 -24920
rect -17192 -24921 -17176 -24887
rect -17000 -24907 -16917 -24887
rect -16856 -24907 -16844 -24708
rect -17000 -24921 -16844 -24907
rect -16928 -24933 -16844 -24921
rect 7298 -24690 7406 -24674
rect 7298 -24702 7372 -24690
rect -17681 -25017 -17665 -24983
rect -17433 -25017 -17417 -24983
rect -17769 -25113 -17665 -25079
rect -17433 -25113 -17417 -25079
rect -17769 -25271 -17750 -25113
rect -17681 -25209 -17665 -25175
rect -17433 -25209 -17417 -25175
rect -12318 -25259 -12302 -25225
rect -11776 -25259 -11262 -25225
rect -11156 -25259 -11140 -25225
rect -17769 -25279 -17665 -25271
rect -17840 -25305 -17665 -25279
rect -17433 -25305 -17417 -25271
rect -17840 -25307 -17750 -25305
rect -12499 -25343 -12373 -25301
rect -12499 -26465 -12471 -25343
rect -12399 -26465 -12373 -25343
rect -12318 -25347 -12302 -25313
rect -11776 -25347 -11760 -25313
rect -12318 -25443 -12302 -25409
rect -11776 -25443 -11760 -25409
rect -12318 -25539 -12302 -25505
rect -11776 -25539 -11760 -25505
rect -12318 -25635 -12302 -25601
rect -11776 -25635 -11760 -25601
rect -11718 -25650 -11641 -25259
rect -11433 -25314 -11337 -25299
rect -11433 -25379 -11411 -25314
rect -11356 -25379 -11337 -25314
rect -11278 -25347 -11262 -25313
rect -11156 -25347 -11140 -25313
rect -11090 -25342 -10999 -25304
rect -11600 -25481 -11494 -25463
rect -11600 -25561 -11582 -25481
rect -11514 -25561 -11494 -25481
rect -11600 -25578 -11494 -25561
rect -11718 -25670 -11501 -25650
rect -12318 -25731 -12302 -25697
rect -11776 -25731 -11760 -25697
rect -12318 -25827 -12302 -25793
rect -11776 -25827 -11760 -25793
rect -11718 -25800 -11700 -25670
rect -11655 -25681 -11501 -25670
rect -11655 -25795 -11583 -25681
rect -11530 -25795 -11501 -25681
rect -11655 -25800 -11501 -25795
rect -11718 -25827 -11501 -25800
rect -11433 -25873 -11337 -25379
rect -11278 -25443 -11277 -25409
rect -11156 -25443 -11140 -25409
rect -11278 -25539 -11262 -25505
rect -11142 -25539 -11140 -25505
rect -11278 -25635 -11277 -25601
rect -11156 -25635 -11140 -25601
rect -11278 -25731 -11262 -25697
rect -11142 -25731 -11140 -25697
rect -11278 -25827 -11277 -25793
rect -11156 -25827 -11140 -25793
rect -11733 -25889 -11303 -25873
rect -12318 -25923 -12302 -25889
rect -11776 -25923 -11262 -25889
rect -11142 -25923 -11140 -25889
rect -11733 -25939 -11303 -25923
rect -12318 -26019 -12302 -25985
rect -11776 -26019 -11760 -25985
rect -11715 -25993 -11314 -25985
rect -11715 -26001 -11376 -25993
rect -12318 -26115 -12302 -26081
rect -11776 -26115 -11760 -26081
rect -11715 -26131 -11705 -26001
rect -11660 -26123 -11376 -26001
rect -11331 -26123 -11314 -25993
rect -11278 -26019 -11276 -25985
rect -11156 -26019 -11140 -25985
rect -11278 -26115 -11262 -26081
rect -11142 -26115 -11140 -26081
rect -11660 -26131 -11314 -26123
rect -11715 -26150 -11314 -26131
rect -12318 -26211 -12302 -26177
rect -11776 -26211 -11760 -26177
rect -12318 -26307 -12302 -26273
rect -11776 -26307 -11760 -26273
rect -12318 -26403 -12302 -26369
rect -11776 -26403 -11760 -26369
rect -12499 -26511 -12373 -26465
rect -12318 -26499 -12302 -26465
rect -11776 -26499 -11760 -26465
rect -11715 -26553 -11646 -26150
rect -11278 -26211 -11277 -26177
rect -11156 -26211 -11140 -26177
rect -11602 -26268 -11312 -26230
rect -11602 -26401 -11575 -26268
rect -11522 -26276 -11312 -26268
rect -11522 -26401 -11384 -26276
rect -11602 -26406 -11384 -26401
rect -11339 -26406 -11312 -26276
rect -11278 -26307 -11262 -26273
rect -11142 -26307 -11140 -26273
rect -11278 -26403 -11277 -26369
rect -11156 -26403 -11140 -26369
rect -11602 -26451 -11312 -26406
rect -11090 -26465 -11068 -25342
rect -11022 -26465 -10999 -25342
rect 7333 -25453 7372 -24702
rect 7298 -25466 7372 -25453
rect 7298 -25482 7406 -25466
rect 7756 -24690 7790 -24674
rect 7756 -25482 7790 -25466
rect 8246 -24690 8354 -24674
rect 8246 -24702 8320 -24690
rect 8281 -25453 8320 -24702
rect 8246 -25466 8320 -25453
rect 8246 -25482 8354 -25466
rect 8704 -24690 8738 -24674
rect 8704 -25482 8738 -25466
rect 9182 -24690 9290 -24674
rect 9182 -24702 9256 -24690
rect 9217 -25453 9256 -24702
rect 9182 -25466 9256 -25453
rect 9182 -25482 9290 -25466
rect 9640 -24690 9674 -24674
rect 9640 -25482 9674 -25466
rect 10113 -24690 10221 -24674
rect 10113 -24702 10187 -24690
rect 10148 -25453 10187 -24702
rect 10113 -25466 10187 -25453
rect 10113 -25482 10221 -25466
rect 10571 -24690 10605 -24674
rect 10571 -25482 10605 -25466
rect 11040 -24690 11148 -24674
rect 11040 -24702 11114 -24690
rect 11075 -25453 11114 -24702
rect 11040 -25466 11114 -25453
rect 11040 -25482 11148 -25466
rect 11498 -24690 11532 -24674
rect 11783 -25016 12203 -24996
rect 11783 -25067 11811 -25016
rect 12168 -25067 12203 -25016
rect 11783 -25086 12203 -25067
rect 11785 -25171 11819 -25086
rect 11785 -25419 11819 -25403
rect 11881 -25171 11915 -25155
rect 11881 -25419 11915 -25403
rect 11977 -25171 12011 -25086
rect 11977 -25419 12011 -25403
rect 12073 -25171 12107 -25155
rect 12073 -25419 12107 -25403
rect 12169 -25171 12203 -25086
rect 12169 -25419 12203 -25403
rect 12265 -25171 12299 -25155
rect 12265 -25419 12299 -25403
rect 12361 -25171 12395 -25155
rect 12361 -25419 12395 -25403
rect 12457 -25171 12491 -25155
rect 12457 -25419 12491 -25403
rect 12553 -25171 12587 -25155
rect 12553 -25419 12587 -25403
rect 12649 -25171 12683 -25155
rect 12649 -25419 12683 -25403
rect 12745 -25171 12779 -25155
rect 12970 -25237 12986 -25203
rect 13077 -25237 13093 -25203
rect 12745 -25419 12779 -25403
rect 12826 -25323 12876 -25306
rect 12919 -25309 12929 -25275
rect 13125 -25309 13141 -25275
rect 11498 -25482 11532 -25466
rect 12154 -25499 12170 -25465
rect 12204 -25499 12220 -25465
rect 12826 -25549 12842 -25323
rect 12919 -25405 12935 -25371
rect 13129 -25405 13147 -25371
rect 12919 -25501 12929 -25467
rect 13125 -25501 13141 -25467
rect 7298 -25618 7406 -25602
rect 7298 -25631 7372 -25618
rect 7333 -26382 7372 -25631
rect 7298 -26394 7372 -26382
rect 7298 -26410 7406 -26394
rect 7756 -25618 7790 -25602
rect 7756 -26410 7790 -26394
rect 8246 -25618 8354 -25602
rect 8246 -25631 8320 -25618
rect 8281 -26382 8320 -25631
rect 8246 -26394 8320 -26382
rect 8246 -26410 8354 -26394
rect 8704 -25618 8738 -25602
rect 8704 -26410 8738 -26394
rect 9182 -25618 9290 -25602
rect 9182 -25631 9256 -25618
rect 9217 -26382 9256 -25631
rect 9182 -26394 9256 -26382
rect 9182 -26410 9290 -26394
rect 9640 -25618 9674 -25602
rect 9640 -26410 9674 -26394
rect 10113 -25617 10221 -25601
rect 10113 -25630 10187 -25617
rect 10148 -26381 10187 -25630
rect 10113 -26393 10187 -26381
rect 10113 -26409 10221 -26393
rect 10571 -25617 10605 -25601
rect 10571 -26409 10605 -26393
rect 11040 -25618 11148 -25602
rect 11040 -25631 11114 -25618
rect 11075 -26382 11114 -25631
rect 11040 -26394 11114 -26382
rect 7298 -26413 7403 -26410
rect 8246 -26413 8351 -26410
rect 9182 -26413 9287 -26410
rect 10113 -26412 10218 -26409
rect 11040 -26410 11148 -26394
rect 11498 -25618 11532 -25602
rect 12297 -25604 12313 -25570
rect 12347 -25604 12363 -25570
rect 12169 -25660 12203 -25644
rect 12169 -25908 12203 -25836
rect 12265 -25660 12299 -25644
rect 12265 -25852 12299 -25836
rect 12361 -25660 12395 -25644
rect 12826 -25769 12876 -25549
rect 12919 -25597 12935 -25563
rect 13129 -25597 13147 -25563
rect 12919 -25759 12935 -25725
rect 13111 -25759 13127 -25725
rect 12826 -25803 12842 -25769
rect 12826 -25819 12876 -25803
rect 12361 -25908 12395 -25836
rect 12919 -25847 12935 -25813
rect 13111 -25847 13127 -25813
rect 12157 -25919 12407 -25908
rect 12157 -25980 12183 -25919
rect 12382 -25980 12407 -25919
rect 12938 -25949 12954 -25915
rect 13086 -25949 13102 -25915
rect 12157 -25992 12407 -25980
rect 11498 -26410 11532 -26394
rect 11040 -26413 11145 -26410
rect -11278 -26499 -11262 -26465
rect -11156 -26499 -11140 -26465
rect -11090 -26506 -10999 -26465
rect -12318 -26587 -12302 -26553
rect -11776 -26587 -11262 -26553
rect -11156 -26587 -11140 -26553
rect -11570 -26810 -11564 -26758
rect -11492 -26810 -11486 -26758
rect 7182 -26766 7198 -26732
rect 7232 -26766 7248 -26732
rect 7374 -26766 7390 -26732
rect 7424 -26766 7440 -26732
rect 7566 -26766 7582 -26732
rect 7616 -26766 7632 -26732
rect 7758 -26766 7774 -26732
rect 7808 -26766 7824 -26732
rect 8130 -26766 8146 -26732
rect 8180 -26766 8196 -26732
rect 8322 -26766 8338 -26732
rect 8372 -26766 8388 -26732
rect 8514 -26766 8530 -26732
rect 8564 -26766 8580 -26732
rect 8706 -26766 8722 -26732
rect 8756 -26766 8772 -26732
rect 9066 -26766 9082 -26732
rect 9116 -26766 9132 -26732
rect 9258 -26766 9274 -26732
rect 9308 -26766 9324 -26732
rect 9450 -26766 9466 -26732
rect 9500 -26766 9516 -26732
rect 9642 -26766 9658 -26732
rect 9692 -26766 9708 -26732
rect 9997 -26765 10013 -26731
rect 10047 -26765 10063 -26731
rect 10189 -26765 10205 -26731
rect 10239 -26765 10255 -26731
rect 10381 -26765 10397 -26731
rect 10431 -26765 10447 -26731
rect 10573 -26765 10589 -26731
rect 10623 -26765 10639 -26731
rect 10924 -26766 10940 -26732
rect 10974 -26766 10990 -26732
rect 11116 -26766 11132 -26732
rect 11166 -26766 11182 -26732
rect 11308 -26766 11324 -26732
rect 11358 -26766 11374 -26732
rect 11500 -26766 11516 -26732
rect 11550 -26766 11566 -26732
rect 7150 -26825 7184 -26809
rect 7246 -26820 7280 -26809
rect 7150 -27139 7184 -27123
rect 7246 -27139 7280 -27123
rect 7342 -26825 7376 -26809
rect 7342 -27139 7376 -27123
rect 7438 -26820 7472 -26809
rect 7534 -26825 7568 -26809
rect 7438 -27139 7472 -27123
rect 7534 -27139 7568 -27123
rect 7630 -26820 7664 -26809
rect 7726 -26825 7760 -26809
rect 7630 -27139 7664 -27123
rect 7726 -27139 7760 -27123
rect 7822 -26820 7856 -26809
rect 7918 -26825 7952 -26809
rect 7822 -27139 7856 -27123
rect 7918 -27139 7952 -27123
rect 8098 -26825 8132 -26809
rect 8194 -26820 8228 -26809
rect 8098 -27139 8132 -27123
rect 8194 -27139 8228 -27123
rect 8290 -26825 8324 -26809
rect 8290 -27139 8324 -27123
rect 8386 -26820 8420 -26809
rect 8482 -26825 8516 -26809
rect 8386 -27139 8420 -27123
rect 8482 -27139 8516 -27123
rect 8578 -26820 8612 -26809
rect 8674 -26825 8708 -26809
rect 8578 -27139 8612 -27123
rect 8674 -27139 8708 -27123
rect 8770 -26820 8804 -26809
rect 8866 -26825 8900 -26809
rect 8770 -27139 8804 -27123
rect 8866 -27139 8900 -27123
rect 9034 -26825 9068 -26809
rect 9130 -26820 9164 -26809
rect 9034 -27139 9068 -27123
rect 9130 -27139 9164 -27123
rect 9226 -26825 9260 -26809
rect 9226 -27139 9260 -27123
rect 9322 -26820 9356 -26809
rect 9418 -26825 9452 -26809
rect 9322 -27139 9356 -27123
rect 9418 -27139 9452 -27123
rect 9514 -26820 9548 -26809
rect 9610 -26825 9644 -26809
rect 9514 -27139 9548 -27123
rect 9610 -27139 9644 -27123
rect 9706 -26820 9740 -26809
rect 9802 -26825 9836 -26809
rect 9706 -27139 9740 -27123
rect 9802 -27139 9836 -27123
rect 9965 -26824 9999 -26808
rect 10061 -26819 10095 -26808
rect 9965 -27138 9999 -27122
rect 10061 -27138 10095 -27122
rect 10157 -26824 10191 -26808
rect 10157 -27138 10191 -27122
rect 10253 -26819 10287 -26808
rect 10349 -26824 10383 -26808
rect 10253 -27138 10287 -27122
rect 10349 -27138 10383 -27122
rect 10445 -26819 10479 -26808
rect 10541 -26824 10575 -26808
rect 10445 -27138 10479 -27122
rect 10541 -27138 10575 -27122
rect 10637 -26819 10671 -26808
rect 10733 -26824 10767 -26808
rect 10637 -27138 10671 -27122
rect 10733 -27138 10767 -27122
rect 10892 -26825 10926 -26809
rect 10988 -26820 11022 -26809
rect 10892 -27139 10926 -27123
rect 10988 -27139 11022 -27123
rect 11084 -26825 11118 -26809
rect 11084 -27139 11118 -27123
rect 11180 -26820 11214 -26809
rect 11276 -26825 11310 -26809
rect 11180 -27139 11214 -27123
rect 11276 -27139 11310 -27123
rect 11372 -26820 11406 -26809
rect 11468 -26825 11502 -26809
rect 11372 -27139 11406 -27123
rect 11468 -27139 11502 -27123
rect 11564 -26820 11598 -26809
rect 11660 -26825 11694 -26809
rect 11564 -27139 11598 -27123
rect 11660 -27139 11694 -27123
rect 7373 -27227 7389 -27192
rect 7677 -27227 7703 -27192
rect 8321 -27227 8337 -27192
rect 8625 -27227 8651 -27192
rect 9257 -27227 9273 -27192
rect 9561 -27227 9587 -27192
rect 10188 -27226 10204 -27191
rect 10492 -27226 10518 -27191
rect 11115 -27227 11131 -27192
rect 11419 -27227 11445 -27192
rect 5705 -27747 5721 -27713
rect 5812 -27747 5828 -27713
rect 6145 -27747 6161 -27713
rect 6252 -27747 6268 -27713
rect 6585 -27747 6601 -27713
rect 6692 -27747 6708 -27713
rect 5561 -27833 5611 -27816
rect 5654 -27819 5664 -27785
rect 5860 -27819 5876 -27785
rect -12318 -27892 -12302 -27858
rect -11776 -27892 -11262 -27858
rect -11156 -27892 -11140 -27858
rect -12499 -27976 -12373 -27934
rect -12499 -29098 -12471 -27976
rect -12399 -29098 -12373 -27976
rect -12318 -27980 -12302 -27946
rect -11776 -27980 -11760 -27946
rect -12318 -28076 -12302 -28042
rect -11776 -28076 -11760 -28042
rect -12318 -28172 -12302 -28138
rect -11776 -28172 -11760 -28138
rect -12318 -28268 -12302 -28234
rect -11776 -28268 -11760 -28234
rect -11718 -28283 -11641 -27892
rect -11433 -27947 -11337 -27932
rect -11433 -28012 -11411 -27947
rect -11356 -28012 -11337 -27947
rect -11278 -27980 -11262 -27946
rect -11156 -27980 -11140 -27946
rect -11090 -27975 -10999 -27937
rect -11600 -28114 -11494 -28096
rect -11600 -28194 -11582 -28114
rect -11514 -28194 -11494 -28114
rect -11600 -28211 -11494 -28194
rect -11718 -28303 -11501 -28283
rect -12318 -28364 -12302 -28330
rect -11776 -28364 -11760 -28330
rect -12318 -28460 -12302 -28426
rect -11776 -28460 -11760 -28426
rect -11718 -28433 -11700 -28303
rect -11655 -28314 -11501 -28303
rect -11655 -28428 -11583 -28314
rect -11530 -28428 -11501 -28314
rect -11655 -28433 -11501 -28428
rect -11718 -28460 -11501 -28433
rect -11433 -28506 -11337 -28012
rect -11278 -28076 -11277 -28042
rect -11156 -28076 -11140 -28042
rect -11278 -28172 -11262 -28138
rect -11142 -28172 -11140 -28138
rect -11278 -28268 -11277 -28234
rect -11156 -28268 -11140 -28234
rect -11278 -28364 -11262 -28330
rect -11142 -28364 -11140 -28330
rect -11278 -28460 -11277 -28426
rect -11156 -28460 -11140 -28426
rect -11733 -28522 -11303 -28506
rect -12318 -28556 -12302 -28522
rect -11776 -28556 -11262 -28522
rect -11142 -28556 -11140 -28522
rect -11733 -28572 -11303 -28556
rect -12318 -28652 -12302 -28618
rect -11776 -28652 -11760 -28618
rect -11715 -28626 -11314 -28618
rect -11715 -28634 -11376 -28626
rect -12318 -28748 -12302 -28714
rect -11776 -28748 -11760 -28714
rect -11715 -28764 -11705 -28634
rect -11660 -28756 -11376 -28634
rect -11331 -28756 -11314 -28626
rect -11278 -28652 -11276 -28618
rect -11156 -28652 -11140 -28618
rect -11278 -28748 -11262 -28714
rect -11142 -28748 -11140 -28714
rect -11660 -28764 -11314 -28756
rect -11715 -28783 -11314 -28764
rect -12318 -28844 -12302 -28810
rect -11776 -28844 -11760 -28810
rect -12318 -28940 -12302 -28906
rect -11776 -28940 -11760 -28906
rect -12318 -29036 -12302 -29002
rect -11776 -29036 -11760 -29002
rect -12499 -29144 -12373 -29098
rect -12318 -29132 -12302 -29098
rect -11776 -29132 -11760 -29098
rect -11715 -29186 -11646 -28783
rect -11278 -28844 -11277 -28810
rect -11156 -28844 -11140 -28810
rect -11602 -28901 -11312 -28863
rect -11602 -29034 -11575 -28901
rect -11522 -28909 -11312 -28901
rect -11522 -29034 -11384 -28909
rect -11602 -29039 -11384 -29034
rect -11339 -29039 -11312 -28909
rect -11278 -28940 -11262 -28906
rect -11142 -28940 -11140 -28906
rect -11278 -29036 -11277 -29002
rect -11156 -29036 -11140 -29002
rect -11602 -29084 -11312 -29039
rect -11090 -29098 -11068 -27975
rect -11022 -29098 -10999 -27975
rect 5561 -28059 5577 -27833
rect 6001 -27833 6051 -27816
rect 6094 -27819 6104 -27785
rect 6300 -27819 6316 -27785
rect 5654 -27915 5670 -27881
rect 5864 -27915 5882 -27881
rect 5654 -28011 5664 -27977
rect 5860 -28011 5876 -27977
rect 5561 -28279 5611 -28059
rect 6001 -28059 6017 -27833
rect 6441 -27833 6491 -27816
rect 6534 -27819 6544 -27785
rect 6740 -27819 6756 -27785
rect 6094 -27915 6110 -27881
rect 6304 -27915 6322 -27881
rect 6094 -28011 6104 -27977
rect 6300 -28011 6316 -27977
rect 5654 -28107 5670 -28073
rect 5864 -28107 5882 -28073
rect 5654 -28269 5670 -28235
rect 5846 -28269 5862 -28235
rect 5561 -28313 5577 -28279
rect 5561 -28329 5611 -28313
rect 6001 -28279 6051 -28059
rect 6441 -28059 6457 -27833
rect 6534 -27915 6550 -27881
rect 6744 -27915 6762 -27881
rect 6534 -28011 6544 -27977
rect 6740 -28011 6756 -27977
rect 6094 -28107 6110 -28073
rect 6304 -28107 6322 -28073
rect 6094 -28269 6110 -28235
rect 6286 -28269 6302 -28235
rect 6001 -28313 6017 -28279
rect 5654 -28357 5670 -28323
rect 5846 -28357 5862 -28323
rect 6001 -28329 6051 -28313
rect 6441 -28279 6491 -28059
rect 6534 -28107 6550 -28073
rect 6744 -28107 6762 -28073
rect 6534 -28269 6550 -28235
rect 6726 -28269 6742 -28235
rect 6441 -28313 6457 -28279
rect 6094 -28357 6110 -28323
rect 6286 -28357 6302 -28323
rect 6441 -28329 6491 -28313
rect 6534 -28357 6550 -28323
rect 6726 -28357 6742 -28323
rect 7373 -28420 7389 -28385
rect 7677 -28420 7703 -28385
rect 8321 -28420 8337 -28385
rect 8625 -28420 8651 -28385
rect 9257 -28420 9273 -28385
rect 9561 -28420 9587 -28385
rect 10188 -28420 10204 -28385
rect 10492 -28420 10518 -28385
rect 11115 -28420 11131 -28385
rect 11419 -28420 11445 -28385
rect 5673 -28459 5689 -28425
rect 5821 -28459 5837 -28425
rect 6113 -28459 6129 -28425
rect 6261 -28459 6277 -28425
rect 6553 -28459 6569 -28425
rect 6701 -28459 6717 -28425
rect 7150 -28489 7184 -28473
rect 7246 -28489 7280 -28473
rect 7150 -28803 7184 -28787
rect 7246 -28803 7280 -28792
rect 7342 -28489 7376 -28473
rect 7342 -28803 7376 -28787
rect 7438 -28489 7472 -28473
rect 7534 -28489 7568 -28473
rect 7438 -28803 7472 -28792
rect 7534 -28803 7568 -28787
rect 7630 -28489 7664 -28473
rect 7726 -28489 7760 -28473
rect 7630 -28803 7664 -28792
rect 7726 -28803 7760 -28787
rect 7822 -28489 7856 -28473
rect 7918 -28489 7952 -28473
rect 7822 -28803 7856 -28792
rect 7918 -28803 7952 -28787
rect 8098 -28489 8132 -28473
rect 8194 -28489 8228 -28473
rect 8098 -28803 8132 -28787
rect 8194 -28803 8228 -28792
rect 8290 -28489 8324 -28473
rect 8290 -28803 8324 -28787
rect 8386 -28489 8420 -28473
rect 8482 -28489 8516 -28473
rect 8386 -28803 8420 -28792
rect 8482 -28803 8516 -28787
rect 8578 -28489 8612 -28473
rect 8674 -28489 8708 -28473
rect 8578 -28803 8612 -28792
rect 8674 -28803 8708 -28787
rect 8770 -28489 8804 -28473
rect 8866 -28489 8900 -28473
rect 8770 -28803 8804 -28792
rect 8866 -28803 8900 -28787
rect 9034 -28489 9068 -28473
rect 9130 -28489 9164 -28473
rect 9034 -28803 9068 -28787
rect 9130 -28803 9164 -28792
rect 9226 -28489 9260 -28473
rect 9226 -28803 9260 -28787
rect 9322 -28489 9356 -28473
rect 9418 -28489 9452 -28473
rect 9322 -28803 9356 -28792
rect 9418 -28803 9452 -28787
rect 9514 -28489 9548 -28473
rect 9610 -28489 9644 -28473
rect 9514 -28803 9548 -28792
rect 9610 -28803 9644 -28787
rect 9706 -28489 9740 -28473
rect 9802 -28489 9836 -28473
rect 9706 -28803 9740 -28792
rect 9802 -28803 9836 -28787
rect 9965 -28489 9999 -28473
rect 10061 -28489 10095 -28473
rect 9965 -28803 9999 -28787
rect 10061 -28803 10095 -28792
rect 10157 -28489 10191 -28473
rect 10157 -28803 10191 -28787
rect 10253 -28489 10287 -28473
rect 10349 -28489 10383 -28473
rect 10253 -28803 10287 -28792
rect 10349 -28803 10383 -28787
rect 10445 -28489 10479 -28473
rect 10541 -28489 10575 -28473
rect 10445 -28803 10479 -28792
rect 10541 -28803 10575 -28787
rect 10637 -28489 10671 -28473
rect 10733 -28489 10767 -28473
rect 10637 -28803 10671 -28792
rect 10733 -28803 10767 -28787
rect 10892 -28489 10926 -28473
rect 10988 -28489 11022 -28473
rect 10892 -28803 10926 -28787
rect 10988 -28803 11022 -28792
rect 11084 -28489 11118 -28473
rect 11084 -28803 11118 -28787
rect 11180 -28489 11214 -28473
rect 11276 -28489 11310 -28473
rect 11180 -28803 11214 -28792
rect 11276 -28803 11310 -28787
rect 11372 -28489 11406 -28473
rect 11468 -28489 11502 -28473
rect 11372 -28803 11406 -28792
rect 11468 -28803 11502 -28787
rect 11564 -28489 11598 -28473
rect 11660 -28489 11694 -28473
rect 11564 -28803 11598 -28792
rect 11660 -28803 11694 -28787
rect 7182 -28880 7198 -28846
rect 7232 -28880 7248 -28846
rect 7374 -28880 7390 -28846
rect 7424 -28880 7440 -28846
rect 7566 -28880 7582 -28846
rect 7616 -28880 7632 -28846
rect 7758 -28880 7774 -28846
rect 7808 -28880 7824 -28846
rect 8130 -28880 8146 -28846
rect 8180 -28880 8196 -28846
rect 8322 -28880 8338 -28846
rect 8372 -28880 8388 -28846
rect 8514 -28880 8530 -28846
rect 8564 -28880 8580 -28846
rect 8706 -28880 8722 -28846
rect 8756 -28880 8772 -28846
rect 9066 -28880 9082 -28846
rect 9116 -28880 9132 -28846
rect 9258 -28880 9274 -28846
rect 9308 -28880 9324 -28846
rect 9450 -28880 9466 -28846
rect 9500 -28880 9516 -28846
rect 9642 -28880 9658 -28846
rect 9692 -28880 9708 -28846
rect 9997 -28880 10013 -28846
rect 10047 -28880 10063 -28846
rect 10189 -28880 10205 -28846
rect 10239 -28880 10255 -28846
rect 10381 -28880 10397 -28846
rect 10431 -28880 10447 -28846
rect 10573 -28880 10589 -28846
rect 10623 -28880 10639 -28846
rect 10924 -28880 10940 -28846
rect 10974 -28880 10990 -28846
rect 11116 -28880 11132 -28846
rect 11166 -28880 11182 -28846
rect 11308 -28880 11324 -28846
rect 11358 -28880 11374 -28846
rect 11500 -28880 11516 -28846
rect 11550 -28880 11566 -28846
rect -11278 -29132 -11262 -29098
rect -11156 -29132 -11140 -29098
rect -11090 -29139 -10999 -29098
rect -12318 -29220 -12302 -29186
rect -11776 -29220 -11262 -29186
rect -11156 -29220 -11140 -29186
rect 7298 -29202 7403 -29199
rect 8246 -29202 8351 -29199
rect 9182 -29202 9287 -29199
rect 10113 -29202 10218 -29199
rect 11040 -29202 11145 -29199
rect 7298 -29218 7406 -29202
rect 7298 -29230 7372 -29218
rect -11568 -29443 -11562 -29395
rect -11494 -29443 -11488 -29395
rect 7333 -29981 7372 -29230
rect 7298 -29994 7372 -29981
rect 7298 -30010 7406 -29994
rect 7756 -29218 7790 -29202
rect 7756 -30010 7790 -29994
rect 8246 -29218 8354 -29202
rect 8246 -29230 8320 -29218
rect 8281 -29981 8320 -29230
rect 8246 -29994 8320 -29981
rect 8246 -30010 8354 -29994
rect 8704 -29218 8738 -29202
rect 8704 -30010 8738 -29994
rect 9182 -29218 9290 -29202
rect 9182 -29230 9256 -29218
rect 9217 -29981 9256 -29230
rect 9182 -29994 9256 -29981
rect 9182 -30010 9290 -29994
rect 9640 -29218 9674 -29202
rect 9640 -30010 9674 -29994
rect 10113 -29218 10221 -29202
rect 10113 -29230 10187 -29218
rect 10148 -29981 10187 -29230
rect 10113 -29994 10187 -29981
rect 10113 -30010 10221 -29994
rect 10571 -29218 10605 -29202
rect 10571 -30010 10605 -29994
rect 11040 -29218 11148 -29202
rect 11040 -29230 11114 -29218
rect 11075 -29981 11114 -29230
rect 11040 -29994 11114 -29981
rect 11040 -30010 11148 -29994
rect 11498 -29218 11532 -29202
rect 11783 -29544 12203 -29524
rect 11783 -29595 11811 -29544
rect 12168 -29595 12203 -29544
rect 11783 -29614 12203 -29595
rect 11785 -29699 11819 -29614
rect 11785 -29947 11819 -29931
rect 11881 -29699 11915 -29683
rect 11881 -29947 11915 -29931
rect 11977 -29699 12011 -29614
rect 11977 -29947 12011 -29931
rect 12073 -29699 12107 -29683
rect 12073 -29947 12107 -29931
rect 12169 -29699 12203 -29614
rect 12169 -29947 12203 -29931
rect 12265 -29699 12299 -29683
rect 12265 -29947 12299 -29931
rect 12361 -29699 12395 -29683
rect 12361 -29947 12395 -29931
rect 12457 -29699 12491 -29683
rect 12457 -29947 12491 -29931
rect 12553 -29699 12587 -29683
rect 12553 -29947 12587 -29931
rect 12649 -29699 12683 -29683
rect 12649 -29947 12683 -29931
rect 12745 -29699 12779 -29683
rect 12970 -29765 12986 -29731
rect 13077 -29765 13093 -29731
rect 12745 -29947 12779 -29931
rect 12826 -29851 12876 -29834
rect 12919 -29837 12929 -29803
rect 13125 -29837 13141 -29803
rect 11498 -30010 11532 -29994
rect 12154 -30027 12170 -29993
rect 12204 -30027 12220 -29993
rect 12826 -30077 12842 -29851
rect 12919 -29933 12935 -29899
rect 13129 -29933 13147 -29899
rect 12919 -30029 12929 -29995
rect 13125 -30029 13141 -29995
rect 7298 -30146 7406 -30130
rect 7298 -30159 7372 -30146
rect -12318 -30501 -12302 -30467
rect -11776 -30501 -11262 -30467
rect -11156 -30501 -11140 -30467
rect -12499 -30585 -12373 -30543
rect -12499 -31707 -12471 -30585
rect -12399 -31707 -12373 -30585
rect -12318 -30589 -12302 -30555
rect -11776 -30589 -11760 -30555
rect -12318 -30685 -12302 -30651
rect -11776 -30685 -11760 -30651
rect -12318 -30781 -12302 -30747
rect -11776 -30781 -11760 -30747
rect -12318 -30877 -12302 -30843
rect -11776 -30877 -11760 -30843
rect -11718 -30892 -11641 -30501
rect -11433 -30556 -11337 -30541
rect -11433 -30621 -11411 -30556
rect -11356 -30621 -11337 -30556
rect -11278 -30589 -11262 -30555
rect -11156 -30589 -11140 -30555
rect -11090 -30584 -10999 -30546
rect -11600 -30723 -11494 -30705
rect -11600 -30803 -11582 -30723
rect -11514 -30803 -11494 -30723
rect -11600 -30820 -11494 -30803
rect -11718 -30912 -11501 -30892
rect -12318 -30973 -12302 -30939
rect -11776 -30973 -11760 -30939
rect -12318 -31069 -12302 -31035
rect -11776 -31069 -11760 -31035
rect -11718 -31042 -11700 -30912
rect -11655 -30923 -11501 -30912
rect -11655 -31037 -11583 -30923
rect -11530 -31037 -11501 -30923
rect -11655 -31042 -11501 -31037
rect -11718 -31069 -11501 -31042
rect -11433 -31115 -11337 -30621
rect -11278 -30685 -11277 -30651
rect -11156 -30685 -11140 -30651
rect -11278 -30781 -11262 -30747
rect -11142 -30781 -11140 -30747
rect -11278 -30877 -11277 -30843
rect -11156 -30877 -11140 -30843
rect -11278 -30973 -11262 -30939
rect -11142 -30973 -11140 -30939
rect -11278 -31069 -11277 -31035
rect -11156 -31069 -11140 -31035
rect -11733 -31131 -11303 -31115
rect -12318 -31165 -12302 -31131
rect -11776 -31165 -11262 -31131
rect -11142 -31165 -11140 -31131
rect -11733 -31181 -11303 -31165
rect -12318 -31261 -12302 -31227
rect -11776 -31261 -11760 -31227
rect -11715 -31235 -11314 -31227
rect -11715 -31243 -11376 -31235
rect -12318 -31357 -12302 -31323
rect -11776 -31357 -11760 -31323
rect -11715 -31373 -11705 -31243
rect -11660 -31365 -11376 -31243
rect -11331 -31365 -11314 -31235
rect -11278 -31261 -11276 -31227
rect -11156 -31261 -11140 -31227
rect -11278 -31357 -11262 -31323
rect -11142 -31357 -11140 -31323
rect -11660 -31373 -11314 -31365
rect -11715 -31392 -11314 -31373
rect -12318 -31453 -12302 -31419
rect -11776 -31453 -11760 -31419
rect -12318 -31549 -12302 -31515
rect -11776 -31549 -11760 -31515
rect -12318 -31645 -12302 -31611
rect -11776 -31645 -11760 -31611
rect -12499 -31753 -12373 -31707
rect -12318 -31741 -12302 -31707
rect -11776 -31741 -11760 -31707
rect -11715 -31795 -11646 -31392
rect -11278 -31453 -11277 -31419
rect -11156 -31453 -11140 -31419
rect -11602 -31510 -11312 -31472
rect -11602 -31643 -11575 -31510
rect -11522 -31518 -11312 -31510
rect -11522 -31643 -11384 -31518
rect -11602 -31648 -11384 -31643
rect -11339 -31648 -11312 -31518
rect -11278 -31549 -11262 -31515
rect -11142 -31549 -11140 -31515
rect -11278 -31645 -11277 -31611
rect -11156 -31645 -11140 -31611
rect -11602 -31693 -11312 -31648
rect -11090 -31707 -11068 -30584
rect -11022 -31707 -10999 -30584
rect 7333 -30910 7372 -30159
rect 7298 -30922 7372 -30910
rect 7298 -30938 7406 -30922
rect 7756 -30146 7790 -30130
rect 7756 -30938 7790 -30922
rect 8246 -30146 8354 -30130
rect 8246 -30159 8320 -30146
rect 8281 -30910 8320 -30159
rect 8246 -30922 8320 -30910
rect 8246 -30938 8354 -30922
rect 8704 -30146 8738 -30130
rect 8704 -30938 8738 -30922
rect 9182 -30146 9290 -30130
rect 9182 -30159 9256 -30146
rect 9217 -30910 9256 -30159
rect 9182 -30922 9256 -30910
rect 9182 -30938 9290 -30922
rect 9640 -30146 9674 -30130
rect 9640 -30938 9674 -30922
rect 10113 -30145 10221 -30129
rect 10113 -30158 10187 -30145
rect 10148 -30909 10187 -30158
rect 10113 -30921 10187 -30909
rect 10113 -30937 10221 -30921
rect 10571 -30145 10605 -30129
rect 10571 -30937 10605 -30921
rect 11040 -30146 11148 -30130
rect 11040 -30159 11114 -30146
rect 11075 -30910 11114 -30159
rect 11040 -30922 11114 -30910
rect 7298 -30941 7403 -30938
rect 8246 -30941 8351 -30938
rect 9182 -30941 9287 -30938
rect 10113 -30940 10218 -30937
rect 11040 -30938 11148 -30922
rect 11498 -30146 11532 -30130
rect 12297 -30132 12313 -30098
rect 12347 -30132 12363 -30098
rect 12169 -30188 12203 -30172
rect 12169 -30436 12203 -30364
rect 12265 -30188 12299 -30172
rect 12265 -30380 12299 -30364
rect 12361 -30188 12395 -30172
rect 12826 -30297 12876 -30077
rect 12919 -30125 12935 -30091
rect 13129 -30125 13147 -30091
rect 12919 -30287 12935 -30253
rect 13111 -30287 13127 -30253
rect 12826 -30331 12842 -30297
rect 12826 -30347 12876 -30331
rect 12361 -30436 12395 -30364
rect 12919 -30375 12935 -30341
rect 13111 -30375 13127 -30341
rect 12157 -30447 12407 -30436
rect 12157 -30508 12183 -30447
rect 12382 -30508 12407 -30447
rect 12938 -30477 12954 -30443
rect 13086 -30477 13102 -30443
rect 12157 -30520 12407 -30508
rect 11498 -30938 11532 -30922
rect 11040 -30941 11145 -30938
rect 7182 -31294 7198 -31260
rect 7232 -31294 7248 -31260
rect 7374 -31294 7390 -31260
rect 7424 -31294 7440 -31260
rect 7566 -31294 7582 -31260
rect 7616 -31294 7632 -31260
rect 7758 -31294 7774 -31260
rect 7808 -31294 7824 -31260
rect 8130 -31294 8146 -31260
rect 8180 -31294 8196 -31260
rect 8322 -31294 8338 -31260
rect 8372 -31294 8388 -31260
rect 8514 -31294 8530 -31260
rect 8564 -31294 8580 -31260
rect 8706 -31294 8722 -31260
rect 8756 -31294 8772 -31260
rect 9066 -31294 9082 -31260
rect 9116 -31294 9132 -31260
rect 9258 -31294 9274 -31260
rect 9308 -31294 9324 -31260
rect 9450 -31294 9466 -31260
rect 9500 -31294 9516 -31260
rect 9642 -31294 9658 -31260
rect 9692 -31294 9708 -31260
rect 9997 -31293 10013 -31259
rect 10047 -31293 10063 -31259
rect 10189 -31293 10205 -31259
rect 10239 -31293 10255 -31259
rect 10381 -31293 10397 -31259
rect 10431 -31293 10447 -31259
rect 10573 -31293 10589 -31259
rect 10623 -31293 10639 -31259
rect 10924 -31294 10940 -31260
rect 10974 -31294 10990 -31260
rect 11116 -31294 11132 -31260
rect 11166 -31294 11182 -31260
rect 11308 -31294 11324 -31260
rect 11358 -31294 11374 -31260
rect 11500 -31294 11516 -31260
rect 11550 -31294 11566 -31260
rect 7150 -31353 7184 -31337
rect 7246 -31348 7280 -31337
rect 7150 -31667 7184 -31651
rect 7246 -31667 7280 -31651
rect 7342 -31353 7376 -31337
rect 7342 -31667 7376 -31651
rect 7438 -31348 7472 -31337
rect 7534 -31353 7568 -31337
rect 7438 -31667 7472 -31651
rect 7534 -31667 7568 -31651
rect 7630 -31348 7664 -31337
rect 7726 -31353 7760 -31337
rect 7630 -31667 7664 -31651
rect 7726 -31667 7760 -31651
rect 7822 -31348 7856 -31337
rect 7918 -31353 7952 -31337
rect 7822 -31667 7856 -31651
rect 7918 -31667 7952 -31651
rect 8098 -31353 8132 -31337
rect 8194 -31348 8228 -31337
rect 8098 -31667 8132 -31651
rect 8194 -31667 8228 -31651
rect 8290 -31353 8324 -31337
rect 8290 -31667 8324 -31651
rect 8386 -31348 8420 -31337
rect 8482 -31353 8516 -31337
rect 8386 -31667 8420 -31651
rect 8482 -31667 8516 -31651
rect 8578 -31348 8612 -31337
rect 8674 -31353 8708 -31337
rect 8578 -31667 8612 -31651
rect 8674 -31667 8708 -31651
rect 8770 -31348 8804 -31337
rect 8866 -31353 8900 -31337
rect 8770 -31667 8804 -31651
rect 8866 -31667 8900 -31651
rect 9034 -31353 9068 -31337
rect 9130 -31348 9164 -31337
rect 9034 -31667 9068 -31651
rect 9130 -31667 9164 -31651
rect 9226 -31353 9260 -31337
rect 9226 -31667 9260 -31651
rect 9322 -31348 9356 -31337
rect 9418 -31353 9452 -31337
rect 9322 -31667 9356 -31651
rect 9418 -31667 9452 -31651
rect 9514 -31348 9548 -31337
rect 9610 -31353 9644 -31337
rect 9514 -31667 9548 -31651
rect 9610 -31667 9644 -31651
rect 9706 -31348 9740 -31337
rect 9802 -31353 9836 -31337
rect 9706 -31667 9740 -31651
rect 9802 -31667 9836 -31651
rect 9965 -31352 9999 -31336
rect 10061 -31347 10095 -31336
rect 9965 -31666 9999 -31650
rect 10061 -31666 10095 -31650
rect 10157 -31352 10191 -31336
rect 10157 -31666 10191 -31650
rect 10253 -31347 10287 -31336
rect 10349 -31352 10383 -31336
rect 10253 -31666 10287 -31650
rect 10349 -31666 10383 -31650
rect 10445 -31347 10479 -31336
rect 10541 -31352 10575 -31336
rect 10445 -31666 10479 -31650
rect 10541 -31666 10575 -31650
rect 10637 -31347 10671 -31336
rect 10733 -31352 10767 -31336
rect 10637 -31666 10671 -31650
rect 10733 -31666 10767 -31650
rect 10892 -31353 10926 -31337
rect 10988 -31348 11022 -31337
rect 10892 -31667 10926 -31651
rect 10988 -31667 11022 -31651
rect 11084 -31353 11118 -31337
rect 11084 -31667 11118 -31651
rect 11180 -31348 11214 -31337
rect 11276 -31353 11310 -31337
rect 11180 -31667 11214 -31651
rect 11276 -31667 11310 -31651
rect 11372 -31348 11406 -31337
rect 11468 -31353 11502 -31337
rect 11372 -31667 11406 -31651
rect 11468 -31667 11502 -31651
rect 11564 -31348 11598 -31337
rect 11660 -31353 11694 -31337
rect 11564 -31667 11598 -31651
rect 11660 -31667 11694 -31651
rect -11278 -31741 -11262 -31707
rect -11156 -31741 -11140 -31707
rect -11090 -31748 -10999 -31707
rect 7373 -31755 7389 -31720
rect 7677 -31755 7703 -31720
rect 8321 -31755 8337 -31720
rect 8625 -31755 8651 -31720
rect 9257 -31755 9273 -31720
rect 9561 -31755 9587 -31720
rect 10188 -31754 10204 -31719
rect 10492 -31754 10518 -31719
rect 11115 -31755 11131 -31720
rect 11419 -31755 11445 -31720
rect -12318 -31829 -12302 -31795
rect -11776 -31829 -11262 -31795
rect -11156 -31829 -11140 -31795
rect -11570 -31988 -11564 -31937
rect -11493 -31988 -11487 -31937
rect 5705 -32275 5721 -32241
rect 5812 -32275 5828 -32241
rect 6145 -32275 6161 -32241
rect 6252 -32275 6268 -32241
rect 6585 -32275 6601 -32241
rect 6692 -32275 6708 -32241
rect 5561 -32361 5611 -32344
rect 5654 -32347 5664 -32313
rect 5860 -32347 5876 -32313
rect 5561 -32587 5577 -32361
rect 6001 -32361 6051 -32344
rect 6094 -32347 6104 -32313
rect 6300 -32347 6316 -32313
rect 5654 -32443 5670 -32409
rect 5864 -32443 5882 -32409
rect 5654 -32539 5664 -32505
rect 5860 -32539 5876 -32505
rect 5561 -32807 5611 -32587
rect 6001 -32587 6017 -32361
rect 6441 -32361 6491 -32344
rect 6534 -32347 6544 -32313
rect 6740 -32347 6756 -32313
rect 6094 -32443 6110 -32409
rect 6304 -32443 6322 -32409
rect 6094 -32539 6104 -32505
rect 6300 -32539 6316 -32505
rect 5654 -32635 5670 -32601
rect 5864 -32635 5882 -32601
rect 5654 -32797 5670 -32763
rect 5846 -32797 5862 -32763
rect 5561 -32841 5577 -32807
rect 5561 -32857 5611 -32841
rect 6001 -32807 6051 -32587
rect 6441 -32587 6457 -32361
rect 6534 -32443 6550 -32409
rect 6744 -32443 6762 -32409
rect 6534 -32539 6544 -32505
rect 6740 -32539 6756 -32505
rect 6094 -32635 6110 -32601
rect 6304 -32635 6322 -32601
rect 6094 -32797 6110 -32763
rect 6286 -32797 6302 -32763
rect 6001 -32841 6017 -32807
rect 5654 -32885 5670 -32851
rect 5846 -32885 5862 -32851
rect 6001 -32857 6051 -32841
rect 6441 -32807 6491 -32587
rect 6534 -32635 6550 -32601
rect 6744 -32635 6762 -32601
rect 6534 -32797 6550 -32763
rect 6726 -32797 6742 -32763
rect 6441 -32841 6457 -32807
rect 6094 -32885 6110 -32851
rect 6286 -32885 6302 -32851
rect 6441 -32857 6491 -32841
rect 6534 -32885 6550 -32851
rect 6726 -32885 6742 -32851
rect 7373 -32948 7389 -32913
rect 7677 -32948 7703 -32913
rect 8321 -32948 8337 -32913
rect 8625 -32948 8651 -32913
rect 9257 -32948 9273 -32913
rect 9561 -32948 9587 -32913
rect 10188 -32948 10204 -32913
rect 10492 -32948 10518 -32913
rect 11115 -32948 11131 -32913
rect 11419 -32948 11445 -32913
rect 5673 -32987 5689 -32953
rect 5821 -32987 5837 -32953
rect 6113 -32987 6129 -32953
rect 6261 -32987 6277 -32953
rect 6553 -32987 6569 -32953
rect 6701 -32987 6717 -32953
rect 7150 -33017 7184 -33001
rect -12320 -33121 -12304 -33087
rect -11778 -33121 -11264 -33087
rect -11158 -33121 -11142 -33087
rect -12501 -33205 -12375 -33163
rect -12501 -34327 -12473 -33205
rect -12401 -34327 -12375 -33205
rect -12320 -33209 -12304 -33175
rect -11778 -33209 -11762 -33175
rect -12320 -33305 -12304 -33271
rect -11778 -33305 -11762 -33271
rect -12320 -33401 -12304 -33367
rect -11778 -33401 -11762 -33367
rect -12320 -33497 -12304 -33463
rect -11778 -33497 -11762 -33463
rect -11720 -33512 -11643 -33121
rect -11435 -33176 -11339 -33161
rect -11435 -33241 -11413 -33176
rect -11358 -33241 -11339 -33176
rect -11280 -33209 -11264 -33175
rect -11158 -33209 -11142 -33175
rect -11092 -33204 -11001 -33166
rect -11602 -33343 -11496 -33325
rect -11602 -33423 -11584 -33343
rect -11516 -33423 -11496 -33343
rect -11602 -33440 -11496 -33423
rect -11720 -33532 -11503 -33512
rect -12320 -33593 -12304 -33559
rect -11778 -33593 -11762 -33559
rect -12320 -33689 -12304 -33655
rect -11778 -33689 -11762 -33655
rect -11720 -33662 -11702 -33532
rect -11657 -33543 -11503 -33532
rect -11657 -33657 -11585 -33543
rect -11532 -33657 -11503 -33543
rect -11657 -33662 -11503 -33657
rect -11720 -33689 -11503 -33662
rect -11435 -33735 -11339 -33241
rect -11280 -33305 -11279 -33271
rect -11158 -33305 -11142 -33271
rect -11280 -33401 -11264 -33367
rect -11144 -33401 -11142 -33367
rect -11280 -33497 -11279 -33463
rect -11158 -33497 -11142 -33463
rect -11280 -33593 -11264 -33559
rect -11144 -33593 -11142 -33559
rect -11280 -33689 -11279 -33655
rect -11158 -33689 -11142 -33655
rect -11735 -33751 -11305 -33735
rect -12320 -33785 -12304 -33751
rect -11778 -33785 -11264 -33751
rect -11144 -33785 -11142 -33751
rect -11735 -33801 -11305 -33785
rect -12320 -33881 -12304 -33847
rect -11778 -33881 -11762 -33847
rect -11717 -33855 -11316 -33847
rect -11717 -33863 -11378 -33855
rect -12320 -33977 -12304 -33943
rect -11778 -33977 -11762 -33943
rect -11717 -33993 -11707 -33863
rect -11662 -33985 -11378 -33863
rect -11333 -33985 -11316 -33855
rect -11280 -33881 -11278 -33847
rect -11158 -33881 -11142 -33847
rect -11280 -33977 -11264 -33943
rect -11144 -33977 -11142 -33943
rect -11662 -33993 -11316 -33985
rect -11717 -34012 -11316 -33993
rect -12320 -34073 -12304 -34039
rect -11778 -34073 -11762 -34039
rect -12320 -34169 -12304 -34135
rect -11778 -34169 -11762 -34135
rect -12320 -34265 -12304 -34231
rect -11778 -34265 -11762 -34231
rect -12501 -34373 -12375 -34327
rect -12320 -34361 -12304 -34327
rect -11778 -34361 -11762 -34327
rect -11717 -34415 -11648 -34012
rect -11280 -34073 -11279 -34039
rect -11158 -34073 -11142 -34039
rect -11604 -34130 -11314 -34092
rect -11604 -34263 -11577 -34130
rect -11524 -34138 -11314 -34130
rect -11524 -34263 -11386 -34138
rect -11604 -34268 -11386 -34263
rect -11341 -34268 -11314 -34138
rect -11280 -34169 -11264 -34135
rect -11144 -34169 -11142 -34135
rect -11280 -34265 -11279 -34231
rect -11158 -34265 -11142 -34231
rect -11604 -34313 -11314 -34268
rect -11092 -34327 -11070 -33204
rect -11024 -34327 -11001 -33204
rect 7246 -33017 7280 -33001
rect 7150 -33331 7184 -33315
rect 7246 -33331 7280 -33320
rect 7342 -33017 7376 -33001
rect 7342 -33331 7376 -33315
rect 7438 -33017 7472 -33001
rect 7534 -33017 7568 -33001
rect 7438 -33331 7472 -33320
rect 7534 -33331 7568 -33315
rect 7630 -33017 7664 -33001
rect 7726 -33017 7760 -33001
rect 7630 -33331 7664 -33320
rect 7726 -33331 7760 -33315
rect 7822 -33017 7856 -33001
rect 7918 -33017 7952 -33001
rect 7822 -33331 7856 -33320
rect 7918 -33331 7952 -33315
rect 8098 -33017 8132 -33001
rect 8194 -33017 8228 -33001
rect 8098 -33331 8132 -33315
rect 8194 -33331 8228 -33320
rect 8290 -33017 8324 -33001
rect 8290 -33331 8324 -33315
rect 8386 -33017 8420 -33001
rect 8482 -33017 8516 -33001
rect 8386 -33331 8420 -33320
rect 8482 -33331 8516 -33315
rect 8578 -33017 8612 -33001
rect 8674 -33017 8708 -33001
rect 8578 -33331 8612 -33320
rect 8674 -33331 8708 -33315
rect 8770 -33017 8804 -33001
rect 8866 -33017 8900 -33001
rect 8770 -33331 8804 -33320
rect 8866 -33331 8900 -33315
rect 9034 -33017 9068 -33001
rect 9130 -33017 9164 -33001
rect 9034 -33331 9068 -33315
rect 9130 -33331 9164 -33320
rect 9226 -33017 9260 -33001
rect 9226 -33331 9260 -33315
rect 9322 -33017 9356 -33001
rect 9418 -33017 9452 -33001
rect 9322 -33331 9356 -33320
rect 9418 -33331 9452 -33315
rect 9514 -33017 9548 -33001
rect 9610 -33017 9644 -33001
rect 9514 -33331 9548 -33320
rect 9610 -33331 9644 -33315
rect 9706 -33017 9740 -33001
rect 9802 -33017 9836 -33001
rect 9706 -33331 9740 -33320
rect 9802 -33331 9836 -33315
rect 9965 -33017 9999 -33001
rect 10061 -33017 10095 -33001
rect 9965 -33331 9999 -33315
rect 10061 -33331 10095 -33320
rect 10157 -33017 10191 -33001
rect 10157 -33331 10191 -33315
rect 10253 -33017 10287 -33001
rect 10349 -33017 10383 -33001
rect 10253 -33331 10287 -33320
rect 10349 -33331 10383 -33315
rect 10445 -33017 10479 -33001
rect 10541 -33017 10575 -33001
rect 10445 -33331 10479 -33320
rect 10541 -33331 10575 -33315
rect 10637 -33017 10671 -33001
rect 10733 -33017 10767 -33001
rect 10637 -33331 10671 -33320
rect 10733 -33331 10767 -33315
rect 10892 -33017 10926 -33001
rect 10988 -33017 11022 -33001
rect 10892 -33331 10926 -33315
rect 10988 -33331 11022 -33320
rect 11084 -33017 11118 -33001
rect 11084 -33331 11118 -33315
rect 11180 -33017 11214 -33001
rect 11276 -33017 11310 -33001
rect 11180 -33331 11214 -33320
rect 11276 -33331 11310 -33315
rect 11372 -33017 11406 -33001
rect 11468 -33017 11502 -33001
rect 11372 -33331 11406 -33320
rect 11468 -33331 11502 -33315
rect 11564 -33017 11598 -33001
rect 11660 -33017 11694 -33001
rect 11564 -33331 11598 -33320
rect 11660 -33331 11694 -33315
rect 7182 -33408 7198 -33374
rect 7232 -33408 7248 -33374
rect 7374 -33408 7390 -33374
rect 7424 -33408 7440 -33374
rect 7566 -33408 7582 -33374
rect 7616 -33408 7632 -33374
rect 7758 -33408 7774 -33374
rect 7808 -33408 7824 -33374
rect 8130 -33408 8146 -33374
rect 8180 -33408 8196 -33374
rect 8322 -33408 8338 -33374
rect 8372 -33408 8388 -33374
rect 8514 -33408 8530 -33374
rect 8564 -33408 8580 -33374
rect 8706 -33408 8722 -33374
rect 8756 -33408 8772 -33374
rect 9066 -33408 9082 -33374
rect 9116 -33408 9132 -33374
rect 9258 -33408 9274 -33374
rect 9308 -33408 9324 -33374
rect 9450 -33408 9466 -33374
rect 9500 -33408 9516 -33374
rect 9642 -33408 9658 -33374
rect 9692 -33408 9708 -33374
rect 9997 -33408 10013 -33374
rect 10047 -33408 10063 -33374
rect 10189 -33408 10205 -33374
rect 10239 -33408 10255 -33374
rect 10381 -33408 10397 -33374
rect 10431 -33408 10447 -33374
rect 10573 -33408 10589 -33374
rect 10623 -33408 10639 -33374
rect 10924 -33408 10940 -33374
rect 10974 -33408 10990 -33374
rect 11116 -33408 11132 -33374
rect 11166 -33408 11182 -33374
rect 11308 -33408 11324 -33374
rect 11358 -33408 11374 -33374
rect 11500 -33408 11516 -33374
rect 11550 -33408 11566 -33374
rect -11280 -34361 -11264 -34327
rect -11158 -34361 -11142 -34327
rect -11092 -34368 -11001 -34327
rect 7298 -33730 7403 -33727
rect 8246 -33730 8351 -33727
rect 9182 -33730 9287 -33727
rect 10113 -33730 10218 -33727
rect 11040 -33730 11145 -33727
rect 7298 -33746 7406 -33730
rect 7298 -33758 7372 -33746
rect -12320 -34449 -12304 -34415
rect -11778 -34449 -11264 -34415
rect -11158 -34449 -11142 -34415
rect 7333 -34509 7372 -33758
rect 7298 -34522 7372 -34509
rect -11564 -34567 -11553 -34533
rect -11510 -34567 -11498 -34533
rect 7298 -34538 7406 -34522
rect 7756 -33746 7790 -33730
rect 7756 -34538 7790 -34522
rect 8246 -33746 8354 -33730
rect 8246 -33758 8320 -33746
rect 8281 -34509 8320 -33758
rect 8246 -34522 8320 -34509
rect 8246 -34538 8354 -34522
rect 8704 -33746 8738 -33730
rect 8704 -34538 8738 -34522
rect 9182 -33746 9290 -33730
rect 9182 -33758 9256 -33746
rect 9217 -34509 9256 -33758
rect 9182 -34522 9256 -34509
rect 9182 -34538 9290 -34522
rect 9640 -33746 9674 -33730
rect 9640 -34538 9674 -34522
rect 10113 -33746 10221 -33730
rect 10113 -33758 10187 -33746
rect 10148 -34509 10187 -33758
rect 10113 -34522 10187 -34509
rect 10113 -34538 10221 -34522
rect 10571 -33746 10605 -33730
rect 10571 -34538 10605 -34522
rect 11040 -33746 11148 -33730
rect 11040 -33758 11114 -33746
rect 11075 -34509 11114 -33758
rect 11040 -34522 11114 -34509
rect 11040 -34538 11148 -34522
rect 11498 -33746 11532 -33730
rect 11783 -34072 12203 -34052
rect 11783 -34123 11811 -34072
rect 12168 -34123 12203 -34072
rect 11783 -34142 12203 -34123
rect 11785 -34227 11819 -34142
rect 11785 -34475 11819 -34459
rect 11881 -34227 11915 -34211
rect 11881 -34475 11915 -34459
rect 11977 -34227 12011 -34142
rect 11977 -34475 12011 -34459
rect 12073 -34227 12107 -34211
rect 12073 -34475 12107 -34459
rect 12169 -34227 12203 -34142
rect 12169 -34475 12203 -34459
rect 12265 -34227 12299 -34211
rect 12265 -34475 12299 -34459
rect 12361 -34227 12395 -34211
rect 12361 -34475 12395 -34459
rect 12457 -34227 12491 -34211
rect 12457 -34475 12491 -34459
rect 12553 -34227 12587 -34211
rect 12553 -34475 12587 -34459
rect 12649 -34227 12683 -34211
rect 12649 -34475 12683 -34459
rect 12745 -34227 12779 -34211
rect 12970 -34293 12986 -34259
rect 13077 -34293 13093 -34259
rect 12745 -34475 12779 -34459
rect 12826 -34379 12876 -34362
rect 12919 -34365 12929 -34331
rect 13125 -34365 13141 -34331
rect 11498 -34538 11532 -34522
rect 12154 -34555 12170 -34521
rect 12204 -34555 12220 -34521
rect 12826 -34605 12842 -34379
rect 12919 -34461 12935 -34427
rect 13129 -34461 13147 -34427
rect 12919 -34557 12929 -34523
rect 13125 -34557 13141 -34523
rect 7298 -34674 7406 -34658
rect 7298 -34687 7372 -34674
rect 7333 -35438 7372 -34687
rect 7298 -35450 7372 -35438
rect 7298 -35466 7406 -35450
rect 7756 -34674 7790 -34658
rect 7756 -35466 7790 -35450
rect 8246 -34674 8354 -34658
rect 8246 -34687 8320 -34674
rect 8281 -35438 8320 -34687
rect 8246 -35450 8320 -35438
rect 8246 -35466 8354 -35450
rect 8704 -34674 8738 -34658
rect 8704 -35466 8738 -35450
rect 9182 -34674 9290 -34658
rect 9182 -34687 9256 -34674
rect 9217 -35438 9256 -34687
rect 9182 -35450 9256 -35438
rect 9182 -35466 9290 -35450
rect 9640 -34674 9674 -34658
rect 9640 -35466 9674 -35450
rect 10113 -34673 10221 -34657
rect 10113 -34686 10187 -34673
rect 10148 -35437 10187 -34686
rect 10113 -35449 10187 -35437
rect 10113 -35465 10221 -35449
rect 10571 -34673 10605 -34657
rect 10571 -35465 10605 -35449
rect 11040 -34674 11148 -34658
rect 11040 -34687 11114 -34674
rect 11075 -35438 11114 -34687
rect 11040 -35450 11114 -35438
rect 7298 -35469 7403 -35466
rect 8246 -35469 8351 -35466
rect 9182 -35469 9287 -35466
rect 10113 -35468 10218 -35465
rect 11040 -35466 11148 -35450
rect 11498 -34674 11532 -34658
rect 12297 -34660 12313 -34626
rect 12347 -34660 12363 -34626
rect 12169 -34716 12203 -34700
rect 12169 -34964 12203 -34892
rect 12265 -34716 12299 -34700
rect 12265 -34908 12299 -34892
rect 12361 -34716 12395 -34700
rect 12826 -34825 12876 -34605
rect 12919 -34653 12935 -34619
rect 13129 -34653 13147 -34619
rect 12919 -34815 12935 -34781
rect 13111 -34815 13127 -34781
rect 12826 -34859 12842 -34825
rect 12826 -34875 12876 -34859
rect 12361 -34964 12395 -34892
rect 12919 -34903 12935 -34869
rect 13111 -34903 13127 -34869
rect 12157 -34975 12407 -34964
rect 12157 -35036 12183 -34975
rect 12382 -35036 12407 -34975
rect 12938 -35005 12954 -34971
rect 13086 -35005 13102 -34971
rect 12157 -35048 12407 -35036
rect 11498 -35466 11532 -35450
rect 11040 -35469 11145 -35466
rect 12914 -35634 13427 -35618
rect 12914 -35668 12930 -35634
rect 12964 -35668 13184 -35634
rect 13410 -35668 13427 -35634
rect 12886 -35727 12920 -35711
rect 12784 -35746 12818 -35730
rect 7182 -35822 7198 -35788
rect 7232 -35822 7248 -35788
rect 7374 -35822 7390 -35788
rect 7424 -35822 7440 -35788
rect 7566 -35822 7582 -35788
rect 7616 -35822 7632 -35788
rect 7758 -35822 7774 -35788
rect 7808 -35822 7824 -35788
rect 8130 -35822 8146 -35788
rect 8180 -35822 8196 -35788
rect 8322 -35822 8338 -35788
rect 8372 -35822 8388 -35788
rect 8514 -35822 8530 -35788
rect 8564 -35822 8580 -35788
rect 8706 -35822 8722 -35788
rect 8756 -35822 8772 -35788
rect 9066 -35822 9082 -35788
rect 9116 -35822 9132 -35788
rect 9258 -35822 9274 -35788
rect 9308 -35822 9324 -35788
rect 9450 -35822 9466 -35788
rect 9500 -35822 9516 -35788
rect 9642 -35822 9658 -35788
rect 9692 -35822 9708 -35788
rect 9997 -35821 10013 -35787
rect 10047 -35821 10063 -35787
rect 10189 -35821 10205 -35787
rect 10239 -35821 10255 -35787
rect 10381 -35821 10397 -35787
rect 10431 -35821 10447 -35787
rect 10573 -35821 10589 -35787
rect 10623 -35821 10639 -35787
rect 10924 -35822 10940 -35788
rect 10974 -35822 10990 -35788
rect 11116 -35822 11132 -35788
rect 11166 -35822 11182 -35788
rect 11308 -35822 11324 -35788
rect 11358 -35822 11374 -35788
rect 11500 -35822 11516 -35788
rect 11550 -35822 11566 -35788
rect 7150 -35881 7184 -35865
rect 7246 -35876 7280 -35865
rect 7150 -36195 7184 -36179
rect 7246 -36195 7280 -36179
rect 7342 -35881 7376 -35865
rect 7342 -36195 7376 -36179
rect 7438 -35876 7472 -35865
rect 7534 -35881 7568 -35865
rect 7438 -36195 7472 -36179
rect 7534 -36195 7568 -36179
rect 7630 -35876 7664 -35865
rect 7726 -35881 7760 -35865
rect 7630 -36195 7664 -36179
rect 7726 -36195 7760 -36179
rect 7822 -35876 7856 -35865
rect 7918 -35881 7952 -35865
rect 7822 -36195 7856 -36179
rect 7918 -36195 7952 -36179
rect 8098 -35881 8132 -35865
rect 8194 -35876 8228 -35865
rect 8098 -36195 8132 -36179
rect 8194 -36195 8228 -36179
rect 8290 -35881 8324 -35865
rect 8290 -36195 8324 -36179
rect 8386 -35876 8420 -35865
rect 8482 -35881 8516 -35865
rect 8386 -36195 8420 -36179
rect 8482 -36195 8516 -36179
rect 8578 -35876 8612 -35865
rect 8674 -35881 8708 -35865
rect 8578 -36195 8612 -36179
rect 8674 -36195 8708 -36179
rect 8770 -35876 8804 -35865
rect 8866 -35881 8900 -35865
rect 8770 -36195 8804 -36179
rect 8866 -36195 8900 -36179
rect 9034 -35881 9068 -35865
rect 9130 -35876 9164 -35865
rect 9034 -36195 9068 -36179
rect 9130 -36195 9164 -36179
rect 9226 -35881 9260 -35865
rect 9226 -36195 9260 -36179
rect 9322 -35876 9356 -35865
rect 9418 -35881 9452 -35865
rect 9322 -36195 9356 -36179
rect 9418 -36195 9452 -36179
rect 9514 -35876 9548 -35865
rect 9610 -35881 9644 -35865
rect 9514 -36195 9548 -36179
rect 9610 -36195 9644 -36179
rect 9706 -35876 9740 -35865
rect 9802 -35881 9836 -35865
rect 9706 -36195 9740 -36179
rect 9802 -36195 9836 -36179
rect 9965 -35880 9999 -35864
rect 10061 -35875 10095 -35864
rect 9965 -36194 9999 -36178
rect 10061 -36194 10095 -36178
rect 10157 -35880 10191 -35864
rect 10157 -36194 10191 -36178
rect 10253 -35875 10287 -35864
rect 10349 -35880 10383 -35864
rect 10253 -36194 10287 -36178
rect 10349 -36194 10383 -36178
rect 10445 -35875 10479 -35864
rect 10541 -35880 10575 -35864
rect 10445 -36194 10479 -36178
rect 10541 -36194 10575 -36178
rect 10637 -35875 10671 -35864
rect 10733 -35880 10767 -35864
rect 10637 -36194 10671 -36178
rect 10733 -36194 10767 -36178
rect 10892 -35881 10926 -35865
rect 10988 -35876 11022 -35865
rect 10892 -36195 10926 -36179
rect 10988 -36195 11022 -36179
rect 11084 -35881 11118 -35865
rect 11084 -36195 11118 -36179
rect 11180 -35876 11214 -35865
rect 11276 -35881 11310 -35865
rect 11180 -36195 11214 -36179
rect 11276 -36195 11310 -36179
rect 11372 -35876 11406 -35865
rect 11468 -35881 11502 -35865
rect 11372 -36195 11406 -36179
rect 11468 -36195 11502 -36179
rect 11564 -35876 11598 -35865
rect 11660 -35881 11694 -35865
rect 11564 -36195 11598 -36179
rect 12784 -35894 12818 -35878
rect 12886 -35919 12920 -35903
rect 12974 -35727 13008 -35711
rect 12974 -35919 13008 -35903
rect 13136 -35727 13170 -35711
rect 13136 -35939 13170 -35921
rect 13232 -35721 13266 -35711
rect 13232 -35933 13266 -35917
rect 13328 -35727 13362 -35711
rect 13328 -35939 13362 -35921
rect 13424 -35721 13458 -35711
rect 13496 -35778 13530 -35762
rect 13496 -35885 13530 -35869
rect 13424 -35933 13458 -35917
rect 12914 -36013 13427 -35997
rect 12914 -36047 12930 -36013
rect 12964 -36047 13184 -36013
rect 13410 -36047 13427 -36013
rect 12886 -36106 12920 -36090
rect 11660 -36195 11694 -36179
rect 12784 -36125 12818 -36109
rect 7373 -36283 7389 -36248
rect 7677 -36283 7703 -36248
rect 8321 -36283 8337 -36248
rect 8625 -36283 8651 -36248
rect 9257 -36283 9273 -36248
rect 9561 -36283 9587 -36248
rect 10188 -36282 10204 -36247
rect 10492 -36282 10518 -36247
rect 11115 -36283 11131 -36248
rect 11419 -36283 11445 -36248
rect 12784 -36273 12818 -36257
rect 12886 -36298 12920 -36282
rect 12974 -36106 13008 -36090
rect 12974 -36298 13008 -36282
rect 13136 -36106 13170 -36090
rect 13136 -36318 13170 -36300
rect 13232 -36100 13266 -36090
rect 13232 -36312 13266 -36296
rect 13328 -36106 13362 -36090
rect 13328 -36318 13362 -36300
rect 13424 -36100 13458 -36090
rect 13496 -36157 13530 -36141
rect 13496 -36264 13530 -36248
rect 13424 -36312 13458 -36296
<< viali >>
rect 1841 6169 2963 6241
rect 3447 6169 4569 6241
rect 5151 6167 6273 6239
rect 1564 5398 1673 5495
rect 1807 5964 1841 6066
rect 1807 5569 1841 5671
rect 1903 5756 1937 5880
rect 1999 5964 2033 6066
rect 1999 5605 2033 5671
rect 2095 5756 2129 5880
rect 2191 5962 2225 6064
rect 2191 5605 2225 5665
rect 2287 5756 2321 5880
rect 2383 5961 2417 6063
rect 2383 5605 2417 5648
rect 2479 5756 2513 5880
rect 2575 5961 2609 6063
rect 2575 5605 2609 5665
rect 2671 5756 2705 5880
rect 2767 5961 2801 6063
rect 2767 5605 2801 5672
rect 2863 5755 2897 5879
rect 2959 5961 2993 6063
rect 2959 5605 2993 5672
rect 1905 5292 2038 5345
rect 3413 5964 3447 6066
rect 3413 5569 3447 5671
rect 3509 5756 3543 5880
rect 3605 5964 3639 6066
rect 3605 5605 3639 5671
rect 3701 5756 3735 5880
rect 3797 5962 3831 6064
rect 3797 5605 3831 5665
rect 3893 5756 3927 5880
rect 3989 5961 4023 6063
rect 3989 5605 4023 5648
rect 4085 5756 4119 5880
rect 4181 5961 4215 6063
rect 4181 5605 4215 5665
rect 4277 5756 4311 5880
rect 4373 5961 4407 6063
rect 4373 5605 4407 5672
rect 4469 5755 4503 5879
rect 4565 5961 4599 6063
rect 4565 5605 4599 5672
rect 2511 5300 2625 5353
rect 2745 5346 2825 5352
rect 2745 5291 2753 5346
rect 2753 5291 2818 5346
rect 2818 5291 2825 5346
rect 2745 5284 2825 5291
rect 2927 5126 2992 5181
rect 1807 4926 1841 5032
rect 1903 5032 1937 5047
rect 1903 5013 1937 5032
rect 1999 4926 2033 4946
rect 1999 4912 2033 4926
rect 2095 5032 2129 5047
rect 2095 5013 2129 5032
rect 2191 4926 2225 4946
rect 2191 4912 2225 4926
rect 2287 5032 2321 5046
rect 2287 5012 2321 5032
rect 2383 4926 2417 4946
rect 2383 4912 2417 4926
rect 2479 5032 2513 5047
rect 2479 5013 2513 5032
rect 2575 4926 2609 4946
rect 2575 4912 2609 4926
rect 2671 5032 2705 5047
rect 2671 5013 2705 5032
rect 2767 4926 2801 4946
rect 2767 4912 2801 4926
rect 2863 5032 2897 5047
rect 2863 5013 2897 5032
rect 2959 4926 2993 5032
rect 3177 5371 3286 5468
rect 3511 5292 3644 5345
rect 4117 5300 4231 5353
rect 4351 5346 4431 5352
rect 4351 5291 4359 5346
rect 4359 5291 4424 5346
rect 4424 5291 4431 5346
rect 4351 5284 4431 5291
rect 4533 5126 4598 5181
rect 3413 4926 3447 5032
rect 3509 5032 3543 5047
rect 3509 5013 3543 5032
rect 3605 4926 3639 4946
rect 3605 4912 3639 4926
rect 3701 5032 3735 5047
rect 3701 5013 3735 5032
rect 3797 4926 3831 4946
rect 3797 4912 3831 4926
rect 3893 5032 3927 5046
rect 3893 5012 3927 5032
rect 3989 4926 4023 4946
rect 3989 4912 4023 4926
rect 4085 5032 4119 5047
rect 4085 5013 4119 5032
rect 4181 4926 4215 4946
rect 4181 4912 4215 4926
rect 4277 5032 4311 5047
rect 4277 5013 4311 5032
rect 4373 4926 4407 4946
rect 4373 4912 4407 4926
rect 4469 5032 4503 5047
rect 4469 5013 4503 5032
rect 4565 4926 4599 5032
rect 4861 5516 4970 5613
rect 5117 5962 5151 6064
rect 5117 5567 5151 5669
rect 5213 5754 5247 5878
rect 5309 5962 5343 6064
rect 5309 5603 5343 5669
rect 5405 5754 5439 5878
rect 5501 5960 5535 6062
rect 5501 5603 5535 5663
rect 5597 5754 5631 5878
rect 5693 5959 5727 6061
rect 5693 5603 5727 5646
rect 5789 5754 5823 5878
rect 5885 5959 5919 6061
rect 5885 5603 5919 5663
rect 5981 5754 6015 5878
rect 6077 5959 6111 6061
rect 6077 5603 6111 5670
rect 6173 5753 6207 5877
rect 6269 5959 6303 6061
rect 6269 5603 6303 5670
rect 5215 5290 5348 5343
rect 6967 5507 7536 5554
rect 7872 5497 7963 5531
rect 5821 5298 5935 5351
rect 6055 5344 6135 5350
rect 6055 5289 6063 5344
rect 6063 5289 6128 5344
rect 6128 5289 6135 5344
rect 6055 5282 6135 5289
rect 6237 5124 6302 5179
rect 5117 4924 5151 5030
rect 5213 5030 5247 5045
rect 5213 5011 5247 5030
rect 5309 4924 5343 4944
rect 5309 4910 5343 4924
rect 5405 5030 5439 5045
rect 5405 5011 5439 5030
rect 5501 4924 5535 4944
rect 5501 4910 5535 4924
rect 5597 5030 5631 5044
rect 5597 5010 5631 5030
rect 5693 4924 5727 4944
rect 5693 4910 5727 4924
rect 5789 5030 5823 5045
rect 5789 5011 5823 5030
rect 5885 4924 5919 4944
rect 5885 4910 5919 4924
rect 5981 5030 6015 5045
rect 5981 5011 6015 5030
rect 6077 4924 6111 4944
rect 6077 4910 6111 4924
rect 6173 5030 6207 5045
rect 6173 5011 6207 5030
rect 6269 4924 6303 5030
rect 6951 5429 6985 5435
rect 6951 5355 6985 5429
rect 7047 5239 7081 5313
rect 7047 5233 7081 5239
rect 7143 5429 7177 5435
rect 7143 5355 7177 5429
rect 7239 5239 7273 5313
rect 7239 5233 7273 5239
rect 7335 5429 7369 5435
rect 7335 5355 7369 5429
rect 7431 5239 7465 5313
rect 7431 5233 7465 5239
rect 7527 5429 7561 5435
rect 7527 5355 7561 5429
rect 7815 5425 7821 5459
rect 7821 5425 7894 5459
rect 7728 5185 7762 5411
rect 7938 5329 8015 5363
rect 7815 5233 7821 5267
rect 7821 5233 7894 5267
rect 7017 5145 7051 5180
rect 7306 5145 7340 5180
rect 7101 5021 7135 5056
rect 7185 5051 7561 5085
rect 7938 5137 8015 5171
rect 7821 4975 7997 5009
rect 7728 4931 7762 4965
rect 1841 4792 2964 4838
rect 7185 4859 7561 4893
rect 7821 4887 7997 4921
rect 3447 4792 4570 4838
rect 5151 4790 6274 4836
rect 7200 4787 7535 4821
rect 7840 4785 7972 4819
rect -24000 4445 -22878 4517
rect -20709 4445 -19587 4517
rect -17418 4445 -16296 4517
rect -14127 4445 -13005 4517
rect -10836 4445 -9714 4517
rect -7546 4445 -6424 4517
rect -4255 4445 -3133 4517
rect -964 4445 158 4517
rect -24030 4237 -23996 4339
rect -24030 3881 -23996 3948
rect -23934 4031 -23900 4155
rect -23838 4237 -23804 4339
rect -23838 3881 -23804 3948
rect -23742 4032 -23708 4156
rect -23646 4237 -23612 4339
rect -23646 3881 -23612 3941
rect -23550 4032 -23516 4156
rect -23454 4237 -23420 4339
rect -23454 3881 -23420 3924
rect -23358 4032 -23324 4156
rect -23262 4238 -23228 4340
rect -23262 3881 -23228 3941
rect -23166 4032 -23132 4156
rect -23070 4240 -23036 4342
rect -23070 3881 -23036 3947
rect -22974 4032 -22940 4156
rect -22878 4240 -22844 4342
rect -22878 3845 -22844 3947
rect -23862 3622 -23782 3628
rect -23862 3567 -23855 3622
rect -23855 3567 -23790 3622
rect -23790 3567 -23782 3622
rect -23862 3560 -23782 3567
rect -23662 3576 -23548 3629
rect -24029 3402 -23964 3457
rect -23075 3568 -22942 3621
rect -24030 3202 -23996 3308
rect -23934 3308 -23900 3323
rect -23934 3289 -23900 3308
rect -23838 3202 -23804 3222
rect -23838 3188 -23804 3202
rect -23742 3308 -23708 3323
rect -23742 3289 -23708 3308
rect -23646 3202 -23612 3222
rect -23646 3188 -23612 3202
rect -23550 3308 -23516 3323
rect -23550 3289 -23516 3308
rect -23454 3202 -23420 3222
rect -23454 3188 -23420 3202
rect -23358 3308 -23324 3322
rect -23358 3288 -23324 3308
rect -23262 3202 -23228 3222
rect -23262 3188 -23228 3202
rect -23166 3308 -23132 3323
rect -23166 3289 -23132 3308
rect -23070 3202 -23036 3222
rect -23070 3188 -23036 3202
rect -22974 3308 -22940 3323
rect -22974 3289 -22940 3308
rect -22878 3202 -22844 3308
rect -22637 3624 -22517 3766
rect -20739 4237 -20705 4339
rect -20739 3881 -20705 3948
rect -20643 4031 -20609 4155
rect -20547 4237 -20513 4339
rect -20547 3881 -20513 3948
rect -20451 4032 -20417 4156
rect -20355 4237 -20321 4339
rect -20355 3881 -20321 3941
rect -20259 4032 -20225 4156
rect -20163 4237 -20129 4339
rect -20163 3881 -20129 3924
rect -20067 4032 -20033 4156
rect -19971 4238 -19937 4340
rect -19971 3881 -19937 3941
rect -19875 4032 -19841 4156
rect -19779 4240 -19745 4342
rect -19779 3881 -19745 3947
rect -19683 4032 -19649 4156
rect -19587 4240 -19553 4342
rect -19587 3845 -19553 3947
rect -20571 3622 -20491 3628
rect -20571 3567 -20564 3622
rect -20564 3567 -20499 3622
rect -20499 3567 -20491 3622
rect -20571 3560 -20491 3567
rect -20371 3576 -20257 3629
rect -20738 3402 -20673 3457
rect -19784 3568 -19651 3621
rect -20739 3202 -20705 3308
rect -20643 3308 -20609 3323
rect -20643 3289 -20609 3308
rect -20547 3202 -20513 3222
rect -20547 3188 -20513 3202
rect -20451 3308 -20417 3323
rect -20451 3289 -20417 3308
rect -20355 3202 -20321 3222
rect -20355 3188 -20321 3202
rect -20259 3308 -20225 3323
rect -20259 3289 -20225 3308
rect -20163 3202 -20129 3222
rect -20163 3188 -20129 3202
rect -20067 3308 -20033 3322
rect -20067 3288 -20033 3308
rect -19971 3202 -19937 3222
rect -19971 3188 -19937 3202
rect -19875 3308 -19841 3323
rect -19875 3289 -19841 3308
rect -19779 3202 -19745 3222
rect -19779 3188 -19745 3202
rect -19683 3308 -19649 3323
rect -19683 3289 -19649 3308
rect -19587 3202 -19553 3308
rect -19346 3624 -19226 3766
rect -17448 4237 -17414 4339
rect -17448 3881 -17414 3948
rect -17352 4031 -17318 4155
rect -17256 4237 -17222 4339
rect -17256 3881 -17222 3948
rect -17160 4032 -17126 4156
rect -17064 4237 -17030 4339
rect -17064 3881 -17030 3941
rect -16968 4032 -16934 4156
rect -16872 4237 -16838 4339
rect -16872 3881 -16838 3924
rect -16776 4032 -16742 4156
rect -16680 4238 -16646 4340
rect -16680 3881 -16646 3941
rect -16584 4032 -16550 4156
rect -16488 4240 -16454 4342
rect -16488 3881 -16454 3947
rect -16392 4032 -16358 4156
rect -16296 4240 -16262 4342
rect -16296 3845 -16262 3947
rect -17280 3622 -17200 3628
rect -17280 3567 -17273 3622
rect -17273 3567 -17208 3622
rect -17208 3567 -17200 3622
rect -17280 3560 -17200 3567
rect -17080 3576 -16966 3629
rect -17447 3402 -17382 3457
rect -16493 3568 -16360 3621
rect -17448 3202 -17414 3308
rect -17352 3308 -17318 3323
rect -17352 3289 -17318 3308
rect -17256 3202 -17222 3222
rect -17256 3188 -17222 3202
rect -17160 3308 -17126 3323
rect -17160 3289 -17126 3308
rect -17064 3202 -17030 3222
rect -17064 3188 -17030 3202
rect -16968 3308 -16934 3323
rect -16968 3289 -16934 3308
rect -16872 3202 -16838 3222
rect -16872 3188 -16838 3202
rect -16776 3308 -16742 3322
rect -16776 3288 -16742 3308
rect -16680 3202 -16646 3222
rect -16680 3188 -16646 3202
rect -16584 3308 -16550 3323
rect -16584 3289 -16550 3308
rect -16488 3202 -16454 3222
rect -16488 3188 -16454 3202
rect -16392 3308 -16358 3323
rect -16392 3289 -16358 3308
rect -16296 3202 -16262 3308
rect -16055 3624 -15935 3766
rect -14157 4237 -14123 4339
rect -14157 3881 -14123 3948
rect -14061 4031 -14027 4155
rect -13965 4237 -13931 4339
rect -13965 3881 -13931 3948
rect -13869 4032 -13835 4156
rect -13773 4237 -13739 4339
rect -13773 3881 -13739 3941
rect -13677 4032 -13643 4156
rect -13581 4237 -13547 4339
rect -13581 3881 -13547 3924
rect -13485 4032 -13451 4156
rect -13389 4238 -13355 4340
rect -13389 3881 -13355 3941
rect -13293 4032 -13259 4156
rect -13197 4240 -13163 4342
rect -13197 3881 -13163 3947
rect -13101 4032 -13067 4156
rect -13005 4240 -12971 4342
rect -13005 3845 -12971 3947
rect -13989 3622 -13909 3628
rect -13989 3567 -13982 3622
rect -13982 3567 -13917 3622
rect -13917 3567 -13909 3622
rect -13989 3560 -13909 3567
rect -13789 3576 -13675 3629
rect -14156 3402 -14091 3457
rect -13202 3568 -13069 3621
rect -14157 3202 -14123 3308
rect -14061 3308 -14027 3323
rect -14061 3289 -14027 3308
rect -13965 3202 -13931 3222
rect -13965 3188 -13931 3202
rect -13869 3308 -13835 3323
rect -13869 3289 -13835 3308
rect -13773 3202 -13739 3222
rect -13773 3188 -13739 3202
rect -13677 3308 -13643 3323
rect -13677 3289 -13643 3308
rect -13581 3202 -13547 3222
rect -13581 3188 -13547 3202
rect -13485 3308 -13451 3322
rect -13485 3288 -13451 3308
rect -13389 3202 -13355 3222
rect -13389 3188 -13355 3202
rect -13293 3308 -13259 3323
rect -13293 3289 -13259 3308
rect -13197 3202 -13163 3222
rect -13197 3188 -13163 3202
rect -13101 3308 -13067 3323
rect -13101 3289 -13067 3308
rect -13005 3202 -12971 3308
rect -12764 3624 -12644 3766
rect -10866 4237 -10832 4339
rect -10866 3881 -10832 3948
rect -10770 4031 -10736 4155
rect -10674 4237 -10640 4339
rect -10674 3881 -10640 3948
rect -10578 4032 -10544 4156
rect -10482 4237 -10448 4339
rect -10482 3881 -10448 3941
rect -10386 4032 -10352 4156
rect -10290 4237 -10256 4339
rect -10290 3881 -10256 3924
rect -10194 4032 -10160 4156
rect -10098 4238 -10064 4340
rect -10098 3881 -10064 3941
rect -10002 4032 -9968 4156
rect -9906 4240 -9872 4342
rect -9906 3881 -9872 3947
rect -9810 4032 -9776 4156
rect -9714 4240 -9680 4342
rect -9714 3845 -9680 3947
rect -10698 3622 -10618 3628
rect -10698 3567 -10691 3622
rect -10691 3567 -10626 3622
rect -10626 3567 -10618 3622
rect -10698 3560 -10618 3567
rect -10498 3576 -10384 3629
rect -10865 3402 -10800 3457
rect -9911 3568 -9778 3621
rect -10866 3202 -10832 3308
rect -10770 3308 -10736 3323
rect -10770 3289 -10736 3308
rect -10674 3202 -10640 3222
rect -10674 3188 -10640 3202
rect -10578 3308 -10544 3323
rect -10578 3289 -10544 3308
rect -10482 3202 -10448 3222
rect -10482 3188 -10448 3202
rect -10386 3308 -10352 3323
rect -10386 3289 -10352 3308
rect -10290 3202 -10256 3222
rect -10290 3188 -10256 3202
rect -10194 3308 -10160 3322
rect -10194 3288 -10160 3308
rect -10098 3202 -10064 3222
rect -10098 3188 -10064 3202
rect -10002 3308 -9968 3323
rect -10002 3289 -9968 3308
rect -9906 3202 -9872 3222
rect -9906 3188 -9872 3202
rect -9810 3308 -9776 3323
rect -9810 3289 -9776 3308
rect -9714 3202 -9680 3308
rect -9473 3624 -9353 3766
rect -7576 4237 -7542 4339
rect -7576 3881 -7542 3948
rect -7480 4031 -7446 4155
rect -7384 4237 -7350 4339
rect -7384 3881 -7350 3948
rect -7288 4032 -7254 4156
rect -7192 4237 -7158 4339
rect -7192 3881 -7158 3941
rect -7096 4032 -7062 4156
rect -7000 4237 -6966 4339
rect -7000 3881 -6966 3924
rect -6904 4032 -6870 4156
rect -6808 4238 -6774 4340
rect -6808 3881 -6774 3941
rect -6712 4032 -6678 4156
rect -6616 4240 -6582 4342
rect -6616 3881 -6582 3947
rect -6520 4032 -6486 4156
rect -6424 4240 -6390 4342
rect -6424 3845 -6390 3947
rect -7408 3622 -7328 3628
rect -7408 3567 -7401 3622
rect -7401 3567 -7336 3622
rect -7336 3567 -7328 3622
rect -7408 3560 -7328 3567
rect -7208 3576 -7094 3629
rect -7575 3402 -7510 3457
rect -6621 3568 -6488 3621
rect -7576 3202 -7542 3308
rect -7480 3308 -7446 3323
rect -7480 3289 -7446 3308
rect -7384 3202 -7350 3222
rect -7384 3188 -7350 3202
rect -7288 3308 -7254 3323
rect -7288 3289 -7254 3308
rect -7192 3202 -7158 3222
rect -7192 3188 -7158 3202
rect -7096 3308 -7062 3323
rect -7096 3289 -7062 3308
rect -7000 3202 -6966 3222
rect -7000 3188 -6966 3202
rect -6904 3308 -6870 3322
rect -6904 3288 -6870 3308
rect -6808 3202 -6774 3222
rect -6808 3188 -6774 3202
rect -6712 3308 -6678 3323
rect -6712 3289 -6678 3308
rect -6616 3202 -6582 3222
rect -6616 3188 -6582 3202
rect -6520 3308 -6486 3323
rect -6520 3289 -6486 3308
rect -6424 3202 -6390 3308
rect -6183 3624 -6063 3766
rect -4285 4237 -4251 4339
rect -4285 3881 -4251 3948
rect -4189 4031 -4155 4155
rect -4093 4237 -4059 4339
rect -4093 3881 -4059 3948
rect -3997 4032 -3963 4156
rect -3901 4237 -3867 4339
rect -3901 3881 -3867 3941
rect -3805 4032 -3771 4156
rect -3709 4237 -3675 4339
rect -3709 3881 -3675 3924
rect -3613 4032 -3579 4156
rect -3517 4238 -3483 4340
rect -3517 3881 -3483 3941
rect -3421 4032 -3387 4156
rect -3325 4240 -3291 4342
rect -3325 3881 -3291 3947
rect -3229 4032 -3195 4156
rect -3133 4240 -3099 4342
rect -3133 3845 -3099 3947
rect -4117 3622 -4037 3628
rect -4117 3567 -4110 3622
rect -4110 3567 -4045 3622
rect -4045 3567 -4037 3622
rect -4117 3560 -4037 3567
rect -3917 3576 -3803 3629
rect -4284 3402 -4219 3457
rect -3330 3568 -3197 3621
rect -4285 3202 -4251 3308
rect -4189 3308 -4155 3323
rect -4189 3289 -4155 3308
rect -4093 3202 -4059 3222
rect -4093 3188 -4059 3202
rect -3997 3308 -3963 3323
rect -3997 3289 -3963 3308
rect -3901 3202 -3867 3222
rect -3901 3188 -3867 3202
rect -3805 3308 -3771 3323
rect -3805 3289 -3771 3308
rect -3709 3202 -3675 3222
rect -3709 3188 -3675 3202
rect -3613 3308 -3579 3322
rect -3613 3288 -3579 3308
rect -3517 3202 -3483 3222
rect -3517 3188 -3483 3202
rect -3421 3308 -3387 3323
rect -3421 3289 -3387 3308
rect -3325 3202 -3291 3222
rect -3325 3188 -3291 3202
rect -3229 3308 -3195 3323
rect -3229 3289 -3195 3308
rect -3133 3202 -3099 3308
rect -2892 3624 -2772 3766
rect -994 4237 -960 4339
rect -994 3881 -960 3948
rect -898 4031 -864 4155
rect -802 4237 -768 4339
rect -802 3881 -768 3948
rect -706 4032 -672 4156
rect -610 4237 -576 4339
rect -610 3881 -576 3941
rect -514 4032 -480 4156
rect -418 4237 -384 4339
rect -418 3881 -384 3924
rect -322 4032 -288 4156
rect -226 4238 -192 4340
rect -226 3881 -192 3941
rect -130 4032 -96 4156
rect -34 4240 0 4342
rect -34 3881 0 3947
rect 62 4032 96 4156
rect 158 4240 192 4342
rect 158 3845 192 3947
rect 5721 3949 5812 3983
rect 6161 3949 6252 3983
rect 6601 3949 6692 3983
rect -826 3622 -746 3628
rect -826 3567 -819 3622
rect -819 3567 -754 3622
rect -754 3567 -746 3622
rect -826 3560 -746 3567
rect -626 3576 -512 3629
rect 5664 3877 5670 3911
rect 5670 3877 5743 3911
rect -993 3402 -928 3457
rect -39 3568 94 3621
rect -994 3202 -960 3308
rect -898 3308 -864 3323
rect -898 3289 -864 3308
rect -802 3202 -768 3222
rect -802 3188 -768 3202
rect -706 3308 -672 3323
rect -706 3289 -672 3308
rect -610 3202 -576 3222
rect -610 3188 -576 3202
rect -514 3308 -480 3323
rect -514 3289 -480 3308
rect -418 3202 -384 3222
rect -418 3188 -384 3202
rect -322 3308 -288 3322
rect -322 3288 -288 3308
rect -226 3202 -192 3222
rect -226 3188 -192 3202
rect -130 3308 -96 3323
rect -130 3289 -96 3308
rect -34 3202 0 3222
rect -34 3188 0 3202
rect 62 3308 96 3323
rect 62 3289 96 3308
rect 158 3202 192 3308
rect 399 3624 519 3766
rect 5577 3637 5611 3863
rect 6104 3877 6110 3911
rect 6110 3877 6183 3911
rect 5787 3781 5864 3815
rect 5664 3685 5670 3719
rect 5670 3685 5743 3719
rect 6017 3637 6051 3863
rect 6544 3877 6550 3911
rect 6550 3877 6623 3911
rect 6227 3781 6304 3815
rect 6104 3685 6110 3719
rect 6110 3685 6183 3719
rect 5787 3589 5864 3623
rect 5670 3427 5846 3461
rect 5577 3383 5611 3417
rect 6457 3637 6491 3863
rect 6667 3781 6744 3815
rect 6544 3685 6550 3719
rect 6550 3685 6623 3719
rect 6227 3589 6304 3623
rect 6110 3427 6286 3461
rect 6017 3383 6051 3417
rect 5670 3339 5846 3373
rect 6667 3589 6744 3623
rect 6550 3427 6726 3461
rect 6457 3383 6491 3417
rect 6110 3339 6286 3373
rect 6550 3339 6726 3373
rect 7389 3276 7677 3311
rect 8337 3276 8625 3311
rect 9273 3276 9561 3311
rect 10204 3276 10492 3311
rect 11131 3276 11419 3311
rect 5689 3237 5821 3271
rect 6129 3237 6261 3271
rect 6569 3237 6701 3271
rect -24001 3068 -22878 3114
rect -20710 3068 -19587 3114
rect -17419 3068 -16296 3114
rect -14128 3068 -13005 3114
rect -10837 3068 -9714 3114
rect -7547 3068 -6424 3114
rect -4256 3068 -3133 3114
rect -965 3068 158 3114
rect 7150 3094 7184 3204
rect 7245 2909 7246 3016
rect 7246 2909 7280 3016
rect 7245 2904 7280 2909
rect 7342 3094 7376 3204
rect 7534 3094 7568 3204
rect 7438 2909 7472 3016
rect 7472 2909 7473 3016
rect 7438 2904 7473 2909
rect 7726 3094 7760 3204
rect 7630 2909 7664 3016
rect 7664 2909 7665 3016
rect 7630 2904 7665 2909
rect 7918 3094 7952 3204
rect 7822 2909 7856 3016
rect 7856 2909 7857 3016
rect 7822 2904 7857 2909
rect 8098 3094 8132 3204
rect 8193 2909 8194 3016
rect 8194 2909 8228 3016
rect 8193 2904 8228 2909
rect 8290 3094 8324 3204
rect 8482 3094 8516 3204
rect 8386 2909 8420 3016
rect 8420 2909 8421 3016
rect 8386 2904 8421 2909
rect 8674 3094 8708 3204
rect 8578 2909 8612 3016
rect 8612 2909 8613 3016
rect 8578 2904 8613 2909
rect 8866 3094 8900 3204
rect 8770 2909 8804 3016
rect 8804 2909 8805 3016
rect 8770 2904 8805 2909
rect 9034 3094 9068 3204
rect 9129 2909 9130 3016
rect 9130 2909 9164 3016
rect 9129 2904 9164 2909
rect 9226 3094 9260 3204
rect 9418 3094 9452 3204
rect 9322 2909 9356 3016
rect 9356 2909 9357 3016
rect 9322 2904 9357 2909
rect 9610 3094 9644 3204
rect 9514 2909 9548 3016
rect 9548 2909 9549 3016
rect 9514 2904 9549 2909
rect 9802 3094 9836 3204
rect 9706 2909 9740 3016
rect 9740 2909 9741 3016
rect 9706 2904 9741 2909
rect 9965 3094 9999 3204
rect 10060 2909 10061 3016
rect 10061 2909 10095 3016
rect 10060 2904 10095 2909
rect 10157 3094 10191 3204
rect 10349 3094 10383 3204
rect 10253 2909 10287 3016
rect 10287 2909 10288 3016
rect 10253 2904 10288 2909
rect 10541 3094 10575 3204
rect 10445 2909 10479 3016
rect 10479 2909 10480 3016
rect 10445 2904 10480 2909
rect 10733 3094 10767 3204
rect 10637 2909 10671 3016
rect 10671 2909 10672 3016
rect 10637 2904 10672 2909
rect 10892 3094 10926 3204
rect 10987 2909 10988 3016
rect 10988 2909 11022 3016
rect 10987 2904 11022 2909
rect 11084 3094 11118 3204
rect 11276 3094 11310 3204
rect 11180 2909 11214 3016
rect 11214 2909 11215 3016
rect 11180 2904 11215 2909
rect 11468 3094 11502 3204
rect 11372 2909 11406 3016
rect 11406 2909 11407 3016
rect 11372 2904 11407 2909
rect 11660 3094 11694 3204
rect 11564 2909 11598 3016
rect 11598 2909 11599 3016
rect 11564 2904 11599 2909
rect 7198 2816 7232 2850
rect 7390 2816 7424 2850
rect 7582 2816 7616 2850
rect 7774 2816 7808 2850
rect 8146 2816 8180 2850
rect 8338 2816 8372 2850
rect 8530 2816 8564 2850
rect 8722 2816 8756 2850
rect 9082 2816 9116 2850
rect 9274 2816 9308 2850
rect 9466 2816 9500 2850
rect 9658 2816 9692 2850
rect 10013 2816 10047 2850
rect 10205 2816 10239 2850
rect 10397 2816 10431 2850
rect 10589 2816 10623 2850
rect 10940 2816 10974 2850
rect 11132 2816 11166 2850
rect 11324 2816 11358 2850
rect 11516 2816 11550 2850
rect -24670 2661 -23548 2733
rect -23111 2661 -21989 2733
rect -21379 2661 -20257 2733
rect -19820 2661 -18698 2733
rect -18088 2661 -16966 2733
rect -16529 2661 -15407 2733
rect -14797 2661 -13675 2733
rect -13238 2661 -12116 2733
rect -11506 2661 -10384 2733
rect -9947 2661 -8825 2733
rect -8216 2661 -7094 2733
rect -6657 2661 -5535 2733
rect -4925 2661 -3803 2733
rect -3366 2661 -2244 2733
rect -1634 2661 -512 2733
rect -75 2661 1047 2733
rect -24704 2456 -24670 2558
rect -24704 2061 -24670 2163
rect -24608 2248 -24574 2372
rect -24512 2456 -24478 2558
rect -24512 2097 -24478 2163
rect -24416 2248 -24382 2372
rect -24320 2454 -24286 2556
rect -24320 2097 -24286 2157
rect -24224 2248 -24190 2372
rect -24128 2453 -24094 2555
rect -24128 2097 -24094 2140
rect -24032 2248 -23998 2372
rect -23936 2453 -23902 2555
rect -23936 2097 -23902 2157
rect -23840 2248 -23806 2372
rect -23744 2453 -23710 2555
rect -23744 2097 -23710 2164
rect -23648 2247 -23614 2371
rect -23552 2453 -23518 2555
rect -23552 2097 -23518 2164
rect -24921 1828 -24874 1938
rect -24606 1784 -24473 1837
rect -23145 2456 -23111 2558
rect -23145 2061 -23111 2163
rect -23049 2248 -23015 2372
rect -22953 2456 -22919 2558
rect -22953 2097 -22919 2163
rect -22857 2248 -22823 2372
rect -22761 2454 -22727 2556
rect -22761 2097 -22727 2157
rect -22665 2248 -22631 2372
rect -22569 2453 -22535 2555
rect -22569 2097 -22535 2140
rect -22473 2248 -22439 2372
rect -22377 2453 -22343 2555
rect -22377 2097 -22343 2157
rect -22281 2248 -22247 2372
rect -22185 2453 -22151 2555
rect -22185 2097 -22151 2164
rect -22089 2247 -22055 2371
rect -21993 2453 -21959 2555
rect -21993 2097 -21959 2164
rect -24000 1792 -23886 1845
rect -23766 1838 -23686 1844
rect -23766 1783 -23758 1838
rect -23758 1783 -23693 1838
rect -23693 1783 -23686 1838
rect -23766 1776 -23686 1783
rect -23584 1618 -23519 1673
rect -24704 1418 -24670 1524
rect -24608 1524 -24574 1539
rect -24608 1505 -24574 1524
rect -24512 1418 -24478 1438
rect -24512 1404 -24478 1418
rect -24416 1524 -24382 1539
rect -24416 1505 -24382 1524
rect -24320 1418 -24286 1438
rect -24320 1404 -24286 1418
rect -24224 1524 -24190 1538
rect -24224 1504 -24190 1524
rect -24128 1418 -24094 1438
rect -24128 1404 -24094 1418
rect -24032 1524 -23998 1539
rect -24032 1505 -23998 1524
rect -23936 1418 -23902 1438
rect -23936 1404 -23902 1418
rect -23840 1524 -23806 1539
rect -23840 1505 -23806 1524
rect -23744 1418 -23710 1438
rect -23744 1404 -23710 1418
rect -23648 1524 -23614 1539
rect -23648 1505 -23614 1524
rect -23552 1418 -23518 1524
rect -23364 1790 -23291 1893
rect -23047 1784 -22914 1837
rect -21413 2456 -21379 2558
rect -21413 2061 -21379 2163
rect -21317 2248 -21283 2372
rect -21221 2456 -21187 2558
rect -21221 2097 -21187 2163
rect -21125 2248 -21091 2372
rect -21029 2454 -20995 2556
rect -21029 2097 -20995 2157
rect -20933 2248 -20899 2372
rect -20837 2453 -20803 2555
rect -20837 2097 -20803 2140
rect -20741 2248 -20707 2372
rect -20645 2453 -20611 2555
rect -20645 2097 -20611 2157
rect -20549 2248 -20515 2372
rect -20453 2453 -20419 2555
rect -20453 2097 -20419 2164
rect -20357 2247 -20323 2371
rect -20261 2453 -20227 2555
rect -20261 2097 -20227 2164
rect -22441 1792 -22327 1845
rect -22207 1838 -22127 1844
rect -22207 1783 -22199 1838
rect -22199 1783 -22134 1838
rect -22134 1783 -22127 1838
rect -22207 1776 -22127 1783
rect -22025 1618 -21960 1673
rect -23145 1418 -23111 1524
rect -23049 1524 -23015 1539
rect -23049 1505 -23015 1524
rect -22953 1418 -22919 1438
rect -22953 1404 -22919 1418
rect -22857 1524 -22823 1539
rect -22857 1505 -22823 1524
rect -22761 1418 -22727 1438
rect -22761 1404 -22727 1418
rect -22665 1524 -22631 1538
rect -22665 1504 -22631 1524
rect -22569 1418 -22535 1438
rect -22569 1404 -22535 1418
rect -22473 1524 -22439 1539
rect -22473 1505 -22439 1524
rect -22377 1418 -22343 1438
rect -22377 1404 -22343 1418
rect -22281 1524 -22247 1539
rect -22281 1505 -22247 1524
rect -22185 1418 -22151 1438
rect -22185 1404 -22151 1418
rect -22089 1524 -22055 1539
rect -22089 1505 -22055 1524
rect -21993 1418 -21959 1524
rect -21630 1828 -21583 1938
rect -21315 1784 -21182 1837
rect -19854 2456 -19820 2558
rect -19854 2061 -19820 2163
rect -19758 2248 -19724 2372
rect -19662 2456 -19628 2558
rect -19662 2097 -19628 2163
rect -19566 2248 -19532 2372
rect -19470 2454 -19436 2556
rect -19470 2097 -19436 2157
rect -19374 2248 -19340 2372
rect -19278 2453 -19244 2555
rect -19278 2097 -19244 2140
rect -19182 2248 -19148 2372
rect -19086 2453 -19052 2555
rect -19086 2097 -19052 2157
rect -18990 2248 -18956 2372
rect -18894 2453 -18860 2555
rect -18894 2097 -18860 2164
rect -18798 2247 -18764 2371
rect -18702 2453 -18668 2555
rect -18702 2097 -18668 2164
rect -20709 1792 -20595 1845
rect -20475 1838 -20395 1844
rect -20475 1783 -20467 1838
rect -20467 1783 -20402 1838
rect -20402 1783 -20395 1838
rect -20475 1776 -20395 1783
rect -20293 1618 -20228 1673
rect -21413 1418 -21379 1524
rect -21317 1524 -21283 1539
rect -21317 1505 -21283 1524
rect -21221 1418 -21187 1438
rect -21221 1404 -21187 1418
rect -21125 1524 -21091 1539
rect -21125 1505 -21091 1524
rect -21029 1418 -20995 1438
rect -21029 1404 -20995 1418
rect -20933 1524 -20899 1538
rect -20933 1504 -20899 1524
rect -20837 1418 -20803 1438
rect -20837 1404 -20803 1418
rect -20741 1524 -20707 1539
rect -20741 1505 -20707 1524
rect -20645 1418 -20611 1438
rect -20645 1404 -20611 1418
rect -20549 1524 -20515 1539
rect -20549 1505 -20515 1524
rect -20453 1418 -20419 1438
rect -20453 1404 -20419 1418
rect -20357 1524 -20323 1539
rect -20357 1505 -20323 1524
rect -20261 1418 -20227 1524
rect -20073 1790 -20000 1893
rect -19756 1784 -19623 1837
rect -18122 2456 -18088 2558
rect -18122 2061 -18088 2163
rect -18026 2248 -17992 2372
rect -17930 2456 -17896 2558
rect -17930 2097 -17896 2163
rect -17834 2248 -17800 2372
rect -17738 2454 -17704 2556
rect -17738 2097 -17704 2157
rect -17642 2248 -17608 2372
rect -17546 2453 -17512 2555
rect -17546 2097 -17512 2140
rect -17450 2248 -17416 2372
rect -17354 2453 -17320 2555
rect -17354 2097 -17320 2157
rect -17258 2248 -17224 2372
rect -17162 2453 -17128 2555
rect -17162 2097 -17128 2164
rect -17066 2247 -17032 2371
rect -16970 2453 -16936 2555
rect -16970 2097 -16936 2164
rect -19150 1792 -19036 1845
rect -18916 1838 -18836 1844
rect -18916 1783 -18908 1838
rect -18908 1783 -18843 1838
rect -18843 1783 -18836 1838
rect -18916 1776 -18836 1783
rect -18734 1618 -18669 1673
rect -19854 1418 -19820 1524
rect -19758 1524 -19724 1539
rect -19758 1505 -19724 1524
rect -19662 1418 -19628 1438
rect -19662 1404 -19628 1418
rect -19566 1524 -19532 1539
rect -19566 1505 -19532 1524
rect -19470 1418 -19436 1438
rect -19470 1404 -19436 1418
rect -19374 1524 -19340 1538
rect -19374 1504 -19340 1524
rect -19278 1418 -19244 1438
rect -19278 1404 -19244 1418
rect -19182 1524 -19148 1539
rect -19182 1505 -19148 1524
rect -19086 1418 -19052 1438
rect -19086 1404 -19052 1418
rect -18990 1524 -18956 1539
rect -18990 1505 -18956 1524
rect -18894 1418 -18860 1438
rect -18894 1404 -18860 1418
rect -18798 1524 -18764 1539
rect -18798 1505 -18764 1524
rect -18702 1418 -18668 1524
rect -18339 1828 -18292 1938
rect -18024 1784 -17891 1837
rect -16563 2456 -16529 2558
rect -16563 2061 -16529 2163
rect -16467 2248 -16433 2372
rect -16371 2456 -16337 2558
rect -16371 2097 -16337 2163
rect -16275 2248 -16241 2372
rect -16179 2454 -16145 2556
rect -16179 2097 -16145 2157
rect -16083 2248 -16049 2372
rect -15987 2453 -15953 2555
rect -15987 2097 -15953 2140
rect -15891 2248 -15857 2372
rect -15795 2453 -15761 2555
rect -15795 2097 -15761 2157
rect -15699 2248 -15665 2372
rect -15603 2453 -15569 2555
rect -15603 2097 -15569 2164
rect -15507 2247 -15473 2371
rect -15411 2453 -15377 2555
rect -15411 2097 -15377 2164
rect -17418 1792 -17304 1845
rect -17184 1838 -17104 1844
rect -17184 1783 -17176 1838
rect -17176 1783 -17111 1838
rect -17111 1783 -17104 1838
rect -17184 1776 -17104 1783
rect -17002 1618 -16937 1673
rect -18122 1418 -18088 1524
rect -18026 1524 -17992 1539
rect -18026 1505 -17992 1524
rect -17930 1418 -17896 1438
rect -17930 1404 -17896 1418
rect -17834 1524 -17800 1539
rect -17834 1505 -17800 1524
rect -17738 1418 -17704 1438
rect -17738 1404 -17704 1418
rect -17642 1524 -17608 1538
rect -17642 1504 -17608 1524
rect -17546 1418 -17512 1438
rect -17546 1404 -17512 1418
rect -17450 1524 -17416 1539
rect -17450 1505 -17416 1524
rect -17354 1418 -17320 1438
rect -17354 1404 -17320 1418
rect -17258 1524 -17224 1539
rect -17258 1505 -17224 1524
rect -17162 1418 -17128 1438
rect -17162 1404 -17128 1418
rect -17066 1524 -17032 1539
rect -17066 1505 -17032 1524
rect -16970 1418 -16936 1524
rect -16782 1790 -16709 1893
rect -16465 1784 -16332 1837
rect -14831 2456 -14797 2558
rect -14831 2061 -14797 2163
rect -14735 2248 -14701 2372
rect -14639 2456 -14605 2558
rect -14639 2097 -14605 2163
rect -14543 2248 -14509 2372
rect -14447 2454 -14413 2556
rect -14447 2097 -14413 2157
rect -14351 2248 -14317 2372
rect -14255 2453 -14221 2555
rect -14255 2097 -14221 2140
rect -14159 2248 -14125 2372
rect -14063 2453 -14029 2555
rect -14063 2097 -14029 2157
rect -13967 2248 -13933 2372
rect -13871 2453 -13837 2555
rect -13871 2097 -13837 2164
rect -13775 2247 -13741 2371
rect -13679 2453 -13645 2555
rect -13679 2097 -13645 2164
rect -15859 1792 -15745 1845
rect -15625 1838 -15545 1844
rect -15625 1783 -15617 1838
rect -15617 1783 -15552 1838
rect -15552 1783 -15545 1838
rect -15625 1776 -15545 1783
rect -15443 1618 -15378 1673
rect -16563 1418 -16529 1524
rect -16467 1524 -16433 1539
rect -16467 1505 -16433 1524
rect -16371 1418 -16337 1438
rect -16371 1404 -16337 1418
rect -16275 1524 -16241 1539
rect -16275 1505 -16241 1524
rect -16179 1418 -16145 1438
rect -16179 1404 -16145 1418
rect -16083 1524 -16049 1538
rect -16083 1504 -16049 1524
rect -15987 1418 -15953 1438
rect -15987 1404 -15953 1418
rect -15891 1524 -15857 1539
rect -15891 1505 -15857 1524
rect -15795 1418 -15761 1438
rect -15795 1404 -15761 1418
rect -15699 1524 -15665 1539
rect -15699 1505 -15665 1524
rect -15603 1418 -15569 1438
rect -15603 1404 -15569 1418
rect -15507 1524 -15473 1539
rect -15507 1505 -15473 1524
rect -15411 1418 -15377 1524
rect -15048 1828 -15001 1938
rect -14733 1784 -14600 1837
rect -13272 2456 -13238 2558
rect -13272 2061 -13238 2163
rect -13176 2248 -13142 2372
rect -13080 2456 -13046 2558
rect -13080 2097 -13046 2163
rect -12984 2248 -12950 2372
rect -12888 2454 -12854 2556
rect -12888 2097 -12854 2157
rect -12792 2248 -12758 2372
rect -12696 2453 -12662 2555
rect -12696 2097 -12662 2140
rect -12600 2248 -12566 2372
rect -12504 2453 -12470 2555
rect -12504 2097 -12470 2157
rect -12408 2248 -12374 2372
rect -12312 2453 -12278 2555
rect -12312 2097 -12278 2164
rect -12216 2247 -12182 2371
rect -12120 2453 -12086 2555
rect -12120 2097 -12086 2164
rect -14127 1792 -14013 1845
rect -13893 1838 -13813 1844
rect -13893 1783 -13885 1838
rect -13885 1783 -13820 1838
rect -13820 1783 -13813 1838
rect -13893 1776 -13813 1783
rect -13711 1618 -13646 1673
rect -14831 1418 -14797 1524
rect -14735 1524 -14701 1539
rect -14735 1505 -14701 1524
rect -14639 1418 -14605 1438
rect -14639 1404 -14605 1418
rect -14543 1524 -14509 1539
rect -14543 1505 -14509 1524
rect -14447 1418 -14413 1438
rect -14447 1404 -14413 1418
rect -14351 1524 -14317 1538
rect -14351 1504 -14317 1524
rect -14255 1418 -14221 1438
rect -14255 1404 -14221 1418
rect -14159 1524 -14125 1539
rect -14159 1505 -14125 1524
rect -14063 1418 -14029 1438
rect -14063 1404 -14029 1418
rect -13967 1524 -13933 1539
rect -13967 1505 -13933 1524
rect -13871 1418 -13837 1438
rect -13871 1404 -13837 1418
rect -13775 1524 -13741 1539
rect -13775 1505 -13741 1524
rect -13679 1418 -13645 1524
rect -13491 1790 -13418 1893
rect -13174 1784 -13041 1837
rect -11540 2456 -11506 2558
rect -11540 2061 -11506 2163
rect -11444 2248 -11410 2372
rect -11348 2456 -11314 2558
rect -11348 2097 -11314 2163
rect -11252 2248 -11218 2372
rect -11156 2454 -11122 2556
rect -11156 2097 -11122 2157
rect -11060 2248 -11026 2372
rect -10964 2453 -10930 2555
rect -10964 2097 -10930 2140
rect -10868 2248 -10834 2372
rect -10772 2453 -10738 2555
rect -10772 2097 -10738 2157
rect -10676 2248 -10642 2372
rect -10580 2453 -10546 2555
rect -10580 2097 -10546 2164
rect -10484 2247 -10450 2371
rect -10388 2453 -10354 2555
rect -10388 2097 -10354 2164
rect -12568 1792 -12454 1845
rect -12334 1838 -12254 1844
rect -12334 1783 -12326 1838
rect -12326 1783 -12261 1838
rect -12261 1783 -12254 1838
rect -12334 1776 -12254 1783
rect -12152 1618 -12087 1673
rect -13272 1418 -13238 1524
rect -13176 1524 -13142 1539
rect -13176 1505 -13142 1524
rect -13080 1418 -13046 1438
rect -13080 1404 -13046 1418
rect -12984 1524 -12950 1539
rect -12984 1505 -12950 1524
rect -12888 1418 -12854 1438
rect -12888 1404 -12854 1418
rect -12792 1524 -12758 1538
rect -12792 1504 -12758 1524
rect -12696 1418 -12662 1438
rect -12696 1404 -12662 1418
rect -12600 1524 -12566 1539
rect -12600 1505 -12566 1524
rect -12504 1418 -12470 1438
rect -12504 1404 -12470 1418
rect -12408 1524 -12374 1539
rect -12408 1505 -12374 1524
rect -12312 1418 -12278 1438
rect -12312 1404 -12278 1418
rect -12216 1524 -12182 1539
rect -12216 1505 -12182 1524
rect -12120 1418 -12086 1524
rect -11757 1828 -11710 1938
rect -11442 1784 -11309 1837
rect -9981 2456 -9947 2558
rect -9981 2061 -9947 2163
rect -9885 2248 -9851 2372
rect -9789 2456 -9755 2558
rect -9789 2097 -9755 2163
rect -9693 2248 -9659 2372
rect -9597 2454 -9563 2556
rect -9597 2097 -9563 2157
rect -9501 2248 -9467 2372
rect -9405 2453 -9371 2555
rect -9405 2097 -9371 2140
rect -9309 2248 -9275 2372
rect -9213 2453 -9179 2555
rect -9213 2097 -9179 2157
rect -9117 2248 -9083 2372
rect -9021 2453 -8987 2555
rect -9021 2097 -8987 2164
rect -8925 2247 -8891 2371
rect -8829 2453 -8795 2555
rect -8829 2097 -8795 2164
rect -10836 1792 -10722 1845
rect -10602 1838 -10522 1844
rect -10602 1783 -10594 1838
rect -10594 1783 -10529 1838
rect -10529 1783 -10522 1838
rect -10602 1776 -10522 1783
rect -10420 1618 -10355 1673
rect -11540 1418 -11506 1524
rect -11444 1524 -11410 1539
rect -11444 1505 -11410 1524
rect -11348 1418 -11314 1438
rect -11348 1404 -11314 1418
rect -11252 1524 -11218 1539
rect -11252 1505 -11218 1524
rect -11156 1418 -11122 1438
rect -11156 1404 -11122 1418
rect -11060 1524 -11026 1538
rect -11060 1504 -11026 1524
rect -10964 1418 -10930 1438
rect -10964 1404 -10930 1418
rect -10868 1524 -10834 1539
rect -10868 1505 -10834 1524
rect -10772 1418 -10738 1438
rect -10772 1404 -10738 1418
rect -10676 1524 -10642 1539
rect -10676 1505 -10642 1524
rect -10580 1418 -10546 1438
rect -10580 1404 -10546 1418
rect -10484 1524 -10450 1539
rect -10484 1505 -10450 1524
rect -10388 1418 -10354 1524
rect -10200 1790 -10127 1893
rect -9883 1784 -9750 1837
rect -8250 2456 -8216 2558
rect -8250 2061 -8216 2163
rect -8154 2248 -8120 2372
rect -8058 2456 -8024 2558
rect -8058 2097 -8024 2163
rect -7962 2248 -7928 2372
rect -7866 2454 -7832 2556
rect -7866 2097 -7832 2157
rect -7770 2248 -7736 2372
rect -7674 2453 -7640 2555
rect -7674 2097 -7640 2140
rect -7578 2248 -7544 2372
rect -7482 2453 -7448 2555
rect -7482 2097 -7448 2157
rect -7386 2248 -7352 2372
rect -7290 2453 -7256 2555
rect -7290 2097 -7256 2164
rect -7194 2247 -7160 2371
rect -7098 2453 -7064 2555
rect -7098 2097 -7064 2164
rect -9277 1792 -9163 1845
rect -9043 1838 -8963 1844
rect -9043 1783 -9035 1838
rect -9035 1783 -8970 1838
rect -8970 1783 -8963 1838
rect -9043 1776 -8963 1783
rect -8861 1618 -8796 1673
rect -9981 1418 -9947 1524
rect -9885 1524 -9851 1539
rect -9885 1505 -9851 1524
rect -9789 1418 -9755 1438
rect -9789 1404 -9755 1418
rect -9693 1524 -9659 1539
rect -9693 1505 -9659 1524
rect -9597 1418 -9563 1438
rect -9597 1404 -9563 1418
rect -9501 1524 -9467 1538
rect -9501 1504 -9467 1524
rect -9405 1418 -9371 1438
rect -9405 1404 -9371 1418
rect -9309 1524 -9275 1539
rect -9309 1505 -9275 1524
rect -9213 1418 -9179 1438
rect -9213 1404 -9179 1418
rect -9117 1524 -9083 1539
rect -9117 1505 -9083 1524
rect -9021 1418 -8987 1438
rect -9021 1404 -8987 1418
rect -8925 1524 -8891 1539
rect -8925 1505 -8891 1524
rect -8829 1418 -8795 1524
rect -8467 1828 -8420 1938
rect -8152 1784 -8019 1837
rect -6691 2456 -6657 2558
rect -6691 2061 -6657 2163
rect -6595 2248 -6561 2372
rect -6499 2456 -6465 2558
rect -6499 2097 -6465 2163
rect -6403 2248 -6369 2372
rect -6307 2454 -6273 2556
rect -6307 2097 -6273 2157
rect -6211 2248 -6177 2372
rect -6115 2453 -6081 2555
rect -6115 2097 -6081 2140
rect -6019 2248 -5985 2372
rect -5923 2453 -5889 2555
rect -5923 2097 -5889 2157
rect -5827 2248 -5793 2372
rect -5731 2453 -5697 2555
rect -5731 2097 -5697 2164
rect -5635 2247 -5601 2371
rect -5539 2453 -5505 2555
rect -5539 2097 -5505 2164
rect -7546 1792 -7432 1845
rect -7312 1838 -7232 1844
rect -7312 1783 -7304 1838
rect -7304 1783 -7239 1838
rect -7239 1783 -7232 1838
rect -7312 1776 -7232 1783
rect -7130 1618 -7065 1673
rect -8250 1418 -8216 1524
rect -8154 1524 -8120 1539
rect -8154 1505 -8120 1524
rect -8058 1418 -8024 1438
rect -8058 1404 -8024 1418
rect -7962 1524 -7928 1539
rect -7962 1505 -7928 1524
rect -7866 1418 -7832 1438
rect -7866 1404 -7832 1418
rect -7770 1524 -7736 1538
rect -7770 1504 -7736 1524
rect -7674 1418 -7640 1438
rect -7674 1404 -7640 1418
rect -7578 1524 -7544 1539
rect -7578 1505 -7544 1524
rect -7482 1418 -7448 1438
rect -7482 1404 -7448 1418
rect -7386 1524 -7352 1539
rect -7386 1505 -7352 1524
rect -7290 1418 -7256 1438
rect -7290 1404 -7256 1418
rect -7194 1524 -7160 1539
rect -7194 1505 -7160 1524
rect -7098 1418 -7064 1524
rect -6910 1790 -6837 1893
rect -6593 1784 -6460 1837
rect -4959 2456 -4925 2558
rect -4959 2061 -4925 2163
rect -4863 2248 -4829 2372
rect -4767 2456 -4733 2558
rect -4767 2097 -4733 2163
rect -4671 2248 -4637 2372
rect -4575 2454 -4541 2556
rect -4575 2097 -4541 2157
rect -4479 2248 -4445 2372
rect -4383 2453 -4349 2555
rect -4383 2097 -4349 2140
rect -4287 2248 -4253 2372
rect -4191 2453 -4157 2555
rect -4191 2097 -4157 2157
rect -4095 2248 -4061 2372
rect -3999 2453 -3965 2555
rect -3999 2097 -3965 2164
rect -3903 2247 -3869 2371
rect -3807 2453 -3773 2555
rect -3807 2097 -3773 2164
rect -5987 1792 -5873 1845
rect -5753 1838 -5673 1844
rect -5753 1783 -5745 1838
rect -5745 1783 -5680 1838
rect -5680 1783 -5673 1838
rect -5753 1776 -5673 1783
rect -5571 1618 -5506 1673
rect -6691 1418 -6657 1524
rect -6595 1524 -6561 1539
rect -6595 1505 -6561 1524
rect -6499 1418 -6465 1438
rect -6499 1404 -6465 1418
rect -6403 1524 -6369 1539
rect -6403 1505 -6369 1524
rect -6307 1418 -6273 1438
rect -6307 1404 -6273 1418
rect -6211 1524 -6177 1538
rect -6211 1504 -6177 1524
rect -6115 1418 -6081 1438
rect -6115 1404 -6081 1418
rect -6019 1524 -5985 1539
rect -6019 1505 -5985 1524
rect -5923 1418 -5889 1438
rect -5923 1404 -5889 1418
rect -5827 1524 -5793 1539
rect -5827 1505 -5793 1524
rect -5731 1418 -5697 1438
rect -5731 1404 -5697 1418
rect -5635 1524 -5601 1539
rect -5635 1505 -5601 1524
rect -5539 1418 -5505 1524
rect -5176 1828 -5129 1938
rect -4861 1784 -4728 1837
rect -3400 2456 -3366 2558
rect -3400 2061 -3366 2163
rect -3304 2248 -3270 2372
rect -3208 2456 -3174 2558
rect -3208 2097 -3174 2163
rect -3112 2248 -3078 2372
rect -3016 2454 -2982 2556
rect -3016 2097 -2982 2157
rect -2920 2248 -2886 2372
rect -2824 2453 -2790 2555
rect -2824 2097 -2790 2140
rect -2728 2248 -2694 2372
rect -2632 2453 -2598 2555
rect -2632 2097 -2598 2157
rect -2536 2248 -2502 2372
rect -2440 2453 -2406 2555
rect -2440 2097 -2406 2164
rect -2344 2247 -2310 2371
rect -2248 2453 -2214 2555
rect -2248 2097 -2214 2164
rect -4255 1792 -4141 1845
rect -4021 1838 -3941 1844
rect -4021 1783 -4013 1838
rect -4013 1783 -3948 1838
rect -3948 1783 -3941 1838
rect -4021 1776 -3941 1783
rect -3839 1618 -3774 1673
rect -4959 1418 -4925 1524
rect -4863 1524 -4829 1539
rect -4863 1505 -4829 1524
rect -4767 1418 -4733 1438
rect -4767 1404 -4733 1418
rect -4671 1524 -4637 1539
rect -4671 1505 -4637 1524
rect -4575 1418 -4541 1438
rect -4575 1404 -4541 1418
rect -4479 1524 -4445 1538
rect -4479 1504 -4445 1524
rect -4383 1418 -4349 1438
rect -4383 1404 -4349 1418
rect -4287 1524 -4253 1539
rect -4287 1505 -4253 1524
rect -4191 1418 -4157 1438
rect -4191 1404 -4157 1418
rect -4095 1524 -4061 1539
rect -4095 1505 -4061 1524
rect -3999 1418 -3965 1438
rect -3999 1404 -3965 1418
rect -3903 1524 -3869 1539
rect -3903 1505 -3869 1524
rect -3807 1418 -3773 1524
rect -3619 1790 -3546 1893
rect -3302 1784 -3169 1837
rect -1668 2456 -1634 2558
rect -1668 2061 -1634 2163
rect -1572 2248 -1538 2372
rect -1476 2456 -1442 2558
rect -1476 2097 -1442 2163
rect -1380 2248 -1346 2372
rect -1284 2454 -1250 2556
rect -1284 2097 -1250 2157
rect -1188 2248 -1154 2372
rect -1092 2453 -1058 2555
rect -1092 2097 -1058 2140
rect -996 2248 -962 2372
rect -900 2453 -866 2555
rect -900 2097 -866 2157
rect -804 2248 -770 2372
rect -708 2453 -674 2555
rect -708 2097 -674 2164
rect -612 2247 -578 2371
rect -516 2453 -482 2555
rect -516 2097 -482 2164
rect -2696 1792 -2582 1845
rect -2462 1838 -2382 1844
rect -2462 1783 -2454 1838
rect -2454 1783 -2389 1838
rect -2389 1783 -2382 1838
rect -2462 1776 -2382 1783
rect -2280 1618 -2215 1673
rect -3400 1418 -3366 1524
rect -3304 1524 -3270 1539
rect -3304 1505 -3270 1524
rect -3208 1418 -3174 1438
rect -3208 1404 -3174 1418
rect -3112 1524 -3078 1539
rect -3112 1505 -3078 1524
rect -3016 1418 -2982 1438
rect -3016 1404 -2982 1418
rect -2920 1524 -2886 1538
rect -2920 1504 -2886 1524
rect -2824 1418 -2790 1438
rect -2824 1404 -2790 1418
rect -2728 1524 -2694 1539
rect -2728 1505 -2694 1524
rect -2632 1418 -2598 1438
rect -2632 1404 -2598 1418
rect -2536 1524 -2502 1539
rect -2536 1505 -2502 1524
rect -2440 1418 -2406 1438
rect -2440 1404 -2406 1418
rect -2344 1524 -2310 1539
rect -2344 1505 -2310 1524
rect -2248 1418 -2214 1524
rect -1885 1828 -1838 1938
rect -1570 1784 -1437 1837
rect -109 2456 -75 2558
rect -109 2061 -75 2163
rect -13 2248 21 2372
rect 83 2456 117 2558
rect 83 2097 117 2163
rect 179 2248 213 2372
rect 275 2454 309 2556
rect 275 2097 309 2157
rect 371 2248 405 2372
rect 467 2453 501 2555
rect 467 2097 501 2140
rect 563 2248 597 2372
rect 659 2453 693 2555
rect 659 2097 693 2157
rect 755 2248 789 2372
rect 851 2453 885 2555
rect 851 2097 885 2164
rect 947 2247 981 2371
rect 1043 2453 1077 2555
rect 1043 2097 1077 2164
rect -964 1792 -850 1845
rect -730 1838 -650 1844
rect -730 1783 -722 1838
rect -722 1783 -657 1838
rect -657 1783 -650 1838
rect -730 1776 -650 1783
rect -548 1618 -483 1673
rect -1668 1418 -1634 1524
rect -1572 1524 -1538 1539
rect -1572 1505 -1538 1524
rect -1476 1418 -1442 1438
rect -1476 1404 -1442 1418
rect -1380 1524 -1346 1539
rect -1380 1505 -1346 1524
rect -1284 1418 -1250 1438
rect -1284 1404 -1250 1418
rect -1188 1524 -1154 1538
rect -1188 1504 -1154 1524
rect -1092 1418 -1058 1438
rect -1092 1404 -1058 1418
rect -996 1524 -962 1539
rect -996 1505 -962 1524
rect -900 1418 -866 1438
rect -900 1404 -866 1418
rect -804 1524 -770 1539
rect -804 1505 -770 1524
rect -708 1418 -674 1438
rect -708 1404 -674 1418
rect -612 1524 -578 1539
rect -612 1505 -578 1524
rect -516 1418 -482 1524
rect -328 1790 -255 1893
rect -11 1784 122 1837
rect 595 1792 709 1845
rect 829 1838 909 1844
rect 829 1783 837 1838
rect 837 1783 902 1838
rect 902 1783 909 1838
rect 829 1776 909 1783
rect 1011 1618 1076 1673
rect -109 1418 -75 1524
rect -13 1524 21 1539
rect -13 1505 21 1524
rect 83 1418 117 1438
rect 83 1404 117 1418
rect 179 1524 213 1539
rect 179 1505 213 1524
rect 275 1418 309 1438
rect 275 1404 309 1418
rect 371 1524 405 1538
rect 371 1504 405 1524
rect 467 1418 501 1438
rect 467 1404 501 1418
rect 563 1524 597 1539
rect 563 1505 597 1524
rect 659 1418 693 1438
rect 659 1404 693 1418
rect 755 1524 789 1539
rect 755 1505 789 1524
rect 851 1418 885 1438
rect 851 1404 885 1418
rect 947 1524 981 1539
rect 947 1505 981 1524
rect 1043 1418 1077 1524
rect 7298 2118 7332 2466
rect 7332 2118 7333 2466
rect 7298 2066 7333 2118
rect 7298 1715 7332 2066
rect 7332 1715 7333 2066
rect 7372 1702 7406 2478
rect 7756 1702 7790 2478
rect 8246 2118 8280 2466
rect 8280 2118 8281 2466
rect 8246 2066 8281 2118
rect 8246 1715 8280 2066
rect 8280 1715 8281 2066
rect 8320 1702 8354 2478
rect 8704 1702 8738 2478
rect 9182 2118 9216 2466
rect 9216 2118 9217 2466
rect 9182 2066 9217 2118
rect 9182 1715 9216 2066
rect 9216 1715 9217 2066
rect 9256 1702 9290 2478
rect 9640 1702 9674 2478
rect 10113 2118 10147 2466
rect 10147 2118 10148 2466
rect 10113 2066 10148 2118
rect 10113 1715 10147 2066
rect 10147 1715 10148 2066
rect 10187 1702 10221 2478
rect 10571 1702 10605 2478
rect 11040 2118 11074 2466
rect 11074 2118 11075 2466
rect 11040 2066 11075 2118
rect 11040 1715 11074 2066
rect 11074 1715 11075 2066
rect 11114 1702 11148 2478
rect 11498 1702 11532 2478
rect 11811 2101 12168 2152
rect 11785 1765 11819 1855
rect 11881 1907 11915 1997
rect 11977 1765 12011 1855
rect 12073 1907 12107 1997
rect 12169 1765 12203 1855
rect 12265 1907 12299 1997
rect 12361 1765 12395 1855
rect 12457 1907 12491 1997
rect 12553 1765 12587 1855
rect 12649 1907 12683 1997
rect 12986 1931 13077 1965
rect 12745 1765 12779 1855
rect 12929 1859 12935 1893
rect 12935 1859 13008 1893
rect 12170 1669 12204 1703
rect 12842 1619 12876 1845
rect 13052 1763 13129 1797
rect 12929 1667 12935 1701
rect 12935 1667 13008 1701
rect -24670 1284 -23547 1330
rect -23111 1284 -21988 1330
rect -21379 1284 -20256 1330
rect -19820 1284 -18697 1330
rect -18088 1284 -16965 1330
rect -16529 1284 -15406 1330
rect -14797 1284 -13674 1330
rect -13238 1284 -12115 1330
rect -11506 1284 -10383 1330
rect -9947 1284 -8824 1330
rect -8216 1284 -7093 1330
rect -6657 1284 -5534 1330
rect -4925 1284 -3802 1330
rect -3366 1284 -2243 1330
rect -1634 1284 -511 1330
rect -75 1284 1048 1330
rect 7298 1186 7332 1537
rect 7332 1186 7333 1537
rect 7298 1134 7333 1186
rect -24569 941 -24000 988
rect -23460 941 -22891 988
rect -22578 941 -22009 988
rect -21278 941 -20709 988
rect -20169 941 -19600 988
rect -19287 941 -18718 988
rect -17987 941 -17418 988
rect -16878 941 -16309 988
rect -15996 941 -15427 988
rect -14696 941 -14127 988
rect -13587 941 -13018 988
rect -12705 941 -12136 988
rect -11405 941 -10836 988
rect -10296 941 -9727 988
rect -9414 941 -8845 988
rect -8115 941 -7546 988
rect -7006 941 -6437 988
rect -6124 941 -5555 988
rect -4824 941 -4255 988
rect -3715 941 -3146 988
rect -2833 941 -2264 988
rect -1533 941 -964 988
rect -424 941 145 988
rect 458 941 1027 988
rect -24585 863 -24551 869
rect -24585 789 -24551 863
rect -24489 673 -24455 747
rect -24489 667 -24455 673
rect -24393 863 -24359 869
rect -24393 789 -24359 863
rect -24297 673 -24263 747
rect -24297 667 -24263 673
rect -24201 863 -24167 869
rect -24201 789 -24167 863
rect -24105 673 -24071 747
rect -24105 667 -24071 673
rect -24009 863 -23975 869
rect -24009 789 -23975 863
rect -23476 863 -23442 869
rect -23476 789 -23442 863
rect -23380 673 -23346 747
rect -23380 667 -23346 673
rect -23284 863 -23250 869
rect -23284 789 -23250 863
rect -23188 673 -23154 747
rect -23188 667 -23154 673
rect -23092 863 -23058 869
rect -23092 789 -23058 863
rect -22996 673 -22962 747
rect -22996 667 -22962 673
rect -22900 863 -22866 869
rect -22900 789 -22866 863
rect -22594 863 -22560 869
rect -22594 789 -22560 863
rect -22498 673 -22464 747
rect -22498 667 -22464 673
rect -22402 863 -22368 869
rect -22402 789 -22368 863
rect -22306 673 -22272 747
rect -22306 667 -22272 673
rect -22210 863 -22176 869
rect -22210 789 -22176 863
rect -22114 673 -22080 747
rect -22114 667 -22080 673
rect -22018 863 -21984 869
rect -22018 789 -21984 863
rect -21294 863 -21260 869
rect -21294 789 -21260 863
rect -21198 673 -21164 747
rect -21198 667 -21164 673
rect -21102 863 -21068 869
rect -21102 789 -21068 863
rect -21006 673 -20972 747
rect -21006 667 -20972 673
rect -20910 863 -20876 869
rect -20910 789 -20876 863
rect -20814 673 -20780 747
rect -20814 667 -20780 673
rect -20718 863 -20684 869
rect -20718 789 -20684 863
rect -20185 863 -20151 869
rect -20185 789 -20151 863
rect -20089 673 -20055 747
rect -20089 667 -20055 673
rect -19993 863 -19959 869
rect -19993 789 -19959 863
rect -19897 673 -19863 747
rect -19897 667 -19863 673
rect -19801 863 -19767 869
rect -19801 789 -19767 863
rect -19705 673 -19671 747
rect -19705 667 -19671 673
rect -19609 863 -19575 869
rect -19609 789 -19575 863
rect -19303 863 -19269 869
rect -19303 789 -19269 863
rect -19207 673 -19173 747
rect -19207 667 -19173 673
rect -19111 863 -19077 869
rect -19111 789 -19077 863
rect -19015 673 -18981 747
rect -19015 667 -18981 673
rect -18919 863 -18885 869
rect -18919 789 -18885 863
rect -18823 673 -18789 747
rect -18823 667 -18789 673
rect -18727 863 -18693 869
rect -18727 789 -18693 863
rect -18003 863 -17969 869
rect -18003 789 -17969 863
rect -17907 673 -17873 747
rect -17907 667 -17873 673
rect -17811 863 -17777 869
rect -17811 789 -17777 863
rect -17715 673 -17681 747
rect -17715 667 -17681 673
rect -17619 863 -17585 869
rect -17619 789 -17585 863
rect -17523 673 -17489 747
rect -17523 667 -17489 673
rect -17427 863 -17393 869
rect -17427 789 -17393 863
rect -16894 863 -16860 869
rect -16894 789 -16860 863
rect -16798 673 -16764 747
rect -16798 667 -16764 673
rect -16702 863 -16668 869
rect -16702 789 -16668 863
rect -16606 673 -16572 747
rect -16606 667 -16572 673
rect -16510 863 -16476 869
rect -16510 789 -16476 863
rect -16414 673 -16380 747
rect -16414 667 -16380 673
rect -16318 863 -16284 869
rect -16318 789 -16284 863
rect -16012 863 -15978 869
rect -16012 789 -15978 863
rect -15916 673 -15882 747
rect -15916 667 -15882 673
rect -15820 863 -15786 869
rect -15820 789 -15786 863
rect -15724 673 -15690 747
rect -15724 667 -15690 673
rect -15628 863 -15594 869
rect -15628 789 -15594 863
rect -15532 673 -15498 747
rect -15532 667 -15498 673
rect -15436 863 -15402 869
rect -15436 789 -15402 863
rect -14712 863 -14678 869
rect -14712 789 -14678 863
rect -14616 673 -14582 747
rect -14616 667 -14582 673
rect -14520 863 -14486 869
rect -14520 789 -14486 863
rect -14424 673 -14390 747
rect -14424 667 -14390 673
rect -14328 863 -14294 869
rect -14328 789 -14294 863
rect -14232 673 -14198 747
rect -14232 667 -14198 673
rect -14136 863 -14102 869
rect -14136 789 -14102 863
rect -13603 863 -13569 869
rect -13603 789 -13569 863
rect -13507 673 -13473 747
rect -13507 667 -13473 673
rect -13411 863 -13377 869
rect -13411 789 -13377 863
rect -13315 673 -13281 747
rect -13315 667 -13281 673
rect -13219 863 -13185 869
rect -13219 789 -13185 863
rect -13123 673 -13089 747
rect -13123 667 -13089 673
rect -13027 863 -12993 869
rect -13027 789 -12993 863
rect -12721 863 -12687 869
rect -12721 789 -12687 863
rect -12625 673 -12591 747
rect -12625 667 -12591 673
rect -12529 863 -12495 869
rect -12529 789 -12495 863
rect -12433 673 -12399 747
rect -12433 667 -12399 673
rect -12337 863 -12303 869
rect -12337 789 -12303 863
rect -12241 673 -12207 747
rect -12241 667 -12207 673
rect -12145 863 -12111 869
rect -12145 789 -12111 863
rect -11421 863 -11387 869
rect -11421 789 -11387 863
rect -11325 673 -11291 747
rect -11325 667 -11291 673
rect -11229 863 -11195 869
rect -11229 789 -11195 863
rect -11133 673 -11099 747
rect -11133 667 -11099 673
rect -11037 863 -11003 869
rect -11037 789 -11003 863
rect -10941 673 -10907 747
rect -10941 667 -10907 673
rect -10845 863 -10811 869
rect -10845 789 -10811 863
rect -10312 863 -10278 869
rect -10312 789 -10278 863
rect -10216 673 -10182 747
rect -10216 667 -10182 673
rect -10120 863 -10086 869
rect -10120 789 -10086 863
rect -10024 673 -9990 747
rect -10024 667 -9990 673
rect -9928 863 -9894 869
rect -9928 789 -9894 863
rect -9832 673 -9798 747
rect -9832 667 -9798 673
rect -9736 863 -9702 869
rect -9736 789 -9702 863
rect -9430 863 -9396 869
rect -9430 789 -9396 863
rect -9334 673 -9300 747
rect -9334 667 -9300 673
rect -9238 863 -9204 869
rect -9238 789 -9204 863
rect -9142 673 -9108 747
rect -9142 667 -9108 673
rect -9046 863 -9012 869
rect -9046 789 -9012 863
rect -8950 673 -8916 747
rect -8950 667 -8916 673
rect -8854 863 -8820 869
rect -8854 789 -8820 863
rect -8131 863 -8097 869
rect -8131 789 -8097 863
rect -8035 673 -8001 747
rect -8035 667 -8001 673
rect -7939 863 -7905 869
rect -7939 789 -7905 863
rect -7843 673 -7809 747
rect -7843 667 -7809 673
rect -7747 863 -7713 869
rect -7747 789 -7713 863
rect -7651 673 -7617 747
rect -7651 667 -7617 673
rect -7555 863 -7521 869
rect -7555 789 -7521 863
rect -7022 863 -6988 869
rect -7022 789 -6988 863
rect -6926 673 -6892 747
rect -6926 667 -6892 673
rect -6830 863 -6796 869
rect -6830 789 -6796 863
rect -6734 673 -6700 747
rect -6734 667 -6700 673
rect -6638 863 -6604 869
rect -6638 789 -6604 863
rect -6542 673 -6508 747
rect -6542 667 -6508 673
rect -6446 863 -6412 869
rect -6446 789 -6412 863
rect -6140 863 -6106 869
rect -6140 789 -6106 863
rect -6044 673 -6010 747
rect -6044 667 -6010 673
rect -5948 863 -5914 869
rect -5948 789 -5914 863
rect -5852 673 -5818 747
rect -5852 667 -5818 673
rect -5756 863 -5722 869
rect -5756 789 -5722 863
rect -5660 673 -5626 747
rect -5660 667 -5626 673
rect -5564 863 -5530 869
rect -5564 789 -5530 863
rect -4840 863 -4806 869
rect -4840 789 -4806 863
rect -4744 673 -4710 747
rect -4744 667 -4710 673
rect -4648 863 -4614 869
rect -4648 789 -4614 863
rect -4552 673 -4518 747
rect -4552 667 -4518 673
rect -4456 863 -4422 869
rect -4456 789 -4422 863
rect -4360 673 -4326 747
rect -4360 667 -4326 673
rect -4264 863 -4230 869
rect -4264 789 -4230 863
rect -3731 863 -3697 869
rect -3731 789 -3697 863
rect -3635 673 -3601 747
rect -3635 667 -3601 673
rect -3539 863 -3505 869
rect -3539 789 -3505 863
rect -3443 673 -3409 747
rect -3443 667 -3409 673
rect -3347 863 -3313 869
rect -3347 789 -3313 863
rect -3251 673 -3217 747
rect -3251 667 -3217 673
rect -3155 863 -3121 869
rect -3155 789 -3121 863
rect -2849 863 -2815 869
rect -2849 789 -2815 863
rect -2753 673 -2719 747
rect -2753 667 -2719 673
rect -2657 863 -2623 869
rect -2657 789 -2623 863
rect -2561 673 -2527 747
rect -2561 667 -2527 673
rect -2465 863 -2431 869
rect -2465 789 -2431 863
rect -2369 673 -2335 747
rect -2369 667 -2335 673
rect -2273 863 -2239 869
rect -2273 789 -2239 863
rect -1549 863 -1515 869
rect -1549 789 -1515 863
rect -1453 673 -1419 747
rect -1453 667 -1419 673
rect -1357 863 -1323 869
rect -1357 789 -1323 863
rect -1261 673 -1227 747
rect -1261 667 -1227 673
rect -1165 863 -1131 869
rect -1165 789 -1131 863
rect -1069 673 -1035 747
rect -1069 667 -1035 673
rect -973 863 -939 869
rect -973 789 -939 863
rect -440 863 -406 869
rect -440 789 -406 863
rect -344 673 -310 747
rect -344 667 -310 673
rect -248 863 -214 869
rect -248 789 -214 863
rect -152 673 -118 747
rect -152 667 -118 673
rect -56 863 -22 869
rect -56 789 -22 863
rect 40 673 74 747
rect 40 667 74 673
rect 136 863 170 869
rect 136 789 170 863
rect 442 863 476 869
rect 442 789 476 863
rect 538 673 572 747
rect 538 667 572 673
rect 634 863 668 869
rect 634 789 668 863
rect 730 673 764 747
rect 730 667 764 673
rect 826 863 860 869
rect 826 789 860 863
rect 922 673 956 747
rect 922 667 956 673
rect 1018 863 1052 869
rect 1018 789 1052 863
rect 7298 786 7332 1134
rect 7332 786 7333 1134
rect 7372 774 7406 1550
rect 7756 774 7790 1550
rect 8246 1186 8280 1537
rect 8280 1186 8281 1537
rect 8246 1134 8281 1186
rect 8246 786 8280 1134
rect 8280 786 8281 1134
rect 8320 774 8354 1550
rect 8704 774 8738 1550
rect 9182 1186 9216 1537
rect 9216 1186 9217 1537
rect 9182 1134 9217 1186
rect 9182 786 9216 1134
rect 9216 786 9217 1134
rect 9256 774 9290 1550
rect 9640 774 9674 1550
rect 10113 1187 10147 1538
rect 10147 1187 10148 1538
rect 10113 1135 10148 1187
rect 10113 787 10147 1135
rect 10147 787 10148 1135
rect 10187 775 10221 1551
rect 10571 775 10605 1551
rect 11040 1186 11074 1537
rect 11074 1186 11075 1537
rect 11040 1134 11075 1186
rect 11040 786 11074 1134
rect 11074 786 11075 1134
rect 11114 774 11148 1550
rect 12313 1564 12347 1598
rect 11498 774 11532 1550
rect 12265 1332 12299 1508
rect 13052 1571 13129 1605
rect 12935 1409 13111 1443
rect 12842 1365 12876 1399
rect 12935 1321 13111 1355
rect 12183 1188 12382 1249
rect 12954 1219 13086 1253
rect -24519 579 -24485 614
rect -24230 579 -24196 614
rect -23410 579 -23376 614
rect -23121 579 -23087 614
rect -24435 455 -24401 490
rect -24351 485 -23975 519
rect -22528 579 -22494 614
rect -22239 579 -22205 614
rect -23326 455 -23292 490
rect -23242 485 -22866 519
rect -21228 579 -21194 614
rect -20939 579 -20905 614
rect -22444 455 -22410 490
rect -22360 485 -21984 519
rect -20119 579 -20085 614
rect -19830 579 -19796 614
rect -21144 455 -21110 490
rect -21060 485 -20684 519
rect -19237 579 -19203 614
rect -18948 579 -18914 614
rect -20035 455 -20001 490
rect -19951 485 -19575 519
rect -17937 579 -17903 614
rect -17648 579 -17614 614
rect -19153 455 -19119 490
rect -19069 485 -18693 519
rect -16828 579 -16794 614
rect -16539 579 -16505 614
rect -17853 455 -17819 490
rect -17769 485 -17393 519
rect -15946 579 -15912 614
rect -15657 579 -15623 614
rect -16744 455 -16710 490
rect -16660 485 -16284 519
rect -14646 579 -14612 614
rect -14357 579 -14323 614
rect -15862 455 -15828 490
rect -15778 485 -15402 519
rect -13537 579 -13503 614
rect -13248 579 -13214 614
rect -14562 455 -14528 490
rect -14478 485 -14102 519
rect -12655 579 -12621 614
rect -12366 579 -12332 614
rect -13453 455 -13419 490
rect -13369 485 -12993 519
rect -11355 579 -11321 614
rect -11066 579 -11032 614
rect -12571 455 -12537 490
rect -12487 485 -12111 519
rect -10246 579 -10212 614
rect -9957 579 -9923 614
rect -11271 455 -11237 490
rect -11187 485 -10811 519
rect -9364 579 -9330 614
rect -9075 579 -9041 614
rect -10162 455 -10128 490
rect -10078 485 -9702 519
rect -8065 579 -8031 614
rect -7776 579 -7742 614
rect -9280 455 -9246 490
rect -9196 485 -8820 519
rect -6956 579 -6922 614
rect -6667 579 -6633 614
rect -7981 455 -7947 490
rect -7897 485 -7521 519
rect -6074 579 -6040 614
rect -5785 579 -5751 614
rect -6872 455 -6838 490
rect -6788 485 -6412 519
rect -4774 579 -4740 614
rect -4485 579 -4451 614
rect -5990 455 -5956 490
rect -5906 485 -5530 519
rect -3665 579 -3631 614
rect -3376 579 -3342 614
rect -4690 455 -4656 490
rect -4606 485 -4230 519
rect -2783 579 -2749 614
rect -2494 579 -2460 614
rect -3581 455 -3547 490
rect -3497 485 -3121 519
rect -1483 579 -1449 614
rect -1194 579 -1160 614
rect -2699 455 -2665 490
rect -2615 485 -2239 519
rect -374 579 -340 614
rect -85 579 -51 614
rect -1399 455 -1365 490
rect -1315 485 -939 519
rect 508 579 542 614
rect 797 579 831 614
rect -290 455 -256 490
rect -206 485 170 519
rect 592 455 626 490
rect 676 485 1052 519
rect 7198 402 7232 436
rect 7390 402 7424 436
rect 7582 402 7616 436
rect 7774 402 7808 436
rect 8146 402 8180 436
rect 8338 402 8372 436
rect 8530 402 8564 436
rect 8722 402 8756 436
rect 9082 402 9116 436
rect 9274 402 9308 436
rect 9466 402 9500 436
rect 9658 402 9692 436
rect 10013 403 10047 437
rect 10205 403 10239 437
rect 10397 403 10431 437
rect 10589 403 10623 437
rect 10940 402 10974 436
rect 11132 402 11166 436
rect 11324 402 11358 436
rect 11516 402 11550 436
rect -24351 293 -23975 327
rect -23242 293 -22866 327
rect -22360 293 -21984 327
rect -21060 293 -20684 327
rect -19951 293 -19575 327
rect -19069 293 -18693 327
rect -17769 293 -17393 327
rect -16660 293 -16284 327
rect -15778 293 -15402 327
rect -14478 293 -14102 327
rect -13369 293 -12993 327
rect -12487 293 -12111 327
rect -11187 293 -10811 327
rect -10078 293 -9702 327
rect -9196 293 -8820 327
rect -7897 293 -7521 327
rect -6788 293 -6412 327
rect -5906 293 -5530 327
rect -4606 293 -4230 327
rect -3497 293 -3121 327
rect -2615 293 -2239 327
rect -1315 293 -939 327
rect -206 293 170 327
rect 676 293 1052 327
rect -24336 221 -24001 255
rect -23227 221 -22892 255
rect -22345 221 -22010 255
rect -21045 221 -20710 255
rect -19936 221 -19601 255
rect -19054 221 -18719 255
rect -17754 221 -17419 255
rect -16645 221 -16310 255
rect -15763 221 -15428 255
rect -14463 221 -14128 255
rect -13354 221 -13019 255
rect -12472 221 -12137 255
rect -11172 221 -10837 255
rect -10063 221 -9728 255
rect -9181 221 -8846 255
rect -7882 221 -7547 255
rect -6773 221 -6438 255
rect -5891 221 -5556 255
rect -4591 221 -4256 255
rect -3482 221 -3147 255
rect -2600 221 -2265 255
rect -1300 221 -965 255
rect -191 221 144 255
rect 691 221 1026 255
rect 7245 343 7280 348
rect 7245 236 7246 343
rect 7246 236 7280 343
rect 7150 48 7184 158
rect 7342 48 7376 158
rect 7438 343 7473 348
rect 7438 236 7472 343
rect 7472 236 7473 343
rect 7534 48 7568 158
rect 7630 343 7665 348
rect 7630 236 7664 343
rect 7664 236 7665 343
rect 7726 48 7760 158
rect 7822 343 7857 348
rect 7822 236 7856 343
rect 7856 236 7857 343
rect 7918 48 7952 158
rect 8193 343 8228 348
rect 8193 236 8194 343
rect 8194 236 8228 343
rect 8098 48 8132 158
rect 8290 48 8324 158
rect 8386 343 8421 348
rect 8386 236 8420 343
rect 8420 236 8421 343
rect 8482 48 8516 158
rect 8578 343 8613 348
rect 8578 236 8612 343
rect 8612 236 8613 343
rect 8674 48 8708 158
rect 8770 343 8805 348
rect 8770 236 8804 343
rect 8804 236 8805 343
rect 8866 48 8900 158
rect 9129 343 9164 348
rect 9129 236 9130 343
rect 9130 236 9164 343
rect 9034 48 9068 158
rect 9226 48 9260 158
rect 9322 343 9357 348
rect 9322 236 9356 343
rect 9356 236 9357 343
rect 9418 48 9452 158
rect 9514 343 9549 348
rect 9514 236 9548 343
rect 9548 236 9549 343
rect 9610 48 9644 158
rect 9706 343 9741 348
rect 9706 236 9740 343
rect 9740 236 9741 343
rect 9802 48 9836 158
rect 10060 344 10095 349
rect 10060 237 10061 344
rect 10061 237 10095 344
rect 9965 49 9999 159
rect 10157 49 10191 159
rect 10253 344 10288 349
rect 10253 237 10287 344
rect 10287 237 10288 344
rect 10349 49 10383 159
rect 10445 344 10480 349
rect 10445 237 10479 344
rect 10479 237 10480 344
rect 10541 49 10575 159
rect 10637 344 10672 349
rect 10637 237 10671 344
rect 10671 237 10672 344
rect 10733 49 10767 159
rect 10987 343 11022 348
rect 10987 236 10988 343
rect 10988 236 11022 343
rect 10892 48 10926 158
rect 11084 48 11118 158
rect 11180 343 11215 348
rect 11180 236 11214 343
rect 11214 236 11215 343
rect 11276 48 11310 158
rect 11372 343 11407 348
rect 11372 236 11406 343
rect 11406 236 11407 343
rect 11468 48 11502 158
rect 11564 343 11599 348
rect 11564 236 11598 343
rect 11598 236 11599 343
rect 11660 48 11694 158
rect 7389 -59 7677 -24
rect 8337 -59 8625 -24
rect 9273 -59 9561 -24
rect 10204 -58 10492 -23
rect 11131 -59 11419 -24
rect 5721 -579 5812 -545
rect 6161 -579 6252 -545
rect 6601 -579 6692 -545
rect 5664 -651 5670 -617
rect 5670 -651 5743 -617
rect 5577 -891 5611 -665
rect 6104 -651 6110 -617
rect 6110 -651 6183 -617
rect 5787 -747 5864 -713
rect 5664 -843 5670 -809
rect 5670 -843 5743 -809
rect 6017 -891 6051 -665
rect 6544 -651 6550 -617
rect 6550 -651 6623 -617
rect 6227 -747 6304 -713
rect 6104 -843 6110 -809
rect 6110 -843 6183 -809
rect 5787 -939 5864 -905
rect 5670 -1101 5846 -1067
rect 5577 -1145 5611 -1111
rect 6457 -891 6491 -665
rect 6667 -747 6744 -713
rect 6544 -843 6550 -809
rect 6550 -843 6623 -809
rect 6227 -939 6304 -905
rect 6110 -1101 6286 -1067
rect 6017 -1145 6051 -1111
rect 5670 -1189 5846 -1155
rect 6667 -939 6744 -905
rect 6550 -1101 6726 -1067
rect 6457 -1145 6491 -1111
rect 6110 -1189 6286 -1155
rect 6550 -1189 6726 -1155
rect 7389 -1252 7677 -1217
rect 8337 -1252 8625 -1217
rect 9273 -1252 9561 -1217
rect 10204 -1252 10492 -1217
rect 11131 -1252 11419 -1217
rect 5689 -1291 5821 -1257
rect 6129 -1291 6261 -1257
rect 6569 -1291 6701 -1257
rect 7150 -1434 7184 -1324
rect 7245 -1619 7246 -1512
rect 7246 -1619 7280 -1512
rect 7245 -1624 7280 -1619
rect 7342 -1434 7376 -1324
rect 7534 -1434 7568 -1324
rect 7438 -1619 7472 -1512
rect 7472 -1619 7473 -1512
rect 7438 -1624 7473 -1619
rect 7726 -1434 7760 -1324
rect 7630 -1619 7664 -1512
rect 7664 -1619 7665 -1512
rect 7630 -1624 7665 -1619
rect 7918 -1434 7952 -1324
rect 7822 -1619 7856 -1512
rect 7856 -1619 7857 -1512
rect 7822 -1624 7857 -1619
rect 8098 -1434 8132 -1324
rect 8193 -1619 8194 -1512
rect 8194 -1619 8228 -1512
rect 8193 -1624 8228 -1619
rect 8290 -1434 8324 -1324
rect 8482 -1434 8516 -1324
rect 8386 -1619 8420 -1512
rect 8420 -1619 8421 -1512
rect 8386 -1624 8421 -1619
rect 8674 -1434 8708 -1324
rect 8578 -1619 8612 -1512
rect 8612 -1619 8613 -1512
rect 8578 -1624 8613 -1619
rect 8866 -1434 8900 -1324
rect 8770 -1619 8804 -1512
rect 8804 -1619 8805 -1512
rect 8770 -1624 8805 -1619
rect 9034 -1434 9068 -1324
rect 9129 -1619 9130 -1512
rect 9130 -1619 9164 -1512
rect 9129 -1624 9164 -1619
rect 9226 -1434 9260 -1324
rect 9418 -1434 9452 -1324
rect 9322 -1619 9356 -1512
rect 9356 -1619 9357 -1512
rect 9322 -1624 9357 -1619
rect 9610 -1434 9644 -1324
rect 9514 -1619 9548 -1512
rect 9548 -1619 9549 -1512
rect 9514 -1624 9549 -1619
rect 9802 -1434 9836 -1324
rect 9706 -1619 9740 -1512
rect 9740 -1619 9741 -1512
rect 9706 -1624 9741 -1619
rect 9965 -1434 9999 -1324
rect 10060 -1619 10061 -1512
rect 10061 -1619 10095 -1512
rect 10060 -1624 10095 -1619
rect 10157 -1434 10191 -1324
rect 10349 -1434 10383 -1324
rect 10253 -1619 10287 -1512
rect 10287 -1619 10288 -1512
rect 10253 -1624 10288 -1619
rect 10541 -1434 10575 -1324
rect 10445 -1619 10479 -1512
rect 10479 -1619 10480 -1512
rect 10445 -1624 10480 -1619
rect 10733 -1434 10767 -1324
rect 10637 -1619 10671 -1512
rect 10671 -1619 10672 -1512
rect 10637 -1624 10672 -1619
rect 10892 -1434 10926 -1324
rect 10987 -1619 10988 -1512
rect 10988 -1619 11022 -1512
rect 10987 -1624 11022 -1619
rect 11084 -1434 11118 -1324
rect 11276 -1434 11310 -1324
rect 11180 -1619 11214 -1512
rect 11214 -1619 11215 -1512
rect 11180 -1624 11215 -1619
rect 11468 -1434 11502 -1324
rect 11372 -1619 11406 -1512
rect 11406 -1619 11407 -1512
rect 11372 -1624 11407 -1619
rect 11660 -1434 11694 -1324
rect 11564 -1619 11598 -1512
rect 11598 -1619 11599 -1512
rect 11564 -1624 11599 -1619
rect 7198 -1712 7232 -1678
rect 7390 -1712 7424 -1678
rect 7582 -1712 7616 -1678
rect 7774 -1712 7808 -1678
rect 8146 -1712 8180 -1678
rect 8338 -1712 8372 -1678
rect 8530 -1712 8564 -1678
rect 8722 -1712 8756 -1678
rect 9082 -1712 9116 -1678
rect 9274 -1712 9308 -1678
rect 9466 -1712 9500 -1678
rect 9658 -1712 9692 -1678
rect 10013 -1712 10047 -1678
rect 10205 -1712 10239 -1678
rect 10397 -1712 10431 -1678
rect 10589 -1712 10623 -1678
rect 10940 -1712 10974 -1678
rect 11132 -1712 11166 -1678
rect 11324 -1712 11358 -1678
rect 11516 -1712 11550 -1678
rect -23565 -2281 -23474 -2247
rect -21545 -2281 -21454 -2247
rect -19804 -2281 -19713 -2247
rect -18025 -2281 -17934 -2247
rect -24419 -2347 -23850 -2300
rect -23622 -2353 -23616 -2319
rect -23616 -2353 -23543 -2319
rect -22382 -2347 -21813 -2300
rect -24435 -2425 -24401 -2419
rect -24435 -2499 -24401 -2425
rect -24339 -2615 -24305 -2541
rect -24339 -2621 -24305 -2615
rect -24243 -2425 -24209 -2419
rect -24243 -2499 -24209 -2425
rect -24147 -2615 -24113 -2541
rect -24147 -2621 -24113 -2615
rect -24051 -2425 -24017 -2419
rect -24051 -2499 -24017 -2425
rect -23955 -2615 -23921 -2541
rect -23955 -2621 -23921 -2615
rect -23859 -2425 -23825 -2419
rect -23859 -2499 -23825 -2425
rect -23709 -2593 -23675 -2367
rect -21602 -2353 -21596 -2319
rect -21596 -2353 -21523 -2319
rect -20652 -2347 -20083 -2300
rect -23499 -2449 -23422 -2415
rect -22398 -2425 -22364 -2419
rect -22398 -2499 -22364 -2425
rect -23622 -2545 -23616 -2511
rect -23616 -2545 -23543 -2511
rect -24369 -2709 -24335 -2674
rect -24080 -2709 -24046 -2674
rect -24285 -2833 -24251 -2798
rect -24201 -2803 -23825 -2769
rect -23499 -2641 -23422 -2607
rect -22302 -2615 -22268 -2541
rect -22302 -2621 -22268 -2615
rect -22206 -2425 -22172 -2419
rect -22206 -2499 -22172 -2425
rect -22110 -2615 -22076 -2541
rect -22110 -2621 -22076 -2615
rect -22014 -2425 -21980 -2419
rect -22014 -2499 -21980 -2425
rect -21918 -2615 -21884 -2541
rect -21918 -2621 -21884 -2615
rect -21822 -2425 -21788 -2419
rect -21822 -2499 -21788 -2425
rect -21689 -2593 -21655 -2367
rect -19861 -2353 -19855 -2319
rect -19855 -2353 -19782 -2319
rect -18892 -2347 -18323 -2300
rect -21479 -2449 -21402 -2415
rect -20668 -2425 -20634 -2419
rect -20668 -2499 -20634 -2425
rect -21602 -2545 -21596 -2511
rect -21596 -2545 -21523 -2511
rect -22332 -2709 -22298 -2674
rect -22043 -2709 -22009 -2674
rect -23616 -2803 -23440 -2769
rect -23709 -2847 -23675 -2813
rect -23616 -2891 -23440 -2857
rect -22248 -2833 -22214 -2798
rect -22164 -2803 -21788 -2769
rect -21479 -2641 -21402 -2607
rect -20572 -2615 -20538 -2541
rect -20572 -2621 -20538 -2615
rect -20476 -2425 -20442 -2419
rect -20476 -2499 -20442 -2425
rect -20380 -2615 -20346 -2541
rect -20380 -2621 -20346 -2615
rect -20284 -2425 -20250 -2419
rect -20284 -2499 -20250 -2425
rect -20188 -2615 -20154 -2541
rect -20188 -2621 -20154 -2615
rect -20092 -2425 -20058 -2419
rect -20092 -2499 -20058 -2425
rect -19948 -2593 -19914 -2367
rect -18082 -2353 -18076 -2319
rect -18076 -2353 -18003 -2319
rect -19738 -2449 -19661 -2415
rect -18908 -2425 -18874 -2419
rect -18908 -2499 -18874 -2425
rect -19861 -2545 -19855 -2511
rect -19855 -2545 -19782 -2511
rect -20602 -2709 -20568 -2674
rect -20313 -2709 -20279 -2674
rect -21596 -2803 -21420 -2769
rect -21689 -2847 -21655 -2813
rect -21596 -2891 -21420 -2857
rect -20518 -2833 -20484 -2798
rect -20434 -2803 -20058 -2769
rect -19738 -2641 -19661 -2607
rect -18812 -2615 -18778 -2541
rect -18812 -2621 -18778 -2615
rect -18716 -2425 -18682 -2419
rect -18716 -2499 -18682 -2425
rect -18620 -2615 -18586 -2541
rect -18620 -2621 -18586 -2615
rect -18524 -2425 -18490 -2419
rect -18524 -2499 -18490 -2425
rect -18428 -2615 -18394 -2541
rect -18428 -2621 -18394 -2615
rect -18332 -2425 -18298 -2419
rect -18332 -2499 -18298 -2425
rect -18169 -2593 -18135 -2367
rect 7298 -2410 7332 -2062
rect 7332 -2410 7333 -2062
rect -17959 -2449 -17882 -2415
rect 7298 -2462 7333 -2410
rect -18082 -2545 -18076 -2511
rect -18076 -2545 -18003 -2511
rect -18842 -2709 -18808 -2674
rect -18553 -2709 -18519 -2674
rect -19855 -2803 -19679 -2769
rect -19948 -2847 -19914 -2813
rect -19855 -2891 -19679 -2857
rect -18758 -2833 -18724 -2798
rect -18674 -2803 -18298 -2769
rect -17959 -2641 -17882 -2607
rect -18076 -2803 -17900 -2769
rect -18169 -2847 -18135 -2813
rect 7298 -2813 7332 -2462
rect 7332 -2813 7333 -2462
rect 7372 -2826 7406 -2050
rect 7756 -2826 7790 -2050
rect 8246 -2410 8280 -2062
rect 8280 -2410 8281 -2062
rect 8246 -2462 8281 -2410
rect 8246 -2813 8280 -2462
rect 8280 -2813 8281 -2462
rect 8320 -2826 8354 -2050
rect 8704 -2826 8738 -2050
rect 9182 -2410 9216 -2062
rect 9216 -2410 9217 -2062
rect 9182 -2462 9217 -2410
rect 9182 -2813 9216 -2462
rect 9216 -2813 9217 -2462
rect 9256 -2826 9290 -2050
rect 9640 -2826 9674 -2050
rect 10113 -2410 10147 -2062
rect 10147 -2410 10148 -2062
rect 10113 -2462 10148 -2410
rect 10113 -2813 10147 -2462
rect 10147 -2813 10148 -2462
rect 10187 -2826 10221 -2050
rect 10571 -2826 10605 -2050
rect 11040 -2410 11074 -2062
rect 11074 -2410 11075 -2062
rect 11040 -2462 11075 -2410
rect 11040 -2813 11074 -2462
rect 11074 -2813 11075 -2462
rect 11114 -2826 11148 -2050
rect 11498 -2826 11532 -2050
rect 11811 -2427 12168 -2376
rect 11785 -2763 11819 -2673
rect 11881 -2621 11915 -2531
rect 11977 -2763 12011 -2673
rect 12073 -2621 12107 -2531
rect 12169 -2763 12203 -2673
rect 12265 -2621 12299 -2531
rect 12361 -2763 12395 -2673
rect 12457 -2621 12491 -2531
rect 12553 -2763 12587 -2673
rect 12649 -2621 12683 -2531
rect 12986 -2597 13077 -2563
rect 12745 -2763 12779 -2673
rect 12929 -2669 12935 -2635
rect 12935 -2669 13008 -2635
rect -18076 -2891 -17900 -2857
rect 12170 -2859 12204 -2825
rect 12842 -2909 12876 -2683
rect 13052 -2765 13129 -2731
rect 12929 -2861 12935 -2827
rect 12935 -2861 13008 -2827
rect -24201 -2995 -23825 -2961
rect -23597 -2993 -23465 -2959
rect -22164 -2995 -21788 -2961
rect -21577 -2993 -21445 -2959
rect -20434 -2995 -20058 -2961
rect -19836 -2993 -19704 -2959
rect -18674 -2995 -18298 -2961
rect -18057 -2993 -17925 -2959
rect -24186 -3067 -23851 -3033
rect -22149 -3067 -21814 -3033
rect -20419 -3067 -20084 -3033
rect -18659 -3067 -18324 -3033
rect 7298 -3342 7332 -2991
rect 7332 -3342 7333 -2991
rect 7298 -3394 7333 -3342
rect 7298 -3742 7332 -3394
rect 7332 -3742 7333 -3394
rect 7372 -3754 7406 -2978
rect 7756 -3754 7790 -2978
rect 8246 -3342 8280 -2991
rect 8280 -3342 8281 -2991
rect 8246 -3394 8281 -3342
rect 8246 -3742 8280 -3394
rect 8280 -3742 8281 -3394
rect 8320 -3754 8354 -2978
rect 8704 -3754 8738 -2978
rect 9182 -3342 9216 -2991
rect 9216 -3342 9217 -2991
rect 9182 -3394 9217 -3342
rect 9182 -3742 9216 -3394
rect 9216 -3742 9217 -3394
rect 9256 -3754 9290 -2978
rect 9640 -3754 9674 -2978
rect 10113 -3341 10147 -2990
rect 10147 -3341 10148 -2990
rect 10113 -3393 10148 -3341
rect 10113 -3741 10147 -3393
rect 10147 -3741 10148 -3393
rect 10187 -3753 10221 -2977
rect 10571 -3753 10605 -2977
rect 11040 -3342 11074 -2991
rect 11074 -3342 11075 -2991
rect 11040 -3394 11075 -3342
rect 11040 -3742 11074 -3394
rect 11074 -3742 11075 -3394
rect 11114 -3754 11148 -2978
rect 12313 -2964 12347 -2930
rect 11498 -3754 11532 -2978
rect 12265 -3196 12299 -3020
rect 13052 -2957 13129 -2923
rect 12935 -3119 13111 -3085
rect 12842 -3163 12876 -3129
rect 12935 -3207 13111 -3173
rect 12183 -3340 12382 -3279
rect 12954 -3309 13086 -3275
rect -20603 -3899 -19481 -3827
rect -19044 -3899 -17922 -3827
rect -17312 -3899 -16190 -3827
rect -15753 -3899 -14631 -3827
rect -14021 -3899 -12899 -3827
rect -12462 -3899 -11340 -3827
rect -10730 -3899 -9608 -3827
rect -9171 -3899 -8049 -3827
rect -23521 -4093 -23430 -4059
rect -21783 -4093 -21692 -4059
rect -24368 -4159 -23799 -4112
rect -23578 -4165 -23572 -4131
rect -23572 -4165 -23499 -4131
rect -22632 -4159 -22063 -4112
rect -24384 -4237 -24350 -4231
rect -24384 -4311 -24350 -4237
rect -24288 -4427 -24254 -4353
rect -24288 -4433 -24254 -4427
rect -24192 -4237 -24158 -4231
rect -24192 -4311 -24158 -4237
rect -24096 -4427 -24062 -4353
rect -24096 -4433 -24062 -4427
rect -24000 -4237 -23966 -4231
rect -24000 -4311 -23966 -4237
rect -23904 -4427 -23870 -4353
rect -23904 -4433 -23870 -4427
rect -23808 -4237 -23774 -4231
rect -23808 -4311 -23774 -4237
rect -23665 -4405 -23631 -4179
rect -21840 -4165 -21834 -4131
rect -21834 -4165 -21761 -4131
rect -23455 -4261 -23378 -4227
rect -22648 -4237 -22614 -4231
rect -22648 -4311 -22614 -4237
rect -23578 -4357 -23572 -4323
rect -23572 -4357 -23499 -4323
rect -24318 -4521 -24284 -4486
rect -24029 -4521 -23995 -4486
rect -24234 -4645 -24200 -4610
rect -24150 -4615 -23774 -4581
rect -23455 -4453 -23378 -4419
rect -22552 -4427 -22518 -4353
rect -22552 -4433 -22518 -4427
rect -22456 -4237 -22422 -4231
rect -22456 -4311 -22422 -4237
rect -22360 -4427 -22326 -4353
rect -22360 -4433 -22326 -4427
rect -22264 -4237 -22230 -4231
rect -22264 -4311 -22230 -4237
rect -22168 -4427 -22134 -4353
rect -22168 -4433 -22134 -4427
rect -22072 -4237 -22038 -4231
rect -22072 -4311 -22038 -4237
rect -21927 -4405 -21893 -4179
rect -21717 -4261 -21640 -4227
rect -21840 -4357 -21834 -4323
rect -21834 -4357 -21761 -4323
rect -22582 -4521 -22548 -4486
rect -22293 -4521 -22259 -4486
rect -23572 -4615 -23396 -4581
rect -23665 -4659 -23631 -4625
rect -23572 -4703 -23396 -4669
rect -22498 -4645 -22464 -4610
rect -22414 -4615 -22038 -4581
rect -21717 -4453 -21640 -4419
rect -21834 -4615 -21658 -4581
rect -20637 -4104 -20603 -4002
rect -20637 -4499 -20603 -4397
rect -20541 -4312 -20507 -4188
rect -20445 -4104 -20411 -4002
rect -20445 -4463 -20411 -4397
rect -20349 -4312 -20315 -4188
rect -20253 -4106 -20219 -4004
rect -20253 -4463 -20219 -4403
rect -20157 -4312 -20123 -4188
rect -20061 -4107 -20027 -4005
rect -20061 -4463 -20027 -4420
rect -19965 -4312 -19931 -4188
rect -19869 -4107 -19835 -4005
rect -19869 -4463 -19835 -4403
rect -19773 -4312 -19739 -4188
rect -19677 -4107 -19643 -4005
rect -19677 -4463 -19643 -4396
rect -19581 -4313 -19547 -4189
rect -19485 -4107 -19451 -4005
rect -19485 -4463 -19451 -4396
rect -21927 -4659 -21893 -4625
rect -21834 -4703 -21658 -4669
rect -24150 -4807 -23774 -4773
rect -23553 -4805 -23421 -4771
rect -20854 -4732 -20807 -4622
rect -22414 -4807 -22038 -4773
rect -21815 -4805 -21683 -4771
rect -24135 -4879 -23800 -4845
rect -22399 -4879 -22064 -4845
rect -20539 -4776 -20406 -4723
rect -19078 -4104 -19044 -4002
rect -19078 -4499 -19044 -4397
rect -18982 -4312 -18948 -4188
rect -18886 -4104 -18852 -4002
rect -18886 -4463 -18852 -4397
rect -18790 -4312 -18756 -4188
rect -18694 -4106 -18660 -4004
rect -18694 -4463 -18660 -4403
rect -18598 -4312 -18564 -4188
rect -18502 -4107 -18468 -4005
rect -18502 -4463 -18468 -4420
rect -18406 -4312 -18372 -4188
rect -18310 -4107 -18276 -4005
rect -18310 -4463 -18276 -4403
rect -18214 -4312 -18180 -4188
rect -18118 -4107 -18084 -4005
rect -18118 -4463 -18084 -4396
rect -18022 -4313 -17988 -4189
rect -17926 -4107 -17892 -4005
rect -17926 -4463 -17892 -4396
rect -19933 -4768 -19819 -4715
rect -19699 -4722 -19619 -4716
rect -19699 -4777 -19691 -4722
rect -19691 -4777 -19626 -4722
rect -19626 -4777 -19619 -4722
rect -19699 -4784 -19619 -4777
rect -19517 -4942 -19452 -4887
rect -20637 -5142 -20603 -5036
rect -20541 -5036 -20507 -5021
rect -20541 -5055 -20507 -5036
rect -20445 -5142 -20411 -5122
rect -20445 -5156 -20411 -5142
rect -20349 -5036 -20315 -5021
rect -20349 -5055 -20315 -5036
rect -20253 -5142 -20219 -5122
rect -20253 -5156 -20219 -5142
rect -20157 -5036 -20123 -5022
rect -20157 -5056 -20123 -5036
rect -20061 -5142 -20027 -5122
rect -20061 -5156 -20027 -5142
rect -19965 -5036 -19931 -5021
rect -19965 -5055 -19931 -5036
rect -19869 -5142 -19835 -5122
rect -19869 -5156 -19835 -5142
rect -19773 -5036 -19739 -5021
rect -19773 -5055 -19739 -5036
rect -19677 -5142 -19643 -5122
rect -19677 -5156 -19643 -5142
rect -19581 -5036 -19547 -5021
rect -19581 -5055 -19547 -5036
rect -19485 -5142 -19451 -5036
rect -19297 -4770 -19224 -4667
rect -18980 -4776 -18847 -4723
rect -17346 -4104 -17312 -4002
rect -17346 -4499 -17312 -4397
rect -17250 -4312 -17216 -4188
rect -17154 -4104 -17120 -4002
rect -17154 -4463 -17120 -4397
rect -17058 -4312 -17024 -4188
rect -16962 -4106 -16928 -4004
rect -16962 -4463 -16928 -4403
rect -16866 -4312 -16832 -4188
rect -16770 -4107 -16736 -4005
rect -16770 -4463 -16736 -4420
rect -16674 -4312 -16640 -4188
rect -16578 -4107 -16544 -4005
rect -16578 -4463 -16544 -4403
rect -16482 -4312 -16448 -4188
rect -16386 -4107 -16352 -4005
rect -16386 -4463 -16352 -4396
rect -16290 -4313 -16256 -4189
rect -16194 -4107 -16160 -4005
rect -16194 -4463 -16160 -4396
rect -18374 -4768 -18260 -4715
rect -18140 -4722 -18060 -4716
rect -18140 -4777 -18132 -4722
rect -18132 -4777 -18067 -4722
rect -18067 -4777 -18060 -4722
rect -18140 -4784 -18060 -4777
rect -17958 -4942 -17893 -4887
rect -19078 -5142 -19044 -5036
rect -18982 -5036 -18948 -5021
rect -18982 -5055 -18948 -5036
rect -18886 -5142 -18852 -5122
rect -18886 -5156 -18852 -5142
rect -18790 -5036 -18756 -5021
rect -18790 -5055 -18756 -5036
rect -18694 -5142 -18660 -5122
rect -18694 -5156 -18660 -5142
rect -18598 -5036 -18564 -5022
rect -18598 -5056 -18564 -5036
rect -18502 -5142 -18468 -5122
rect -18502 -5156 -18468 -5142
rect -18406 -5036 -18372 -5021
rect -18406 -5055 -18372 -5036
rect -18310 -5142 -18276 -5122
rect -18310 -5156 -18276 -5142
rect -18214 -5036 -18180 -5021
rect -18214 -5055 -18180 -5036
rect -18118 -5142 -18084 -5122
rect -18118 -5156 -18084 -5142
rect -18022 -5036 -17988 -5021
rect -18022 -5055 -17988 -5036
rect -17926 -5142 -17892 -5036
rect -17563 -4732 -17516 -4622
rect -17248 -4776 -17115 -4723
rect -15787 -4104 -15753 -4002
rect -15787 -4499 -15753 -4397
rect -15691 -4312 -15657 -4188
rect -15595 -4104 -15561 -4002
rect -15595 -4463 -15561 -4397
rect -15499 -4312 -15465 -4188
rect -15403 -4106 -15369 -4004
rect -15403 -4463 -15369 -4403
rect -15307 -4312 -15273 -4188
rect -15211 -4107 -15177 -4005
rect -15211 -4463 -15177 -4420
rect -15115 -4312 -15081 -4188
rect -15019 -4107 -14985 -4005
rect -15019 -4463 -14985 -4403
rect -14923 -4312 -14889 -4188
rect -14827 -4107 -14793 -4005
rect -14827 -4463 -14793 -4396
rect -14731 -4313 -14697 -4189
rect -14635 -4107 -14601 -4005
rect -14635 -4463 -14601 -4396
rect -16642 -4768 -16528 -4715
rect -16408 -4722 -16328 -4716
rect -16408 -4777 -16400 -4722
rect -16400 -4777 -16335 -4722
rect -16335 -4777 -16328 -4722
rect -16408 -4784 -16328 -4777
rect -16226 -4942 -16161 -4887
rect -17346 -5142 -17312 -5036
rect -17250 -5036 -17216 -5021
rect -17250 -5055 -17216 -5036
rect -17154 -5142 -17120 -5122
rect -17154 -5156 -17120 -5142
rect -17058 -5036 -17024 -5021
rect -17058 -5055 -17024 -5036
rect -16962 -5142 -16928 -5122
rect -16962 -5156 -16928 -5142
rect -16866 -5036 -16832 -5022
rect -16866 -5056 -16832 -5036
rect -16770 -5142 -16736 -5122
rect -16770 -5156 -16736 -5142
rect -16674 -5036 -16640 -5021
rect -16674 -5055 -16640 -5036
rect -16578 -5142 -16544 -5122
rect -16578 -5156 -16544 -5142
rect -16482 -5036 -16448 -5021
rect -16482 -5055 -16448 -5036
rect -16386 -5142 -16352 -5122
rect -16386 -5156 -16352 -5142
rect -16290 -5036 -16256 -5021
rect -16290 -5055 -16256 -5036
rect -16194 -5142 -16160 -5036
rect -16006 -4770 -15933 -4667
rect -15689 -4776 -15556 -4723
rect -14055 -4104 -14021 -4002
rect -14055 -4499 -14021 -4397
rect -13959 -4312 -13925 -4188
rect -13863 -4104 -13829 -4002
rect -13863 -4463 -13829 -4397
rect -13767 -4312 -13733 -4188
rect -13671 -4106 -13637 -4004
rect -13671 -4463 -13637 -4403
rect -13575 -4312 -13541 -4188
rect -13479 -4107 -13445 -4005
rect -13479 -4463 -13445 -4420
rect -13383 -4312 -13349 -4188
rect -13287 -4107 -13253 -4005
rect -13287 -4463 -13253 -4403
rect -13191 -4312 -13157 -4188
rect -13095 -4107 -13061 -4005
rect -13095 -4463 -13061 -4396
rect -12999 -4313 -12965 -4189
rect -12903 -4107 -12869 -4005
rect -12903 -4463 -12869 -4396
rect -15083 -4768 -14969 -4715
rect -14849 -4722 -14769 -4716
rect -14849 -4777 -14841 -4722
rect -14841 -4777 -14776 -4722
rect -14776 -4777 -14769 -4722
rect -14849 -4784 -14769 -4777
rect -14667 -4942 -14602 -4887
rect -15787 -5142 -15753 -5036
rect -15691 -5036 -15657 -5021
rect -15691 -5055 -15657 -5036
rect -15595 -5142 -15561 -5122
rect -15595 -5156 -15561 -5142
rect -15499 -5036 -15465 -5021
rect -15499 -5055 -15465 -5036
rect -15403 -5142 -15369 -5122
rect -15403 -5156 -15369 -5142
rect -15307 -5036 -15273 -5022
rect -15307 -5056 -15273 -5036
rect -15211 -5142 -15177 -5122
rect -15211 -5156 -15177 -5142
rect -15115 -5036 -15081 -5021
rect -15115 -5055 -15081 -5036
rect -15019 -5142 -14985 -5122
rect -15019 -5156 -14985 -5142
rect -14923 -5036 -14889 -5021
rect -14923 -5055 -14889 -5036
rect -14827 -5142 -14793 -5122
rect -14827 -5156 -14793 -5142
rect -14731 -5036 -14697 -5021
rect -14731 -5055 -14697 -5036
rect -14635 -5142 -14601 -5036
rect -14272 -4732 -14225 -4622
rect -13957 -4776 -13824 -4723
rect -12496 -4104 -12462 -4002
rect -12496 -4499 -12462 -4397
rect -12400 -4312 -12366 -4188
rect -12304 -4104 -12270 -4002
rect -12304 -4463 -12270 -4397
rect -12208 -4312 -12174 -4188
rect -12112 -4106 -12078 -4004
rect -12112 -4463 -12078 -4403
rect -12016 -4312 -11982 -4188
rect -11920 -4107 -11886 -4005
rect -11920 -4463 -11886 -4420
rect -11824 -4312 -11790 -4188
rect -11728 -4107 -11694 -4005
rect -11728 -4463 -11694 -4403
rect -11632 -4312 -11598 -4188
rect -11536 -4107 -11502 -4005
rect -11536 -4463 -11502 -4396
rect -11440 -4313 -11406 -4189
rect -11344 -4107 -11310 -4005
rect -11344 -4463 -11310 -4396
rect -13351 -4768 -13237 -4715
rect -13117 -4722 -13037 -4716
rect -13117 -4777 -13109 -4722
rect -13109 -4777 -13044 -4722
rect -13044 -4777 -13037 -4722
rect -13117 -4784 -13037 -4777
rect -12935 -4942 -12870 -4887
rect -14055 -5142 -14021 -5036
rect -13959 -5036 -13925 -5021
rect -13959 -5055 -13925 -5036
rect -13863 -5142 -13829 -5122
rect -13863 -5156 -13829 -5142
rect -13767 -5036 -13733 -5021
rect -13767 -5055 -13733 -5036
rect -13671 -5142 -13637 -5122
rect -13671 -5156 -13637 -5142
rect -13575 -5036 -13541 -5022
rect -13575 -5056 -13541 -5036
rect -13479 -5142 -13445 -5122
rect -13479 -5156 -13445 -5142
rect -13383 -5036 -13349 -5021
rect -13383 -5055 -13349 -5036
rect -13287 -5142 -13253 -5122
rect -13287 -5156 -13253 -5142
rect -13191 -5036 -13157 -5021
rect -13191 -5055 -13157 -5036
rect -13095 -5142 -13061 -5122
rect -13095 -5156 -13061 -5142
rect -12999 -5036 -12965 -5021
rect -12999 -5055 -12965 -5036
rect -12903 -5142 -12869 -5036
rect -12715 -4770 -12642 -4667
rect -12398 -4776 -12265 -4723
rect -10764 -4104 -10730 -4002
rect -10764 -4499 -10730 -4397
rect -10668 -4312 -10634 -4188
rect -10572 -4104 -10538 -4002
rect -10572 -4463 -10538 -4397
rect -10476 -4312 -10442 -4188
rect -10380 -4106 -10346 -4004
rect -10380 -4463 -10346 -4403
rect -10284 -4312 -10250 -4188
rect -10188 -4107 -10154 -4005
rect -10188 -4463 -10154 -4420
rect -10092 -4312 -10058 -4188
rect -9996 -4107 -9962 -4005
rect -9996 -4463 -9962 -4403
rect -9900 -4312 -9866 -4188
rect -9804 -4107 -9770 -4005
rect -9804 -4463 -9770 -4396
rect -9708 -4313 -9674 -4189
rect -9612 -4107 -9578 -4005
rect -9612 -4463 -9578 -4396
rect -11792 -4768 -11678 -4715
rect -11558 -4722 -11478 -4716
rect -11558 -4777 -11550 -4722
rect -11550 -4777 -11485 -4722
rect -11485 -4777 -11478 -4722
rect -11558 -4784 -11478 -4777
rect -11376 -4942 -11311 -4887
rect -12496 -5142 -12462 -5036
rect -12400 -5036 -12366 -5021
rect -12400 -5055 -12366 -5036
rect -12304 -5142 -12270 -5122
rect -12304 -5156 -12270 -5142
rect -12208 -5036 -12174 -5021
rect -12208 -5055 -12174 -5036
rect -12112 -5142 -12078 -5122
rect -12112 -5156 -12078 -5142
rect -12016 -5036 -11982 -5022
rect -12016 -5056 -11982 -5036
rect -11920 -5142 -11886 -5122
rect -11920 -5156 -11886 -5142
rect -11824 -5036 -11790 -5021
rect -11824 -5055 -11790 -5036
rect -11728 -5142 -11694 -5122
rect -11728 -5156 -11694 -5142
rect -11632 -5036 -11598 -5021
rect -11632 -5055 -11598 -5036
rect -11536 -5142 -11502 -5122
rect -11536 -5156 -11502 -5142
rect -11440 -5036 -11406 -5021
rect -11440 -5055 -11406 -5036
rect -11344 -5142 -11310 -5036
rect -10981 -4732 -10934 -4622
rect -10666 -4776 -10533 -4723
rect -9205 -4104 -9171 -4002
rect -9205 -4499 -9171 -4397
rect -9109 -4312 -9075 -4188
rect -9013 -4104 -8979 -4002
rect -9013 -4463 -8979 -4397
rect -8917 -4312 -8883 -4188
rect -8821 -4106 -8787 -4004
rect -8821 -4463 -8787 -4403
rect -8725 -4312 -8691 -4188
rect -8629 -4107 -8595 -4005
rect -8629 -4463 -8595 -4420
rect -8533 -4312 -8499 -4188
rect -8437 -4107 -8403 -4005
rect -8437 -4463 -8403 -4403
rect -8341 -4312 -8307 -4188
rect -8245 -4107 -8211 -4005
rect -8245 -4463 -8211 -4396
rect -8149 -4313 -8115 -4189
rect -8053 -4107 -8019 -4005
rect -8053 -4463 -8019 -4396
rect 7198 -4126 7232 -4092
rect 7390 -4126 7424 -4092
rect 7582 -4126 7616 -4092
rect 7774 -4126 7808 -4092
rect 8146 -4126 8180 -4092
rect 8338 -4126 8372 -4092
rect 8530 -4126 8564 -4092
rect 8722 -4126 8756 -4092
rect 9082 -4126 9116 -4092
rect 9274 -4126 9308 -4092
rect 9466 -4126 9500 -4092
rect 9658 -4126 9692 -4092
rect 10013 -4125 10047 -4091
rect 10205 -4125 10239 -4091
rect 10397 -4125 10431 -4091
rect 10589 -4125 10623 -4091
rect 10940 -4126 10974 -4092
rect 11132 -4126 11166 -4092
rect 11324 -4126 11358 -4092
rect 11516 -4126 11550 -4092
rect 7245 -4185 7280 -4180
rect 7245 -4292 7246 -4185
rect 7246 -4292 7280 -4185
rect 7150 -4480 7184 -4370
rect 7342 -4480 7376 -4370
rect 7438 -4185 7473 -4180
rect 7438 -4292 7472 -4185
rect 7472 -4292 7473 -4185
rect 7534 -4480 7568 -4370
rect 7630 -4185 7665 -4180
rect 7630 -4292 7664 -4185
rect 7664 -4292 7665 -4185
rect 7726 -4480 7760 -4370
rect 7822 -4185 7857 -4180
rect 7822 -4292 7856 -4185
rect 7856 -4292 7857 -4185
rect 7918 -4480 7952 -4370
rect 8193 -4185 8228 -4180
rect 8193 -4292 8194 -4185
rect 8194 -4292 8228 -4185
rect 8098 -4480 8132 -4370
rect 8290 -4480 8324 -4370
rect 8386 -4185 8421 -4180
rect 8386 -4292 8420 -4185
rect 8420 -4292 8421 -4185
rect 8482 -4480 8516 -4370
rect 8578 -4185 8613 -4180
rect 8578 -4292 8612 -4185
rect 8612 -4292 8613 -4185
rect 8674 -4480 8708 -4370
rect 8770 -4185 8805 -4180
rect 8770 -4292 8804 -4185
rect 8804 -4292 8805 -4185
rect 8866 -4480 8900 -4370
rect 9129 -4185 9164 -4180
rect 9129 -4292 9130 -4185
rect 9130 -4292 9164 -4185
rect 9034 -4480 9068 -4370
rect 9226 -4480 9260 -4370
rect 9322 -4185 9357 -4180
rect 9322 -4292 9356 -4185
rect 9356 -4292 9357 -4185
rect 9418 -4480 9452 -4370
rect 9514 -4185 9549 -4180
rect 9514 -4292 9548 -4185
rect 9548 -4292 9549 -4185
rect 9610 -4480 9644 -4370
rect 9706 -4185 9741 -4180
rect 9706 -4292 9740 -4185
rect 9740 -4292 9741 -4185
rect 9802 -4480 9836 -4370
rect 10060 -4184 10095 -4179
rect 10060 -4291 10061 -4184
rect 10061 -4291 10095 -4184
rect 9965 -4479 9999 -4369
rect 10157 -4479 10191 -4369
rect 10253 -4184 10288 -4179
rect 10253 -4291 10287 -4184
rect 10287 -4291 10288 -4184
rect 10349 -4479 10383 -4369
rect 10445 -4184 10480 -4179
rect 10445 -4291 10479 -4184
rect 10479 -4291 10480 -4184
rect 10541 -4479 10575 -4369
rect 10637 -4184 10672 -4179
rect 10637 -4291 10671 -4184
rect 10671 -4291 10672 -4184
rect 10733 -4479 10767 -4369
rect 10987 -4185 11022 -4180
rect 10987 -4292 10988 -4185
rect 10988 -4292 11022 -4185
rect 10892 -4480 10926 -4370
rect 11084 -4480 11118 -4370
rect 11180 -4185 11215 -4180
rect 11180 -4292 11214 -4185
rect 11214 -4292 11215 -4185
rect 11276 -4480 11310 -4370
rect 11372 -4185 11407 -4180
rect 11372 -4292 11406 -4185
rect 11406 -4292 11407 -4185
rect 11468 -4480 11502 -4370
rect 11564 -4185 11599 -4180
rect 11564 -4292 11598 -4185
rect 11598 -4292 11599 -4185
rect 11660 -4480 11694 -4370
rect -10060 -4768 -9946 -4715
rect -9826 -4722 -9746 -4716
rect -9826 -4777 -9818 -4722
rect -9818 -4777 -9753 -4722
rect -9753 -4777 -9746 -4722
rect -9826 -4784 -9746 -4777
rect -9644 -4942 -9579 -4887
rect -10764 -5142 -10730 -5036
rect -10668 -5036 -10634 -5021
rect -10668 -5055 -10634 -5036
rect -10572 -5142 -10538 -5122
rect -10572 -5156 -10538 -5142
rect -10476 -5036 -10442 -5021
rect -10476 -5055 -10442 -5036
rect -10380 -5142 -10346 -5122
rect -10380 -5156 -10346 -5142
rect -10284 -5036 -10250 -5022
rect -10284 -5056 -10250 -5036
rect -10188 -5142 -10154 -5122
rect -10188 -5156 -10154 -5142
rect -10092 -5036 -10058 -5021
rect -10092 -5055 -10058 -5036
rect -9996 -5142 -9962 -5122
rect -9996 -5156 -9962 -5142
rect -9900 -5036 -9866 -5021
rect -9900 -5055 -9866 -5036
rect -9804 -5142 -9770 -5122
rect -9804 -5156 -9770 -5142
rect -9708 -5036 -9674 -5021
rect -9708 -5055 -9674 -5036
rect -9612 -5142 -9578 -5036
rect -9424 -4770 -9351 -4667
rect -9107 -4776 -8974 -4723
rect 7389 -4587 7677 -4552
rect 8337 -4587 8625 -4552
rect 9273 -4587 9561 -4552
rect 10204 -4586 10492 -4551
rect 11131 -4587 11419 -4552
rect -8501 -4768 -8387 -4715
rect -8267 -4722 -8187 -4716
rect -8267 -4777 -8259 -4722
rect -8259 -4777 -8194 -4722
rect -8194 -4777 -8187 -4722
rect -8267 -4784 -8187 -4777
rect -8085 -4942 -8020 -4887
rect -9205 -5142 -9171 -5036
rect -9109 -5036 -9075 -5021
rect -9109 -5055 -9075 -5036
rect -9013 -5142 -8979 -5122
rect -9013 -5156 -8979 -5142
rect -8917 -5036 -8883 -5021
rect -8917 -5055 -8883 -5036
rect -8821 -5142 -8787 -5122
rect -8821 -5156 -8787 -5142
rect -8725 -5036 -8691 -5022
rect -8725 -5056 -8691 -5036
rect -8629 -5142 -8595 -5122
rect -8629 -5156 -8595 -5142
rect -8533 -5036 -8499 -5021
rect -8533 -5055 -8499 -5036
rect -8437 -5142 -8403 -5122
rect -8437 -5156 -8403 -5142
rect -8341 -5036 -8307 -5021
rect -8341 -5055 -8307 -5036
rect -8245 -5142 -8211 -5122
rect -8245 -5156 -8211 -5142
rect -8149 -5036 -8115 -5021
rect -8149 -5055 -8115 -5036
rect -8053 -5142 -8019 -5036
rect 5721 -5007 5812 -4973
rect 6161 -5007 6252 -4973
rect 6601 -5007 6692 -4973
rect 5664 -5079 5670 -5045
rect 5670 -5079 5743 -5045
rect -20603 -5276 -19480 -5230
rect -19044 -5276 -17921 -5230
rect -17312 -5276 -16189 -5230
rect -15753 -5276 -14630 -5230
rect -14021 -5276 -12898 -5230
rect -12462 -5276 -11339 -5230
rect -10730 -5276 -9607 -5230
rect -9171 -5276 -8048 -5230
rect 5577 -5319 5611 -5093
rect 6104 -5079 6110 -5045
rect 6110 -5079 6183 -5045
rect 5787 -5175 5864 -5141
rect 5664 -5271 5670 -5237
rect 5670 -5271 5743 -5237
rect -23523 -5385 -23432 -5351
rect -21789 -5385 -21698 -5351
rect -24368 -5451 -23799 -5404
rect -23580 -5457 -23574 -5423
rect -23574 -5457 -23501 -5423
rect -22632 -5451 -22063 -5404
rect -24384 -5529 -24350 -5523
rect -24384 -5603 -24350 -5529
rect -24288 -5719 -24254 -5645
rect -24288 -5725 -24254 -5719
rect -24192 -5529 -24158 -5523
rect -24192 -5603 -24158 -5529
rect -24096 -5719 -24062 -5645
rect -24096 -5725 -24062 -5719
rect -24000 -5529 -23966 -5523
rect -24000 -5603 -23966 -5529
rect -23904 -5719 -23870 -5645
rect -23904 -5725 -23870 -5719
rect -23808 -5529 -23774 -5523
rect -23808 -5603 -23774 -5529
rect -23667 -5697 -23633 -5471
rect -21846 -5457 -21840 -5423
rect -21840 -5457 -21767 -5423
rect -23457 -5553 -23380 -5519
rect -22648 -5529 -22614 -5523
rect -22648 -5603 -22614 -5529
rect -23580 -5649 -23574 -5615
rect -23574 -5649 -23501 -5615
rect -24318 -5813 -24284 -5778
rect -24029 -5813 -23995 -5778
rect -24234 -5937 -24200 -5902
rect -24150 -5907 -23774 -5873
rect -23457 -5745 -23380 -5711
rect -22552 -5719 -22518 -5645
rect -22552 -5725 -22518 -5719
rect -22456 -5529 -22422 -5523
rect -22456 -5603 -22422 -5529
rect -22360 -5719 -22326 -5645
rect -22360 -5725 -22326 -5719
rect -22264 -5529 -22230 -5523
rect -22264 -5603 -22230 -5529
rect -22168 -5719 -22134 -5645
rect -22168 -5725 -22134 -5719
rect -22072 -5529 -22038 -5523
rect -22072 -5603 -22038 -5529
rect -21933 -5697 -21899 -5471
rect -21723 -5553 -21646 -5519
rect 6017 -5319 6051 -5093
rect 6544 -5079 6550 -5045
rect 6550 -5079 6623 -5045
rect 6227 -5175 6304 -5141
rect 6104 -5271 6110 -5237
rect 6110 -5271 6183 -5237
rect 5787 -5367 5864 -5333
rect 5670 -5529 5846 -5495
rect -21846 -5649 -21840 -5615
rect -21840 -5649 -21767 -5615
rect -20502 -5619 -19933 -5572
rect -19393 -5619 -18824 -5572
rect -18511 -5619 -17942 -5572
rect -17211 -5619 -16642 -5572
rect -16102 -5619 -15533 -5572
rect -15220 -5619 -14651 -5572
rect -13920 -5619 -13351 -5572
rect -12811 -5619 -12242 -5572
rect -11929 -5619 -11360 -5572
rect -10629 -5619 -10060 -5572
rect -9520 -5619 -8951 -5572
rect -8638 -5619 -8069 -5572
rect 5577 -5573 5611 -5539
rect 6457 -5319 6491 -5093
rect 6667 -5175 6744 -5141
rect 6544 -5271 6550 -5237
rect 6550 -5271 6623 -5237
rect 6227 -5367 6304 -5333
rect 6110 -5529 6286 -5495
rect 6017 -5573 6051 -5539
rect 5670 -5617 5846 -5583
rect 6667 -5367 6744 -5333
rect 6550 -5529 6726 -5495
rect 6457 -5573 6491 -5539
rect 6110 -5617 6286 -5583
rect 6550 -5617 6726 -5583
rect 7389 -5680 7677 -5645
rect 8337 -5680 8625 -5645
rect 9273 -5680 9561 -5645
rect 10204 -5680 10492 -5645
rect 11131 -5680 11419 -5645
rect -22582 -5813 -22548 -5778
rect -22293 -5813 -22259 -5778
rect -23574 -5907 -23398 -5873
rect -23667 -5951 -23633 -5917
rect -23574 -5995 -23398 -5961
rect -22498 -5937 -22464 -5902
rect -22414 -5907 -22038 -5873
rect -20518 -5697 -20484 -5691
rect -21723 -5745 -21646 -5711
rect -20518 -5771 -20484 -5697
rect -21840 -5907 -21664 -5873
rect -20422 -5887 -20388 -5813
rect -20422 -5893 -20388 -5887
rect -20326 -5697 -20292 -5691
rect -20326 -5771 -20292 -5697
rect -20230 -5887 -20196 -5813
rect -20230 -5893 -20196 -5887
rect -20134 -5697 -20100 -5691
rect -20134 -5771 -20100 -5697
rect -20038 -5887 -20004 -5813
rect -20038 -5893 -20004 -5887
rect -19942 -5697 -19908 -5691
rect -19942 -5771 -19908 -5697
rect -19409 -5697 -19375 -5691
rect -19409 -5771 -19375 -5697
rect -19313 -5887 -19279 -5813
rect -19313 -5893 -19279 -5887
rect -19217 -5697 -19183 -5691
rect -19217 -5771 -19183 -5697
rect -19121 -5887 -19087 -5813
rect -19121 -5893 -19087 -5887
rect -19025 -5697 -18991 -5691
rect -19025 -5771 -18991 -5697
rect -18929 -5887 -18895 -5813
rect -18929 -5893 -18895 -5887
rect -18833 -5697 -18799 -5691
rect -18833 -5771 -18799 -5697
rect -18527 -5697 -18493 -5691
rect -18527 -5771 -18493 -5697
rect -18431 -5887 -18397 -5813
rect -18431 -5893 -18397 -5887
rect -18335 -5697 -18301 -5691
rect -18335 -5771 -18301 -5697
rect -18239 -5887 -18205 -5813
rect -18239 -5893 -18205 -5887
rect -18143 -5697 -18109 -5691
rect -18143 -5771 -18109 -5697
rect -18047 -5887 -18013 -5813
rect -18047 -5893 -18013 -5887
rect -17951 -5697 -17917 -5691
rect -17951 -5771 -17917 -5697
rect -17227 -5697 -17193 -5691
rect -17227 -5771 -17193 -5697
rect -17131 -5887 -17097 -5813
rect -17131 -5893 -17097 -5887
rect -17035 -5697 -17001 -5691
rect -17035 -5771 -17001 -5697
rect -16939 -5887 -16905 -5813
rect -16939 -5893 -16905 -5887
rect -16843 -5697 -16809 -5691
rect -16843 -5771 -16809 -5697
rect -16747 -5887 -16713 -5813
rect -16747 -5893 -16713 -5887
rect -16651 -5697 -16617 -5691
rect -16651 -5771 -16617 -5697
rect -16118 -5697 -16084 -5691
rect -16118 -5771 -16084 -5697
rect -16022 -5887 -15988 -5813
rect -16022 -5893 -15988 -5887
rect -15926 -5697 -15892 -5691
rect -15926 -5771 -15892 -5697
rect -15830 -5887 -15796 -5813
rect -15830 -5893 -15796 -5887
rect -15734 -5697 -15700 -5691
rect -15734 -5771 -15700 -5697
rect -15638 -5887 -15604 -5813
rect -15638 -5893 -15604 -5887
rect -15542 -5697 -15508 -5691
rect -15542 -5771 -15508 -5697
rect -15236 -5697 -15202 -5691
rect -15236 -5771 -15202 -5697
rect -15140 -5887 -15106 -5813
rect -15140 -5893 -15106 -5887
rect -15044 -5697 -15010 -5691
rect -15044 -5771 -15010 -5697
rect -14948 -5887 -14914 -5813
rect -14948 -5893 -14914 -5887
rect -14852 -5697 -14818 -5691
rect -14852 -5771 -14818 -5697
rect -14756 -5887 -14722 -5813
rect -14756 -5893 -14722 -5887
rect -14660 -5697 -14626 -5691
rect -14660 -5771 -14626 -5697
rect -13936 -5697 -13902 -5691
rect -13936 -5771 -13902 -5697
rect -13840 -5887 -13806 -5813
rect -13840 -5893 -13806 -5887
rect -13744 -5697 -13710 -5691
rect -13744 -5771 -13710 -5697
rect -13648 -5887 -13614 -5813
rect -13648 -5893 -13614 -5887
rect -13552 -5697 -13518 -5691
rect -13552 -5771 -13518 -5697
rect -13456 -5887 -13422 -5813
rect -13456 -5893 -13422 -5887
rect -13360 -5697 -13326 -5691
rect -13360 -5771 -13326 -5697
rect -12827 -5697 -12793 -5691
rect -12827 -5771 -12793 -5697
rect -12731 -5887 -12697 -5813
rect -12731 -5893 -12697 -5887
rect -12635 -5697 -12601 -5691
rect -12635 -5771 -12601 -5697
rect -12539 -5887 -12505 -5813
rect -12539 -5893 -12505 -5887
rect -12443 -5697 -12409 -5691
rect -12443 -5771 -12409 -5697
rect -12347 -5887 -12313 -5813
rect -12347 -5893 -12313 -5887
rect -12251 -5697 -12217 -5691
rect -12251 -5771 -12217 -5697
rect -11945 -5697 -11911 -5691
rect -11945 -5771 -11911 -5697
rect -11849 -5887 -11815 -5813
rect -11849 -5893 -11815 -5887
rect -11753 -5697 -11719 -5691
rect -11753 -5771 -11719 -5697
rect -11657 -5887 -11623 -5813
rect -11657 -5893 -11623 -5887
rect -11561 -5697 -11527 -5691
rect -11561 -5771 -11527 -5697
rect -11465 -5887 -11431 -5813
rect -11465 -5893 -11431 -5887
rect -11369 -5697 -11335 -5691
rect -11369 -5771 -11335 -5697
rect -10645 -5697 -10611 -5691
rect -10645 -5771 -10611 -5697
rect -10549 -5887 -10515 -5813
rect -10549 -5893 -10515 -5887
rect -10453 -5697 -10419 -5691
rect -10453 -5771 -10419 -5697
rect -10357 -5887 -10323 -5813
rect -10357 -5893 -10323 -5887
rect -10261 -5697 -10227 -5691
rect -10261 -5771 -10227 -5697
rect -10165 -5887 -10131 -5813
rect -10165 -5893 -10131 -5887
rect -10069 -5697 -10035 -5691
rect -10069 -5771 -10035 -5697
rect -9536 -5697 -9502 -5691
rect -9536 -5771 -9502 -5697
rect -9440 -5887 -9406 -5813
rect -9440 -5893 -9406 -5887
rect -9344 -5697 -9310 -5691
rect -9344 -5771 -9310 -5697
rect -9248 -5887 -9214 -5813
rect -9248 -5893 -9214 -5887
rect -9152 -5697 -9118 -5691
rect -9152 -5771 -9118 -5697
rect -9056 -5887 -9022 -5813
rect -9056 -5893 -9022 -5887
rect -8960 -5697 -8926 -5691
rect -8960 -5771 -8926 -5697
rect -8654 -5697 -8620 -5691
rect -8654 -5771 -8620 -5697
rect -8558 -5887 -8524 -5813
rect -8558 -5893 -8524 -5887
rect -8462 -5697 -8428 -5691
rect -8462 -5771 -8428 -5697
rect -8366 -5887 -8332 -5813
rect -8366 -5893 -8332 -5887
rect -8270 -5697 -8236 -5691
rect -8270 -5771 -8236 -5697
rect -8174 -5887 -8140 -5813
rect -8174 -5893 -8140 -5887
rect -8078 -5697 -8044 -5691
rect -8078 -5771 -8044 -5697
rect 5689 -5719 5821 -5685
rect 6129 -5719 6261 -5685
rect 6569 -5719 6701 -5685
rect 7150 -5862 7184 -5752
rect -21933 -5951 -21899 -5917
rect -21840 -5995 -21664 -5961
rect -20452 -5981 -20418 -5946
rect -20163 -5981 -20129 -5946
rect -24150 -6099 -23774 -6065
rect -23555 -6097 -23423 -6063
rect -22414 -6099 -22038 -6065
rect -21821 -6097 -21689 -6063
rect -24135 -6171 -23800 -6137
rect -22399 -6171 -22064 -6137
rect -19343 -5981 -19309 -5946
rect -19054 -5981 -19020 -5946
rect -20368 -6105 -20334 -6070
rect -20284 -6075 -19908 -6041
rect -18461 -5981 -18427 -5946
rect -18172 -5981 -18138 -5946
rect -19259 -6105 -19225 -6070
rect -19175 -6075 -18799 -6041
rect -17161 -5981 -17127 -5946
rect -16872 -5981 -16838 -5946
rect -18377 -6105 -18343 -6070
rect -18293 -6075 -17917 -6041
rect -16052 -5981 -16018 -5946
rect -15763 -5981 -15729 -5946
rect -17077 -6105 -17043 -6070
rect -16993 -6075 -16617 -6041
rect -15170 -5981 -15136 -5946
rect -14881 -5981 -14847 -5946
rect -15968 -6105 -15934 -6070
rect -15884 -6075 -15508 -6041
rect -13870 -5981 -13836 -5946
rect -13581 -5981 -13547 -5946
rect -15086 -6105 -15052 -6070
rect -15002 -6075 -14626 -6041
rect -12761 -5981 -12727 -5946
rect -12472 -5981 -12438 -5946
rect -13786 -6105 -13752 -6070
rect -13702 -6075 -13326 -6041
rect -11879 -5981 -11845 -5946
rect -11590 -5981 -11556 -5946
rect -12677 -6105 -12643 -6070
rect -12593 -6075 -12217 -6041
rect -10579 -5981 -10545 -5946
rect -10290 -5981 -10256 -5946
rect -11795 -6105 -11761 -6070
rect -11711 -6075 -11335 -6041
rect -9470 -5981 -9436 -5946
rect -9181 -5981 -9147 -5946
rect -10495 -6105 -10461 -6070
rect -10411 -6075 -10035 -6041
rect -8588 -5981 -8554 -5946
rect -8299 -5981 -8265 -5946
rect -9386 -6105 -9352 -6070
rect -9302 -6075 -8926 -6041
rect -8504 -6105 -8470 -6070
rect -8420 -6075 -8044 -6041
rect 7245 -6047 7246 -5940
rect 7246 -6047 7280 -5940
rect 7245 -6052 7280 -6047
rect 7342 -5862 7376 -5752
rect 7534 -5862 7568 -5752
rect 7438 -6047 7472 -5940
rect 7472 -6047 7473 -5940
rect 7438 -6052 7473 -6047
rect 7726 -5862 7760 -5752
rect 7630 -6047 7664 -5940
rect 7664 -6047 7665 -5940
rect 7630 -6052 7665 -6047
rect 7918 -5862 7952 -5752
rect 7822 -6047 7856 -5940
rect 7856 -6047 7857 -5940
rect 7822 -6052 7857 -6047
rect 8098 -5862 8132 -5752
rect 8193 -6047 8194 -5940
rect 8194 -6047 8228 -5940
rect 8193 -6052 8228 -6047
rect 8290 -5862 8324 -5752
rect 8482 -5862 8516 -5752
rect 8386 -6047 8420 -5940
rect 8420 -6047 8421 -5940
rect 8386 -6052 8421 -6047
rect 8674 -5862 8708 -5752
rect 8578 -6047 8612 -5940
rect 8612 -6047 8613 -5940
rect 8578 -6052 8613 -6047
rect 8866 -5862 8900 -5752
rect 8770 -6047 8804 -5940
rect 8804 -6047 8805 -5940
rect 8770 -6052 8805 -6047
rect 9034 -5862 9068 -5752
rect 9129 -6047 9130 -5940
rect 9130 -6047 9164 -5940
rect 9129 -6052 9164 -6047
rect 9226 -5862 9260 -5752
rect 9418 -5862 9452 -5752
rect 9322 -6047 9356 -5940
rect 9356 -6047 9357 -5940
rect 9322 -6052 9357 -6047
rect 9610 -5862 9644 -5752
rect 9514 -6047 9548 -5940
rect 9548 -6047 9549 -5940
rect 9514 -6052 9549 -6047
rect 9802 -5862 9836 -5752
rect 9706 -6047 9740 -5940
rect 9740 -6047 9741 -5940
rect 9706 -6052 9741 -6047
rect 9965 -5862 9999 -5752
rect 10060 -6047 10061 -5940
rect 10061 -6047 10095 -5940
rect 10060 -6052 10095 -6047
rect 10157 -5862 10191 -5752
rect 10349 -5862 10383 -5752
rect 10253 -6047 10287 -5940
rect 10287 -6047 10288 -5940
rect 10253 -6052 10288 -6047
rect 10541 -5862 10575 -5752
rect 10445 -6047 10479 -5940
rect 10479 -6047 10480 -5940
rect 10445 -6052 10480 -6047
rect 10733 -5862 10767 -5752
rect 10637 -6047 10671 -5940
rect 10671 -6047 10672 -5940
rect 10637 -6052 10672 -6047
rect 10892 -5862 10926 -5752
rect 10987 -6047 10988 -5940
rect 10988 -6047 11022 -5940
rect 10987 -6052 11022 -6047
rect 11084 -5862 11118 -5752
rect 11276 -5862 11310 -5752
rect 11180 -6047 11214 -5940
rect 11214 -6047 11215 -5940
rect 11180 -6052 11215 -6047
rect 11468 -5862 11502 -5752
rect 11372 -6047 11406 -5940
rect 11406 -6047 11407 -5940
rect 11372 -6052 11407 -6047
rect 11660 -5862 11694 -5752
rect 11564 -6047 11598 -5940
rect 11598 -6047 11599 -5940
rect 11564 -6052 11599 -6047
rect 7198 -6140 7232 -6106
rect 7390 -6140 7424 -6106
rect 7582 -6140 7616 -6106
rect 7774 -6140 7808 -6106
rect 8146 -6140 8180 -6106
rect 8338 -6140 8372 -6106
rect 8530 -6140 8564 -6106
rect 8722 -6140 8756 -6106
rect 9082 -6140 9116 -6106
rect 9274 -6140 9308 -6106
rect 9466 -6140 9500 -6106
rect 9658 -6140 9692 -6106
rect 10013 -6140 10047 -6106
rect 10205 -6140 10239 -6106
rect 10397 -6140 10431 -6106
rect 10589 -6140 10623 -6106
rect 10940 -6140 10974 -6106
rect 11132 -6140 11166 -6106
rect 11324 -6140 11358 -6106
rect 11516 -6140 11550 -6106
rect -20284 -6267 -19908 -6233
rect -19175 -6267 -18799 -6233
rect -18293 -6267 -17917 -6233
rect -16993 -6267 -16617 -6233
rect -15884 -6267 -15508 -6233
rect -15002 -6267 -14626 -6233
rect -13702 -6267 -13326 -6233
rect -12593 -6267 -12217 -6233
rect -11711 -6267 -11335 -6233
rect -10411 -6267 -10035 -6233
rect -9302 -6267 -8926 -6233
rect -8420 -6267 -8044 -6233
rect -20269 -6339 -19934 -6305
rect -19160 -6339 -18825 -6305
rect -18278 -6339 -17943 -6305
rect -16978 -6339 -16643 -6305
rect -15869 -6339 -15534 -6305
rect -14987 -6339 -14652 -6305
rect -13687 -6339 -13352 -6305
rect -12578 -6339 -12243 -6305
rect -11696 -6339 -11361 -6305
rect -10396 -6339 -10061 -6305
rect -9287 -6339 -8952 -6305
rect -8405 -6339 -8070 -6305
rect 7298 -6838 7332 -6490
rect 7332 -6838 7333 -6490
rect 7298 -6890 7333 -6838
rect -20603 -7164 -19481 -7092
rect -19044 -7164 -17922 -7092
rect -17312 -7164 -16190 -7092
rect -15753 -7164 -14631 -7092
rect -14021 -7164 -12899 -7092
rect -12462 -7164 -11340 -7092
rect -10730 -7164 -9608 -7092
rect -9171 -7164 -8049 -7092
rect 7298 -7241 7332 -6890
rect 7332 -7241 7333 -6890
rect -23521 -7358 -23430 -7324
rect -21787 -7358 -21696 -7324
rect -24368 -7424 -23799 -7377
rect -23578 -7430 -23572 -7396
rect -23572 -7430 -23499 -7396
rect -22631 -7424 -22062 -7377
rect -24384 -7502 -24350 -7496
rect -24384 -7576 -24350 -7502
rect -24288 -7692 -24254 -7618
rect -24288 -7698 -24254 -7692
rect -24192 -7502 -24158 -7496
rect -24192 -7576 -24158 -7502
rect -24096 -7692 -24062 -7618
rect -24096 -7698 -24062 -7692
rect -24000 -7502 -23966 -7496
rect -24000 -7576 -23966 -7502
rect -23904 -7692 -23870 -7618
rect -23904 -7698 -23870 -7692
rect -23808 -7502 -23774 -7496
rect -23808 -7576 -23774 -7502
rect -23665 -7670 -23631 -7444
rect -21844 -7430 -21838 -7396
rect -21838 -7430 -21765 -7396
rect -23455 -7526 -23378 -7492
rect -22647 -7502 -22613 -7496
rect -22647 -7576 -22613 -7502
rect -23578 -7622 -23572 -7588
rect -23572 -7622 -23499 -7588
rect -24318 -7786 -24284 -7751
rect -24029 -7786 -23995 -7751
rect -24234 -7910 -24200 -7875
rect -24150 -7880 -23774 -7846
rect -23455 -7718 -23378 -7684
rect -22551 -7692 -22517 -7618
rect -22551 -7698 -22517 -7692
rect -22455 -7502 -22421 -7496
rect -22455 -7576 -22421 -7502
rect -22359 -7692 -22325 -7618
rect -22359 -7698 -22325 -7692
rect -22263 -7502 -22229 -7496
rect -22263 -7576 -22229 -7502
rect -22167 -7692 -22133 -7618
rect -22167 -7698 -22133 -7692
rect -22071 -7502 -22037 -7496
rect -22071 -7576 -22037 -7502
rect -21931 -7670 -21897 -7444
rect -21721 -7526 -21644 -7492
rect -21844 -7622 -21838 -7588
rect -21838 -7622 -21765 -7588
rect -22581 -7786 -22547 -7751
rect -22292 -7786 -22258 -7751
rect -23572 -7880 -23396 -7846
rect -23665 -7924 -23631 -7890
rect -23572 -7968 -23396 -7934
rect -22497 -7910 -22463 -7875
rect -22413 -7880 -22037 -7846
rect -21721 -7718 -21644 -7684
rect -21838 -7880 -21662 -7846
rect -20637 -7369 -20603 -7267
rect -20637 -7764 -20603 -7662
rect -20541 -7577 -20507 -7453
rect -20445 -7369 -20411 -7267
rect -20445 -7728 -20411 -7662
rect -20349 -7577 -20315 -7453
rect -20253 -7371 -20219 -7269
rect -20253 -7728 -20219 -7668
rect -20157 -7577 -20123 -7453
rect -20061 -7372 -20027 -7270
rect -20061 -7728 -20027 -7685
rect -19965 -7577 -19931 -7453
rect -19869 -7372 -19835 -7270
rect -19869 -7728 -19835 -7668
rect -19773 -7577 -19739 -7453
rect -19677 -7372 -19643 -7270
rect -19677 -7728 -19643 -7661
rect -19581 -7578 -19547 -7454
rect -19485 -7372 -19451 -7270
rect -19485 -7728 -19451 -7661
rect -21931 -7924 -21897 -7890
rect -21838 -7968 -21662 -7934
rect -24150 -8072 -23774 -8038
rect -23553 -8070 -23421 -8036
rect -20854 -7997 -20807 -7887
rect -22413 -8072 -22037 -8038
rect -21819 -8070 -21687 -8036
rect -24135 -8144 -23800 -8110
rect -22398 -8144 -22063 -8110
rect -20539 -8041 -20406 -7988
rect -19078 -7369 -19044 -7267
rect -19078 -7764 -19044 -7662
rect -18982 -7577 -18948 -7453
rect -18886 -7369 -18852 -7267
rect -18886 -7728 -18852 -7662
rect -18790 -7577 -18756 -7453
rect -18694 -7371 -18660 -7269
rect -18694 -7728 -18660 -7668
rect -18598 -7577 -18564 -7453
rect -18502 -7372 -18468 -7270
rect -18502 -7728 -18468 -7685
rect -18406 -7577 -18372 -7453
rect -18310 -7372 -18276 -7270
rect -18310 -7728 -18276 -7668
rect -18214 -7577 -18180 -7453
rect -18118 -7372 -18084 -7270
rect -18118 -7728 -18084 -7661
rect -18022 -7578 -17988 -7454
rect -17926 -7372 -17892 -7270
rect -17926 -7728 -17892 -7661
rect -19933 -8033 -19819 -7980
rect -19699 -7987 -19619 -7981
rect -19699 -8042 -19691 -7987
rect -19691 -8042 -19626 -7987
rect -19626 -8042 -19619 -7987
rect -19699 -8049 -19619 -8042
rect -19517 -8207 -19452 -8152
rect -20637 -8407 -20603 -8301
rect -20541 -8301 -20507 -8286
rect -20541 -8320 -20507 -8301
rect -20445 -8407 -20411 -8387
rect -20445 -8421 -20411 -8407
rect -20349 -8301 -20315 -8286
rect -20349 -8320 -20315 -8301
rect -20253 -8407 -20219 -8387
rect -20253 -8421 -20219 -8407
rect -20157 -8301 -20123 -8287
rect -20157 -8321 -20123 -8301
rect -20061 -8407 -20027 -8387
rect -20061 -8421 -20027 -8407
rect -19965 -8301 -19931 -8286
rect -19965 -8320 -19931 -8301
rect -19869 -8407 -19835 -8387
rect -19869 -8421 -19835 -8407
rect -19773 -8301 -19739 -8286
rect -19773 -8320 -19739 -8301
rect -19677 -8407 -19643 -8387
rect -19677 -8421 -19643 -8407
rect -19581 -8301 -19547 -8286
rect -19581 -8320 -19547 -8301
rect -19485 -8407 -19451 -8301
rect -19297 -8035 -19224 -7932
rect -18980 -8041 -18847 -7988
rect -17346 -7369 -17312 -7267
rect -17346 -7764 -17312 -7662
rect -17250 -7577 -17216 -7453
rect -17154 -7369 -17120 -7267
rect -17154 -7728 -17120 -7662
rect -17058 -7577 -17024 -7453
rect -16962 -7371 -16928 -7269
rect -16962 -7728 -16928 -7668
rect -16866 -7577 -16832 -7453
rect -16770 -7372 -16736 -7270
rect -16770 -7728 -16736 -7685
rect -16674 -7577 -16640 -7453
rect -16578 -7372 -16544 -7270
rect -16578 -7728 -16544 -7668
rect -16482 -7577 -16448 -7453
rect -16386 -7372 -16352 -7270
rect -16386 -7728 -16352 -7661
rect -16290 -7578 -16256 -7454
rect -16194 -7372 -16160 -7270
rect -16194 -7728 -16160 -7661
rect -18374 -8033 -18260 -7980
rect -18140 -7987 -18060 -7981
rect -18140 -8042 -18132 -7987
rect -18132 -8042 -18067 -7987
rect -18067 -8042 -18060 -7987
rect -18140 -8049 -18060 -8042
rect -17958 -8207 -17893 -8152
rect -19078 -8407 -19044 -8301
rect -18982 -8301 -18948 -8286
rect -18982 -8320 -18948 -8301
rect -18886 -8407 -18852 -8387
rect -18886 -8421 -18852 -8407
rect -18790 -8301 -18756 -8286
rect -18790 -8320 -18756 -8301
rect -18694 -8407 -18660 -8387
rect -18694 -8421 -18660 -8407
rect -18598 -8301 -18564 -8287
rect -18598 -8321 -18564 -8301
rect -18502 -8407 -18468 -8387
rect -18502 -8421 -18468 -8407
rect -18406 -8301 -18372 -8286
rect -18406 -8320 -18372 -8301
rect -18310 -8407 -18276 -8387
rect -18310 -8421 -18276 -8407
rect -18214 -8301 -18180 -8286
rect -18214 -8320 -18180 -8301
rect -18118 -8407 -18084 -8387
rect -18118 -8421 -18084 -8407
rect -18022 -8301 -17988 -8286
rect -18022 -8320 -17988 -8301
rect -17926 -8407 -17892 -8301
rect -17563 -7997 -17516 -7887
rect -17248 -8041 -17115 -7988
rect -15787 -7369 -15753 -7267
rect -15787 -7764 -15753 -7662
rect -15691 -7577 -15657 -7453
rect -15595 -7369 -15561 -7267
rect -15595 -7728 -15561 -7662
rect -15499 -7577 -15465 -7453
rect -15403 -7371 -15369 -7269
rect -15403 -7728 -15369 -7668
rect -15307 -7577 -15273 -7453
rect -15211 -7372 -15177 -7270
rect -15211 -7728 -15177 -7685
rect -15115 -7577 -15081 -7453
rect -15019 -7372 -14985 -7270
rect -15019 -7728 -14985 -7668
rect -14923 -7577 -14889 -7453
rect -14827 -7372 -14793 -7270
rect -14827 -7728 -14793 -7661
rect -14731 -7578 -14697 -7454
rect -14635 -7372 -14601 -7270
rect -14635 -7728 -14601 -7661
rect -16642 -8033 -16528 -7980
rect -16408 -7987 -16328 -7981
rect -16408 -8042 -16400 -7987
rect -16400 -8042 -16335 -7987
rect -16335 -8042 -16328 -7987
rect -16408 -8049 -16328 -8042
rect -16226 -8207 -16161 -8152
rect -17346 -8407 -17312 -8301
rect -17250 -8301 -17216 -8286
rect -17250 -8320 -17216 -8301
rect -17154 -8407 -17120 -8387
rect -17154 -8421 -17120 -8407
rect -17058 -8301 -17024 -8286
rect -17058 -8320 -17024 -8301
rect -16962 -8407 -16928 -8387
rect -16962 -8421 -16928 -8407
rect -16866 -8301 -16832 -8287
rect -16866 -8321 -16832 -8301
rect -16770 -8407 -16736 -8387
rect -16770 -8421 -16736 -8407
rect -16674 -8301 -16640 -8286
rect -16674 -8320 -16640 -8301
rect -16578 -8407 -16544 -8387
rect -16578 -8421 -16544 -8407
rect -16482 -8301 -16448 -8286
rect -16482 -8320 -16448 -8301
rect -16386 -8407 -16352 -8387
rect -16386 -8421 -16352 -8407
rect -16290 -8301 -16256 -8286
rect -16290 -8320 -16256 -8301
rect -16194 -8407 -16160 -8301
rect -16006 -8035 -15933 -7932
rect -15689 -8041 -15556 -7988
rect -14055 -7369 -14021 -7267
rect -14055 -7764 -14021 -7662
rect -13959 -7577 -13925 -7453
rect -13863 -7369 -13829 -7267
rect -13863 -7728 -13829 -7662
rect -13767 -7577 -13733 -7453
rect -13671 -7371 -13637 -7269
rect -13671 -7728 -13637 -7668
rect -13575 -7577 -13541 -7453
rect -13479 -7372 -13445 -7270
rect -13479 -7728 -13445 -7685
rect -13383 -7577 -13349 -7453
rect -13287 -7372 -13253 -7270
rect -13287 -7728 -13253 -7668
rect -13191 -7577 -13157 -7453
rect -13095 -7372 -13061 -7270
rect -13095 -7728 -13061 -7661
rect -12999 -7578 -12965 -7454
rect -12903 -7372 -12869 -7270
rect -12903 -7728 -12869 -7661
rect -15083 -8033 -14969 -7980
rect -14849 -7987 -14769 -7981
rect -14849 -8042 -14841 -7987
rect -14841 -8042 -14776 -7987
rect -14776 -8042 -14769 -7987
rect -14849 -8049 -14769 -8042
rect -14667 -8207 -14602 -8152
rect -15787 -8407 -15753 -8301
rect -15691 -8301 -15657 -8286
rect -15691 -8320 -15657 -8301
rect -15595 -8407 -15561 -8387
rect -15595 -8421 -15561 -8407
rect -15499 -8301 -15465 -8286
rect -15499 -8320 -15465 -8301
rect -15403 -8407 -15369 -8387
rect -15403 -8421 -15369 -8407
rect -15307 -8301 -15273 -8287
rect -15307 -8321 -15273 -8301
rect -15211 -8407 -15177 -8387
rect -15211 -8421 -15177 -8407
rect -15115 -8301 -15081 -8286
rect -15115 -8320 -15081 -8301
rect -15019 -8407 -14985 -8387
rect -15019 -8421 -14985 -8407
rect -14923 -8301 -14889 -8286
rect -14923 -8320 -14889 -8301
rect -14827 -8407 -14793 -8387
rect -14827 -8421 -14793 -8407
rect -14731 -8301 -14697 -8286
rect -14731 -8320 -14697 -8301
rect -14635 -8407 -14601 -8301
rect -14272 -7997 -14225 -7887
rect -13957 -8041 -13824 -7988
rect -12496 -7369 -12462 -7267
rect -12496 -7764 -12462 -7662
rect -12400 -7577 -12366 -7453
rect -12304 -7369 -12270 -7267
rect -12304 -7728 -12270 -7662
rect -12208 -7577 -12174 -7453
rect -12112 -7371 -12078 -7269
rect -12112 -7728 -12078 -7668
rect -12016 -7577 -11982 -7453
rect -11920 -7372 -11886 -7270
rect -11920 -7728 -11886 -7685
rect -11824 -7577 -11790 -7453
rect -11728 -7372 -11694 -7270
rect -11728 -7728 -11694 -7668
rect -11632 -7577 -11598 -7453
rect -11536 -7372 -11502 -7270
rect -11536 -7728 -11502 -7661
rect -11440 -7578 -11406 -7454
rect -11344 -7372 -11310 -7270
rect -11344 -7728 -11310 -7661
rect -13351 -8033 -13237 -7980
rect -13117 -7987 -13037 -7981
rect -13117 -8042 -13109 -7987
rect -13109 -8042 -13044 -7987
rect -13044 -8042 -13037 -7987
rect -13117 -8049 -13037 -8042
rect -12935 -8207 -12870 -8152
rect -14055 -8407 -14021 -8301
rect -13959 -8301 -13925 -8286
rect -13959 -8320 -13925 -8301
rect -13863 -8407 -13829 -8387
rect -13863 -8421 -13829 -8407
rect -13767 -8301 -13733 -8286
rect -13767 -8320 -13733 -8301
rect -13671 -8407 -13637 -8387
rect -13671 -8421 -13637 -8407
rect -13575 -8301 -13541 -8287
rect -13575 -8321 -13541 -8301
rect -13479 -8407 -13445 -8387
rect -13479 -8421 -13445 -8407
rect -13383 -8301 -13349 -8286
rect -13383 -8320 -13349 -8301
rect -13287 -8407 -13253 -8387
rect -13287 -8421 -13253 -8407
rect -13191 -8301 -13157 -8286
rect -13191 -8320 -13157 -8301
rect -13095 -8407 -13061 -8387
rect -13095 -8421 -13061 -8407
rect -12999 -8301 -12965 -8286
rect -12999 -8320 -12965 -8301
rect -12903 -8407 -12869 -8301
rect -12715 -8035 -12642 -7932
rect -12398 -8041 -12265 -7988
rect -10764 -7369 -10730 -7267
rect -10764 -7764 -10730 -7662
rect -10668 -7577 -10634 -7453
rect -10572 -7369 -10538 -7267
rect -10572 -7728 -10538 -7662
rect -10476 -7577 -10442 -7453
rect -10380 -7371 -10346 -7269
rect -10380 -7728 -10346 -7668
rect -10284 -7577 -10250 -7453
rect -10188 -7372 -10154 -7270
rect -10188 -7728 -10154 -7685
rect -10092 -7577 -10058 -7453
rect -9996 -7372 -9962 -7270
rect -9996 -7728 -9962 -7668
rect -9900 -7577 -9866 -7453
rect -9804 -7372 -9770 -7270
rect -9804 -7728 -9770 -7661
rect -9708 -7578 -9674 -7454
rect -9612 -7372 -9578 -7270
rect -9612 -7728 -9578 -7661
rect -11792 -8033 -11678 -7980
rect -11558 -7987 -11478 -7981
rect -11558 -8042 -11550 -7987
rect -11550 -8042 -11485 -7987
rect -11485 -8042 -11478 -7987
rect -11558 -8049 -11478 -8042
rect -11376 -8207 -11311 -8152
rect -12496 -8407 -12462 -8301
rect -12400 -8301 -12366 -8286
rect -12400 -8320 -12366 -8301
rect -12304 -8407 -12270 -8387
rect -12304 -8421 -12270 -8407
rect -12208 -8301 -12174 -8286
rect -12208 -8320 -12174 -8301
rect -12112 -8407 -12078 -8387
rect -12112 -8421 -12078 -8407
rect -12016 -8301 -11982 -8287
rect -12016 -8321 -11982 -8301
rect -11920 -8407 -11886 -8387
rect -11920 -8421 -11886 -8407
rect -11824 -8301 -11790 -8286
rect -11824 -8320 -11790 -8301
rect -11728 -8407 -11694 -8387
rect -11728 -8421 -11694 -8407
rect -11632 -8301 -11598 -8286
rect -11632 -8320 -11598 -8301
rect -11536 -8407 -11502 -8387
rect -11536 -8421 -11502 -8407
rect -11440 -8301 -11406 -8286
rect -11440 -8320 -11406 -8301
rect -11344 -8407 -11310 -8301
rect -10981 -7997 -10934 -7887
rect -10666 -8041 -10533 -7988
rect -9205 -7369 -9171 -7267
rect -9205 -7764 -9171 -7662
rect -9109 -7577 -9075 -7453
rect -9013 -7369 -8979 -7267
rect -9013 -7728 -8979 -7662
rect -8917 -7577 -8883 -7453
rect -8821 -7371 -8787 -7269
rect -8821 -7728 -8787 -7668
rect -8725 -7577 -8691 -7453
rect -8629 -7372 -8595 -7270
rect -8629 -7728 -8595 -7685
rect -8533 -7577 -8499 -7453
rect -8437 -7372 -8403 -7270
rect -8437 -7728 -8403 -7668
rect -8341 -7577 -8307 -7453
rect -8245 -7372 -8211 -7270
rect -8245 -7728 -8211 -7661
rect -8149 -7578 -8115 -7454
rect -8053 -7372 -8019 -7270
rect -8053 -7728 -8019 -7661
rect 7372 -7254 7406 -6478
rect 7756 -7254 7790 -6478
rect 8246 -6838 8280 -6490
rect 8280 -6838 8281 -6490
rect 8246 -6890 8281 -6838
rect 8246 -7241 8280 -6890
rect 8280 -7241 8281 -6890
rect 8320 -7254 8354 -6478
rect 8704 -7254 8738 -6478
rect 9182 -6838 9216 -6490
rect 9216 -6838 9217 -6490
rect 9182 -6890 9217 -6838
rect 9182 -7241 9216 -6890
rect 9216 -7241 9217 -6890
rect 9256 -7254 9290 -6478
rect 9640 -7254 9674 -6478
rect 10113 -6838 10147 -6490
rect 10147 -6838 10148 -6490
rect 10113 -6890 10148 -6838
rect 10113 -7241 10147 -6890
rect 10147 -7241 10148 -6890
rect 10187 -7254 10221 -6478
rect 10571 -7254 10605 -6478
rect 11040 -6838 11074 -6490
rect 11074 -6838 11075 -6490
rect 11040 -6890 11075 -6838
rect 11040 -7241 11074 -6890
rect 11074 -7241 11075 -6890
rect 11114 -7254 11148 -6478
rect 11498 -7254 11532 -6478
rect 11811 -6855 12168 -6804
rect 11785 -7191 11819 -7101
rect 11881 -7049 11915 -6959
rect 11977 -7191 12011 -7101
rect 12073 -7049 12107 -6959
rect 12169 -7191 12203 -7101
rect 12265 -7049 12299 -6959
rect 12361 -7191 12395 -7101
rect 12457 -7049 12491 -6959
rect 12553 -7191 12587 -7101
rect 12649 -7049 12683 -6959
rect 12986 -7025 13077 -6991
rect 12745 -7191 12779 -7101
rect 12929 -7097 12935 -7063
rect 12935 -7097 13008 -7063
rect 12170 -7287 12204 -7253
rect 12842 -7337 12876 -7111
rect 13052 -7193 13129 -7159
rect 12929 -7289 12935 -7255
rect 12935 -7289 13008 -7255
rect -10060 -8033 -9946 -7980
rect -9826 -7987 -9746 -7981
rect -9826 -8042 -9818 -7987
rect -9818 -8042 -9753 -7987
rect -9753 -8042 -9746 -7987
rect -9826 -8049 -9746 -8042
rect -9644 -8207 -9579 -8152
rect -10764 -8407 -10730 -8301
rect -10668 -8301 -10634 -8286
rect -10668 -8320 -10634 -8301
rect -10572 -8407 -10538 -8387
rect -10572 -8421 -10538 -8407
rect -10476 -8301 -10442 -8286
rect -10476 -8320 -10442 -8301
rect -10380 -8407 -10346 -8387
rect -10380 -8421 -10346 -8407
rect -10284 -8301 -10250 -8287
rect -10284 -8321 -10250 -8301
rect -10188 -8407 -10154 -8387
rect -10188 -8421 -10154 -8407
rect -10092 -8301 -10058 -8286
rect -10092 -8320 -10058 -8301
rect -9996 -8407 -9962 -8387
rect -9996 -8421 -9962 -8407
rect -9900 -8301 -9866 -8286
rect -9900 -8320 -9866 -8301
rect -9804 -8407 -9770 -8387
rect -9804 -8421 -9770 -8407
rect -9708 -8301 -9674 -8286
rect -9708 -8320 -9674 -8301
rect -9612 -8407 -9578 -8301
rect -9424 -8035 -9351 -7932
rect -9107 -8041 -8974 -7988
rect -8501 -8033 -8387 -7980
rect -8267 -7987 -8187 -7981
rect -8267 -8042 -8259 -7987
rect -8259 -8042 -8194 -7987
rect -8194 -8042 -8187 -7987
rect -8267 -8049 -8187 -8042
rect -8085 -8207 -8020 -8152
rect -9205 -8407 -9171 -8301
rect -9109 -8301 -9075 -8286
rect -9109 -8320 -9075 -8301
rect -9013 -8407 -8979 -8387
rect -9013 -8421 -8979 -8407
rect -8917 -8301 -8883 -8286
rect -8917 -8320 -8883 -8301
rect -8821 -8407 -8787 -8387
rect -8821 -8421 -8787 -8407
rect -8725 -8301 -8691 -8287
rect -8725 -8321 -8691 -8301
rect -8629 -8407 -8595 -8387
rect -8629 -8421 -8595 -8407
rect -8533 -8301 -8499 -8286
rect -8533 -8320 -8499 -8301
rect -8437 -8407 -8403 -8387
rect -8437 -8421 -8403 -8407
rect -8341 -8301 -8307 -8286
rect -8341 -8320 -8307 -8301
rect -8245 -8407 -8211 -8387
rect -8245 -8421 -8211 -8407
rect -8149 -8301 -8115 -8286
rect -8149 -8320 -8115 -8301
rect -8053 -8407 -8019 -8301
rect 7298 -7770 7332 -7419
rect 7332 -7770 7333 -7419
rect 7298 -7822 7333 -7770
rect 7298 -8170 7332 -7822
rect 7332 -8170 7333 -7822
rect 7372 -8182 7406 -7406
rect 7756 -8182 7790 -7406
rect 8246 -7770 8280 -7419
rect 8280 -7770 8281 -7419
rect 8246 -7822 8281 -7770
rect 8246 -8170 8280 -7822
rect 8280 -8170 8281 -7822
rect 8320 -8182 8354 -7406
rect 8704 -8182 8738 -7406
rect 9182 -7770 9216 -7419
rect 9216 -7770 9217 -7419
rect 9182 -7822 9217 -7770
rect 9182 -8170 9216 -7822
rect 9216 -8170 9217 -7822
rect 9256 -8182 9290 -7406
rect 9640 -8182 9674 -7406
rect 10113 -7769 10147 -7418
rect 10147 -7769 10148 -7418
rect 10113 -7821 10148 -7769
rect 10113 -8169 10147 -7821
rect 10147 -8169 10148 -7821
rect 10187 -8181 10221 -7405
rect 10571 -8181 10605 -7405
rect 11040 -7770 11074 -7419
rect 11074 -7770 11075 -7419
rect 11040 -7822 11075 -7770
rect 11040 -8170 11074 -7822
rect 11074 -8170 11075 -7822
rect 11114 -8182 11148 -7406
rect 12313 -7392 12347 -7358
rect 11498 -8182 11532 -7406
rect 12265 -7624 12299 -7448
rect 13052 -7385 13129 -7351
rect 12935 -7547 13111 -7513
rect 12842 -7591 12876 -7557
rect 12935 -7635 13111 -7601
rect 12183 -7768 12382 -7707
rect 12954 -7737 13086 -7703
rect -20603 -8541 -19480 -8495
rect -19044 -8541 -17921 -8495
rect -17312 -8541 -16189 -8495
rect -15753 -8541 -14630 -8495
rect -14021 -8541 -12898 -8495
rect -12462 -8541 -11339 -8495
rect -10730 -8541 -9607 -8495
rect -9171 -8541 -8048 -8495
rect 7198 -8554 7232 -8520
rect 7390 -8554 7424 -8520
rect 7582 -8554 7616 -8520
rect 7774 -8554 7808 -8520
rect 8146 -8554 8180 -8520
rect 8338 -8554 8372 -8520
rect 8530 -8554 8564 -8520
rect 8722 -8554 8756 -8520
rect 9082 -8554 9116 -8520
rect 9274 -8554 9308 -8520
rect 9466 -8554 9500 -8520
rect 9658 -8554 9692 -8520
rect 10013 -8553 10047 -8519
rect 10205 -8553 10239 -8519
rect 10397 -8553 10431 -8519
rect 10589 -8553 10623 -8519
rect 10940 -8554 10974 -8520
rect 11132 -8554 11166 -8520
rect 11324 -8554 11358 -8520
rect 11516 -8554 11550 -8520
rect -23520 -8650 -23429 -8616
rect -21783 -8650 -21692 -8616
rect -24368 -8716 -23799 -8669
rect -23577 -8722 -23571 -8688
rect -23571 -8722 -23498 -8688
rect -22632 -8716 -22063 -8669
rect -24384 -8794 -24350 -8788
rect -24384 -8868 -24350 -8794
rect -24288 -8984 -24254 -8910
rect -24288 -8990 -24254 -8984
rect -24192 -8794 -24158 -8788
rect -24192 -8868 -24158 -8794
rect -24096 -8984 -24062 -8910
rect -24096 -8990 -24062 -8984
rect -24000 -8794 -23966 -8788
rect -24000 -8868 -23966 -8794
rect -23904 -8984 -23870 -8910
rect -23904 -8990 -23870 -8984
rect -23808 -8794 -23774 -8788
rect -23808 -8868 -23774 -8794
rect -23664 -8962 -23630 -8736
rect -21840 -8722 -21834 -8688
rect -21834 -8722 -21761 -8688
rect -23454 -8818 -23377 -8784
rect -22648 -8794 -22614 -8788
rect -22648 -8868 -22614 -8794
rect -23577 -8914 -23571 -8880
rect -23571 -8914 -23498 -8880
rect -24318 -9078 -24284 -9043
rect -24029 -9078 -23995 -9043
rect -24234 -9202 -24200 -9167
rect -24150 -9172 -23774 -9138
rect -23454 -9010 -23377 -8976
rect -22552 -8984 -22518 -8910
rect -22552 -8990 -22518 -8984
rect -22456 -8794 -22422 -8788
rect -22456 -8868 -22422 -8794
rect -22360 -8984 -22326 -8910
rect -22360 -8990 -22326 -8984
rect -22264 -8794 -22230 -8788
rect -22264 -8868 -22230 -8794
rect -22168 -8984 -22134 -8910
rect -22168 -8990 -22134 -8984
rect -22072 -8794 -22038 -8788
rect -22072 -8868 -22038 -8794
rect -21927 -8962 -21893 -8736
rect -21717 -8818 -21640 -8784
rect 7245 -8613 7280 -8608
rect 7245 -8720 7246 -8613
rect 7246 -8720 7280 -8613
rect -21840 -8914 -21834 -8880
rect -21834 -8914 -21761 -8880
rect -20502 -8884 -19933 -8837
rect -19393 -8884 -18824 -8837
rect -18511 -8884 -17942 -8837
rect -17211 -8884 -16642 -8837
rect -16102 -8884 -15533 -8837
rect -15220 -8884 -14651 -8837
rect -13920 -8884 -13351 -8837
rect -12811 -8884 -12242 -8837
rect -11929 -8884 -11360 -8837
rect -10629 -8884 -10060 -8837
rect -9520 -8884 -8951 -8837
rect -8638 -8884 -8069 -8837
rect 7150 -8908 7184 -8798
rect 7342 -8908 7376 -8798
rect 7438 -8613 7473 -8608
rect 7438 -8720 7472 -8613
rect 7472 -8720 7473 -8613
rect 7534 -8908 7568 -8798
rect 7630 -8613 7665 -8608
rect 7630 -8720 7664 -8613
rect 7664 -8720 7665 -8613
rect 7726 -8908 7760 -8798
rect 7822 -8613 7857 -8608
rect 7822 -8720 7856 -8613
rect 7856 -8720 7857 -8613
rect 7918 -8908 7952 -8798
rect 8193 -8613 8228 -8608
rect 8193 -8720 8194 -8613
rect 8194 -8720 8228 -8613
rect 8098 -8908 8132 -8798
rect 8290 -8908 8324 -8798
rect 8386 -8613 8421 -8608
rect 8386 -8720 8420 -8613
rect 8420 -8720 8421 -8613
rect 8482 -8908 8516 -8798
rect 8578 -8613 8613 -8608
rect 8578 -8720 8612 -8613
rect 8612 -8720 8613 -8613
rect 8674 -8908 8708 -8798
rect 8770 -8613 8805 -8608
rect 8770 -8720 8804 -8613
rect 8804 -8720 8805 -8613
rect 8866 -8908 8900 -8798
rect 9129 -8613 9164 -8608
rect 9129 -8720 9130 -8613
rect 9130 -8720 9164 -8613
rect 9034 -8908 9068 -8798
rect 9226 -8908 9260 -8798
rect 9322 -8613 9357 -8608
rect 9322 -8720 9356 -8613
rect 9356 -8720 9357 -8613
rect 9418 -8908 9452 -8798
rect 9514 -8613 9549 -8608
rect 9514 -8720 9548 -8613
rect 9548 -8720 9549 -8613
rect 9610 -8908 9644 -8798
rect 9706 -8613 9741 -8608
rect 9706 -8720 9740 -8613
rect 9740 -8720 9741 -8613
rect 9802 -8908 9836 -8798
rect 10060 -8612 10095 -8607
rect 10060 -8719 10061 -8612
rect 10061 -8719 10095 -8612
rect 9965 -8907 9999 -8797
rect 10157 -8907 10191 -8797
rect 10253 -8612 10288 -8607
rect 10253 -8719 10287 -8612
rect 10287 -8719 10288 -8612
rect 10349 -8907 10383 -8797
rect 10445 -8612 10480 -8607
rect 10445 -8719 10479 -8612
rect 10479 -8719 10480 -8612
rect 10541 -8907 10575 -8797
rect 10637 -8612 10672 -8607
rect 10637 -8719 10671 -8612
rect 10671 -8719 10672 -8612
rect 10733 -8907 10767 -8797
rect 10987 -8613 11022 -8608
rect 10987 -8720 10988 -8613
rect 10988 -8720 11022 -8613
rect 10892 -8908 10926 -8798
rect 11084 -8908 11118 -8798
rect 11180 -8613 11215 -8608
rect 11180 -8720 11214 -8613
rect 11214 -8720 11215 -8613
rect 11276 -8908 11310 -8798
rect 11372 -8613 11407 -8608
rect 11372 -8720 11406 -8613
rect 11406 -8720 11407 -8613
rect 11468 -8908 11502 -8798
rect 11564 -8613 11599 -8608
rect 11564 -8720 11598 -8613
rect 11598 -8720 11599 -8613
rect 11660 -8908 11694 -8798
rect -22582 -9078 -22548 -9043
rect -22293 -9078 -22259 -9043
rect -23571 -9172 -23395 -9138
rect -23664 -9216 -23630 -9182
rect -23571 -9260 -23395 -9226
rect -22498 -9202 -22464 -9167
rect -22414 -9172 -22038 -9138
rect -20518 -8962 -20484 -8956
rect -21717 -9010 -21640 -8976
rect -20518 -9036 -20484 -8962
rect -21834 -9172 -21658 -9138
rect -20422 -9152 -20388 -9078
rect -20422 -9158 -20388 -9152
rect -20326 -8962 -20292 -8956
rect -20326 -9036 -20292 -8962
rect -20230 -9152 -20196 -9078
rect -20230 -9158 -20196 -9152
rect -20134 -8962 -20100 -8956
rect -20134 -9036 -20100 -8962
rect -20038 -9152 -20004 -9078
rect -20038 -9158 -20004 -9152
rect -19942 -8962 -19908 -8956
rect -19942 -9036 -19908 -8962
rect -19409 -8962 -19375 -8956
rect -19409 -9036 -19375 -8962
rect -19313 -9152 -19279 -9078
rect -19313 -9158 -19279 -9152
rect -19217 -8962 -19183 -8956
rect -19217 -9036 -19183 -8962
rect -19121 -9152 -19087 -9078
rect -19121 -9158 -19087 -9152
rect -19025 -8962 -18991 -8956
rect -19025 -9036 -18991 -8962
rect -18929 -9152 -18895 -9078
rect -18929 -9158 -18895 -9152
rect -18833 -8962 -18799 -8956
rect -18833 -9036 -18799 -8962
rect -18527 -8962 -18493 -8956
rect -18527 -9036 -18493 -8962
rect -18431 -9152 -18397 -9078
rect -18431 -9158 -18397 -9152
rect -18335 -8962 -18301 -8956
rect -18335 -9036 -18301 -8962
rect -18239 -9152 -18205 -9078
rect -18239 -9158 -18205 -9152
rect -18143 -8962 -18109 -8956
rect -18143 -9036 -18109 -8962
rect -18047 -9152 -18013 -9078
rect -18047 -9158 -18013 -9152
rect -17951 -8962 -17917 -8956
rect -17951 -9036 -17917 -8962
rect -17227 -8962 -17193 -8956
rect -17227 -9036 -17193 -8962
rect -17131 -9152 -17097 -9078
rect -17131 -9158 -17097 -9152
rect -17035 -8962 -17001 -8956
rect -17035 -9036 -17001 -8962
rect -16939 -9152 -16905 -9078
rect -16939 -9158 -16905 -9152
rect -16843 -8962 -16809 -8956
rect -16843 -9036 -16809 -8962
rect -16747 -9152 -16713 -9078
rect -16747 -9158 -16713 -9152
rect -16651 -8962 -16617 -8956
rect -16651 -9036 -16617 -8962
rect -16118 -8962 -16084 -8956
rect -16118 -9036 -16084 -8962
rect -16022 -9152 -15988 -9078
rect -16022 -9158 -15988 -9152
rect -15926 -8962 -15892 -8956
rect -15926 -9036 -15892 -8962
rect -15830 -9152 -15796 -9078
rect -15830 -9158 -15796 -9152
rect -15734 -8962 -15700 -8956
rect -15734 -9036 -15700 -8962
rect -15638 -9152 -15604 -9078
rect -15638 -9158 -15604 -9152
rect -15542 -8962 -15508 -8956
rect -15542 -9036 -15508 -8962
rect -15236 -8962 -15202 -8956
rect -15236 -9036 -15202 -8962
rect -15140 -9152 -15106 -9078
rect -15140 -9158 -15106 -9152
rect -15044 -8962 -15010 -8956
rect -15044 -9036 -15010 -8962
rect -14948 -9152 -14914 -9078
rect -14948 -9158 -14914 -9152
rect -14852 -8962 -14818 -8956
rect -14852 -9036 -14818 -8962
rect -14756 -9152 -14722 -9078
rect -14756 -9158 -14722 -9152
rect -14660 -8962 -14626 -8956
rect -14660 -9036 -14626 -8962
rect -13936 -8962 -13902 -8956
rect -13936 -9036 -13902 -8962
rect -13840 -9152 -13806 -9078
rect -13840 -9158 -13806 -9152
rect -13744 -8962 -13710 -8956
rect -13744 -9036 -13710 -8962
rect -13648 -9152 -13614 -9078
rect -13648 -9158 -13614 -9152
rect -13552 -8962 -13518 -8956
rect -13552 -9036 -13518 -8962
rect -13456 -9152 -13422 -9078
rect -13456 -9158 -13422 -9152
rect -13360 -8962 -13326 -8956
rect -13360 -9036 -13326 -8962
rect -12827 -8962 -12793 -8956
rect -12827 -9036 -12793 -8962
rect -12731 -9152 -12697 -9078
rect -12731 -9158 -12697 -9152
rect -12635 -8962 -12601 -8956
rect -12635 -9036 -12601 -8962
rect -12539 -9152 -12505 -9078
rect -12539 -9158 -12505 -9152
rect -12443 -8962 -12409 -8956
rect -12443 -9036 -12409 -8962
rect -12347 -9152 -12313 -9078
rect -12347 -9158 -12313 -9152
rect -12251 -8962 -12217 -8956
rect -12251 -9036 -12217 -8962
rect -11945 -8962 -11911 -8956
rect -11945 -9036 -11911 -8962
rect -11849 -9152 -11815 -9078
rect -11849 -9158 -11815 -9152
rect -11753 -8962 -11719 -8956
rect -11753 -9036 -11719 -8962
rect -11657 -9152 -11623 -9078
rect -11657 -9158 -11623 -9152
rect -11561 -8962 -11527 -8956
rect -11561 -9036 -11527 -8962
rect -11465 -9152 -11431 -9078
rect -11465 -9158 -11431 -9152
rect -11369 -8962 -11335 -8956
rect -11369 -9036 -11335 -8962
rect -10645 -8962 -10611 -8956
rect -10645 -9036 -10611 -8962
rect -10549 -9152 -10515 -9078
rect -10549 -9158 -10515 -9152
rect -10453 -8962 -10419 -8956
rect -10453 -9036 -10419 -8962
rect -10357 -9152 -10323 -9078
rect -10357 -9158 -10323 -9152
rect -10261 -8962 -10227 -8956
rect -10261 -9036 -10227 -8962
rect -10165 -9152 -10131 -9078
rect -10165 -9158 -10131 -9152
rect -10069 -8962 -10035 -8956
rect -10069 -9036 -10035 -8962
rect -9536 -8962 -9502 -8956
rect -9536 -9036 -9502 -8962
rect -9440 -9152 -9406 -9078
rect -9440 -9158 -9406 -9152
rect -9344 -8962 -9310 -8956
rect -9344 -9036 -9310 -8962
rect -9248 -9152 -9214 -9078
rect -9248 -9158 -9214 -9152
rect -9152 -8962 -9118 -8956
rect -9152 -9036 -9118 -8962
rect -9056 -9152 -9022 -9078
rect -9056 -9158 -9022 -9152
rect -8960 -8962 -8926 -8956
rect -8960 -9036 -8926 -8962
rect -8654 -8962 -8620 -8956
rect -8654 -9036 -8620 -8962
rect -8558 -9152 -8524 -9078
rect -8558 -9158 -8524 -9152
rect -8462 -8962 -8428 -8956
rect -8462 -9036 -8428 -8962
rect -8366 -9152 -8332 -9078
rect -8366 -9158 -8332 -9152
rect -8270 -8962 -8236 -8956
rect -8270 -9036 -8236 -8962
rect -8174 -9152 -8140 -9078
rect -8174 -9158 -8140 -9152
rect -8078 -8962 -8044 -8956
rect -8078 -9036 -8044 -8962
rect 7389 -9015 7677 -8980
rect 8337 -9015 8625 -8980
rect 9273 -9015 9561 -8980
rect 10204 -9014 10492 -8979
rect 11131 -9015 11419 -8980
rect -21927 -9216 -21893 -9182
rect -21834 -9260 -21658 -9226
rect -20452 -9246 -20418 -9211
rect -20163 -9246 -20129 -9211
rect -24150 -9364 -23774 -9330
rect -23552 -9362 -23420 -9328
rect -22414 -9364 -22038 -9330
rect -21815 -9362 -21683 -9328
rect -24135 -9436 -23800 -9402
rect -22399 -9436 -22064 -9402
rect -19343 -9246 -19309 -9211
rect -19054 -9246 -19020 -9211
rect -20368 -9370 -20334 -9335
rect -20284 -9340 -19908 -9306
rect -18461 -9246 -18427 -9211
rect -18172 -9246 -18138 -9211
rect -19259 -9370 -19225 -9335
rect -19175 -9340 -18799 -9306
rect -17161 -9246 -17127 -9211
rect -16872 -9246 -16838 -9211
rect -18377 -9370 -18343 -9335
rect -18293 -9340 -17917 -9306
rect -16052 -9246 -16018 -9211
rect -15763 -9246 -15729 -9211
rect -17077 -9370 -17043 -9335
rect -16993 -9340 -16617 -9306
rect -15170 -9246 -15136 -9211
rect -14881 -9246 -14847 -9211
rect -15968 -9370 -15934 -9335
rect -15884 -9340 -15508 -9306
rect -13870 -9246 -13836 -9211
rect -13581 -9246 -13547 -9211
rect -15086 -9370 -15052 -9335
rect -15002 -9340 -14626 -9306
rect -12761 -9246 -12727 -9211
rect -12472 -9246 -12438 -9211
rect -13786 -9370 -13752 -9335
rect -13702 -9340 -13326 -9306
rect -11879 -9246 -11845 -9211
rect -11590 -9246 -11556 -9211
rect -12677 -9370 -12643 -9335
rect -12593 -9340 -12217 -9306
rect -10579 -9246 -10545 -9211
rect -10290 -9246 -10256 -9211
rect -11795 -9370 -11761 -9335
rect -11711 -9340 -11335 -9306
rect -9470 -9246 -9436 -9211
rect -9181 -9246 -9147 -9211
rect -10495 -9370 -10461 -9335
rect -10411 -9340 -10035 -9306
rect -8588 -9246 -8554 -9211
rect -8299 -9246 -8265 -9211
rect -9386 -9370 -9352 -9335
rect -9302 -9340 -8926 -9306
rect -8504 -9370 -8470 -9335
rect -8420 -9340 -8044 -9306
rect -20284 -9532 -19908 -9498
rect -19175 -9532 -18799 -9498
rect -18293 -9532 -17917 -9498
rect -16993 -9532 -16617 -9498
rect -15884 -9532 -15508 -9498
rect -15002 -9532 -14626 -9498
rect -13702 -9532 -13326 -9498
rect -12593 -9532 -12217 -9498
rect -11711 -9532 -11335 -9498
rect -10411 -9532 -10035 -9498
rect -9302 -9532 -8926 -9498
rect -8420 -9532 -8044 -9498
rect -20269 -9604 -19934 -9570
rect -19160 -9604 -18825 -9570
rect -18278 -9604 -17943 -9570
rect -16978 -9604 -16643 -9570
rect -15869 -9604 -15534 -9570
rect -14987 -9604 -14652 -9570
rect -13687 -9604 -13352 -9570
rect -12578 -9604 -12243 -9570
rect -11696 -9604 -11361 -9570
rect -10396 -9604 -10061 -9570
rect -9287 -9604 -8952 -9570
rect -8405 -9604 -8070 -9570
rect 5721 -9635 5812 -9601
rect 6161 -9635 6252 -9601
rect 6601 -9635 6692 -9601
rect 5664 -9707 5670 -9673
rect 5670 -9707 5743 -9673
rect 5577 -9947 5611 -9721
rect 6104 -9707 6110 -9673
rect 6110 -9707 6183 -9673
rect 5787 -9803 5864 -9769
rect 5664 -9899 5670 -9865
rect 5670 -9899 5743 -9865
rect 6017 -9947 6051 -9721
rect 6544 -9707 6550 -9673
rect 6550 -9707 6623 -9673
rect 6227 -9803 6304 -9769
rect 6104 -9899 6110 -9865
rect 6110 -9899 6183 -9865
rect 5787 -9995 5864 -9961
rect 5670 -10157 5846 -10123
rect 5577 -10201 5611 -10167
rect 6457 -9947 6491 -9721
rect 6667 -9803 6744 -9769
rect 6544 -9899 6550 -9865
rect 6550 -9899 6623 -9865
rect 6227 -9995 6304 -9961
rect 6110 -10157 6286 -10123
rect 6017 -10201 6051 -10167
rect 5670 -10245 5846 -10211
rect 6667 -9995 6744 -9961
rect 6550 -10157 6726 -10123
rect 6457 -10201 6491 -10167
rect 6110 -10245 6286 -10211
rect 6550 -10245 6726 -10211
rect 7389 -10308 7677 -10273
rect 8337 -10308 8625 -10273
rect 9273 -10308 9561 -10273
rect 10204 -10308 10492 -10273
rect 11131 -10308 11419 -10273
rect -20603 -10428 -19481 -10356
rect -19044 -10428 -17922 -10356
rect -17312 -10428 -16190 -10356
rect -15753 -10428 -14631 -10356
rect -14021 -10428 -12899 -10356
rect -12462 -10428 -11340 -10356
rect -10730 -10428 -9608 -10356
rect 5689 -10347 5821 -10313
rect 6129 -10347 6261 -10313
rect 6569 -10347 6701 -10313
rect -9171 -10428 -8049 -10356
rect 7150 -10490 7184 -10380
rect -23520 -10622 -23429 -10588
rect -21787 -10622 -21696 -10588
rect -24368 -10688 -23799 -10641
rect -23577 -10694 -23571 -10660
rect -23571 -10694 -23498 -10660
rect -22631 -10688 -22062 -10641
rect -24384 -10766 -24350 -10760
rect -24384 -10840 -24350 -10766
rect -24288 -10956 -24254 -10882
rect -24288 -10962 -24254 -10956
rect -24192 -10766 -24158 -10760
rect -24192 -10840 -24158 -10766
rect -24096 -10956 -24062 -10882
rect -24096 -10962 -24062 -10956
rect -24000 -10766 -23966 -10760
rect -24000 -10840 -23966 -10766
rect -23904 -10956 -23870 -10882
rect -23904 -10962 -23870 -10956
rect -23808 -10766 -23774 -10760
rect -23808 -10840 -23774 -10766
rect -23664 -10934 -23630 -10708
rect -21844 -10694 -21838 -10660
rect -21838 -10694 -21765 -10660
rect -23454 -10790 -23377 -10756
rect -22647 -10766 -22613 -10760
rect -22647 -10840 -22613 -10766
rect -23577 -10886 -23571 -10852
rect -23571 -10886 -23498 -10852
rect -24318 -11050 -24284 -11015
rect -24029 -11050 -23995 -11015
rect -24234 -11174 -24200 -11139
rect -24150 -11144 -23774 -11110
rect -23454 -10982 -23377 -10948
rect -22551 -10956 -22517 -10882
rect -22551 -10962 -22517 -10956
rect -22455 -10766 -22421 -10760
rect -22455 -10840 -22421 -10766
rect -22359 -10956 -22325 -10882
rect -22359 -10962 -22325 -10956
rect -22263 -10766 -22229 -10760
rect -22263 -10840 -22229 -10766
rect -22167 -10956 -22133 -10882
rect -22167 -10962 -22133 -10956
rect -22071 -10766 -22037 -10760
rect -22071 -10840 -22037 -10766
rect -21931 -10934 -21897 -10708
rect -21721 -10790 -21644 -10756
rect -21844 -10886 -21838 -10852
rect -21838 -10886 -21765 -10852
rect -22581 -11050 -22547 -11015
rect -22292 -11050 -22258 -11015
rect -23571 -11144 -23395 -11110
rect -23664 -11188 -23630 -11154
rect -23571 -11232 -23395 -11198
rect -22497 -11174 -22463 -11139
rect -22413 -11144 -22037 -11110
rect -21721 -10982 -21644 -10948
rect -21838 -11144 -21662 -11110
rect -20637 -10633 -20603 -10531
rect -20637 -11028 -20603 -10926
rect -20541 -10841 -20507 -10717
rect -20445 -10633 -20411 -10531
rect -20445 -10992 -20411 -10926
rect -20349 -10841 -20315 -10717
rect -20253 -10635 -20219 -10533
rect -20253 -10992 -20219 -10932
rect -20157 -10841 -20123 -10717
rect -20061 -10636 -20027 -10534
rect -20061 -10992 -20027 -10949
rect -19965 -10841 -19931 -10717
rect -19869 -10636 -19835 -10534
rect -19869 -10992 -19835 -10932
rect -19773 -10841 -19739 -10717
rect -19677 -10636 -19643 -10534
rect -19677 -10992 -19643 -10925
rect -19581 -10842 -19547 -10718
rect -19485 -10636 -19451 -10534
rect -19485 -10992 -19451 -10925
rect -21931 -11188 -21897 -11154
rect -21838 -11232 -21662 -11198
rect -24150 -11336 -23774 -11302
rect -23552 -11334 -23420 -11300
rect -20854 -11261 -20807 -11151
rect -22413 -11336 -22037 -11302
rect -21819 -11334 -21687 -11300
rect -24135 -11408 -23800 -11374
rect -22398 -11408 -22063 -11374
rect -20539 -11305 -20406 -11252
rect -19078 -10633 -19044 -10531
rect -19078 -11028 -19044 -10926
rect -18982 -10841 -18948 -10717
rect -18886 -10633 -18852 -10531
rect -18886 -10992 -18852 -10926
rect -18790 -10841 -18756 -10717
rect -18694 -10635 -18660 -10533
rect -18694 -10992 -18660 -10932
rect -18598 -10841 -18564 -10717
rect -18502 -10636 -18468 -10534
rect -18502 -10992 -18468 -10949
rect -18406 -10841 -18372 -10717
rect -18310 -10636 -18276 -10534
rect -18310 -10992 -18276 -10932
rect -18214 -10841 -18180 -10717
rect -18118 -10636 -18084 -10534
rect -18118 -10992 -18084 -10925
rect -18022 -10842 -17988 -10718
rect -17926 -10636 -17892 -10534
rect -17926 -10992 -17892 -10925
rect -19933 -11297 -19819 -11244
rect -19699 -11251 -19619 -11245
rect -19699 -11306 -19691 -11251
rect -19691 -11306 -19626 -11251
rect -19626 -11306 -19619 -11251
rect -19699 -11313 -19619 -11306
rect -19517 -11471 -19452 -11416
rect -20637 -11671 -20603 -11565
rect -20541 -11565 -20507 -11550
rect -20541 -11584 -20507 -11565
rect -20445 -11671 -20411 -11651
rect -20445 -11685 -20411 -11671
rect -20349 -11565 -20315 -11550
rect -20349 -11584 -20315 -11565
rect -20253 -11671 -20219 -11651
rect -20253 -11685 -20219 -11671
rect -20157 -11565 -20123 -11551
rect -20157 -11585 -20123 -11565
rect -20061 -11671 -20027 -11651
rect -20061 -11685 -20027 -11671
rect -19965 -11565 -19931 -11550
rect -19965 -11584 -19931 -11565
rect -19869 -11671 -19835 -11651
rect -19869 -11685 -19835 -11671
rect -19773 -11565 -19739 -11550
rect -19773 -11584 -19739 -11565
rect -19677 -11671 -19643 -11651
rect -19677 -11685 -19643 -11671
rect -19581 -11565 -19547 -11550
rect -19581 -11584 -19547 -11565
rect -19485 -11671 -19451 -11565
rect -19297 -11299 -19224 -11196
rect -18980 -11305 -18847 -11252
rect -17346 -10633 -17312 -10531
rect -17346 -11028 -17312 -10926
rect -17250 -10841 -17216 -10717
rect -17154 -10633 -17120 -10531
rect -17154 -10992 -17120 -10926
rect -17058 -10841 -17024 -10717
rect -16962 -10635 -16928 -10533
rect -16962 -10992 -16928 -10932
rect -16866 -10841 -16832 -10717
rect -16770 -10636 -16736 -10534
rect -16770 -10992 -16736 -10949
rect -16674 -10841 -16640 -10717
rect -16578 -10636 -16544 -10534
rect -16578 -10992 -16544 -10932
rect -16482 -10841 -16448 -10717
rect -16386 -10636 -16352 -10534
rect -16386 -10992 -16352 -10925
rect -16290 -10842 -16256 -10718
rect -16194 -10636 -16160 -10534
rect -16194 -10992 -16160 -10925
rect -18374 -11297 -18260 -11244
rect -18140 -11251 -18060 -11245
rect -18140 -11306 -18132 -11251
rect -18132 -11306 -18067 -11251
rect -18067 -11306 -18060 -11251
rect -18140 -11313 -18060 -11306
rect -17958 -11471 -17893 -11416
rect -19078 -11671 -19044 -11565
rect -18982 -11565 -18948 -11550
rect -18982 -11584 -18948 -11565
rect -18886 -11671 -18852 -11651
rect -18886 -11685 -18852 -11671
rect -18790 -11565 -18756 -11550
rect -18790 -11584 -18756 -11565
rect -18694 -11671 -18660 -11651
rect -18694 -11685 -18660 -11671
rect -18598 -11565 -18564 -11551
rect -18598 -11585 -18564 -11565
rect -18502 -11671 -18468 -11651
rect -18502 -11685 -18468 -11671
rect -18406 -11565 -18372 -11550
rect -18406 -11584 -18372 -11565
rect -18310 -11671 -18276 -11651
rect -18310 -11685 -18276 -11671
rect -18214 -11565 -18180 -11550
rect -18214 -11584 -18180 -11565
rect -18118 -11671 -18084 -11651
rect -18118 -11685 -18084 -11671
rect -18022 -11565 -17988 -11550
rect -18022 -11584 -17988 -11565
rect -17926 -11671 -17892 -11565
rect -17563 -11261 -17516 -11151
rect -17248 -11305 -17115 -11252
rect -15787 -10633 -15753 -10531
rect -15787 -11028 -15753 -10926
rect -15691 -10841 -15657 -10717
rect -15595 -10633 -15561 -10531
rect -15595 -10992 -15561 -10926
rect -15499 -10841 -15465 -10717
rect -15403 -10635 -15369 -10533
rect -15403 -10992 -15369 -10932
rect -15307 -10841 -15273 -10717
rect -15211 -10636 -15177 -10534
rect -15211 -10992 -15177 -10949
rect -15115 -10841 -15081 -10717
rect -15019 -10636 -14985 -10534
rect -15019 -10992 -14985 -10932
rect -14923 -10841 -14889 -10717
rect -14827 -10636 -14793 -10534
rect -14827 -10992 -14793 -10925
rect -14731 -10842 -14697 -10718
rect -14635 -10636 -14601 -10534
rect -14635 -10992 -14601 -10925
rect -16642 -11297 -16528 -11244
rect -16408 -11251 -16328 -11245
rect -16408 -11306 -16400 -11251
rect -16400 -11306 -16335 -11251
rect -16335 -11306 -16328 -11251
rect -16408 -11313 -16328 -11306
rect -16226 -11471 -16161 -11416
rect -17346 -11671 -17312 -11565
rect -17250 -11565 -17216 -11550
rect -17250 -11584 -17216 -11565
rect -17154 -11671 -17120 -11651
rect -17154 -11685 -17120 -11671
rect -17058 -11565 -17024 -11550
rect -17058 -11584 -17024 -11565
rect -16962 -11671 -16928 -11651
rect -16962 -11685 -16928 -11671
rect -16866 -11565 -16832 -11551
rect -16866 -11585 -16832 -11565
rect -16770 -11671 -16736 -11651
rect -16770 -11685 -16736 -11671
rect -16674 -11565 -16640 -11550
rect -16674 -11584 -16640 -11565
rect -16578 -11671 -16544 -11651
rect -16578 -11685 -16544 -11671
rect -16482 -11565 -16448 -11550
rect -16482 -11584 -16448 -11565
rect -16386 -11671 -16352 -11651
rect -16386 -11685 -16352 -11671
rect -16290 -11565 -16256 -11550
rect -16290 -11584 -16256 -11565
rect -16194 -11671 -16160 -11565
rect -16006 -11299 -15933 -11196
rect -15689 -11305 -15556 -11252
rect -14055 -10633 -14021 -10531
rect -14055 -11028 -14021 -10926
rect -13959 -10841 -13925 -10717
rect -13863 -10633 -13829 -10531
rect -13863 -10992 -13829 -10926
rect -13767 -10841 -13733 -10717
rect -13671 -10635 -13637 -10533
rect -13671 -10992 -13637 -10932
rect -13575 -10841 -13541 -10717
rect -13479 -10636 -13445 -10534
rect -13479 -10992 -13445 -10949
rect -13383 -10841 -13349 -10717
rect -13287 -10636 -13253 -10534
rect -13287 -10992 -13253 -10932
rect -13191 -10841 -13157 -10717
rect -13095 -10636 -13061 -10534
rect -13095 -10992 -13061 -10925
rect -12999 -10842 -12965 -10718
rect -12903 -10636 -12869 -10534
rect -12903 -10992 -12869 -10925
rect -15083 -11297 -14969 -11244
rect -14849 -11251 -14769 -11245
rect -14849 -11306 -14841 -11251
rect -14841 -11306 -14776 -11251
rect -14776 -11306 -14769 -11251
rect -14849 -11313 -14769 -11306
rect -14667 -11471 -14602 -11416
rect -15787 -11671 -15753 -11565
rect -15691 -11565 -15657 -11550
rect -15691 -11584 -15657 -11565
rect -15595 -11671 -15561 -11651
rect -15595 -11685 -15561 -11671
rect -15499 -11565 -15465 -11550
rect -15499 -11584 -15465 -11565
rect -15403 -11671 -15369 -11651
rect -15403 -11685 -15369 -11671
rect -15307 -11565 -15273 -11551
rect -15307 -11585 -15273 -11565
rect -15211 -11671 -15177 -11651
rect -15211 -11685 -15177 -11671
rect -15115 -11565 -15081 -11550
rect -15115 -11584 -15081 -11565
rect -15019 -11671 -14985 -11651
rect -15019 -11685 -14985 -11671
rect -14923 -11565 -14889 -11550
rect -14923 -11584 -14889 -11565
rect -14827 -11671 -14793 -11651
rect -14827 -11685 -14793 -11671
rect -14731 -11565 -14697 -11550
rect -14731 -11584 -14697 -11565
rect -14635 -11671 -14601 -11565
rect -14272 -11261 -14225 -11151
rect -13957 -11305 -13824 -11252
rect -12496 -10633 -12462 -10531
rect -12496 -11028 -12462 -10926
rect -12400 -10841 -12366 -10717
rect -12304 -10633 -12270 -10531
rect -12304 -10992 -12270 -10926
rect -12208 -10841 -12174 -10717
rect -12112 -10635 -12078 -10533
rect -12112 -10992 -12078 -10932
rect -12016 -10841 -11982 -10717
rect -11920 -10636 -11886 -10534
rect -11920 -10992 -11886 -10949
rect -11824 -10841 -11790 -10717
rect -11728 -10636 -11694 -10534
rect -11728 -10992 -11694 -10932
rect -11632 -10841 -11598 -10717
rect -11536 -10636 -11502 -10534
rect -11536 -10992 -11502 -10925
rect -11440 -10842 -11406 -10718
rect -11344 -10636 -11310 -10534
rect -11344 -10992 -11310 -10925
rect -13351 -11297 -13237 -11244
rect -13117 -11251 -13037 -11245
rect -13117 -11306 -13109 -11251
rect -13109 -11306 -13044 -11251
rect -13044 -11306 -13037 -11251
rect -13117 -11313 -13037 -11306
rect -12935 -11471 -12870 -11416
rect -14055 -11671 -14021 -11565
rect -13959 -11565 -13925 -11550
rect -13959 -11584 -13925 -11565
rect -13863 -11671 -13829 -11651
rect -13863 -11685 -13829 -11671
rect -13767 -11565 -13733 -11550
rect -13767 -11584 -13733 -11565
rect -13671 -11671 -13637 -11651
rect -13671 -11685 -13637 -11671
rect -13575 -11565 -13541 -11551
rect -13575 -11585 -13541 -11565
rect -13479 -11671 -13445 -11651
rect -13479 -11685 -13445 -11671
rect -13383 -11565 -13349 -11550
rect -13383 -11584 -13349 -11565
rect -13287 -11671 -13253 -11651
rect -13287 -11685 -13253 -11671
rect -13191 -11565 -13157 -11550
rect -13191 -11584 -13157 -11565
rect -13095 -11671 -13061 -11651
rect -13095 -11685 -13061 -11671
rect -12999 -11565 -12965 -11550
rect -12999 -11584 -12965 -11565
rect -12903 -11671 -12869 -11565
rect -12715 -11299 -12642 -11196
rect -12398 -11305 -12265 -11252
rect -10764 -10633 -10730 -10531
rect -10764 -11028 -10730 -10926
rect -10668 -10841 -10634 -10717
rect -10572 -10633 -10538 -10531
rect -10572 -10992 -10538 -10926
rect -10476 -10841 -10442 -10717
rect -10380 -10635 -10346 -10533
rect -10380 -10992 -10346 -10932
rect -10284 -10841 -10250 -10717
rect -10188 -10636 -10154 -10534
rect -10188 -10992 -10154 -10949
rect -10092 -10841 -10058 -10717
rect -9996 -10636 -9962 -10534
rect -9996 -10992 -9962 -10932
rect -9900 -10841 -9866 -10717
rect -9804 -10636 -9770 -10534
rect -9804 -10992 -9770 -10925
rect -9708 -10842 -9674 -10718
rect -9612 -10636 -9578 -10534
rect -9612 -10992 -9578 -10925
rect -11792 -11297 -11678 -11244
rect -11558 -11251 -11478 -11245
rect -11558 -11306 -11550 -11251
rect -11550 -11306 -11485 -11251
rect -11485 -11306 -11478 -11251
rect -11558 -11313 -11478 -11306
rect -11376 -11471 -11311 -11416
rect -12496 -11671 -12462 -11565
rect -12400 -11565 -12366 -11550
rect -12400 -11584 -12366 -11565
rect -12304 -11671 -12270 -11651
rect -12304 -11685 -12270 -11671
rect -12208 -11565 -12174 -11550
rect -12208 -11584 -12174 -11565
rect -12112 -11671 -12078 -11651
rect -12112 -11685 -12078 -11671
rect -12016 -11565 -11982 -11551
rect -12016 -11585 -11982 -11565
rect -11920 -11671 -11886 -11651
rect -11920 -11685 -11886 -11671
rect -11824 -11565 -11790 -11550
rect -11824 -11584 -11790 -11565
rect -11728 -11671 -11694 -11651
rect -11728 -11685 -11694 -11671
rect -11632 -11565 -11598 -11550
rect -11632 -11584 -11598 -11565
rect -11536 -11671 -11502 -11651
rect -11536 -11685 -11502 -11671
rect -11440 -11565 -11406 -11550
rect -11440 -11584 -11406 -11565
rect -11344 -11671 -11310 -11565
rect -10981 -11261 -10934 -11151
rect -10666 -11305 -10533 -11252
rect -9205 -10633 -9171 -10531
rect -9205 -11028 -9171 -10926
rect -9109 -10841 -9075 -10717
rect -9013 -10633 -8979 -10531
rect -9013 -10992 -8979 -10926
rect -8917 -10841 -8883 -10717
rect -8821 -10635 -8787 -10533
rect -8821 -10992 -8787 -10932
rect -8725 -10841 -8691 -10717
rect -8629 -10636 -8595 -10534
rect -8629 -10992 -8595 -10949
rect -8533 -10841 -8499 -10717
rect -8437 -10636 -8403 -10534
rect -8437 -10992 -8403 -10932
rect -8341 -10841 -8307 -10717
rect -8245 -10636 -8211 -10534
rect -8245 -10992 -8211 -10925
rect -8149 -10842 -8115 -10718
rect -8053 -10636 -8019 -10534
rect -8053 -10992 -8019 -10925
rect 7245 -10675 7246 -10568
rect 7246 -10675 7280 -10568
rect 7245 -10680 7280 -10675
rect 7342 -10490 7376 -10380
rect 7534 -10490 7568 -10380
rect 7438 -10675 7472 -10568
rect 7472 -10675 7473 -10568
rect 7438 -10680 7473 -10675
rect 7726 -10490 7760 -10380
rect 7630 -10675 7664 -10568
rect 7664 -10675 7665 -10568
rect 7630 -10680 7665 -10675
rect 7918 -10490 7952 -10380
rect 7822 -10675 7856 -10568
rect 7856 -10675 7857 -10568
rect 7822 -10680 7857 -10675
rect 8098 -10490 8132 -10380
rect 8193 -10675 8194 -10568
rect 8194 -10675 8228 -10568
rect 8193 -10680 8228 -10675
rect 8290 -10490 8324 -10380
rect 8482 -10490 8516 -10380
rect 8386 -10675 8420 -10568
rect 8420 -10675 8421 -10568
rect 8386 -10680 8421 -10675
rect 8674 -10490 8708 -10380
rect 8578 -10675 8612 -10568
rect 8612 -10675 8613 -10568
rect 8578 -10680 8613 -10675
rect 8866 -10490 8900 -10380
rect 8770 -10675 8804 -10568
rect 8804 -10675 8805 -10568
rect 8770 -10680 8805 -10675
rect 9034 -10490 9068 -10380
rect 9129 -10675 9130 -10568
rect 9130 -10675 9164 -10568
rect 9129 -10680 9164 -10675
rect 9226 -10490 9260 -10380
rect 9418 -10490 9452 -10380
rect 9322 -10675 9356 -10568
rect 9356 -10675 9357 -10568
rect 9322 -10680 9357 -10675
rect 9610 -10490 9644 -10380
rect 9514 -10675 9548 -10568
rect 9548 -10675 9549 -10568
rect 9514 -10680 9549 -10675
rect 9802 -10490 9836 -10380
rect 9706 -10675 9740 -10568
rect 9740 -10675 9741 -10568
rect 9706 -10680 9741 -10675
rect 9965 -10490 9999 -10380
rect 10060 -10675 10061 -10568
rect 10061 -10675 10095 -10568
rect 10060 -10680 10095 -10675
rect 10157 -10490 10191 -10380
rect 10349 -10490 10383 -10380
rect 10253 -10675 10287 -10568
rect 10287 -10675 10288 -10568
rect 10253 -10680 10288 -10675
rect 10541 -10490 10575 -10380
rect 10445 -10675 10479 -10568
rect 10479 -10675 10480 -10568
rect 10445 -10680 10480 -10675
rect 10733 -10490 10767 -10380
rect 10637 -10675 10671 -10568
rect 10671 -10675 10672 -10568
rect 10637 -10680 10672 -10675
rect 10892 -10490 10926 -10380
rect 10987 -10675 10988 -10568
rect 10988 -10675 11022 -10568
rect 10987 -10680 11022 -10675
rect 11084 -10490 11118 -10380
rect 11276 -10490 11310 -10380
rect 11180 -10675 11214 -10568
rect 11214 -10675 11215 -10568
rect 11180 -10680 11215 -10675
rect 11468 -10490 11502 -10380
rect 11372 -10675 11406 -10568
rect 11406 -10675 11407 -10568
rect 11372 -10680 11407 -10675
rect 11660 -10490 11694 -10380
rect 11564 -10675 11598 -10568
rect 11598 -10675 11599 -10568
rect 11564 -10680 11599 -10675
rect 7198 -10768 7232 -10734
rect 7390 -10768 7424 -10734
rect 7582 -10768 7616 -10734
rect 7774 -10768 7808 -10734
rect 8146 -10768 8180 -10734
rect 8338 -10768 8372 -10734
rect 8530 -10768 8564 -10734
rect 8722 -10768 8756 -10734
rect 9082 -10768 9116 -10734
rect 9274 -10768 9308 -10734
rect 9466 -10768 9500 -10734
rect 9658 -10768 9692 -10734
rect 10013 -10768 10047 -10734
rect 10205 -10768 10239 -10734
rect 10397 -10768 10431 -10734
rect 10589 -10768 10623 -10734
rect 10940 -10768 10974 -10734
rect 11132 -10768 11166 -10734
rect 11324 -10768 11358 -10734
rect 11516 -10768 11550 -10734
rect -10060 -11297 -9946 -11244
rect -9826 -11251 -9746 -11245
rect -9826 -11306 -9818 -11251
rect -9818 -11306 -9753 -11251
rect -9753 -11306 -9746 -11251
rect -9826 -11313 -9746 -11306
rect -9644 -11471 -9579 -11416
rect -10764 -11671 -10730 -11565
rect -10668 -11565 -10634 -11550
rect -10668 -11584 -10634 -11565
rect -10572 -11671 -10538 -11651
rect -10572 -11685 -10538 -11671
rect -10476 -11565 -10442 -11550
rect -10476 -11584 -10442 -11565
rect -10380 -11671 -10346 -11651
rect -10380 -11685 -10346 -11671
rect -10284 -11565 -10250 -11551
rect -10284 -11585 -10250 -11565
rect -10188 -11671 -10154 -11651
rect -10188 -11685 -10154 -11671
rect -10092 -11565 -10058 -11550
rect -10092 -11584 -10058 -11565
rect -9996 -11671 -9962 -11651
rect -9996 -11685 -9962 -11671
rect -9900 -11565 -9866 -11550
rect -9900 -11584 -9866 -11565
rect -9804 -11671 -9770 -11651
rect -9804 -11685 -9770 -11671
rect -9708 -11565 -9674 -11550
rect -9708 -11584 -9674 -11565
rect -9612 -11671 -9578 -11565
rect -9424 -11299 -9351 -11196
rect -9107 -11305 -8974 -11252
rect -8501 -11297 -8387 -11244
rect -8267 -11251 -8187 -11245
rect -8267 -11306 -8259 -11251
rect -8259 -11306 -8194 -11251
rect -8194 -11306 -8187 -11251
rect -8267 -11313 -8187 -11306
rect -8085 -11471 -8020 -11416
rect -9205 -11671 -9171 -11565
rect -9109 -11565 -9075 -11550
rect -9109 -11584 -9075 -11565
rect -9013 -11671 -8979 -11651
rect -9013 -11685 -8979 -11671
rect -8917 -11565 -8883 -11550
rect -8917 -11584 -8883 -11565
rect -8821 -11671 -8787 -11651
rect -8821 -11685 -8787 -11671
rect -8725 -11565 -8691 -11551
rect -8725 -11585 -8691 -11565
rect -8629 -11671 -8595 -11651
rect -8629 -11685 -8595 -11671
rect -8533 -11565 -8499 -11550
rect -8533 -11584 -8499 -11565
rect -8437 -11671 -8403 -11651
rect -8437 -11685 -8403 -11671
rect -8341 -11565 -8307 -11550
rect -8341 -11584 -8307 -11565
rect -8245 -11671 -8211 -11651
rect -8245 -11685 -8211 -11671
rect -8149 -11565 -8115 -11550
rect -8149 -11584 -8115 -11565
rect -8053 -11671 -8019 -11565
rect 7298 -11466 7332 -11118
rect 7332 -11466 7333 -11118
rect 7298 -11518 7333 -11466
rect -20603 -11805 -19480 -11759
rect -19044 -11805 -17921 -11759
rect -17312 -11805 -16189 -11759
rect -15753 -11805 -14630 -11759
rect -14021 -11805 -12898 -11759
rect -12462 -11805 -11339 -11759
rect -10730 -11805 -9607 -11759
rect -9171 -11805 -8048 -11759
rect 7298 -11869 7332 -11518
rect 7332 -11869 7333 -11518
rect -23520 -11914 -23429 -11880
rect -21791 -11914 -21700 -11880
rect 7372 -11882 7406 -11106
rect 7756 -11882 7790 -11106
rect 8246 -11466 8280 -11118
rect 8280 -11466 8281 -11118
rect 8246 -11518 8281 -11466
rect 8246 -11869 8280 -11518
rect 8280 -11869 8281 -11518
rect 8320 -11882 8354 -11106
rect 8704 -11882 8738 -11106
rect 9182 -11466 9216 -11118
rect 9216 -11466 9217 -11118
rect 9182 -11518 9217 -11466
rect 9182 -11869 9216 -11518
rect 9216 -11869 9217 -11518
rect 9256 -11882 9290 -11106
rect 9640 -11882 9674 -11106
rect 10113 -11466 10147 -11118
rect 10147 -11466 10148 -11118
rect 10113 -11518 10148 -11466
rect 10113 -11869 10147 -11518
rect 10147 -11869 10148 -11518
rect 10187 -11882 10221 -11106
rect 10571 -11882 10605 -11106
rect 11040 -11466 11074 -11118
rect 11074 -11466 11075 -11118
rect 11040 -11518 11075 -11466
rect 11040 -11869 11074 -11518
rect 11074 -11869 11075 -11518
rect 11114 -11882 11148 -11106
rect 11498 -11882 11532 -11106
rect 11811 -11483 12168 -11432
rect 11785 -11819 11819 -11729
rect 11881 -11677 11915 -11587
rect 11977 -11819 12011 -11729
rect 12073 -11677 12107 -11587
rect 12169 -11819 12203 -11729
rect 12265 -11677 12299 -11587
rect 12361 -11819 12395 -11729
rect 12457 -11677 12491 -11587
rect 12553 -11819 12587 -11729
rect 12649 -11677 12683 -11587
rect 12986 -11653 13077 -11619
rect 12745 -11819 12779 -11729
rect 12929 -11725 12935 -11691
rect 12935 -11725 13008 -11691
rect 12170 -11915 12204 -11881
rect -24368 -11980 -23799 -11933
rect -23577 -11986 -23571 -11952
rect -23571 -11986 -23498 -11952
rect -22631 -11980 -22062 -11933
rect -24384 -12058 -24350 -12052
rect -24384 -12132 -24350 -12058
rect -24288 -12248 -24254 -12174
rect -24288 -12254 -24254 -12248
rect -24192 -12058 -24158 -12052
rect -24192 -12132 -24158 -12058
rect -24096 -12248 -24062 -12174
rect -24096 -12254 -24062 -12248
rect -24000 -12058 -23966 -12052
rect -24000 -12132 -23966 -12058
rect -23904 -12248 -23870 -12174
rect -23904 -12254 -23870 -12248
rect -23808 -12058 -23774 -12052
rect -23808 -12132 -23774 -12058
rect -23664 -12226 -23630 -12000
rect -21848 -11986 -21842 -11952
rect -21842 -11986 -21769 -11952
rect 12842 -11965 12876 -11739
rect 13052 -11821 13129 -11787
rect 12929 -11917 12935 -11883
rect 12935 -11917 13008 -11883
rect -23454 -12082 -23377 -12048
rect -22647 -12058 -22613 -12052
rect -22647 -12132 -22613 -12058
rect -23577 -12178 -23571 -12144
rect -23571 -12178 -23498 -12144
rect -24318 -12342 -24284 -12307
rect -24029 -12342 -23995 -12307
rect -24234 -12466 -24200 -12431
rect -24150 -12436 -23774 -12402
rect -23454 -12274 -23377 -12240
rect -22551 -12248 -22517 -12174
rect -22551 -12254 -22517 -12248
rect -22455 -12058 -22421 -12052
rect -22455 -12132 -22421 -12058
rect -22359 -12248 -22325 -12174
rect -22359 -12254 -22325 -12248
rect -22263 -12058 -22229 -12052
rect -22263 -12132 -22229 -12058
rect -22167 -12248 -22133 -12174
rect -22167 -12254 -22133 -12248
rect -22071 -12058 -22037 -12052
rect -22071 -12132 -22037 -12058
rect -21935 -12226 -21901 -12000
rect -21725 -12082 -21648 -12048
rect -21848 -12178 -21842 -12144
rect -21842 -12178 -21769 -12144
rect -20502 -12148 -19933 -12101
rect -19393 -12148 -18824 -12101
rect -18511 -12148 -17942 -12101
rect -17211 -12148 -16642 -12101
rect -16102 -12148 -15533 -12101
rect -15220 -12148 -14651 -12101
rect -13920 -12148 -13351 -12101
rect -12811 -12148 -12242 -12101
rect -11929 -12148 -11360 -12101
rect -10629 -12148 -10060 -12101
rect -9520 -12148 -8951 -12101
rect -8638 -12148 -8069 -12101
rect -22581 -12342 -22547 -12307
rect -22292 -12342 -22258 -12307
rect -23571 -12436 -23395 -12402
rect -23664 -12480 -23630 -12446
rect -23571 -12524 -23395 -12490
rect -22497 -12466 -22463 -12431
rect -22413 -12436 -22037 -12402
rect -20518 -12226 -20484 -12220
rect -21725 -12274 -21648 -12240
rect -20518 -12300 -20484 -12226
rect -21842 -12436 -21666 -12402
rect -20422 -12416 -20388 -12342
rect -20422 -12422 -20388 -12416
rect -20326 -12226 -20292 -12220
rect -20326 -12300 -20292 -12226
rect -20230 -12416 -20196 -12342
rect -20230 -12422 -20196 -12416
rect -20134 -12226 -20100 -12220
rect -20134 -12300 -20100 -12226
rect -20038 -12416 -20004 -12342
rect -20038 -12422 -20004 -12416
rect -19942 -12226 -19908 -12220
rect -19942 -12300 -19908 -12226
rect -19409 -12226 -19375 -12220
rect -19409 -12300 -19375 -12226
rect -19313 -12416 -19279 -12342
rect -19313 -12422 -19279 -12416
rect -19217 -12226 -19183 -12220
rect -19217 -12300 -19183 -12226
rect -19121 -12416 -19087 -12342
rect -19121 -12422 -19087 -12416
rect -19025 -12226 -18991 -12220
rect -19025 -12300 -18991 -12226
rect -18929 -12416 -18895 -12342
rect -18929 -12422 -18895 -12416
rect -18833 -12226 -18799 -12220
rect -18833 -12300 -18799 -12226
rect -18527 -12226 -18493 -12220
rect -18527 -12300 -18493 -12226
rect -18431 -12416 -18397 -12342
rect -18431 -12422 -18397 -12416
rect -18335 -12226 -18301 -12220
rect -18335 -12300 -18301 -12226
rect -18239 -12416 -18205 -12342
rect -18239 -12422 -18205 -12416
rect -18143 -12226 -18109 -12220
rect -18143 -12300 -18109 -12226
rect -18047 -12416 -18013 -12342
rect -18047 -12422 -18013 -12416
rect -17951 -12226 -17917 -12220
rect -17951 -12300 -17917 -12226
rect -17227 -12226 -17193 -12220
rect -17227 -12300 -17193 -12226
rect -17131 -12416 -17097 -12342
rect -17131 -12422 -17097 -12416
rect -17035 -12226 -17001 -12220
rect -17035 -12300 -17001 -12226
rect -16939 -12416 -16905 -12342
rect -16939 -12422 -16905 -12416
rect -16843 -12226 -16809 -12220
rect -16843 -12300 -16809 -12226
rect -16747 -12416 -16713 -12342
rect -16747 -12422 -16713 -12416
rect -16651 -12226 -16617 -12220
rect -16651 -12300 -16617 -12226
rect -16118 -12226 -16084 -12220
rect -16118 -12300 -16084 -12226
rect -16022 -12416 -15988 -12342
rect -16022 -12422 -15988 -12416
rect -15926 -12226 -15892 -12220
rect -15926 -12300 -15892 -12226
rect -15830 -12416 -15796 -12342
rect -15830 -12422 -15796 -12416
rect -15734 -12226 -15700 -12220
rect -15734 -12300 -15700 -12226
rect -15638 -12416 -15604 -12342
rect -15638 -12422 -15604 -12416
rect -15542 -12226 -15508 -12220
rect -15542 -12300 -15508 -12226
rect -15236 -12226 -15202 -12220
rect -15236 -12300 -15202 -12226
rect -15140 -12416 -15106 -12342
rect -15140 -12422 -15106 -12416
rect -15044 -12226 -15010 -12220
rect -15044 -12300 -15010 -12226
rect -14948 -12416 -14914 -12342
rect -14948 -12422 -14914 -12416
rect -14852 -12226 -14818 -12220
rect -14852 -12300 -14818 -12226
rect -14756 -12416 -14722 -12342
rect -14756 -12422 -14722 -12416
rect -14660 -12226 -14626 -12220
rect -14660 -12300 -14626 -12226
rect -13936 -12226 -13902 -12220
rect -13936 -12300 -13902 -12226
rect -13840 -12416 -13806 -12342
rect -13840 -12422 -13806 -12416
rect -13744 -12226 -13710 -12220
rect -13744 -12300 -13710 -12226
rect -13648 -12416 -13614 -12342
rect -13648 -12422 -13614 -12416
rect -13552 -12226 -13518 -12220
rect -13552 -12300 -13518 -12226
rect -13456 -12416 -13422 -12342
rect -13456 -12422 -13422 -12416
rect -13360 -12226 -13326 -12220
rect -13360 -12300 -13326 -12226
rect -12827 -12226 -12793 -12220
rect -12827 -12300 -12793 -12226
rect -12731 -12416 -12697 -12342
rect -12731 -12422 -12697 -12416
rect -12635 -12226 -12601 -12220
rect -12635 -12300 -12601 -12226
rect -12539 -12416 -12505 -12342
rect -12539 -12422 -12505 -12416
rect -12443 -12226 -12409 -12220
rect -12443 -12300 -12409 -12226
rect -12347 -12416 -12313 -12342
rect -12347 -12422 -12313 -12416
rect -12251 -12226 -12217 -12220
rect -12251 -12300 -12217 -12226
rect -11945 -12226 -11911 -12220
rect -11945 -12300 -11911 -12226
rect -11849 -12416 -11815 -12342
rect -11849 -12422 -11815 -12416
rect -11753 -12226 -11719 -12220
rect -11753 -12300 -11719 -12226
rect -11657 -12416 -11623 -12342
rect -11657 -12422 -11623 -12416
rect -11561 -12226 -11527 -12220
rect -11561 -12300 -11527 -12226
rect -11465 -12416 -11431 -12342
rect -11465 -12422 -11431 -12416
rect -11369 -12226 -11335 -12220
rect -11369 -12300 -11335 -12226
rect -10645 -12226 -10611 -12220
rect -10645 -12300 -10611 -12226
rect -10549 -12416 -10515 -12342
rect -10549 -12422 -10515 -12416
rect -10453 -12226 -10419 -12220
rect -10453 -12300 -10419 -12226
rect -10357 -12416 -10323 -12342
rect -10357 -12422 -10323 -12416
rect -10261 -12226 -10227 -12220
rect -10261 -12300 -10227 -12226
rect -10165 -12416 -10131 -12342
rect -10165 -12422 -10131 -12416
rect -10069 -12226 -10035 -12220
rect -10069 -12300 -10035 -12226
rect -9536 -12226 -9502 -12220
rect -9536 -12300 -9502 -12226
rect -9440 -12416 -9406 -12342
rect -9440 -12422 -9406 -12416
rect -9344 -12226 -9310 -12220
rect -9344 -12300 -9310 -12226
rect -9248 -12416 -9214 -12342
rect -9248 -12422 -9214 -12416
rect -9152 -12226 -9118 -12220
rect -9152 -12300 -9118 -12226
rect -9056 -12416 -9022 -12342
rect -9056 -12422 -9022 -12416
rect -8960 -12226 -8926 -12220
rect -8960 -12300 -8926 -12226
rect -8654 -12226 -8620 -12220
rect -8654 -12300 -8620 -12226
rect -8558 -12416 -8524 -12342
rect -8558 -12422 -8524 -12416
rect -8462 -12226 -8428 -12220
rect -8462 -12300 -8428 -12226
rect -8366 -12416 -8332 -12342
rect -8366 -12422 -8332 -12416
rect -8270 -12226 -8236 -12220
rect -8270 -12300 -8236 -12226
rect -8174 -12416 -8140 -12342
rect -8174 -12422 -8140 -12416
rect -8078 -12226 -8044 -12220
rect -8078 -12300 -8044 -12226
rect 7298 -12398 7332 -12047
rect 7332 -12398 7333 -12047
rect -21935 -12480 -21901 -12446
rect 7298 -12450 7333 -12398
rect -21842 -12524 -21666 -12490
rect -20452 -12510 -20418 -12475
rect -20163 -12510 -20129 -12475
rect -24150 -12628 -23774 -12594
rect -23552 -12626 -23420 -12592
rect -22413 -12628 -22037 -12594
rect -21823 -12626 -21691 -12592
rect -24135 -12700 -23800 -12666
rect -22398 -12700 -22063 -12666
rect -19343 -12510 -19309 -12475
rect -19054 -12510 -19020 -12475
rect -20368 -12634 -20334 -12599
rect -20284 -12604 -19908 -12570
rect -18461 -12510 -18427 -12475
rect -18172 -12510 -18138 -12475
rect -19259 -12634 -19225 -12599
rect -19175 -12604 -18799 -12570
rect -17161 -12510 -17127 -12475
rect -16872 -12510 -16838 -12475
rect -18377 -12634 -18343 -12599
rect -18293 -12604 -17917 -12570
rect -16052 -12510 -16018 -12475
rect -15763 -12510 -15729 -12475
rect -17077 -12634 -17043 -12599
rect -16993 -12604 -16617 -12570
rect -15170 -12510 -15136 -12475
rect -14881 -12510 -14847 -12475
rect -15968 -12634 -15934 -12599
rect -15884 -12604 -15508 -12570
rect -13870 -12510 -13836 -12475
rect -13581 -12510 -13547 -12475
rect -15086 -12634 -15052 -12599
rect -15002 -12604 -14626 -12570
rect -12761 -12510 -12727 -12475
rect -12472 -12510 -12438 -12475
rect -13786 -12634 -13752 -12599
rect -13702 -12604 -13326 -12570
rect -11879 -12510 -11845 -12475
rect -11590 -12510 -11556 -12475
rect -12677 -12634 -12643 -12599
rect -12593 -12604 -12217 -12570
rect -10579 -12510 -10545 -12475
rect -10290 -12510 -10256 -12475
rect -11795 -12634 -11761 -12599
rect -11711 -12604 -11335 -12570
rect -9470 -12510 -9436 -12475
rect -9181 -12510 -9147 -12475
rect -10495 -12634 -10461 -12599
rect -10411 -12604 -10035 -12570
rect -8588 -12510 -8554 -12475
rect -8299 -12510 -8265 -12475
rect -9386 -12634 -9352 -12599
rect -9302 -12604 -8926 -12570
rect -8504 -12634 -8470 -12599
rect -8420 -12604 -8044 -12570
rect -20284 -12796 -19908 -12762
rect -19175 -12796 -18799 -12762
rect -18293 -12796 -17917 -12762
rect -16993 -12796 -16617 -12762
rect -15884 -12796 -15508 -12762
rect -15002 -12796 -14626 -12762
rect -13702 -12796 -13326 -12762
rect -12593 -12796 -12217 -12762
rect -11711 -12796 -11335 -12762
rect -10411 -12796 -10035 -12762
rect -9302 -12796 -8926 -12762
rect -8420 -12796 -8044 -12762
rect 7298 -12798 7332 -12450
rect 7332 -12798 7333 -12450
rect 7372 -12810 7406 -12034
rect 7756 -12810 7790 -12034
rect 8246 -12398 8280 -12047
rect 8280 -12398 8281 -12047
rect 8246 -12450 8281 -12398
rect 8246 -12798 8280 -12450
rect 8280 -12798 8281 -12450
rect 8320 -12810 8354 -12034
rect 8704 -12810 8738 -12034
rect 9182 -12398 9216 -12047
rect 9216 -12398 9217 -12047
rect 9182 -12450 9217 -12398
rect 9182 -12798 9216 -12450
rect 9216 -12798 9217 -12450
rect 9256 -12810 9290 -12034
rect 9640 -12810 9674 -12034
rect 10113 -12397 10147 -12046
rect 10147 -12397 10148 -12046
rect 10113 -12449 10148 -12397
rect 10113 -12797 10147 -12449
rect 10147 -12797 10148 -12449
rect 10187 -12809 10221 -12033
rect 10571 -12809 10605 -12033
rect 11040 -12398 11074 -12047
rect 11074 -12398 11075 -12047
rect 11040 -12450 11075 -12398
rect 11040 -12798 11074 -12450
rect 11074 -12798 11075 -12450
rect 11114 -12810 11148 -12034
rect 12313 -12020 12347 -11986
rect 11498 -12810 11532 -12034
rect 12265 -12252 12299 -12076
rect 13052 -12013 13129 -11979
rect 12935 -12175 13111 -12141
rect 12842 -12219 12876 -12185
rect 12935 -12263 13111 -12229
rect 12183 -12396 12382 -12335
rect 12954 -12365 13086 -12331
rect -20269 -12868 -19934 -12834
rect -19160 -12868 -18825 -12834
rect -18278 -12868 -17943 -12834
rect -16978 -12868 -16643 -12834
rect -15869 -12868 -15534 -12834
rect -14987 -12868 -14652 -12834
rect -13687 -12868 -13352 -12834
rect -12578 -12868 -12243 -12834
rect -11696 -12868 -11361 -12834
rect -10396 -12868 -10061 -12834
rect -9287 -12868 -8952 -12834
rect -8405 -12868 -8070 -12834
rect 7198 -13182 7232 -13148
rect 7390 -13182 7424 -13148
rect 7582 -13182 7616 -13148
rect 7774 -13182 7808 -13148
rect 8146 -13182 8180 -13148
rect 8338 -13182 8372 -13148
rect 8530 -13182 8564 -13148
rect 8722 -13182 8756 -13148
rect 9082 -13182 9116 -13148
rect 9274 -13182 9308 -13148
rect 9466 -13182 9500 -13148
rect 9658 -13182 9692 -13148
rect 10013 -13181 10047 -13147
rect 10205 -13181 10239 -13147
rect 10397 -13181 10431 -13147
rect 10589 -13181 10623 -13147
rect 10940 -13182 10974 -13148
rect 11132 -13182 11166 -13148
rect 11324 -13182 11358 -13148
rect 11516 -13182 11550 -13148
rect 7245 -13241 7280 -13236
rect 7245 -13348 7246 -13241
rect 7246 -13348 7280 -13241
rect 7150 -13536 7184 -13426
rect 7342 -13536 7376 -13426
rect 7438 -13241 7473 -13236
rect 7438 -13348 7472 -13241
rect 7472 -13348 7473 -13241
rect 7534 -13536 7568 -13426
rect 7630 -13241 7665 -13236
rect 7630 -13348 7664 -13241
rect 7664 -13348 7665 -13241
rect 7726 -13536 7760 -13426
rect 7822 -13241 7857 -13236
rect 7822 -13348 7856 -13241
rect 7856 -13348 7857 -13241
rect 7918 -13536 7952 -13426
rect 8193 -13241 8228 -13236
rect 8193 -13348 8194 -13241
rect 8194 -13348 8228 -13241
rect 8098 -13536 8132 -13426
rect 8290 -13536 8324 -13426
rect 8386 -13241 8421 -13236
rect 8386 -13348 8420 -13241
rect 8420 -13348 8421 -13241
rect 8482 -13536 8516 -13426
rect 8578 -13241 8613 -13236
rect 8578 -13348 8612 -13241
rect 8612 -13348 8613 -13241
rect 8674 -13536 8708 -13426
rect 8770 -13241 8805 -13236
rect 8770 -13348 8804 -13241
rect 8804 -13348 8805 -13241
rect 8866 -13536 8900 -13426
rect 9129 -13241 9164 -13236
rect 9129 -13348 9130 -13241
rect 9130 -13348 9164 -13241
rect 9034 -13536 9068 -13426
rect 9226 -13536 9260 -13426
rect 9322 -13241 9357 -13236
rect 9322 -13348 9356 -13241
rect 9356 -13348 9357 -13241
rect 9418 -13536 9452 -13426
rect 9514 -13241 9549 -13236
rect 9514 -13348 9548 -13241
rect 9548 -13348 9549 -13241
rect 9610 -13536 9644 -13426
rect 9706 -13241 9741 -13236
rect 9706 -13348 9740 -13241
rect 9740 -13348 9741 -13241
rect 9802 -13536 9836 -13426
rect 10060 -13240 10095 -13235
rect 10060 -13347 10061 -13240
rect 10061 -13347 10095 -13240
rect 9965 -13535 9999 -13425
rect 10157 -13535 10191 -13425
rect 10253 -13240 10288 -13235
rect 10253 -13347 10287 -13240
rect 10287 -13347 10288 -13240
rect 10349 -13535 10383 -13425
rect 10445 -13240 10480 -13235
rect 10445 -13347 10479 -13240
rect 10479 -13347 10480 -13240
rect 10541 -13535 10575 -13425
rect 10637 -13240 10672 -13235
rect 10637 -13347 10671 -13240
rect 10671 -13347 10672 -13240
rect 10733 -13535 10767 -13425
rect 10987 -13241 11022 -13236
rect 10987 -13348 10988 -13241
rect 10988 -13348 11022 -13241
rect 10892 -13536 10926 -13426
rect 11084 -13536 11118 -13426
rect 11180 -13241 11215 -13236
rect 11180 -13348 11214 -13241
rect 11214 -13348 11215 -13241
rect 11276 -13536 11310 -13426
rect 11372 -13241 11407 -13236
rect 11372 -13348 11406 -13241
rect 11406 -13348 11407 -13241
rect 11468 -13536 11502 -13426
rect 11564 -13241 11599 -13236
rect 11564 -13348 11598 -13241
rect 11598 -13348 11599 -13241
rect 11660 -13536 11694 -13426
rect 7389 -13643 7677 -13608
rect 8337 -13643 8625 -13608
rect 9273 -13643 9561 -13608
rect 10204 -13642 10492 -13607
rect 11131 -13643 11419 -13608
rect -2172 -13969 -2138 -13878
rect -2100 -14020 -2066 -13947
rect -2100 -14026 -2066 -14020
rect -2004 -13903 -1970 -13826
rect -1908 -14020 -1874 -13947
rect -1908 -14026 -1874 -14020
rect -1812 -13903 -1778 -13826
rect -1650 -14020 -1616 -13844
rect -1562 -14020 -1528 -13844
rect -1460 -14001 -1426 -13869
rect -17523 -14545 -17433 -14511
rect -17665 -14641 -17575 -14607
rect -17523 -14737 -17433 -14703
rect -17665 -14833 -17575 -14799
rect -24562 -15522 -24515 -14953
rect -24443 -14962 -24437 -14928
rect -24437 -14962 -24363 -14928
rect -24321 -15058 -24247 -15024
rect -24247 -15058 -24241 -15024
rect -24443 -15154 -24437 -15120
rect -24437 -15154 -24363 -15120
rect -24188 -15183 -24153 -15149
rect -24321 -15250 -24247 -15216
rect -24247 -15250 -24241 -15216
rect -24443 -15346 -24437 -15312
rect -24437 -15346 -24363 -15312
rect -24093 -15304 -24059 -14928
rect -23901 -15304 -23867 -14928
rect -17523 -14929 -17433 -14895
rect -23829 -15289 -23795 -14954
rect -17266 -14977 -17232 -14943
rect -17665 -15025 -17575 -14991
rect -17176 -15025 -17000 -14991
rect -17523 -15121 -17433 -15087
rect -17371 -15120 -17337 -15086
rect -24064 -15388 -24029 -15354
rect -24321 -15442 -24247 -15408
rect -24247 -15442 -24241 -15408
rect -24188 -15472 -24153 -15438
rect -17820 -15479 -17769 -15122
rect -16917 -15107 -16856 -14908
rect -17665 -15217 -17575 -15183
rect -17523 -15313 -17433 -15279
rect -12473 -15345 -12401 -14223
rect -12295 -14227 -12193 -14193
rect -11904 -14227 -11837 -14193
rect -12111 -14323 -11987 -14289
rect -12295 -14419 -12193 -14385
rect -11904 -14419 -11837 -14385
rect -12112 -14515 -11988 -14481
rect -4768 -14156 -4542 -14122
rect -4322 -14156 -4288 -14122
rect -2052 -14113 -1826 -14079
rect -1606 -14113 -1572 -14079
rect 5721 -14163 5812 -14129
rect 6161 -14163 6252 -14129
rect 6601 -14163 6692 -14129
rect -11413 -14259 -11358 -14194
rect -11264 -14227 -11158 -14193
rect -11584 -14368 -11516 -14361
rect -11584 -14433 -11578 -14368
rect -11578 -14433 -11523 -14368
rect -11523 -14433 -11516 -14368
rect -11584 -14441 -11516 -14433
rect -12295 -14611 -12193 -14577
rect -11897 -14611 -11837 -14577
rect -12112 -14707 -11988 -14673
rect -11585 -14675 -11532 -14561
rect -11279 -14323 -11264 -14289
rect -11264 -14323 -11245 -14289
rect -11178 -14419 -11158 -14385
rect -11158 -14419 -11144 -14385
rect -11279 -14515 -11264 -14481
rect -11264 -14515 -11245 -14481
rect -11178 -14611 -11158 -14577
rect -11158 -14611 -11144 -14577
rect -11279 -14707 -11264 -14673
rect -11264 -14707 -11245 -14673
rect -12295 -14803 -12193 -14769
rect -11880 -14803 -11837 -14769
rect -11178 -14803 -11158 -14769
rect -11158 -14803 -11144 -14769
rect -12112 -14899 -11988 -14865
rect -12296 -14995 -12194 -14961
rect -11897 -14995 -11837 -14961
rect -11278 -14899 -11264 -14865
rect -11264 -14899 -11244 -14865
rect -11178 -14995 -11158 -14961
rect -11158 -14995 -11144 -14961
rect -12112 -15091 -11988 -15057
rect -12298 -15187 -12196 -15153
rect -11903 -15187 -11837 -15153
rect -12112 -15283 -11988 -15249
rect -17665 -15409 -17575 -15375
rect -12298 -15379 -12196 -15345
rect -11903 -15379 -11801 -15345
rect -11279 -15091 -11264 -15057
rect -11264 -15091 -11245 -15057
rect -11577 -15281 -11524 -15148
rect -11178 -15187 -11158 -15153
rect -11158 -15187 -11144 -15153
rect -11279 -15283 -11264 -15249
rect -11264 -15283 -11245 -15249
rect -11070 -15345 -11024 -14222
rect -4816 -14215 -4782 -14209
rect -4888 -14357 -4854 -14266
rect -4816 -14288 -4782 -14215
rect -4720 -14409 -4686 -14332
rect -4624 -14215 -4590 -14209
rect -4624 -14288 -4590 -14215
rect -4528 -14409 -4494 -14332
rect -4366 -14391 -4332 -14215
rect -4278 -14391 -4244 -14215
rect -4176 -14366 -4142 -14234
rect -2172 -14348 -2138 -14257
rect -2100 -14399 -2066 -14326
rect -2100 -14405 -2066 -14399
rect -2004 -14282 -1970 -14205
rect -1908 -14399 -1874 -14326
rect -1908 -14405 -1874 -14399
rect -1812 -14282 -1778 -14205
rect -1650 -14399 -1616 -14223
rect -1562 -14399 -1528 -14223
rect -1460 -14380 -1426 -14248
rect 5664 -14235 5670 -14201
rect 5670 -14235 5743 -14201
rect -2052 -14492 -1826 -14458
rect -1606 -14492 -1572 -14458
rect 5577 -14475 5611 -14249
rect 6104 -14235 6110 -14201
rect 6110 -14235 6183 -14201
rect 5787 -14331 5864 -14297
rect 5664 -14427 5670 -14393
rect 5670 -14427 5743 -14393
rect -4768 -14596 -4542 -14562
rect -4322 -14596 -4288 -14562
rect -4816 -14655 -4782 -14649
rect -4888 -14797 -4854 -14706
rect -4816 -14728 -4782 -14655
rect -4720 -14849 -4686 -14772
rect -4624 -14655 -4590 -14649
rect -4624 -14728 -4590 -14655
rect -4528 -14849 -4494 -14772
rect -4366 -14831 -4332 -14655
rect -4278 -14831 -4244 -14655
rect -4176 -14806 -4142 -14674
rect -2172 -14788 -2138 -14697
rect -2100 -14839 -2066 -14766
rect -2100 -14845 -2066 -14839
rect -2004 -14722 -1970 -14645
rect -1908 -14839 -1874 -14766
rect -1908 -14845 -1874 -14839
rect -1812 -14722 -1778 -14645
rect -1650 -14839 -1616 -14663
rect -1562 -14839 -1528 -14663
rect -1460 -14820 -1426 -14688
rect 6017 -14475 6051 -14249
rect 6544 -14235 6550 -14201
rect 6550 -14235 6623 -14201
rect 6227 -14331 6304 -14297
rect 6104 -14427 6110 -14393
rect 6110 -14427 6183 -14393
rect 5787 -14523 5864 -14489
rect 5670 -14685 5846 -14651
rect 5577 -14729 5611 -14695
rect 6457 -14475 6491 -14249
rect 6667 -14331 6744 -14297
rect 6544 -14427 6550 -14393
rect 6550 -14427 6623 -14393
rect 6227 -14523 6304 -14489
rect 6110 -14685 6286 -14651
rect 6017 -14729 6051 -14695
rect 5670 -14773 5846 -14739
rect 6667 -14523 6744 -14489
rect 6550 -14685 6726 -14651
rect 6457 -14729 6491 -14695
rect 6110 -14773 6286 -14739
rect 6550 -14773 6726 -14739
rect 7389 -14836 7677 -14801
rect 8337 -14836 8625 -14801
rect 9273 -14836 9561 -14801
rect 10204 -14836 10492 -14801
rect 11131 -14836 11419 -14801
rect 5689 -14875 5821 -14841
rect 6129 -14875 6261 -14841
rect 6569 -14875 6701 -14841
rect -4768 -14975 -4542 -14941
rect -4322 -14975 -4288 -14941
rect -2052 -14932 -1826 -14898
rect -1606 -14932 -1572 -14898
rect -4816 -15034 -4782 -15028
rect -4888 -15176 -4854 -15085
rect -4816 -15107 -4782 -15034
rect -4720 -15228 -4686 -15151
rect -4624 -15034 -4590 -15028
rect -4624 -15107 -4590 -15034
rect -4528 -15228 -4494 -15151
rect -4366 -15210 -4332 -15034
rect -4278 -15210 -4244 -15034
rect -4176 -15185 -4142 -15053
rect -2172 -15167 -2138 -15076
rect -2100 -15218 -2066 -15145
rect -2100 -15224 -2066 -15218
rect -2004 -15101 -1970 -15024
rect -1908 -15218 -1874 -15145
rect -1908 -15224 -1874 -15218
rect -1812 -15101 -1778 -15024
rect 7150 -15018 7184 -14908
rect -1650 -15218 -1616 -15042
rect -1562 -15218 -1528 -15042
rect -1460 -15199 -1426 -15067
rect 7245 -15203 7246 -15096
rect 7246 -15203 7280 -15096
rect 7245 -15208 7280 -15203
rect 7342 -15018 7376 -14908
rect 7534 -15018 7568 -14908
rect 7438 -15203 7472 -15096
rect 7472 -15203 7473 -15096
rect 7438 -15208 7473 -15203
rect 7726 -15018 7760 -14908
rect 7630 -15203 7664 -15096
rect 7664 -15203 7665 -15096
rect 7630 -15208 7665 -15203
rect 7918 -15018 7952 -14908
rect 7822 -15203 7856 -15096
rect 7856 -15203 7857 -15096
rect 7822 -15208 7857 -15203
rect 8098 -15018 8132 -14908
rect 8193 -15203 8194 -15096
rect 8194 -15203 8228 -15096
rect 8193 -15208 8228 -15203
rect 8290 -15018 8324 -14908
rect 8482 -15018 8516 -14908
rect 8386 -15203 8420 -15096
rect 8420 -15203 8421 -15096
rect 8386 -15208 8421 -15203
rect 8674 -15018 8708 -14908
rect 8578 -15203 8612 -15096
rect 8612 -15203 8613 -15096
rect 8578 -15208 8613 -15203
rect 8866 -15018 8900 -14908
rect 8770 -15203 8804 -15096
rect 8804 -15203 8805 -15096
rect 8770 -15208 8805 -15203
rect 9034 -15018 9068 -14908
rect 9129 -15203 9130 -15096
rect 9130 -15203 9164 -15096
rect 9129 -15208 9164 -15203
rect 9226 -15018 9260 -14908
rect 9418 -15018 9452 -14908
rect 9322 -15203 9356 -15096
rect 9356 -15203 9357 -15096
rect 9322 -15208 9357 -15203
rect 9610 -15018 9644 -14908
rect 9514 -15203 9548 -15096
rect 9548 -15203 9549 -15096
rect 9514 -15208 9549 -15203
rect 9802 -15018 9836 -14908
rect 9706 -15203 9740 -15096
rect 9740 -15203 9741 -15096
rect 9706 -15208 9741 -15203
rect 9965 -15018 9999 -14908
rect 10060 -15203 10061 -15096
rect 10061 -15203 10095 -15096
rect 10060 -15208 10095 -15203
rect 10157 -15018 10191 -14908
rect 10349 -15018 10383 -14908
rect 10253 -15203 10287 -15096
rect 10287 -15203 10288 -15096
rect 10253 -15208 10288 -15203
rect 10541 -15018 10575 -14908
rect 10445 -15203 10479 -15096
rect 10479 -15203 10480 -15096
rect 10445 -15208 10480 -15203
rect 10733 -15018 10767 -14908
rect 10637 -15203 10671 -15096
rect 10671 -15203 10672 -15096
rect 10637 -15208 10672 -15203
rect 10892 -15018 10926 -14908
rect 10987 -15203 10988 -15096
rect 10988 -15203 11022 -15096
rect 10987 -15208 11022 -15203
rect 11084 -15018 11118 -14908
rect 11276 -15018 11310 -14908
rect 11180 -15203 11214 -15096
rect 11214 -15203 11215 -15096
rect 11180 -15208 11215 -15203
rect 11468 -15018 11502 -14908
rect 11372 -15203 11406 -15096
rect 11406 -15203 11407 -15096
rect 11372 -15208 11407 -15203
rect 11660 -15018 11694 -14908
rect 11564 -15203 11598 -15096
rect 11598 -15203 11599 -15096
rect 11564 -15208 11599 -15203
rect -2052 -15311 -1826 -15277
rect -1606 -15311 -1572 -15277
rect 7198 -15296 7232 -15262
rect 7390 -15296 7424 -15262
rect 7582 -15296 7616 -15262
rect 7774 -15296 7808 -15262
rect 8146 -15296 8180 -15262
rect 8338 -15296 8372 -15262
rect 8530 -15296 8564 -15262
rect 8722 -15296 8756 -15262
rect 9082 -15296 9116 -15262
rect 9274 -15296 9308 -15262
rect 9466 -15296 9500 -15262
rect 9658 -15296 9692 -15262
rect 10013 -15296 10047 -15262
rect 10205 -15296 10239 -15262
rect 10397 -15296 10431 -15262
rect 10589 -15296 10623 -15262
rect 10940 -15296 10974 -15262
rect 11132 -15296 11166 -15262
rect 11324 -15296 11358 -15262
rect 11516 -15296 11550 -15262
rect -11264 -15379 -11158 -15345
rect -24443 -15538 -24437 -15504
rect -24437 -15538 -24363 -15504
rect -17523 -15505 -17433 -15471
rect -8239 -15497 -8205 -15406
rect -8167 -15548 -8133 -15475
rect -8167 -15554 -8133 -15548
rect -8071 -15431 -8037 -15354
rect -7975 -15548 -7941 -15475
rect -7975 -15554 -7941 -15548
rect -7879 -15431 -7845 -15354
rect -7717 -15548 -7683 -15372
rect -7629 -15548 -7595 -15372
rect -7527 -15529 -7493 -15397
rect -4768 -15415 -4542 -15381
rect -4322 -15415 -4288 -15381
rect -4816 -15474 -4782 -15468
rect -11567 -15604 -11493 -15594
rect -11567 -15658 -11557 -15604
rect -11557 -15658 -11503 -15604
rect -11503 -15658 -11493 -15604
rect -8119 -15641 -7893 -15607
rect -7673 -15641 -7639 -15607
rect -4888 -15616 -4854 -15525
rect -4816 -15547 -4782 -15474
rect -11567 -15668 -11493 -15658
rect -4720 -15668 -4686 -15591
rect -4624 -15474 -4590 -15468
rect -4624 -15547 -4590 -15474
rect -4528 -15668 -4494 -15591
rect -4366 -15650 -4332 -15474
rect -4278 -15650 -4244 -15474
rect -4176 -15625 -4142 -15493
rect -2172 -15607 -2138 -15516
rect -2100 -15658 -2066 -15585
rect -2100 -15664 -2066 -15658
rect -2004 -15541 -1970 -15464
rect -1908 -15658 -1874 -15585
rect -1908 -15664 -1874 -15658
rect -1812 -15541 -1778 -15464
rect -1650 -15658 -1616 -15482
rect -1562 -15658 -1528 -15482
rect -1460 -15639 -1426 -15507
rect -4768 -15794 -4542 -15760
rect -4322 -15794 -4288 -15760
rect -2052 -15751 -1826 -15717
rect -1606 -15751 -1572 -15717
rect -17523 -15945 -17433 -15911
rect -8238 -15997 -8204 -15906
rect -17665 -16041 -17575 -16007
rect -8166 -16048 -8132 -15975
rect -8166 -16054 -8132 -16048
rect -8070 -15931 -8036 -15854
rect -7974 -16048 -7940 -15975
rect -7974 -16054 -7940 -16048
rect -7878 -15931 -7844 -15854
rect -4816 -15853 -4782 -15847
rect -7716 -16048 -7682 -15872
rect -7628 -16048 -7594 -15872
rect -7526 -16029 -7492 -15897
rect -4888 -15995 -4854 -15904
rect -4816 -15926 -4782 -15853
rect -4720 -16047 -4686 -15970
rect -4624 -15853 -4590 -15847
rect -4624 -15926 -4590 -15853
rect -4528 -16047 -4494 -15970
rect -4366 -16029 -4332 -15853
rect -4278 -16029 -4244 -15853
rect -4176 -16004 -4142 -15872
rect -2172 -15986 -2138 -15895
rect -2100 -16037 -2066 -15964
rect -2100 -16043 -2066 -16037
rect -2004 -15920 -1970 -15843
rect -1908 -16037 -1874 -15964
rect -1908 -16043 -1874 -16037
rect -1812 -15920 -1778 -15843
rect -1650 -16037 -1616 -15861
rect -1562 -16037 -1528 -15861
rect -1460 -16018 -1426 -15886
rect 7298 -15994 7332 -15646
rect 7332 -15994 7333 -15646
rect 7298 -16046 7333 -15994
rect -24561 -16707 -24514 -16138
rect -24442 -16147 -24436 -16113
rect -24436 -16147 -24362 -16113
rect -24320 -16243 -24246 -16209
rect -24246 -16243 -24240 -16209
rect -24442 -16339 -24436 -16305
rect -24436 -16339 -24362 -16305
rect -24187 -16368 -24152 -16334
rect -24320 -16435 -24246 -16401
rect -24246 -16435 -24240 -16401
rect -24442 -16531 -24436 -16497
rect -24436 -16531 -24362 -16497
rect -24092 -16489 -24058 -16113
rect -23900 -16489 -23866 -16113
rect -17523 -16137 -17433 -16103
rect -23828 -16474 -23794 -16139
rect -8118 -16141 -7892 -16107
rect -7672 -16141 -7638 -16107
rect -2052 -16130 -1826 -16096
rect -1606 -16130 -1572 -16096
rect -17665 -16233 -17575 -16199
rect -4768 -16234 -4542 -16200
rect -4322 -16234 -4288 -16200
rect -17523 -16329 -17433 -16295
rect -17266 -16377 -17232 -16343
rect -17665 -16425 -17575 -16391
rect -17176 -16425 -17000 -16391
rect -17523 -16521 -17433 -16487
rect -17371 -16520 -17337 -16486
rect -24063 -16573 -24028 -16539
rect -24320 -16627 -24246 -16593
rect -24246 -16627 -24240 -16593
rect -24187 -16657 -24152 -16623
rect -24442 -16723 -24436 -16689
rect -24436 -16723 -24362 -16689
rect -17820 -16879 -17769 -16522
rect -16917 -16507 -16856 -16308
rect -4816 -16293 -4782 -16287
rect -8239 -16477 -8205 -16386
rect -8167 -16528 -8133 -16455
rect -8167 -16534 -8133 -16528
rect -8071 -16411 -8037 -16334
rect -7975 -16528 -7941 -16455
rect -7975 -16534 -7941 -16528
rect -7879 -16411 -7845 -16334
rect -7717 -16528 -7683 -16352
rect -7629 -16528 -7595 -16352
rect -7527 -16509 -7493 -16377
rect -4888 -16435 -4854 -16344
rect -4816 -16366 -4782 -16293
rect -4720 -16487 -4686 -16410
rect -4624 -16293 -4590 -16287
rect -4624 -16366 -4590 -16293
rect -4528 -16487 -4494 -16410
rect -4366 -16469 -4332 -16293
rect -4278 -16469 -4244 -16293
rect -4176 -16444 -4142 -16312
rect -2172 -16426 -2138 -16335
rect -2100 -16477 -2066 -16404
rect -2100 -16483 -2066 -16477
rect -2004 -16360 -1970 -16283
rect -1908 -16477 -1874 -16404
rect -1908 -16483 -1874 -16477
rect -1812 -16360 -1778 -16283
rect -1650 -16477 -1616 -16301
rect -1562 -16477 -1528 -16301
rect -1460 -16458 -1426 -16326
rect 7298 -16397 7332 -16046
rect 7332 -16397 7333 -16046
rect 7372 -16410 7406 -15634
rect 7756 -16410 7790 -15634
rect 8246 -15994 8280 -15646
rect 8280 -15994 8281 -15646
rect 8246 -16046 8281 -15994
rect 8246 -16397 8280 -16046
rect 8280 -16397 8281 -16046
rect 8320 -16410 8354 -15634
rect 8704 -16410 8738 -15634
rect 9182 -15994 9216 -15646
rect 9216 -15994 9217 -15646
rect 9182 -16046 9217 -15994
rect 9182 -16397 9216 -16046
rect 9216 -16397 9217 -16046
rect 9256 -16410 9290 -15634
rect 9640 -16410 9674 -15634
rect 10113 -15994 10147 -15646
rect 10147 -15994 10148 -15646
rect 10113 -16046 10148 -15994
rect 10113 -16397 10147 -16046
rect 10147 -16397 10148 -16046
rect 10187 -16410 10221 -15634
rect 10571 -16410 10605 -15634
rect 11040 -15994 11074 -15646
rect 11074 -15994 11075 -15646
rect 11040 -16046 11075 -15994
rect 11040 -16397 11074 -16046
rect 11074 -16397 11075 -16046
rect 11114 -16410 11148 -15634
rect 11498 -16410 11532 -15634
rect 11811 -16011 12168 -15960
rect 11785 -16347 11819 -16257
rect 11881 -16205 11915 -16115
rect 11977 -16347 12011 -16257
rect 12073 -16205 12107 -16115
rect 12169 -16347 12203 -16257
rect 12265 -16205 12299 -16115
rect 12361 -16347 12395 -16257
rect 12457 -16205 12491 -16115
rect 12553 -16347 12587 -16257
rect 12649 -16205 12683 -16115
rect 12986 -16181 13077 -16147
rect 12745 -16347 12779 -16257
rect 12929 -16253 12935 -16219
rect 12935 -16253 13008 -16219
rect 12170 -16443 12204 -16409
rect 12842 -16493 12876 -16267
rect 13052 -16349 13129 -16315
rect 12929 -16445 12935 -16411
rect 12935 -16445 13008 -16411
rect -17665 -16617 -17575 -16583
rect -8119 -16621 -7893 -16587
rect -7673 -16621 -7639 -16587
rect -4768 -16613 -4542 -16579
rect -4322 -16613 -4288 -16579
rect -2052 -16570 -1826 -16536
rect -1606 -16570 -1572 -16536
rect -4816 -16672 -4782 -16666
rect -17523 -16713 -17433 -16679
rect -17665 -16809 -17575 -16775
rect -4888 -16814 -4854 -16723
rect -17523 -16905 -17433 -16871
rect -24556 -17920 -24509 -17351
rect -24437 -17360 -24431 -17326
rect -24431 -17360 -24357 -17326
rect -24315 -17456 -24241 -17422
rect -24241 -17456 -24235 -17422
rect -24437 -17552 -24431 -17518
rect -24431 -17552 -24357 -17518
rect -24182 -17581 -24147 -17547
rect -24315 -17648 -24241 -17614
rect -24241 -17648 -24235 -17614
rect -24437 -17744 -24431 -17710
rect -24431 -17744 -24357 -17710
rect -24087 -17702 -24053 -17326
rect -23895 -17702 -23861 -17326
rect -17523 -17345 -17433 -17311
rect -23823 -17687 -23789 -17352
rect -17665 -17441 -17575 -17407
rect -17523 -17537 -17433 -17503
rect -17665 -17633 -17575 -17599
rect -17523 -17729 -17433 -17695
rect -24058 -17786 -24023 -17752
rect -24315 -17840 -24241 -17806
rect -24241 -17840 -24235 -17806
rect -24182 -17870 -24147 -17836
rect -17266 -17777 -17232 -17743
rect -17665 -17825 -17575 -17791
rect -17176 -17825 -17000 -17791
rect -24437 -17936 -24431 -17902
rect -24431 -17936 -24357 -17902
rect -17523 -17921 -17433 -17887
rect -17371 -17920 -17337 -17886
rect -21678 -18185 -21644 -18094
rect -21606 -18236 -21572 -18163
rect -21606 -18242 -21572 -18236
rect -21510 -18119 -21476 -18042
rect -21414 -18236 -21380 -18163
rect -21414 -18242 -21380 -18236
rect -21318 -18119 -21284 -18042
rect -21156 -18236 -21122 -18060
rect -21068 -18236 -21034 -18060
rect -20966 -18217 -20932 -18085
rect -17820 -18279 -17769 -17922
rect -16917 -17907 -16856 -17708
rect -17665 -18017 -17575 -17983
rect -16087 -18056 -16053 -17965
rect -17523 -18113 -17433 -18079
rect -16015 -18107 -15981 -18034
rect -16015 -18113 -15981 -18107
rect -15919 -17990 -15885 -17913
rect -15823 -18107 -15789 -18034
rect -15823 -18113 -15789 -18107
rect -15727 -17990 -15693 -17913
rect -15565 -18107 -15531 -17931
rect -15477 -18107 -15443 -17931
rect -15375 -18088 -15341 -17956
rect -12471 -18161 -12399 -17039
rect -12293 -17043 -12191 -17009
rect -11902 -17043 -11835 -17009
rect -12109 -17139 -11985 -17105
rect -12293 -17235 -12191 -17201
rect -11902 -17235 -11835 -17201
rect -12110 -17331 -11986 -17297
rect -8239 -16977 -8205 -16886
rect -11411 -17075 -11356 -17010
rect -11262 -17043 -11156 -17009
rect -11582 -17184 -11514 -17177
rect -11582 -17249 -11576 -17184
rect -11576 -17249 -11521 -17184
rect -11521 -17249 -11514 -17184
rect -11582 -17257 -11514 -17249
rect -12293 -17427 -12191 -17393
rect -11895 -17427 -11835 -17393
rect -12110 -17523 -11986 -17489
rect -11583 -17491 -11530 -17377
rect -11277 -17139 -11262 -17105
rect -11262 -17139 -11243 -17105
rect -11176 -17235 -11156 -17201
rect -11156 -17235 -11142 -17201
rect -11277 -17331 -11262 -17297
rect -11262 -17331 -11243 -17297
rect -11176 -17427 -11156 -17393
rect -11156 -17427 -11142 -17393
rect -11277 -17523 -11262 -17489
rect -11262 -17523 -11243 -17489
rect -12293 -17619 -12191 -17585
rect -11878 -17619 -11835 -17585
rect -11176 -17619 -11156 -17585
rect -11156 -17619 -11142 -17585
rect -12110 -17715 -11986 -17681
rect -12294 -17811 -12192 -17777
rect -11895 -17811 -11835 -17777
rect -11276 -17715 -11262 -17681
rect -11262 -17715 -11242 -17681
rect -11176 -17811 -11156 -17777
rect -11156 -17811 -11142 -17777
rect -12110 -17907 -11986 -17873
rect -12296 -18003 -12194 -17969
rect -11901 -18003 -11835 -17969
rect -12110 -18099 -11986 -18065
rect -17665 -18209 -17575 -18175
rect -15967 -18200 -15741 -18166
rect -15521 -18200 -15487 -18166
rect -12296 -18195 -12194 -18161
rect -11901 -18195 -11799 -18161
rect -11277 -17907 -11262 -17873
rect -11262 -17907 -11243 -17873
rect -11575 -18097 -11522 -17964
rect -11176 -18003 -11156 -17969
rect -11156 -18003 -11142 -17969
rect -11277 -18099 -11262 -18065
rect -11262 -18099 -11243 -18065
rect -11068 -18161 -11022 -17038
rect -8167 -17028 -8133 -16955
rect -8167 -17034 -8133 -17028
rect -8071 -16911 -8037 -16834
rect -7975 -17028 -7941 -16955
rect -7975 -17034 -7941 -17028
rect -4816 -16745 -4782 -16672
rect -7879 -16911 -7845 -16834
rect -7717 -17028 -7683 -16852
rect -7629 -17028 -7595 -16852
rect -7527 -17009 -7493 -16877
rect -4720 -16866 -4686 -16789
rect -4624 -16672 -4590 -16666
rect -4624 -16745 -4590 -16672
rect -4528 -16866 -4494 -16789
rect -4366 -16848 -4332 -16672
rect -4278 -16848 -4244 -16672
rect -4176 -16823 -4142 -16691
rect -2172 -16805 -2138 -16714
rect -2100 -16856 -2066 -16783
rect -2100 -16862 -2066 -16856
rect -2004 -16739 -1970 -16662
rect -1908 -16856 -1874 -16783
rect -1908 -16862 -1874 -16856
rect -1812 -16739 -1778 -16662
rect -1650 -16856 -1616 -16680
rect -1562 -16856 -1528 -16680
rect -1460 -16837 -1426 -16705
rect -2052 -16949 -1826 -16915
rect -1606 -16949 -1572 -16915
rect 7298 -16926 7332 -16575
rect 7332 -16926 7333 -16575
rect 7298 -16978 7333 -16926
rect -4768 -17053 -4542 -17019
rect -4322 -17053 -4288 -17019
rect -8119 -17121 -7893 -17087
rect -7673 -17121 -7639 -17087
rect -4816 -17112 -4782 -17106
rect -4888 -17254 -4854 -17163
rect -4816 -17185 -4782 -17112
rect -8239 -17457 -8205 -17366
rect -8167 -17508 -8133 -17435
rect -8167 -17514 -8133 -17508
rect -8071 -17391 -8037 -17314
rect -7975 -17508 -7941 -17435
rect -7975 -17514 -7941 -17508
rect -7879 -17391 -7845 -17314
rect -7717 -17508 -7683 -17332
rect -4720 -17306 -4686 -17229
rect -4624 -17112 -4590 -17106
rect -4624 -17185 -4590 -17112
rect -4528 -17306 -4494 -17229
rect -4366 -17288 -4332 -17112
rect -4278 -17288 -4244 -17112
rect -4176 -17263 -4142 -17131
rect -2172 -17245 -2138 -17154
rect -2100 -17296 -2066 -17223
rect -2100 -17302 -2066 -17296
rect -2004 -17179 -1970 -17102
rect -1908 -17296 -1874 -17223
rect -1908 -17302 -1874 -17296
rect -1812 -17179 -1778 -17102
rect -1650 -17296 -1616 -17120
rect -1562 -17296 -1528 -17120
rect -1460 -17277 -1426 -17145
rect -7629 -17508 -7595 -17332
rect 7298 -17326 7332 -16978
rect 7332 -17326 7333 -16978
rect 7372 -17338 7406 -16562
rect 7756 -17338 7790 -16562
rect 8246 -16926 8280 -16575
rect 8280 -16926 8281 -16575
rect 8246 -16978 8281 -16926
rect 8246 -17326 8280 -16978
rect 8280 -17326 8281 -16978
rect 8320 -17338 8354 -16562
rect 8704 -17338 8738 -16562
rect 9182 -16926 9216 -16575
rect 9216 -16926 9217 -16575
rect 9182 -16978 9217 -16926
rect 9182 -17326 9216 -16978
rect 9216 -17326 9217 -16978
rect 9256 -17338 9290 -16562
rect 9640 -17338 9674 -16562
rect 10113 -16925 10147 -16574
rect 10147 -16925 10148 -16574
rect 10113 -16977 10148 -16925
rect 10113 -17325 10147 -16977
rect 10147 -17325 10148 -16977
rect 10187 -17337 10221 -16561
rect 10571 -17337 10605 -16561
rect 11040 -16926 11074 -16575
rect 11074 -16926 11075 -16575
rect 11040 -16978 11075 -16926
rect 11040 -17326 11074 -16978
rect 11074 -17326 11075 -16978
rect 11114 -17338 11148 -16562
rect -7527 -17489 -7493 -17357
rect -4768 -17432 -4542 -17398
rect -4322 -17432 -4288 -17398
rect -2052 -17389 -1826 -17355
rect -1606 -17389 -1572 -17355
rect 12313 -16548 12347 -16514
rect 11498 -17338 11532 -16562
rect 12265 -16780 12299 -16604
rect 13052 -16541 13129 -16507
rect 12935 -16703 13111 -16669
rect 12842 -16747 12876 -16713
rect 12935 -16791 13111 -16757
rect 12183 -16924 12382 -16863
rect 12954 -16893 13086 -16859
rect 16211 -16927 16541 -16814
rect 16255 -17237 16289 -17061
rect 16447 -17237 16481 -17061
rect 16669 -17338 16703 -17304
rect -4816 -17491 -4782 -17485
rect -8119 -17601 -7893 -17567
rect -7673 -17601 -7639 -17567
rect -4888 -17633 -4854 -17542
rect -4816 -17564 -4782 -17491
rect -4720 -17685 -4686 -17608
rect -4624 -17491 -4590 -17485
rect -4624 -17564 -4590 -17491
rect -4528 -17685 -4494 -17608
rect -4366 -17667 -4332 -17491
rect -4278 -17667 -4244 -17491
rect -4176 -17642 -4142 -17510
rect -2172 -17624 -2138 -17533
rect -2100 -17675 -2066 -17602
rect -2100 -17681 -2066 -17675
rect -2004 -17558 -1970 -17481
rect -1908 -17675 -1874 -17602
rect -1908 -17681 -1874 -17675
rect -1812 -17558 -1778 -17481
rect -1650 -17675 -1616 -17499
rect -1562 -17675 -1528 -17499
rect -1460 -17656 -1426 -17524
rect 15997 -17620 16031 -17586
rect 16285 -17620 16319 -17586
rect 16417 -17620 16451 -17586
rect 7198 -17710 7232 -17676
rect 7390 -17710 7424 -17676
rect 7582 -17710 7616 -17676
rect 7774 -17710 7808 -17676
rect 8146 -17710 8180 -17676
rect 8338 -17710 8372 -17676
rect 8530 -17710 8564 -17676
rect 8722 -17710 8756 -17676
rect 9082 -17710 9116 -17676
rect 9274 -17710 9308 -17676
rect 9466 -17710 9500 -17676
rect 9658 -17710 9692 -17676
rect 10013 -17709 10047 -17675
rect 10205 -17709 10239 -17675
rect 10397 -17709 10431 -17675
rect 10589 -17709 10623 -17675
rect 10940 -17710 10974 -17676
rect 11132 -17710 11166 -17676
rect 11324 -17710 11358 -17676
rect 11516 -17710 11550 -17676
rect -8239 -17917 -8205 -17826
rect -8167 -17968 -8133 -17895
rect -8167 -17974 -8133 -17968
rect -8071 -17851 -8037 -17774
rect -7975 -17968 -7941 -17895
rect -7975 -17974 -7941 -17968
rect -7879 -17851 -7845 -17774
rect -2052 -17768 -1826 -17734
rect -1606 -17768 -1572 -17734
rect -7717 -17968 -7683 -17792
rect -7629 -17968 -7595 -17792
rect -7527 -17949 -7493 -17817
rect -4768 -17872 -4542 -17838
rect -4322 -17872 -4288 -17838
rect -4816 -17931 -4782 -17925
rect -8119 -18061 -7893 -18027
rect -7673 -18061 -7639 -18027
rect -4888 -18073 -4854 -17982
rect -4816 -18004 -4782 -17931
rect -4720 -18125 -4686 -18048
rect -4624 -17931 -4590 -17925
rect -4624 -18004 -4590 -17931
rect -4528 -18125 -4494 -18048
rect -4366 -18107 -4332 -17931
rect -4278 -18107 -4244 -17931
rect -4176 -18082 -4142 -17950
rect -2172 -18064 -2138 -17973
rect -2100 -18115 -2066 -18042
rect -2100 -18121 -2066 -18115
rect -2004 -17998 -1970 -17921
rect -1908 -18115 -1874 -18042
rect -1908 -18121 -1874 -18115
rect -1812 -17998 -1778 -17921
rect -1650 -18115 -1616 -17939
rect -1562 -18115 -1528 -17939
rect -1460 -18096 -1426 -17964
rect 7245 -17769 7280 -17764
rect 7245 -17876 7246 -17769
rect 7246 -17876 7280 -17769
rect 7150 -18064 7184 -17954
rect 7342 -18064 7376 -17954
rect 7438 -17769 7473 -17764
rect 7438 -17876 7472 -17769
rect 7472 -17876 7473 -17769
rect 7534 -18064 7568 -17954
rect 7630 -17769 7665 -17764
rect 7630 -17876 7664 -17769
rect 7664 -17876 7665 -17769
rect 7726 -18064 7760 -17954
rect 7822 -17769 7857 -17764
rect 7822 -17876 7856 -17769
rect 7856 -17876 7857 -17769
rect 7918 -18064 7952 -17954
rect 8193 -17769 8228 -17764
rect 8193 -17876 8194 -17769
rect 8194 -17876 8228 -17769
rect 8098 -18064 8132 -17954
rect 8290 -18064 8324 -17954
rect 8386 -17769 8421 -17764
rect 8386 -17876 8420 -17769
rect 8420 -17876 8421 -17769
rect 8482 -18064 8516 -17954
rect 8578 -17769 8613 -17764
rect 8578 -17876 8612 -17769
rect 8612 -17876 8613 -17769
rect 8674 -18064 8708 -17954
rect 8770 -17769 8805 -17764
rect 8770 -17876 8804 -17769
rect 8804 -17876 8805 -17769
rect 8866 -18064 8900 -17954
rect 9129 -17769 9164 -17764
rect 9129 -17876 9130 -17769
rect 9130 -17876 9164 -17769
rect 9034 -18064 9068 -17954
rect 9226 -18064 9260 -17954
rect 9322 -17769 9357 -17764
rect 9322 -17876 9356 -17769
rect 9356 -17876 9357 -17769
rect 9418 -18064 9452 -17954
rect 9514 -17769 9549 -17764
rect 9514 -17876 9548 -17769
rect 9548 -17876 9549 -17769
rect 9610 -18064 9644 -17954
rect 9706 -17769 9741 -17764
rect 9706 -17876 9740 -17769
rect 9740 -17876 9741 -17769
rect 9802 -18064 9836 -17954
rect 10060 -17768 10095 -17763
rect 10060 -17875 10061 -17768
rect 10061 -17875 10095 -17768
rect 9965 -18063 9999 -17953
rect 10157 -18063 10191 -17953
rect 10253 -17768 10288 -17763
rect 10253 -17875 10287 -17768
rect 10287 -17875 10288 -17768
rect 10349 -18063 10383 -17953
rect 10445 -17768 10480 -17763
rect 10445 -17875 10479 -17768
rect 10479 -17875 10480 -17768
rect 10541 -18063 10575 -17953
rect 10637 -17768 10672 -17763
rect 10637 -17875 10671 -17768
rect 10671 -17875 10672 -17768
rect 10733 -18063 10767 -17953
rect 10987 -17769 11022 -17764
rect 10987 -17876 10988 -17769
rect 10988 -17876 11022 -17769
rect 10892 -18064 10926 -17954
rect 11084 -18064 11118 -17954
rect 11180 -17769 11215 -17764
rect 11180 -17876 11214 -17769
rect 11214 -17876 11215 -17769
rect 11276 -18064 11310 -17954
rect 11372 -17769 11407 -17764
rect 11372 -17876 11406 -17769
rect 11406 -17876 11407 -17769
rect 11468 -18064 11502 -17954
rect 11564 -17769 11599 -17764
rect 11564 -17876 11598 -17769
rect 11598 -17876 11599 -17769
rect 11660 -18064 11694 -17954
rect 15703 -18033 15737 -17679
rect 15775 -18033 15809 -17679
rect -11262 -18195 -11156 -18161
rect 7389 -18171 7677 -18136
rect 8337 -18171 8625 -18136
rect 9273 -18171 9561 -18136
rect 10204 -18170 10492 -18135
rect 11131 -18171 11419 -18136
rect -21558 -18329 -21332 -18295
rect -21112 -18329 -21078 -18295
rect -17523 -18305 -17433 -18271
rect -8253 -18377 -8219 -18286
rect -24541 -19039 -24494 -18470
rect -24422 -18479 -24416 -18445
rect -24416 -18479 -24342 -18445
rect -24300 -18575 -24226 -18541
rect -24226 -18575 -24220 -18541
rect -24422 -18671 -24416 -18637
rect -24416 -18671 -24342 -18637
rect -24167 -18700 -24132 -18666
rect -24300 -18767 -24226 -18733
rect -24226 -18767 -24220 -18733
rect -24422 -18863 -24416 -18829
rect -24416 -18863 -24342 -18829
rect -24072 -18821 -24038 -18445
rect -23880 -18821 -23846 -18445
rect -23808 -18806 -23774 -18471
rect -21677 -18685 -21643 -18594
rect -21605 -18736 -21571 -18663
rect -21605 -18742 -21571 -18736
rect -21509 -18619 -21475 -18542
rect -21413 -18736 -21379 -18663
rect -21413 -18742 -21379 -18736
rect -21317 -18619 -21283 -18542
rect -21155 -18736 -21121 -18560
rect -21067 -18736 -21033 -18560
rect -16086 -18556 -16052 -18465
rect -20965 -18717 -20931 -18585
rect -16014 -18607 -15980 -18534
rect -16014 -18613 -15980 -18607
rect -15918 -18490 -15884 -18413
rect -15822 -18607 -15788 -18534
rect -15822 -18613 -15788 -18607
rect -11565 -18413 -11491 -18403
rect -15726 -18490 -15692 -18413
rect -15564 -18607 -15530 -18431
rect -15476 -18607 -15442 -18431
rect -15374 -18588 -15340 -18456
rect -11565 -18467 -11555 -18413
rect -11555 -18467 -11501 -18413
rect -11501 -18467 -11491 -18413
rect -8181 -18428 -8147 -18355
rect -8181 -18434 -8147 -18428
rect -8085 -18311 -8051 -18234
rect -7989 -18428 -7955 -18355
rect -7989 -18434 -7955 -18428
rect -7893 -18311 -7859 -18234
rect -7731 -18428 -7697 -18252
rect -4768 -18251 -4542 -18217
rect -4322 -18251 -4288 -18217
rect -2052 -18208 -1826 -18174
rect -1606 -18208 -1572 -18174
rect -7643 -18428 -7609 -18252
rect -7541 -18409 -7507 -18277
rect -4816 -18310 -4782 -18304
rect -4888 -18452 -4854 -18361
rect -11565 -18477 -11491 -18467
rect -4816 -18383 -4782 -18310
rect -8133 -18521 -7907 -18487
rect -7687 -18521 -7653 -18487
rect -4720 -18504 -4686 -18427
rect -4624 -18310 -4590 -18304
rect -4624 -18383 -4590 -18310
rect -4528 -18504 -4494 -18427
rect -4366 -18486 -4332 -18310
rect -4278 -18486 -4244 -18310
rect -4176 -18461 -4142 -18329
rect -2172 -18443 -2138 -18352
rect -2100 -18494 -2066 -18421
rect -2100 -18500 -2066 -18494
rect -2004 -18377 -1970 -18300
rect -1908 -18494 -1874 -18421
rect -1908 -18500 -1874 -18494
rect -1812 -18377 -1778 -18300
rect -1650 -18494 -1616 -18318
rect -1562 -18494 -1528 -18318
rect -1460 -18475 -1426 -18343
rect 15871 -18511 15905 -18155
rect 15967 -18033 16001 -17679
rect 16063 -18511 16097 -18155
rect 16159 -18033 16193 -17679
rect 16255 -18511 16289 -18155
rect 16351 -18033 16385 -17679
rect 16447 -18511 16481 -18155
rect 16543 -18033 16577 -17679
rect 16639 -18511 16673 -18155
rect 16735 -18033 16769 -17679
rect 16831 -18511 16865 -18155
rect 16927 -18033 16961 -17679
rect 17322 -18209 17891 -18162
rect 18159 -18221 18250 -18187
rect 17306 -18287 17340 -18281
rect 17306 -18361 17340 -18287
rect 17402 -18477 17436 -18403
rect 17402 -18483 17436 -18477
rect 17498 -18287 17532 -18281
rect 17498 -18361 17532 -18287
rect 17594 -18477 17628 -18403
rect 17594 -18483 17628 -18477
rect 17690 -18287 17724 -18281
rect 17690 -18361 17724 -18287
rect 17786 -18477 17820 -18403
rect 17786 -18483 17820 -18477
rect 17882 -18287 17916 -18281
rect 17882 -18361 17916 -18287
rect 18102 -18293 18108 -18259
rect 18108 -18293 18181 -18259
rect 18015 -18533 18049 -18307
rect 18225 -18389 18302 -18355
rect 18102 -18485 18108 -18451
rect 18108 -18485 18181 -18451
rect -2052 -18587 -1826 -18553
rect -1606 -18587 -1572 -18553
rect 17372 -18571 17406 -18536
rect 17661 -18571 17695 -18536
rect -15966 -18700 -15740 -18666
rect -15520 -18700 -15486 -18666
rect -4768 -18691 -4542 -18657
rect -4322 -18691 -4288 -18657
rect 5721 -18691 5812 -18657
rect 6161 -18691 6252 -18657
rect 6601 -18691 6692 -18657
rect -17523 -18745 -17433 -18711
rect -21557 -18829 -21331 -18795
rect -21111 -18829 -21077 -18795
rect -17665 -18841 -17575 -18807
rect -8251 -18857 -8217 -18766
rect -24043 -18905 -24008 -18871
rect -24300 -18959 -24226 -18925
rect -24226 -18959 -24220 -18925
rect -24167 -18989 -24132 -18955
rect -17523 -18937 -17433 -18903
rect -24422 -19055 -24416 -19021
rect -24416 -19055 -24342 -19021
rect -21678 -19165 -21644 -19074
rect -21606 -19216 -21572 -19143
rect -21606 -19222 -21572 -19216
rect -21510 -19099 -21476 -19022
rect -21414 -19216 -21380 -19143
rect -21414 -19222 -21380 -19216
rect -21318 -19099 -21284 -19022
rect -21156 -19216 -21122 -19040
rect -17665 -19033 -17575 -18999
rect -21068 -19216 -21034 -19040
rect -16087 -19036 -16053 -18945
rect -20966 -19197 -20932 -19065
rect -17523 -19129 -17433 -19095
rect -16015 -19087 -15981 -19014
rect -16015 -19093 -15981 -19087
rect -15919 -18970 -15885 -18893
rect -15823 -19087 -15789 -19014
rect -15823 -19093 -15789 -19087
rect -15727 -18970 -15693 -18893
rect -15565 -19087 -15531 -18911
rect -15477 -19087 -15443 -18911
rect -8179 -18908 -8145 -18835
rect -8179 -18914 -8145 -18908
rect -8083 -18791 -8049 -18714
rect -7987 -18908 -7953 -18835
rect -7987 -18914 -7953 -18908
rect -7891 -18791 -7857 -18714
rect -7729 -18908 -7695 -18732
rect -7641 -18908 -7607 -18732
rect -7539 -18889 -7505 -18757
rect -4816 -18750 -4782 -18744
rect -4888 -18892 -4854 -18801
rect -4816 -18823 -4782 -18750
rect -15375 -19068 -15341 -18936
rect -4720 -18944 -4686 -18867
rect -4624 -18750 -4590 -18744
rect -4624 -18823 -4590 -18750
rect -4528 -18944 -4494 -18867
rect -4366 -18926 -4332 -18750
rect -4278 -18926 -4244 -18750
rect -4176 -18901 -4142 -18769
rect -2172 -18883 -2138 -18792
rect -2100 -18934 -2066 -18861
rect -2100 -18940 -2066 -18934
rect -2004 -18817 -1970 -18740
rect -1908 -18934 -1874 -18861
rect -1908 -18940 -1874 -18934
rect -1812 -18817 -1778 -18740
rect -1650 -18934 -1616 -18758
rect -1562 -18934 -1528 -18758
rect -1460 -18915 -1426 -18783
rect 5664 -18763 5670 -18729
rect 5670 -18763 5743 -18729
rect -8131 -19001 -7905 -18967
rect -7685 -19001 -7651 -18967
rect -4768 -19070 -4542 -19036
rect -4322 -19070 -4288 -19036
rect -2052 -19027 -1826 -18993
rect -1606 -19027 -1572 -18993
rect 5577 -19003 5611 -18777
rect 6104 -18763 6110 -18729
rect 6110 -18763 6183 -18729
rect 5787 -18859 5864 -18825
rect 5664 -18955 5670 -18921
rect 5670 -18955 5743 -18921
rect -17266 -19177 -17232 -19143
rect -17665 -19225 -17575 -19191
rect -17176 -19225 -17000 -19191
rect -21558 -19309 -21332 -19275
rect -21112 -19309 -21078 -19275
rect -17523 -19321 -17433 -19287
rect -17371 -19320 -17337 -19286
rect -24539 -20233 -24492 -19664
rect -24420 -19673 -24414 -19639
rect -24414 -19673 -24340 -19639
rect -24298 -19769 -24224 -19735
rect -24224 -19769 -24218 -19735
rect -24420 -19865 -24414 -19831
rect -24414 -19865 -24340 -19831
rect -24165 -19894 -24130 -19860
rect -24298 -19961 -24224 -19927
rect -24224 -19961 -24218 -19927
rect -24420 -20057 -24414 -20023
rect -24414 -20057 -24340 -20023
rect -24070 -20015 -24036 -19639
rect -23878 -20015 -23844 -19639
rect -23806 -20000 -23772 -19665
rect -21678 -19665 -21644 -19574
rect -21606 -19716 -21572 -19643
rect -21606 -19722 -21572 -19716
rect -21510 -19599 -21476 -19522
rect -21414 -19716 -21380 -19643
rect -21414 -19722 -21380 -19716
rect -21318 -19599 -21284 -19522
rect -21156 -19716 -21122 -19540
rect -21068 -19716 -21034 -19540
rect -20966 -19697 -20932 -19565
rect -17820 -19679 -17769 -19322
rect -16917 -19307 -16856 -19108
rect -4816 -19129 -4782 -19123
rect -15967 -19180 -15741 -19146
rect -15521 -19180 -15487 -19146
rect -4888 -19271 -4854 -19180
rect -4816 -19202 -4782 -19129
rect -4720 -19323 -4686 -19246
rect -4624 -19129 -4590 -19123
rect -4624 -19202 -4590 -19129
rect -4528 -19323 -4494 -19246
rect -4366 -19305 -4332 -19129
rect -4278 -19305 -4244 -19129
rect -4176 -19280 -4142 -19148
rect -2172 -19262 -2138 -19171
rect -2100 -19313 -2066 -19240
rect -2100 -19319 -2066 -19313
rect -2004 -19196 -1970 -19119
rect -1908 -19313 -1874 -19240
rect -1908 -19319 -1874 -19313
rect -1812 -19196 -1778 -19119
rect -1650 -19313 -1616 -19137
rect -1562 -19313 -1528 -19137
rect -1460 -19294 -1426 -19162
rect 6017 -19003 6051 -18777
rect 6544 -18763 6550 -18729
rect 6550 -18763 6623 -18729
rect 6227 -18859 6304 -18825
rect 6104 -18955 6110 -18921
rect 6110 -18955 6183 -18921
rect 5787 -19051 5864 -19017
rect 5670 -19213 5846 -19179
rect 5577 -19257 5611 -19223
rect 6457 -19003 6491 -18777
rect 6667 -18859 6744 -18825
rect 6544 -18955 6550 -18921
rect 6550 -18955 6623 -18921
rect 6227 -19051 6304 -19017
rect 6110 -19213 6286 -19179
rect 6017 -19257 6051 -19223
rect 5670 -19301 5846 -19267
rect 6667 -19051 6744 -19017
rect 6550 -19213 6726 -19179
rect 6457 -19257 6491 -19223
rect 6110 -19301 6286 -19267
rect 6550 -19301 6726 -19267
rect 7389 -19364 7677 -19329
rect 8337 -19364 8625 -19329
rect 9273 -19364 9561 -19329
rect 10204 -19364 10492 -19329
rect 11131 -19364 11419 -19329
rect -17665 -19417 -17575 -19383
rect -17523 -19513 -17433 -19479
rect -16087 -19536 -16053 -19445
rect -17665 -19609 -17575 -19575
rect -16015 -19587 -15981 -19514
rect -16015 -19593 -15981 -19587
rect -15919 -19470 -15885 -19393
rect -15823 -19587 -15789 -19514
rect -15823 -19593 -15789 -19587
rect -15727 -19470 -15693 -19393
rect -15565 -19587 -15531 -19411
rect -15477 -19587 -15443 -19411
rect -2052 -19406 -1826 -19372
rect -1606 -19406 -1572 -19372
rect 5689 -19403 5821 -19369
rect 6129 -19403 6261 -19369
rect 6569 -19403 6701 -19369
rect -15375 -19568 -15341 -19436
rect -4768 -19510 -4542 -19476
rect -4322 -19510 -4288 -19476
rect -4816 -19569 -4782 -19563
rect -17523 -19705 -17433 -19671
rect -15967 -19680 -15741 -19646
rect -15521 -19680 -15487 -19646
rect -4888 -19711 -4854 -19620
rect -4816 -19642 -4782 -19569
rect -4720 -19763 -4686 -19686
rect -21558 -19809 -21332 -19775
rect -21112 -19809 -21078 -19775
rect -4624 -19569 -4590 -19563
rect -4624 -19642 -4590 -19569
rect -4528 -19763 -4494 -19686
rect -4366 -19745 -4332 -19569
rect -4278 -19745 -4244 -19569
rect -4176 -19720 -4142 -19588
rect -2172 -19702 -2138 -19611
rect -2100 -19753 -2066 -19680
rect -2100 -19759 -2066 -19753
rect -2004 -19636 -1970 -19559
rect -1908 -19753 -1874 -19680
rect -1908 -19759 -1874 -19753
rect -1812 -19636 -1778 -19559
rect 7150 -19546 7184 -19436
rect -1650 -19753 -1616 -19577
rect -1562 -19753 -1528 -19577
rect -1460 -19734 -1426 -19602
rect 7245 -19731 7246 -19624
rect 7246 -19731 7280 -19624
rect 7245 -19736 7280 -19731
rect 7342 -19546 7376 -19436
rect 7534 -19546 7568 -19436
rect 7438 -19731 7472 -19624
rect 7472 -19731 7473 -19624
rect 7438 -19736 7473 -19731
rect 7726 -19546 7760 -19436
rect 7630 -19731 7664 -19624
rect 7664 -19731 7665 -19624
rect 7630 -19736 7665 -19731
rect 7918 -19546 7952 -19436
rect 7822 -19731 7856 -19624
rect 7856 -19731 7857 -19624
rect 7822 -19736 7857 -19731
rect 8098 -19546 8132 -19436
rect 8193 -19731 8194 -19624
rect 8194 -19731 8228 -19624
rect 8193 -19736 8228 -19731
rect 8290 -19546 8324 -19436
rect 8482 -19546 8516 -19436
rect 8386 -19731 8420 -19624
rect 8420 -19731 8421 -19624
rect 8386 -19736 8421 -19731
rect 8674 -19546 8708 -19436
rect 8578 -19731 8612 -19624
rect 8612 -19731 8613 -19624
rect 8578 -19736 8613 -19731
rect 8866 -19546 8900 -19436
rect 8770 -19731 8804 -19624
rect 8804 -19731 8805 -19624
rect 8770 -19736 8805 -19731
rect 9034 -19546 9068 -19436
rect 9129 -19731 9130 -19624
rect 9130 -19731 9164 -19624
rect 9129 -19736 9164 -19731
rect 9226 -19546 9260 -19436
rect 9418 -19546 9452 -19436
rect 9322 -19731 9356 -19624
rect 9356 -19731 9357 -19624
rect 9322 -19736 9357 -19731
rect 9610 -19546 9644 -19436
rect 9514 -19731 9548 -19624
rect 9548 -19731 9549 -19624
rect 9514 -19736 9549 -19731
rect 9802 -19546 9836 -19436
rect 9706 -19731 9740 -19624
rect 9740 -19731 9741 -19624
rect 9706 -19736 9741 -19731
rect 9965 -19546 9999 -19436
rect 10060 -19731 10061 -19624
rect 10061 -19731 10095 -19624
rect 10060 -19736 10095 -19731
rect 10157 -19546 10191 -19436
rect 10349 -19546 10383 -19436
rect 10253 -19731 10287 -19624
rect 10287 -19731 10288 -19624
rect 10253 -19736 10288 -19731
rect 10541 -19546 10575 -19436
rect 10445 -19731 10479 -19624
rect 10479 -19731 10480 -19624
rect 10445 -19736 10480 -19731
rect 10733 -19546 10767 -19436
rect 10637 -19731 10671 -19624
rect 10671 -19731 10672 -19624
rect 10637 -19736 10672 -19731
rect 10892 -19546 10926 -19436
rect 10987 -19731 10988 -19624
rect 10988 -19731 11022 -19624
rect 10987 -19736 11022 -19731
rect 11084 -19546 11118 -19436
rect 11276 -19546 11310 -19436
rect 11180 -19731 11214 -19624
rect 11214 -19731 11215 -19624
rect 11180 -19736 11215 -19731
rect 11468 -19546 11502 -19436
rect 11372 -19731 11406 -19624
rect 11406 -19731 11407 -19624
rect 11372 -19736 11407 -19731
rect 11660 -19546 11694 -19436
rect 15703 -19493 15737 -19139
rect 15775 -19493 15809 -19139
rect 15871 -19017 15905 -18661
rect 15967 -19493 16001 -19139
rect 16063 -19017 16097 -18661
rect 16159 -19493 16193 -19139
rect 16255 -19017 16289 -18661
rect 16351 -19493 16385 -19139
rect 16447 -19017 16481 -18661
rect 16543 -19493 16577 -19139
rect 16639 -19017 16673 -18661
rect 16735 -19493 16769 -19139
rect 16831 -19017 16865 -18661
rect 17456 -18695 17490 -18660
rect 17540 -18665 17916 -18631
rect 18225 -18581 18302 -18547
rect 18108 -18743 18284 -18709
rect 18015 -18787 18049 -18753
rect 17540 -18857 17916 -18823
rect 18108 -18831 18284 -18797
rect 17555 -18929 17890 -18895
rect 18127 -18933 18259 -18899
rect 16927 -19493 16961 -19139
rect 11564 -19731 11598 -19624
rect 11598 -19731 11599 -19624
rect 11564 -19736 11599 -19731
rect 15997 -19586 16031 -19552
rect 16285 -19586 16319 -19552
rect 16417 -19586 16451 -19552
rect -24041 -20099 -24006 -20065
rect -24298 -20153 -24224 -20119
rect -24224 -20153 -24218 -20119
rect -24165 -20183 -24130 -20149
rect -21678 -20145 -21644 -20054
rect -21606 -20196 -21572 -20123
rect -21606 -20202 -21572 -20196
rect -21510 -20079 -21476 -20002
rect -21414 -20196 -21380 -20123
rect -21414 -20202 -21380 -20196
rect -21318 -20079 -21284 -20002
rect -21156 -20196 -21122 -20020
rect -21068 -20196 -21034 -20020
rect -16087 -20016 -16053 -19925
rect -20966 -20177 -20932 -20045
rect -16015 -20067 -15981 -19994
rect -16015 -20073 -15981 -20067
rect -15919 -19950 -15885 -19873
rect -15823 -20067 -15789 -19994
rect -15823 -20073 -15789 -20067
rect -15727 -19950 -15693 -19873
rect -15565 -20067 -15531 -19891
rect -15477 -20067 -15443 -19891
rect -4768 -19889 -4542 -19855
rect -4322 -19889 -4288 -19855
rect -2052 -19846 -1826 -19812
rect -1606 -19846 -1572 -19812
rect 7198 -19824 7232 -19790
rect 7390 -19824 7424 -19790
rect 7582 -19824 7616 -19790
rect 7774 -19824 7808 -19790
rect 8146 -19824 8180 -19790
rect 8338 -19824 8372 -19790
rect 8530 -19824 8564 -19790
rect 8722 -19824 8756 -19790
rect 9082 -19824 9116 -19790
rect 9274 -19824 9308 -19790
rect 9466 -19824 9500 -19790
rect 9658 -19824 9692 -19790
rect 10013 -19824 10047 -19790
rect 10205 -19824 10239 -19790
rect 10397 -19824 10431 -19790
rect 10589 -19824 10623 -19790
rect 10940 -19824 10974 -19790
rect 11132 -19824 11166 -19790
rect 11324 -19824 11358 -19790
rect 11516 -19824 11550 -19790
rect 16669 -19868 16703 -19834
rect -15375 -20048 -15341 -19916
rect -17523 -20145 -17433 -20111
rect -15967 -20160 -15741 -20126
rect -15521 -20160 -15487 -20126
rect -24420 -20249 -24414 -20215
rect -24414 -20249 -24340 -20215
rect -17665 -20241 -17575 -20207
rect -21558 -20289 -21332 -20255
rect -21112 -20289 -21078 -20255
rect -17523 -20337 -17433 -20303
rect -17665 -20433 -17575 -20399
rect -21678 -20605 -21644 -20514
rect -21606 -20656 -21572 -20583
rect -21606 -20662 -21572 -20656
rect -21510 -20539 -21476 -20462
rect -21414 -20656 -21380 -20583
rect -21414 -20662 -21380 -20656
rect -21318 -20539 -21284 -20462
rect -21156 -20656 -21122 -20480
rect -21068 -20656 -21034 -20480
rect -16087 -20476 -16053 -20385
rect -20966 -20637 -20932 -20505
rect -17523 -20529 -17433 -20495
rect -17266 -20577 -17232 -20543
rect -17665 -20625 -17575 -20591
rect -17176 -20625 -17000 -20591
rect -21558 -20749 -21332 -20715
rect -21112 -20749 -21078 -20715
rect -17523 -20721 -17433 -20687
rect -17371 -20720 -17337 -20686
rect -24508 -21433 -24461 -20864
rect -24389 -20873 -24383 -20839
rect -24383 -20873 -24309 -20839
rect -24267 -20969 -24193 -20935
rect -24193 -20969 -24187 -20935
rect -24389 -21065 -24383 -21031
rect -24383 -21065 -24309 -21031
rect -24134 -21094 -24099 -21060
rect -24267 -21161 -24193 -21127
rect -24193 -21161 -24187 -21127
rect -24389 -21257 -24383 -21223
rect -24383 -21257 -24309 -21223
rect -24039 -21215 -24005 -20839
rect -23847 -21215 -23813 -20839
rect -23775 -21200 -23741 -20865
rect -21692 -21065 -21658 -20974
rect -21620 -21116 -21586 -21043
rect -21620 -21122 -21586 -21116
rect -21524 -20999 -21490 -20922
rect -21428 -21116 -21394 -21043
rect -21428 -21122 -21394 -21116
rect -21332 -20999 -21298 -20922
rect -21170 -21116 -21136 -20940
rect -21082 -21116 -21048 -20940
rect -20980 -21097 -20946 -20965
rect -17820 -21079 -17769 -20722
rect -16917 -20707 -16856 -20508
rect -16015 -20527 -15981 -20454
rect -16015 -20533 -15981 -20527
rect -15919 -20410 -15885 -20333
rect -15823 -20527 -15789 -20454
rect -15823 -20533 -15789 -20527
rect -15727 -20410 -15693 -20333
rect -15565 -20527 -15531 -20351
rect -15477 -20527 -15443 -20351
rect -15375 -20508 -15341 -20376
rect -15967 -20620 -15741 -20586
rect -15521 -20620 -15487 -20586
rect -17665 -20817 -17575 -20783
rect -17523 -20913 -17433 -20879
rect -16101 -20936 -16067 -20845
rect -17665 -21009 -17575 -20975
rect -16029 -20987 -15995 -20914
rect -16029 -20993 -15995 -20987
rect -15933 -20870 -15899 -20793
rect -15837 -20987 -15803 -20914
rect -15837 -20993 -15803 -20987
rect -15741 -20870 -15707 -20793
rect -15579 -20987 -15545 -20811
rect -15491 -20987 -15457 -20811
rect -15389 -20968 -15355 -20836
rect -17523 -21105 -17433 -21071
rect -15981 -21080 -15755 -21046
rect -15535 -21080 -15501 -21046
rect -12471 -21118 -12399 -19996
rect -12293 -20000 -12191 -19966
rect -11902 -20000 -11835 -19966
rect -12109 -20096 -11985 -20062
rect -12293 -20192 -12191 -20158
rect -11902 -20192 -11835 -20158
rect -12110 -20288 -11986 -20254
rect -4816 -19948 -4782 -19942
rect -11411 -20032 -11356 -19967
rect -11262 -20000 -11156 -19966
rect -11582 -20141 -11514 -20134
rect -11582 -20206 -11576 -20141
rect -11576 -20206 -11521 -20141
rect -11521 -20206 -11514 -20141
rect -11582 -20214 -11514 -20206
rect -12293 -20384 -12191 -20350
rect -11895 -20384 -11835 -20350
rect -12110 -20480 -11986 -20446
rect -11583 -20448 -11530 -20334
rect -11277 -20096 -11262 -20062
rect -11262 -20096 -11243 -20062
rect -11176 -20192 -11156 -20158
rect -11156 -20192 -11142 -20158
rect -11277 -20288 -11262 -20254
rect -11262 -20288 -11243 -20254
rect -11176 -20384 -11156 -20350
rect -11156 -20384 -11142 -20350
rect -11277 -20480 -11262 -20446
rect -11262 -20480 -11243 -20446
rect -12293 -20576 -12191 -20542
rect -11878 -20576 -11835 -20542
rect -11176 -20576 -11156 -20542
rect -11156 -20576 -11142 -20542
rect -12110 -20672 -11986 -20638
rect -12294 -20768 -12192 -20734
rect -11895 -20768 -11835 -20734
rect -11276 -20672 -11262 -20638
rect -11262 -20672 -11242 -20638
rect -11176 -20768 -11156 -20734
rect -11156 -20768 -11142 -20734
rect -12110 -20864 -11986 -20830
rect -12296 -20960 -12194 -20926
rect -11901 -20960 -11835 -20926
rect -12110 -21056 -11986 -21022
rect -12296 -21152 -12194 -21118
rect -11901 -21152 -11799 -21118
rect -21572 -21209 -21346 -21175
rect -21126 -21209 -21092 -21175
rect -11277 -20864 -11262 -20830
rect -11262 -20864 -11243 -20830
rect -11575 -21054 -11522 -20921
rect -11176 -20960 -11156 -20926
rect -11156 -20960 -11142 -20926
rect -11277 -21056 -11262 -21022
rect -11262 -21056 -11243 -21022
rect -11068 -21118 -11022 -19995
rect -4888 -20090 -4854 -19999
rect -4816 -20021 -4782 -19948
rect -4720 -20142 -4686 -20065
rect -4624 -19948 -4590 -19942
rect -4624 -20021 -4590 -19948
rect -4528 -20142 -4494 -20065
rect -4366 -20124 -4332 -19948
rect -4278 -20124 -4244 -19948
rect -4176 -20099 -4142 -19967
rect -2172 -20081 -2138 -19990
rect -2100 -20132 -2066 -20059
rect -2100 -20138 -2066 -20132
rect -2004 -20015 -1970 -19938
rect -1908 -20132 -1874 -20059
rect -1908 -20138 -1874 -20132
rect -1812 -20015 -1778 -19938
rect -1650 -20132 -1616 -19956
rect -1562 -20132 -1528 -19956
rect -1460 -20113 -1426 -19981
rect -2052 -20225 -1826 -20191
rect -1606 -20225 -1572 -20191
rect -4768 -20329 -4542 -20295
rect -4322 -20329 -4288 -20295
rect -4816 -20388 -4782 -20382
rect -4888 -20530 -4854 -20439
rect -4816 -20461 -4782 -20388
rect -4720 -20582 -4686 -20505
rect -4624 -20388 -4590 -20382
rect -4624 -20461 -4590 -20388
rect -4528 -20582 -4494 -20505
rect -4366 -20564 -4332 -20388
rect -4278 -20564 -4244 -20388
rect -4176 -20539 -4142 -20407
rect -2172 -20521 -2138 -20430
rect -2100 -20572 -2066 -20499
rect -2100 -20578 -2066 -20572
rect -2004 -20455 -1970 -20378
rect -1908 -20572 -1874 -20499
rect -1908 -20578 -1874 -20572
rect -1812 -20455 -1778 -20378
rect -1650 -20572 -1616 -20396
rect -1562 -20572 -1528 -20396
rect -1460 -20553 -1426 -20421
rect 7298 -20522 7332 -20174
rect 7332 -20522 7333 -20174
rect 7298 -20574 7333 -20522
rect -4768 -20708 -4542 -20674
rect -4322 -20708 -4288 -20674
rect -2052 -20665 -1826 -20631
rect -1606 -20665 -1572 -20631
rect -4816 -20767 -4782 -20761
rect -4888 -20909 -4854 -20818
rect -4816 -20840 -4782 -20767
rect -4720 -20961 -4686 -20884
rect -4624 -20767 -4590 -20761
rect -4624 -20840 -4590 -20767
rect -4528 -20961 -4494 -20884
rect -4366 -20943 -4332 -20767
rect -4278 -20943 -4244 -20767
rect -4176 -20918 -4142 -20786
rect 7298 -20925 7332 -20574
rect 7332 -20925 7333 -20574
rect 7372 -20938 7406 -20162
rect 7756 -20938 7790 -20162
rect 8246 -20522 8280 -20174
rect 8280 -20522 8281 -20174
rect 8246 -20574 8281 -20522
rect 8246 -20925 8280 -20574
rect 8280 -20925 8281 -20574
rect 8320 -20938 8354 -20162
rect 8704 -20938 8738 -20162
rect 9182 -20522 9216 -20174
rect 9216 -20522 9217 -20174
rect 9182 -20574 9217 -20522
rect 9182 -20925 9216 -20574
rect 9216 -20925 9217 -20574
rect 9256 -20938 9290 -20162
rect 9640 -20938 9674 -20162
rect 10113 -20522 10147 -20174
rect 10147 -20522 10148 -20174
rect 10113 -20574 10148 -20522
rect 10113 -20925 10147 -20574
rect 10147 -20925 10148 -20574
rect 10187 -20938 10221 -20162
rect 10571 -20938 10605 -20162
rect 11040 -20522 11074 -20174
rect 11074 -20522 11075 -20174
rect 11040 -20574 11075 -20522
rect 11040 -20925 11074 -20574
rect 11074 -20925 11075 -20574
rect 11114 -20938 11148 -20162
rect 11498 -20938 11532 -20162
rect 16255 -20111 16289 -19935
rect 16447 -20111 16481 -19935
rect 16211 -20358 16541 -20245
rect 11811 -20539 12168 -20488
rect 11785 -20875 11819 -20785
rect 11881 -20733 11915 -20643
rect 11977 -20875 12011 -20785
rect 12073 -20733 12107 -20643
rect 12169 -20875 12203 -20785
rect 12265 -20733 12299 -20643
rect 12361 -20875 12395 -20785
rect 12457 -20733 12491 -20643
rect 12553 -20875 12587 -20785
rect 12649 -20733 12683 -20643
rect 12986 -20709 13077 -20675
rect 12745 -20875 12779 -20785
rect 12929 -20781 12935 -20747
rect 12935 -20781 13008 -20747
rect 12170 -20971 12204 -20937
rect 12842 -21021 12876 -20795
rect 13052 -20877 13129 -20843
rect 12929 -20973 12935 -20939
rect 12935 -20973 13008 -20939
rect -11262 -21152 -11156 -21118
rect -24010 -21299 -23975 -21265
rect -24267 -21353 -24193 -21319
rect -24193 -21353 -24187 -21319
rect -24134 -21383 -24099 -21349
rect -24389 -21449 -24383 -21415
rect -24383 -21449 -24309 -21415
rect -21690 -21545 -21656 -21454
rect -21618 -21596 -21584 -21523
rect -21618 -21602 -21584 -21596
rect -21522 -21479 -21488 -21402
rect -21426 -21596 -21392 -21523
rect -21426 -21602 -21392 -21596
rect -21330 -21479 -21296 -21402
rect -21168 -21596 -21134 -21420
rect -21080 -21596 -21046 -21420
rect -16099 -21416 -16065 -21325
rect -20978 -21577 -20944 -21445
rect -16027 -21467 -15993 -21394
rect -16027 -21473 -15993 -21467
rect -15931 -21350 -15897 -21273
rect -15835 -21467 -15801 -21394
rect -15835 -21473 -15801 -21467
rect -15739 -21350 -15705 -21273
rect -15577 -21467 -15543 -21291
rect -15489 -21467 -15455 -21291
rect -15387 -21448 -15353 -21316
rect -11559 -21389 -11497 -21379
rect -11559 -21431 -11549 -21389
rect -11549 -21431 -11507 -21389
rect -11507 -21431 -11497 -21389
rect -11559 -21441 -11497 -21431
rect 7298 -21454 7332 -21103
rect 7332 -21454 7333 -21103
rect 7298 -21506 7333 -21454
rect -17523 -21545 -17433 -21511
rect -15979 -21560 -15753 -21526
rect -15533 -21560 -15499 -21526
rect -17665 -21641 -17575 -21607
rect -21570 -21689 -21344 -21655
rect -21124 -21689 -21090 -21655
rect -17523 -21737 -17433 -21703
rect -17665 -21833 -17575 -21799
rect 7298 -21854 7332 -21506
rect 7332 -21854 7333 -21506
rect 7372 -21866 7406 -21090
rect 7756 -21866 7790 -21090
rect 8246 -21454 8280 -21103
rect 8280 -21454 8281 -21103
rect 8246 -21506 8281 -21454
rect 8246 -21854 8280 -21506
rect 8280 -21854 8281 -21506
rect 8320 -21866 8354 -21090
rect 8704 -21866 8738 -21090
rect 9182 -21454 9216 -21103
rect 9216 -21454 9217 -21103
rect 9182 -21506 9217 -21454
rect 9182 -21854 9216 -21506
rect 9216 -21854 9217 -21506
rect 9256 -21866 9290 -21090
rect 9640 -21866 9674 -21090
rect 10113 -21453 10147 -21102
rect 10147 -21453 10148 -21102
rect 10113 -21505 10148 -21453
rect 10113 -21853 10147 -21505
rect 10147 -21853 10148 -21505
rect 10187 -21865 10221 -21089
rect 10571 -21865 10605 -21089
rect 11040 -21454 11074 -21103
rect 11074 -21454 11075 -21103
rect 11040 -21506 11075 -21454
rect 11040 -21854 11074 -21506
rect 11074 -21854 11075 -21506
rect 11114 -21866 11148 -21090
rect 12313 -21076 12347 -21042
rect 11498 -21866 11532 -21090
rect 12265 -21308 12299 -21132
rect 13052 -21069 13129 -21035
rect 12935 -21231 13111 -21197
rect 12842 -21275 12876 -21241
rect 12935 -21319 13111 -21285
rect 12183 -21452 12382 -21391
rect 12954 -21421 13086 -21387
rect -17523 -21929 -17433 -21895
rect -17266 -21977 -17232 -21943
rect -17665 -22025 -17575 -21991
rect -17176 -22025 -17000 -21991
rect -17523 -22121 -17433 -22087
rect -17371 -22120 -17337 -22086
rect -24509 -22736 -24462 -22167
rect -24390 -22176 -24384 -22142
rect -24384 -22176 -24310 -22142
rect -24268 -22272 -24194 -22238
rect -24194 -22272 -24188 -22238
rect -24390 -22368 -24384 -22334
rect -24384 -22368 -24310 -22334
rect -24135 -22397 -24100 -22363
rect -24268 -22464 -24194 -22430
rect -24194 -22464 -24188 -22430
rect -24390 -22560 -24384 -22526
rect -24384 -22560 -24310 -22526
rect -24040 -22518 -24006 -22142
rect -23848 -22518 -23814 -22142
rect -23776 -22503 -23742 -22168
rect -17820 -22479 -17769 -22122
rect -16917 -22107 -16856 -21908
rect -17665 -22217 -17575 -22183
rect 7198 -22238 7232 -22204
rect 7390 -22238 7424 -22204
rect 7582 -22238 7616 -22204
rect 7774 -22238 7808 -22204
rect 8146 -22238 8180 -22204
rect 8338 -22238 8372 -22204
rect 8530 -22238 8564 -22204
rect 8722 -22238 8756 -22204
rect 9082 -22238 9116 -22204
rect 9274 -22238 9308 -22204
rect 9466 -22238 9500 -22204
rect 9658 -22238 9692 -22204
rect 10013 -22237 10047 -22203
rect 10205 -22237 10239 -22203
rect 10397 -22237 10431 -22203
rect 10589 -22237 10623 -22203
rect 10940 -22238 10974 -22204
rect 11132 -22238 11166 -22204
rect 11324 -22238 11358 -22204
rect 11516 -22238 11550 -22204
rect -17523 -22313 -17433 -22279
rect -17665 -22409 -17575 -22375
rect -17523 -22505 -17433 -22471
rect 7245 -22297 7280 -22292
rect 7245 -22404 7246 -22297
rect 7246 -22404 7280 -22297
rect -24011 -22602 -23976 -22568
rect -24268 -22656 -24194 -22622
rect -24194 -22656 -24188 -22622
rect -24135 -22686 -24100 -22652
rect -24390 -22752 -24384 -22718
rect -24384 -22752 -24310 -22718
rect -17523 -22945 -17433 -22911
rect -17665 -23041 -17575 -23007
rect -17523 -23137 -17433 -23103
rect -17665 -23233 -17575 -23199
rect -17523 -23329 -17433 -23295
rect -17266 -23377 -17232 -23343
rect -17665 -23425 -17575 -23391
rect -17176 -23425 -17000 -23391
rect -24509 -24045 -24462 -23476
rect -24390 -23485 -24384 -23451
rect -24384 -23485 -24310 -23451
rect -24268 -23581 -24194 -23547
rect -24194 -23581 -24188 -23547
rect -24390 -23677 -24384 -23643
rect -24384 -23677 -24310 -23643
rect -24135 -23706 -24100 -23672
rect -24268 -23773 -24194 -23739
rect -24194 -23773 -24188 -23739
rect -24390 -23869 -24384 -23835
rect -24384 -23869 -24310 -23835
rect -24040 -23827 -24006 -23451
rect -23848 -23827 -23814 -23451
rect -23776 -23812 -23742 -23477
rect -17523 -23521 -17433 -23487
rect -17371 -23520 -17337 -23486
rect -24011 -23911 -23976 -23877
rect -17820 -23879 -17769 -23522
rect -16917 -23507 -16856 -23308
rect -17665 -23617 -17575 -23583
rect -17523 -23713 -17433 -23679
rect -12471 -23697 -12399 -22575
rect -12293 -22579 -12191 -22545
rect -11902 -22579 -11835 -22545
rect -12109 -22675 -11985 -22641
rect -12293 -22771 -12191 -22737
rect -11902 -22771 -11835 -22737
rect -12110 -22867 -11986 -22833
rect -11411 -22611 -11356 -22546
rect -11262 -22579 -11156 -22545
rect -11582 -22720 -11514 -22713
rect -11582 -22785 -11576 -22720
rect -11576 -22785 -11521 -22720
rect -11521 -22785 -11514 -22720
rect -11582 -22793 -11514 -22785
rect -12293 -22963 -12191 -22929
rect -11895 -22963 -11835 -22929
rect -12110 -23059 -11986 -23025
rect -11583 -23027 -11530 -22913
rect -11277 -22675 -11262 -22641
rect -11262 -22675 -11243 -22641
rect -11176 -22771 -11156 -22737
rect -11156 -22771 -11142 -22737
rect -11277 -22867 -11262 -22833
rect -11262 -22867 -11243 -22833
rect -11176 -22963 -11156 -22929
rect -11156 -22963 -11142 -22929
rect -11277 -23059 -11262 -23025
rect -11262 -23059 -11243 -23025
rect -12293 -23155 -12191 -23121
rect -11878 -23155 -11835 -23121
rect -11176 -23155 -11156 -23121
rect -11156 -23155 -11142 -23121
rect -12110 -23251 -11986 -23217
rect -12294 -23347 -12192 -23313
rect -11895 -23347 -11835 -23313
rect -11276 -23251 -11262 -23217
rect -11262 -23251 -11242 -23217
rect -11176 -23347 -11156 -23313
rect -11156 -23347 -11142 -23313
rect -12110 -23443 -11986 -23409
rect -12296 -23539 -12194 -23505
rect -11901 -23539 -11835 -23505
rect -12110 -23635 -11986 -23601
rect -12296 -23731 -12194 -23697
rect -11901 -23731 -11799 -23697
rect -17665 -23809 -17575 -23775
rect -11277 -23443 -11262 -23409
rect -11262 -23443 -11243 -23409
rect -11575 -23633 -11522 -23500
rect -11176 -23539 -11156 -23505
rect -11156 -23539 -11142 -23505
rect -11277 -23635 -11262 -23601
rect -11262 -23635 -11243 -23601
rect -11068 -23697 -11022 -22574
rect 7150 -22592 7184 -22482
rect 7342 -22592 7376 -22482
rect 7438 -22297 7473 -22292
rect 7438 -22404 7472 -22297
rect 7472 -22404 7473 -22297
rect 7534 -22592 7568 -22482
rect 7630 -22297 7665 -22292
rect 7630 -22404 7664 -22297
rect 7664 -22404 7665 -22297
rect 7726 -22592 7760 -22482
rect 7822 -22297 7857 -22292
rect 7822 -22404 7856 -22297
rect 7856 -22404 7857 -22297
rect 7918 -22592 7952 -22482
rect 8193 -22297 8228 -22292
rect 8193 -22404 8194 -22297
rect 8194 -22404 8228 -22297
rect 8098 -22592 8132 -22482
rect 8290 -22592 8324 -22482
rect 8386 -22297 8421 -22292
rect 8386 -22404 8420 -22297
rect 8420 -22404 8421 -22297
rect 8482 -22592 8516 -22482
rect 8578 -22297 8613 -22292
rect 8578 -22404 8612 -22297
rect 8612 -22404 8613 -22297
rect 8674 -22592 8708 -22482
rect 8770 -22297 8805 -22292
rect 8770 -22404 8804 -22297
rect 8804 -22404 8805 -22297
rect 8866 -22592 8900 -22482
rect 9129 -22297 9164 -22292
rect 9129 -22404 9130 -22297
rect 9130 -22404 9164 -22297
rect 9034 -22592 9068 -22482
rect 9226 -22592 9260 -22482
rect 9322 -22297 9357 -22292
rect 9322 -22404 9356 -22297
rect 9356 -22404 9357 -22297
rect 9418 -22592 9452 -22482
rect 9514 -22297 9549 -22292
rect 9514 -22404 9548 -22297
rect 9548 -22404 9549 -22297
rect 9610 -22592 9644 -22482
rect 9706 -22297 9741 -22292
rect 9706 -22404 9740 -22297
rect 9740 -22404 9741 -22297
rect 9802 -22592 9836 -22482
rect 10060 -22296 10095 -22291
rect 10060 -22403 10061 -22296
rect 10061 -22403 10095 -22296
rect 9965 -22591 9999 -22481
rect 10157 -22591 10191 -22481
rect 10253 -22296 10288 -22291
rect 10253 -22403 10287 -22296
rect 10287 -22403 10288 -22296
rect 10349 -22591 10383 -22481
rect 10445 -22296 10480 -22291
rect 10445 -22403 10479 -22296
rect 10479 -22403 10480 -22296
rect 10541 -22591 10575 -22481
rect 10637 -22296 10672 -22291
rect 10637 -22403 10671 -22296
rect 10671 -22403 10672 -22296
rect 10733 -22591 10767 -22481
rect 10987 -22297 11022 -22292
rect 10987 -22404 10988 -22297
rect 10988 -22404 11022 -22297
rect 10892 -22592 10926 -22482
rect 11084 -22592 11118 -22482
rect 11180 -22297 11215 -22292
rect 11180 -22404 11214 -22297
rect 11214 -22404 11215 -22297
rect 11276 -22592 11310 -22482
rect 11372 -22297 11407 -22292
rect 11372 -22404 11406 -22297
rect 11406 -22404 11407 -22297
rect 11468 -22592 11502 -22482
rect 11564 -22297 11599 -22292
rect 11564 -22404 11598 -22297
rect 11598 -22404 11599 -22297
rect 11660 -22592 11694 -22482
rect 7389 -22699 7677 -22664
rect 8337 -22699 8625 -22664
rect 9273 -22699 9561 -22664
rect 10204 -22698 10492 -22663
rect 11131 -22699 11419 -22664
rect 5721 -23219 5812 -23185
rect 6161 -23219 6252 -23185
rect 6601 -23219 6692 -23185
rect -11262 -23731 -11156 -23697
rect 5664 -23291 5670 -23257
rect 5670 -23291 5743 -23257
rect 5577 -23531 5611 -23305
rect 6104 -23291 6110 -23257
rect 6110 -23291 6183 -23257
rect 5787 -23387 5864 -23353
rect 5664 -23483 5670 -23449
rect 5670 -23483 5743 -23449
rect 6017 -23531 6051 -23305
rect 6544 -23291 6550 -23257
rect 6550 -23291 6623 -23257
rect 6227 -23387 6304 -23353
rect 6104 -23483 6110 -23449
rect 6110 -23483 6183 -23449
rect 5787 -23579 5864 -23545
rect 5670 -23741 5846 -23707
rect 5577 -23785 5611 -23751
rect 6457 -23531 6491 -23305
rect 6667 -23387 6744 -23353
rect 6544 -23483 6550 -23449
rect 6550 -23483 6623 -23449
rect 6227 -23579 6304 -23545
rect 6110 -23741 6286 -23707
rect 6017 -23785 6051 -23751
rect 5670 -23829 5846 -23795
rect 6667 -23579 6744 -23545
rect 6550 -23741 6726 -23707
rect 6457 -23785 6491 -23751
rect 6110 -23829 6286 -23795
rect 6550 -23829 6726 -23795
rect -17523 -23905 -17433 -23871
rect 7389 -23892 7677 -23857
rect 8337 -23892 8625 -23857
rect 9273 -23892 9561 -23857
rect 10204 -23892 10492 -23857
rect 11131 -23892 11419 -23857
rect -24268 -23965 -24194 -23931
rect -24194 -23965 -24188 -23931
rect -24135 -23995 -24100 -23961
rect 5689 -23931 5821 -23897
rect 6129 -23931 6261 -23897
rect 6569 -23931 6701 -23897
rect -11563 -23970 -11494 -23960
rect -11563 -24019 -11553 -23970
rect -11553 -24019 -11504 -23970
rect -11504 -24019 -11494 -23970
rect -24390 -24061 -24384 -24027
rect -24384 -24061 -24310 -24027
rect -11563 -24029 -11494 -24019
rect 7150 -24074 7184 -23964
rect 7245 -24259 7246 -24152
rect 7246 -24259 7280 -24152
rect 7245 -24264 7280 -24259
rect 7342 -24074 7376 -23964
rect 7534 -24074 7568 -23964
rect 7438 -24259 7472 -24152
rect 7472 -24259 7473 -24152
rect 7438 -24264 7473 -24259
rect 7726 -24074 7760 -23964
rect 7630 -24259 7664 -24152
rect 7664 -24259 7665 -24152
rect 7630 -24264 7665 -24259
rect 7918 -24074 7952 -23964
rect 7822 -24259 7856 -24152
rect 7856 -24259 7857 -24152
rect 7822 -24264 7857 -24259
rect 8098 -24074 8132 -23964
rect 8193 -24259 8194 -24152
rect 8194 -24259 8228 -24152
rect 8193 -24264 8228 -24259
rect 8290 -24074 8324 -23964
rect 8482 -24074 8516 -23964
rect 8386 -24259 8420 -24152
rect 8420 -24259 8421 -24152
rect 8386 -24264 8421 -24259
rect 8674 -24074 8708 -23964
rect 8578 -24259 8612 -24152
rect 8612 -24259 8613 -24152
rect 8578 -24264 8613 -24259
rect 8866 -24074 8900 -23964
rect 8770 -24259 8804 -24152
rect 8804 -24259 8805 -24152
rect 8770 -24264 8805 -24259
rect 9034 -24074 9068 -23964
rect 9129 -24259 9130 -24152
rect 9130 -24259 9164 -24152
rect 9129 -24264 9164 -24259
rect 9226 -24074 9260 -23964
rect 9418 -24074 9452 -23964
rect 9322 -24259 9356 -24152
rect 9356 -24259 9357 -24152
rect 9322 -24264 9357 -24259
rect 9610 -24074 9644 -23964
rect 9514 -24259 9548 -24152
rect 9548 -24259 9549 -24152
rect 9514 -24264 9549 -24259
rect 9802 -24074 9836 -23964
rect 9706 -24259 9740 -24152
rect 9740 -24259 9741 -24152
rect 9706 -24264 9741 -24259
rect 9965 -24074 9999 -23964
rect 10060 -24259 10061 -24152
rect 10061 -24259 10095 -24152
rect 10060 -24264 10095 -24259
rect 10157 -24074 10191 -23964
rect 10349 -24074 10383 -23964
rect 10253 -24259 10287 -24152
rect 10287 -24259 10288 -24152
rect 10253 -24264 10288 -24259
rect 10541 -24074 10575 -23964
rect 10445 -24259 10479 -24152
rect 10479 -24259 10480 -24152
rect 10445 -24264 10480 -24259
rect 10733 -24074 10767 -23964
rect 10637 -24259 10671 -24152
rect 10671 -24259 10672 -24152
rect 10637 -24264 10672 -24259
rect 10892 -24074 10926 -23964
rect 10987 -24259 10988 -24152
rect 10988 -24259 11022 -24152
rect 10987 -24264 11022 -24259
rect 11084 -24074 11118 -23964
rect 11276 -24074 11310 -23964
rect 11180 -24259 11214 -24152
rect 11214 -24259 11215 -24152
rect 11180 -24264 11215 -24259
rect 11468 -24074 11502 -23964
rect 11372 -24259 11406 -24152
rect 11406 -24259 11407 -24152
rect 11372 -24264 11407 -24259
rect 11660 -24074 11694 -23964
rect 11564 -24259 11598 -24152
rect 11598 -24259 11599 -24152
rect 11564 -24264 11599 -24259
rect -17523 -24345 -17433 -24311
rect 7198 -24352 7232 -24318
rect 7390 -24352 7424 -24318
rect 7582 -24352 7616 -24318
rect 7774 -24352 7808 -24318
rect 8146 -24352 8180 -24318
rect 8338 -24352 8372 -24318
rect 8530 -24352 8564 -24318
rect 8722 -24352 8756 -24318
rect 9082 -24352 9116 -24318
rect 9274 -24352 9308 -24318
rect 9466 -24352 9500 -24318
rect 9658 -24352 9692 -24318
rect 10013 -24352 10047 -24318
rect 10205 -24352 10239 -24318
rect 10397 -24352 10431 -24318
rect 10589 -24352 10623 -24318
rect 10940 -24352 10974 -24318
rect 11132 -24352 11166 -24318
rect 11324 -24352 11358 -24318
rect 11516 -24352 11550 -24318
rect -17665 -24441 -17575 -24407
rect -17523 -24537 -17433 -24503
rect -17665 -24633 -17575 -24599
rect -17523 -24729 -17433 -24695
rect -17266 -24777 -17232 -24743
rect -17665 -24825 -17575 -24791
rect -17176 -24825 -17000 -24791
rect -17523 -24921 -17433 -24887
rect -17371 -24920 -17337 -24886
rect -17820 -25279 -17769 -24922
rect -16917 -24907 -16856 -24708
rect -17665 -25017 -17575 -24983
rect 7298 -25050 7332 -24702
rect 7332 -25050 7333 -24702
rect -17523 -25113 -17433 -25079
rect 7298 -25102 7333 -25050
rect -17665 -25209 -17575 -25175
rect -17523 -25305 -17433 -25271
rect -12471 -26465 -12399 -25343
rect -12293 -25347 -12191 -25313
rect -11902 -25347 -11835 -25313
rect -12109 -25443 -11985 -25409
rect -12293 -25539 -12191 -25505
rect -11902 -25539 -11835 -25505
rect -12110 -25635 -11986 -25601
rect -11411 -25379 -11356 -25314
rect -11262 -25347 -11156 -25313
rect -11582 -25488 -11514 -25481
rect -11582 -25553 -11576 -25488
rect -11576 -25553 -11521 -25488
rect -11521 -25553 -11514 -25488
rect -11582 -25561 -11514 -25553
rect -12293 -25731 -12191 -25697
rect -11895 -25731 -11835 -25697
rect -12110 -25827 -11986 -25793
rect -11583 -25795 -11530 -25681
rect -11277 -25443 -11262 -25409
rect -11262 -25443 -11243 -25409
rect -11176 -25539 -11156 -25505
rect -11156 -25539 -11142 -25505
rect -11277 -25635 -11262 -25601
rect -11262 -25635 -11243 -25601
rect -11176 -25731 -11156 -25697
rect -11156 -25731 -11142 -25697
rect -11277 -25827 -11262 -25793
rect -11262 -25827 -11243 -25793
rect -12293 -25923 -12191 -25889
rect -11878 -25923 -11835 -25889
rect -11176 -25923 -11156 -25889
rect -11156 -25923 -11142 -25889
rect -12110 -26019 -11986 -25985
rect -12294 -26115 -12192 -26081
rect -11895 -26115 -11835 -26081
rect -11276 -26019 -11262 -25985
rect -11262 -26019 -11242 -25985
rect -11176 -26115 -11156 -26081
rect -11156 -26115 -11142 -26081
rect -12110 -26211 -11986 -26177
rect -12296 -26307 -12194 -26273
rect -11901 -26307 -11835 -26273
rect -12110 -26403 -11986 -26369
rect -12296 -26499 -12194 -26465
rect -11901 -26499 -11799 -26465
rect -11277 -26211 -11262 -26177
rect -11262 -26211 -11243 -26177
rect -11575 -26401 -11522 -26268
rect -11176 -26307 -11156 -26273
rect -11156 -26307 -11142 -26273
rect -11277 -26403 -11262 -26369
rect -11262 -26403 -11243 -26369
rect -11068 -26465 -11022 -25342
rect 7298 -25453 7332 -25102
rect 7332 -25453 7333 -25102
rect 7372 -25466 7406 -24690
rect 7756 -25466 7790 -24690
rect 8246 -25050 8280 -24702
rect 8280 -25050 8281 -24702
rect 8246 -25102 8281 -25050
rect 8246 -25453 8280 -25102
rect 8280 -25453 8281 -25102
rect 8320 -25466 8354 -24690
rect 8704 -25466 8738 -24690
rect 9182 -25050 9216 -24702
rect 9216 -25050 9217 -24702
rect 9182 -25102 9217 -25050
rect 9182 -25453 9216 -25102
rect 9216 -25453 9217 -25102
rect 9256 -25466 9290 -24690
rect 9640 -25466 9674 -24690
rect 10113 -25050 10147 -24702
rect 10147 -25050 10148 -24702
rect 10113 -25102 10148 -25050
rect 10113 -25453 10147 -25102
rect 10147 -25453 10148 -25102
rect 10187 -25466 10221 -24690
rect 10571 -25466 10605 -24690
rect 11040 -25050 11074 -24702
rect 11074 -25050 11075 -24702
rect 11040 -25102 11075 -25050
rect 11040 -25453 11074 -25102
rect 11074 -25453 11075 -25102
rect 11114 -25466 11148 -24690
rect 11498 -25466 11532 -24690
rect 11811 -25067 12168 -25016
rect 11785 -25403 11819 -25313
rect 11881 -25261 11915 -25171
rect 11977 -25403 12011 -25313
rect 12073 -25261 12107 -25171
rect 12169 -25403 12203 -25313
rect 12265 -25261 12299 -25171
rect 12361 -25403 12395 -25313
rect 12457 -25261 12491 -25171
rect 12553 -25403 12587 -25313
rect 12649 -25261 12683 -25171
rect 12986 -25237 13077 -25203
rect 12745 -25403 12779 -25313
rect 12929 -25309 12935 -25275
rect 12935 -25309 13008 -25275
rect 12170 -25499 12204 -25465
rect 12842 -25549 12876 -25323
rect 13052 -25405 13129 -25371
rect 12929 -25501 12935 -25467
rect 12935 -25501 13008 -25467
rect 7298 -25982 7332 -25631
rect 7332 -25982 7333 -25631
rect 7298 -26034 7333 -25982
rect 7298 -26382 7332 -26034
rect 7332 -26382 7333 -26034
rect 7372 -26394 7406 -25618
rect 7756 -26394 7790 -25618
rect 8246 -25982 8280 -25631
rect 8280 -25982 8281 -25631
rect 8246 -26034 8281 -25982
rect 8246 -26382 8280 -26034
rect 8280 -26382 8281 -26034
rect 8320 -26394 8354 -25618
rect 8704 -26394 8738 -25618
rect 9182 -25982 9216 -25631
rect 9216 -25982 9217 -25631
rect 9182 -26034 9217 -25982
rect 9182 -26382 9216 -26034
rect 9216 -26382 9217 -26034
rect 9256 -26394 9290 -25618
rect 9640 -26394 9674 -25618
rect 10113 -25981 10147 -25630
rect 10147 -25981 10148 -25630
rect 10113 -26033 10148 -25981
rect 10113 -26381 10147 -26033
rect 10147 -26381 10148 -26033
rect 10187 -26393 10221 -25617
rect 10571 -26393 10605 -25617
rect 11040 -25982 11074 -25631
rect 11074 -25982 11075 -25631
rect 11040 -26034 11075 -25982
rect 11040 -26382 11074 -26034
rect 11074 -26382 11075 -26034
rect 11114 -26394 11148 -25618
rect 12313 -25604 12347 -25570
rect 11498 -26394 11532 -25618
rect 12265 -25836 12299 -25660
rect 13052 -25597 13129 -25563
rect 12935 -25759 13111 -25725
rect 12842 -25803 12876 -25769
rect 12935 -25847 13111 -25813
rect 12183 -25980 12382 -25919
rect 12954 -25949 13086 -25915
rect -11262 -26499 -11156 -26465
rect -11564 -26758 -11492 -26748
rect -11564 -26810 -11554 -26758
rect -11554 -26810 -11502 -26758
rect -11502 -26810 -11492 -26758
rect 7198 -26766 7232 -26732
rect 7390 -26766 7424 -26732
rect 7582 -26766 7616 -26732
rect 7774 -26766 7808 -26732
rect 8146 -26766 8180 -26732
rect 8338 -26766 8372 -26732
rect 8530 -26766 8564 -26732
rect 8722 -26766 8756 -26732
rect 9082 -26766 9116 -26732
rect 9274 -26766 9308 -26732
rect 9466 -26766 9500 -26732
rect 9658 -26766 9692 -26732
rect 10013 -26765 10047 -26731
rect 10205 -26765 10239 -26731
rect 10397 -26765 10431 -26731
rect 10589 -26765 10623 -26731
rect 10940 -26766 10974 -26732
rect 11132 -26766 11166 -26732
rect 11324 -26766 11358 -26732
rect 11516 -26766 11550 -26732
rect -11564 -26820 -11492 -26810
rect 7245 -26825 7280 -26820
rect 7245 -26932 7246 -26825
rect 7246 -26932 7280 -26825
rect 7150 -27120 7184 -27010
rect 7342 -27120 7376 -27010
rect 7438 -26825 7473 -26820
rect 7438 -26932 7472 -26825
rect 7472 -26932 7473 -26825
rect 7534 -27120 7568 -27010
rect 7630 -26825 7665 -26820
rect 7630 -26932 7664 -26825
rect 7664 -26932 7665 -26825
rect 7726 -27120 7760 -27010
rect 7822 -26825 7857 -26820
rect 7822 -26932 7856 -26825
rect 7856 -26932 7857 -26825
rect 7918 -27120 7952 -27010
rect 8193 -26825 8228 -26820
rect 8193 -26932 8194 -26825
rect 8194 -26932 8228 -26825
rect 8098 -27120 8132 -27010
rect 8290 -27120 8324 -27010
rect 8386 -26825 8421 -26820
rect 8386 -26932 8420 -26825
rect 8420 -26932 8421 -26825
rect 8482 -27120 8516 -27010
rect 8578 -26825 8613 -26820
rect 8578 -26932 8612 -26825
rect 8612 -26932 8613 -26825
rect 8674 -27120 8708 -27010
rect 8770 -26825 8805 -26820
rect 8770 -26932 8804 -26825
rect 8804 -26932 8805 -26825
rect 8866 -27120 8900 -27010
rect 9129 -26825 9164 -26820
rect 9129 -26932 9130 -26825
rect 9130 -26932 9164 -26825
rect 9034 -27120 9068 -27010
rect 9226 -27120 9260 -27010
rect 9322 -26825 9357 -26820
rect 9322 -26932 9356 -26825
rect 9356 -26932 9357 -26825
rect 9418 -27120 9452 -27010
rect 9514 -26825 9549 -26820
rect 9514 -26932 9548 -26825
rect 9548 -26932 9549 -26825
rect 9610 -27120 9644 -27010
rect 9706 -26825 9741 -26820
rect 9706 -26932 9740 -26825
rect 9740 -26932 9741 -26825
rect 9802 -27120 9836 -27010
rect 10060 -26824 10095 -26819
rect 10060 -26931 10061 -26824
rect 10061 -26931 10095 -26824
rect 9965 -27119 9999 -27009
rect 10157 -27119 10191 -27009
rect 10253 -26824 10288 -26819
rect 10253 -26931 10287 -26824
rect 10287 -26931 10288 -26824
rect 10349 -27119 10383 -27009
rect 10445 -26824 10480 -26819
rect 10445 -26931 10479 -26824
rect 10479 -26931 10480 -26824
rect 10541 -27119 10575 -27009
rect 10637 -26824 10672 -26819
rect 10637 -26931 10671 -26824
rect 10671 -26931 10672 -26824
rect 10733 -27119 10767 -27009
rect 10987 -26825 11022 -26820
rect 10987 -26932 10988 -26825
rect 10988 -26932 11022 -26825
rect 10892 -27120 10926 -27010
rect 11084 -27120 11118 -27010
rect 11180 -26825 11215 -26820
rect 11180 -26932 11214 -26825
rect 11214 -26932 11215 -26825
rect 11276 -27120 11310 -27010
rect 11372 -26825 11407 -26820
rect 11372 -26932 11406 -26825
rect 11406 -26932 11407 -26825
rect 11468 -27120 11502 -27010
rect 11564 -26825 11599 -26820
rect 11564 -26932 11598 -26825
rect 11598 -26932 11599 -26825
rect 11660 -27120 11694 -27010
rect 7389 -27227 7677 -27192
rect 8337 -27227 8625 -27192
rect 9273 -27227 9561 -27192
rect 10204 -27226 10492 -27191
rect 11131 -27227 11419 -27192
rect 5721 -27747 5812 -27713
rect 6161 -27747 6252 -27713
rect 6601 -27747 6692 -27713
rect 5664 -27819 5670 -27785
rect 5670 -27819 5743 -27785
rect -12471 -29098 -12399 -27976
rect -12293 -27980 -12191 -27946
rect -11902 -27980 -11835 -27946
rect -12109 -28076 -11985 -28042
rect -12293 -28172 -12191 -28138
rect -11902 -28172 -11835 -28138
rect -12110 -28268 -11986 -28234
rect -11411 -28012 -11356 -27947
rect -11262 -27980 -11156 -27946
rect -11582 -28121 -11514 -28114
rect -11582 -28186 -11576 -28121
rect -11576 -28186 -11521 -28121
rect -11521 -28186 -11514 -28121
rect -11582 -28194 -11514 -28186
rect -12293 -28364 -12191 -28330
rect -11895 -28364 -11835 -28330
rect -12110 -28460 -11986 -28426
rect -11583 -28428 -11530 -28314
rect -11277 -28076 -11262 -28042
rect -11262 -28076 -11243 -28042
rect -11176 -28172 -11156 -28138
rect -11156 -28172 -11142 -28138
rect -11277 -28268 -11262 -28234
rect -11262 -28268 -11243 -28234
rect -11176 -28364 -11156 -28330
rect -11156 -28364 -11142 -28330
rect -11277 -28460 -11262 -28426
rect -11262 -28460 -11243 -28426
rect -12293 -28556 -12191 -28522
rect -11878 -28556 -11835 -28522
rect -11176 -28556 -11156 -28522
rect -11156 -28556 -11142 -28522
rect -12110 -28652 -11986 -28618
rect -12294 -28748 -12192 -28714
rect -11895 -28748 -11835 -28714
rect -11276 -28652 -11262 -28618
rect -11262 -28652 -11242 -28618
rect -11176 -28748 -11156 -28714
rect -11156 -28748 -11142 -28714
rect -12110 -28844 -11986 -28810
rect -12296 -28940 -12194 -28906
rect -11901 -28940 -11835 -28906
rect -12110 -29036 -11986 -29002
rect -12296 -29132 -12194 -29098
rect -11901 -29132 -11799 -29098
rect -11277 -28844 -11262 -28810
rect -11262 -28844 -11243 -28810
rect -11575 -29034 -11522 -28901
rect -11176 -28940 -11156 -28906
rect -11156 -28940 -11142 -28906
rect -11277 -29036 -11262 -29002
rect -11262 -29036 -11243 -29002
rect -11068 -29098 -11022 -27975
rect 5577 -28059 5611 -27833
rect 6104 -27819 6110 -27785
rect 6110 -27819 6183 -27785
rect 5787 -27915 5864 -27881
rect 5664 -28011 5670 -27977
rect 5670 -28011 5743 -27977
rect 6017 -28059 6051 -27833
rect 6544 -27819 6550 -27785
rect 6550 -27819 6623 -27785
rect 6227 -27915 6304 -27881
rect 6104 -28011 6110 -27977
rect 6110 -28011 6183 -27977
rect 5787 -28107 5864 -28073
rect 5670 -28269 5846 -28235
rect 5577 -28313 5611 -28279
rect 6457 -28059 6491 -27833
rect 6667 -27915 6744 -27881
rect 6544 -28011 6550 -27977
rect 6550 -28011 6623 -27977
rect 6227 -28107 6304 -28073
rect 6110 -28269 6286 -28235
rect 6017 -28313 6051 -28279
rect 5670 -28357 5846 -28323
rect 6667 -28107 6744 -28073
rect 6550 -28269 6726 -28235
rect 6457 -28313 6491 -28279
rect 6110 -28357 6286 -28323
rect 6550 -28357 6726 -28323
rect 7389 -28420 7677 -28385
rect 8337 -28420 8625 -28385
rect 9273 -28420 9561 -28385
rect 10204 -28420 10492 -28385
rect 11131 -28420 11419 -28385
rect 5689 -28459 5821 -28425
rect 6129 -28459 6261 -28425
rect 6569 -28459 6701 -28425
rect 7150 -28602 7184 -28492
rect 7245 -28787 7246 -28680
rect 7246 -28787 7280 -28680
rect 7245 -28792 7280 -28787
rect 7342 -28602 7376 -28492
rect 7534 -28602 7568 -28492
rect 7438 -28787 7472 -28680
rect 7472 -28787 7473 -28680
rect 7438 -28792 7473 -28787
rect 7726 -28602 7760 -28492
rect 7630 -28787 7664 -28680
rect 7664 -28787 7665 -28680
rect 7630 -28792 7665 -28787
rect 7918 -28602 7952 -28492
rect 7822 -28787 7856 -28680
rect 7856 -28787 7857 -28680
rect 7822 -28792 7857 -28787
rect 8098 -28602 8132 -28492
rect 8193 -28787 8194 -28680
rect 8194 -28787 8228 -28680
rect 8193 -28792 8228 -28787
rect 8290 -28602 8324 -28492
rect 8482 -28602 8516 -28492
rect 8386 -28787 8420 -28680
rect 8420 -28787 8421 -28680
rect 8386 -28792 8421 -28787
rect 8674 -28602 8708 -28492
rect 8578 -28787 8612 -28680
rect 8612 -28787 8613 -28680
rect 8578 -28792 8613 -28787
rect 8866 -28602 8900 -28492
rect 8770 -28787 8804 -28680
rect 8804 -28787 8805 -28680
rect 8770 -28792 8805 -28787
rect 9034 -28602 9068 -28492
rect 9129 -28787 9130 -28680
rect 9130 -28787 9164 -28680
rect 9129 -28792 9164 -28787
rect 9226 -28602 9260 -28492
rect 9418 -28602 9452 -28492
rect 9322 -28787 9356 -28680
rect 9356 -28787 9357 -28680
rect 9322 -28792 9357 -28787
rect 9610 -28602 9644 -28492
rect 9514 -28787 9548 -28680
rect 9548 -28787 9549 -28680
rect 9514 -28792 9549 -28787
rect 9802 -28602 9836 -28492
rect 9706 -28787 9740 -28680
rect 9740 -28787 9741 -28680
rect 9706 -28792 9741 -28787
rect 9965 -28602 9999 -28492
rect 10060 -28787 10061 -28680
rect 10061 -28787 10095 -28680
rect 10060 -28792 10095 -28787
rect 10157 -28602 10191 -28492
rect 10349 -28602 10383 -28492
rect 10253 -28787 10287 -28680
rect 10287 -28787 10288 -28680
rect 10253 -28792 10288 -28787
rect 10541 -28602 10575 -28492
rect 10445 -28787 10479 -28680
rect 10479 -28787 10480 -28680
rect 10445 -28792 10480 -28787
rect 10733 -28602 10767 -28492
rect 10637 -28787 10671 -28680
rect 10671 -28787 10672 -28680
rect 10637 -28792 10672 -28787
rect 10892 -28602 10926 -28492
rect 10987 -28787 10988 -28680
rect 10988 -28787 11022 -28680
rect 10987 -28792 11022 -28787
rect 11084 -28602 11118 -28492
rect 11276 -28602 11310 -28492
rect 11180 -28787 11214 -28680
rect 11214 -28787 11215 -28680
rect 11180 -28792 11215 -28787
rect 11468 -28602 11502 -28492
rect 11372 -28787 11406 -28680
rect 11406 -28787 11407 -28680
rect 11372 -28792 11407 -28787
rect 11660 -28602 11694 -28492
rect 11564 -28787 11598 -28680
rect 11598 -28787 11599 -28680
rect 11564 -28792 11599 -28787
rect 7198 -28880 7232 -28846
rect 7390 -28880 7424 -28846
rect 7582 -28880 7616 -28846
rect 7774 -28880 7808 -28846
rect 8146 -28880 8180 -28846
rect 8338 -28880 8372 -28846
rect 8530 -28880 8564 -28846
rect 8722 -28880 8756 -28846
rect 9082 -28880 9116 -28846
rect 9274 -28880 9308 -28846
rect 9466 -28880 9500 -28846
rect 9658 -28880 9692 -28846
rect 10013 -28880 10047 -28846
rect 10205 -28880 10239 -28846
rect 10397 -28880 10431 -28846
rect 10589 -28880 10623 -28846
rect 10940 -28880 10974 -28846
rect 11132 -28880 11166 -28846
rect 11324 -28880 11358 -28846
rect 11516 -28880 11550 -28846
rect -11262 -29132 -11156 -29098
rect -11562 -29395 -11494 -29385
rect -11562 -29443 -11552 -29395
rect -11552 -29443 -11504 -29395
rect -11504 -29443 -11494 -29395
rect -11562 -29453 -11494 -29443
rect 7298 -29578 7332 -29230
rect 7332 -29578 7333 -29230
rect 7298 -29630 7333 -29578
rect 7298 -29981 7332 -29630
rect 7332 -29981 7333 -29630
rect 7372 -29994 7406 -29218
rect 7756 -29994 7790 -29218
rect 8246 -29578 8280 -29230
rect 8280 -29578 8281 -29230
rect 8246 -29630 8281 -29578
rect 8246 -29981 8280 -29630
rect 8280 -29981 8281 -29630
rect 8320 -29994 8354 -29218
rect 8704 -29994 8738 -29218
rect 9182 -29578 9216 -29230
rect 9216 -29578 9217 -29230
rect 9182 -29630 9217 -29578
rect 9182 -29981 9216 -29630
rect 9216 -29981 9217 -29630
rect 9256 -29994 9290 -29218
rect 9640 -29994 9674 -29218
rect 10113 -29578 10147 -29230
rect 10147 -29578 10148 -29230
rect 10113 -29630 10148 -29578
rect 10113 -29981 10147 -29630
rect 10147 -29981 10148 -29630
rect 10187 -29994 10221 -29218
rect 10571 -29994 10605 -29218
rect 11040 -29578 11074 -29230
rect 11074 -29578 11075 -29230
rect 11040 -29630 11075 -29578
rect 11040 -29981 11074 -29630
rect 11074 -29981 11075 -29630
rect 11114 -29994 11148 -29218
rect 11498 -29994 11532 -29218
rect 11811 -29595 12168 -29544
rect 11785 -29931 11819 -29841
rect 11881 -29789 11915 -29699
rect 11977 -29931 12011 -29841
rect 12073 -29789 12107 -29699
rect 12169 -29931 12203 -29841
rect 12265 -29789 12299 -29699
rect 12361 -29931 12395 -29841
rect 12457 -29789 12491 -29699
rect 12553 -29931 12587 -29841
rect 12649 -29789 12683 -29699
rect 12986 -29765 13077 -29731
rect 12745 -29931 12779 -29841
rect 12929 -29837 12935 -29803
rect 12935 -29837 13008 -29803
rect 12170 -30027 12204 -29993
rect 12842 -30077 12876 -29851
rect 13052 -29933 13129 -29899
rect 12929 -30029 12935 -29995
rect 12935 -30029 13008 -29995
rect -12471 -31707 -12399 -30585
rect -12293 -30589 -12191 -30555
rect -11902 -30589 -11835 -30555
rect -12109 -30685 -11985 -30651
rect -12293 -30781 -12191 -30747
rect -11902 -30781 -11835 -30747
rect -12110 -30877 -11986 -30843
rect 7298 -30510 7332 -30159
rect 7332 -30510 7333 -30159
rect -11411 -30621 -11356 -30556
rect -11262 -30589 -11156 -30555
rect -11582 -30730 -11514 -30723
rect -11582 -30795 -11576 -30730
rect -11576 -30795 -11521 -30730
rect -11521 -30795 -11514 -30730
rect -11582 -30803 -11514 -30795
rect -12293 -30973 -12191 -30939
rect -11895 -30973 -11835 -30939
rect -12110 -31069 -11986 -31035
rect -11583 -31037 -11530 -30923
rect -11277 -30685 -11262 -30651
rect -11262 -30685 -11243 -30651
rect -11176 -30781 -11156 -30747
rect -11156 -30781 -11142 -30747
rect -11277 -30877 -11262 -30843
rect -11262 -30877 -11243 -30843
rect -11176 -30973 -11156 -30939
rect -11156 -30973 -11142 -30939
rect -11277 -31069 -11262 -31035
rect -11262 -31069 -11243 -31035
rect -12293 -31165 -12191 -31131
rect -11878 -31165 -11835 -31131
rect -11176 -31165 -11156 -31131
rect -11156 -31165 -11142 -31131
rect -12110 -31261 -11986 -31227
rect -12294 -31357 -12192 -31323
rect -11895 -31357 -11835 -31323
rect -11276 -31261 -11262 -31227
rect -11262 -31261 -11242 -31227
rect -11176 -31357 -11156 -31323
rect -11156 -31357 -11142 -31323
rect -12110 -31453 -11986 -31419
rect -12296 -31549 -12194 -31515
rect -11901 -31549 -11835 -31515
rect -12110 -31645 -11986 -31611
rect -12296 -31741 -12194 -31707
rect -11901 -31741 -11799 -31707
rect -11277 -31453 -11262 -31419
rect -11262 -31453 -11243 -31419
rect -11575 -31643 -11522 -31510
rect -11176 -31549 -11156 -31515
rect -11156 -31549 -11142 -31515
rect -11277 -31645 -11262 -31611
rect -11262 -31645 -11243 -31611
rect -11068 -31707 -11022 -30584
rect 7298 -30562 7333 -30510
rect 7298 -30910 7332 -30562
rect 7332 -30910 7333 -30562
rect 7372 -30922 7406 -30146
rect 7756 -30922 7790 -30146
rect 8246 -30510 8280 -30159
rect 8280 -30510 8281 -30159
rect 8246 -30562 8281 -30510
rect 8246 -30910 8280 -30562
rect 8280 -30910 8281 -30562
rect 8320 -30922 8354 -30146
rect 8704 -30922 8738 -30146
rect 9182 -30510 9216 -30159
rect 9216 -30510 9217 -30159
rect 9182 -30562 9217 -30510
rect 9182 -30910 9216 -30562
rect 9216 -30910 9217 -30562
rect 9256 -30922 9290 -30146
rect 9640 -30922 9674 -30146
rect 10113 -30509 10147 -30158
rect 10147 -30509 10148 -30158
rect 10113 -30561 10148 -30509
rect 10113 -30909 10147 -30561
rect 10147 -30909 10148 -30561
rect 10187 -30921 10221 -30145
rect 10571 -30921 10605 -30145
rect 11040 -30510 11074 -30159
rect 11074 -30510 11075 -30159
rect 11040 -30562 11075 -30510
rect 11040 -30910 11074 -30562
rect 11074 -30910 11075 -30562
rect 11114 -30922 11148 -30146
rect 12313 -30132 12347 -30098
rect 11498 -30922 11532 -30146
rect 12265 -30364 12299 -30188
rect 13052 -30125 13129 -30091
rect 12935 -30287 13111 -30253
rect 12842 -30331 12876 -30297
rect 12935 -30375 13111 -30341
rect 12183 -30508 12382 -30447
rect 12954 -30477 13086 -30443
rect 7198 -31294 7232 -31260
rect 7390 -31294 7424 -31260
rect 7582 -31294 7616 -31260
rect 7774 -31294 7808 -31260
rect 8146 -31294 8180 -31260
rect 8338 -31294 8372 -31260
rect 8530 -31294 8564 -31260
rect 8722 -31294 8756 -31260
rect 9082 -31294 9116 -31260
rect 9274 -31294 9308 -31260
rect 9466 -31294 9500 -31260
rect 9658 -31294 9692 -31260
rect 10013 -31293 10047 -31259
rect 10205 -31293 10239 -31259
rect 10397 -31293 10431 -31259
rect 10589 -31293 10623 -31259
rect 10940 -31294 10974 -31260
rect 11132 -31294 11166 -31260
rect 11324 -31294 11358 -31260
rect 11516 -31294 11550 -31260
rect 7245 -31353 7280 -31348
rect 7245 -31460 7246 -31353
rect 7246 -31460 7280 -31353
rect 7150 -31648 7184 -31538
rect 7342 -31648 7376 -31538
rect 7438 -31353 7473 -31348
rect 7438 -31460 7472 -31353
rect 7472 -31460 7473 -31353
rect 7534 -31648 7568 -31538
rect 7630 -31353 7665 -31348
rect 7630 -31460 7664 -31353
rect 7664 -31460 7665 -31353
rect 7726 -31648 7760 -31538
rect 7822 -31353 7857 -31348
rect 7822 -31460 7856 -31353
rect 7856 -31460 7857 -31353
rect 7918 -31648 7952 -31538
rect 8193 -31353 8228 -31348
rect 8193 -31460 8194 -31353
rect 8194 -31460 8228 -31353
rect 8098 -31648 8132 -31538
rect 8290 -31648 8324 -31538
rect 8386 -31353 8421 -31348
rect 8386 -31460 8420 -31353
rect 8420 -31460 8421 -31353
rect 8482 -31648 8516 -31538
rect 8578 -31353 8613 -31348
rect 8578 -31460 8612 -31353
rect 8612 -31460 8613 -31353
rect 8674 -31648 8708 -31538
rect 8770 -31353 8805 -31348
rect 8770 -31460 8804 -31353
rect 8804 -31460 8805 -31353
rect 8866 -31648 8900 -31538
rect 9129 -31353 9164 -31348
rect 9129 -31460 9130 -31353
rect 9130 -31460 9164 -31353
rect 9034 -31648 9068 -31538
rect 9226 -31648 9260 -31538
rect 9322 -31353 9357 -31348
rect 9322 -31460 9356 -31353
rect 9356 -31460 9357 -31353
rect 9418 -31648 9452 -31538
rect 9514 -31353 9549 -31348
rect 9514 -31460 9548 -31353
rect 9548 -31460 9549 -31353
rect 9610 -31648 9644 -31538
rect 9706 -31353 9741 -31348
rect 9706 -31460 9740 -31353
rect 9740 -31460 9741 -31353
rect 9802 -31648 9836 -31538
rect 10060 -31352 10095 -31347
rect 10060 -31459 10061 -31352
rect 10061 -31459 10095 -31352
rect 9965 -31647 9999 -31537
rect 10157 -31647 10191 -31537
rect 10253 -31352 10288 -31347
rect 10253 -31459 10287 -31352
rect 10287 -31459 10288 -31352
rect 10349 -31647 10383 -31537
rect 10445 -31352 10480 -31347
rect 10445 -31459 10479 -31352
rect 10479 -31459 10480 -31352
rect 10541 -31647 10575 -31537
rect 10637 -31352 10672 -31347
rect 10637 -31459 10671 -31352
rect 10671 -31459 10672 -31352
rect 10733 -31647 10767 -31537
rect 10987 -31353 11022 -31348
rect 10987 -31460 10988 -31353
rect 10988 -31460 11022 -31353
rect 10892 -31648 10926 -31538
rect 11084 -31648 11118 -31538
rect 11180 -31353 11215 -31348
rect 11180 -31460 11214 -31353
rect 11214 -31460 11215 -31353
rect 11276 -31648 11310 -31538
rect 11372 -31353 11407 -31348
rect 11372 -31460 11406 -31353
rect 11406 -31460 11407 -31353
rect 11468 -31648 11502 -31538
rect 11564 -31353 11599 -31348
rect 11564 -31460 11598 -31353
rect 11598 -31460 11599 -31353
rect 11660 -31648 11694 -31538
rect -11262 -31741 -11156 -31707
rect 7389 -31755 7677 -31720
rect 8337 -31755 8625 -31720
rect 9273 -31755 9561 -31720
rect 10204 -31754 10492 -31719
rect 11131 -31755 11419 -31720
rect -11564 -31937 -11493 -31927
rect -11564 -31988 -11554 -31937
rect -11554 -31988 -11503 -31937
rect -11503 -31988 -11493 -31937
rect -11564 -31998 -11493 -31988
rect 5721 -32275 5812 -32241
rect 6161 -32275 6252 -32241
rect 6601 -32275 6692 -32241
rect 5664 -32347 5670 -32313
rect 5670 -32347 5743 -32313
rect 5577 -32587 5611 -32361
rect 6104 -32347 6110 -32313
rect 6110 -32347 6183 -32313
rect 5787 -32443 5864 -32409
rect 5664 -32539 5670 -32505
rect 5670 -32539 5743 -32505
rect 6017 -32587 6051 -32361
rect 6544 -32347 6550 -32313
rect 6550 -32347 6623 -32313
rect 6227 -32443 6304 -32409
rect 6104 -32539 6110 -32505
rect 6110 -32539 6183 -32505
rect 5787 -32635 5864 -32601
rect 5670 -32797 5846 -32763
rect 5577 -32841 5611 -32807
rect 6457 -32587 6491 -32361
rect 6667 -32443 6744 -32409
rect 6544 -32539 6550 -32505
rect 6550 -32539 6623 -32505
rect 6227 -32635 6304 -32601
rect 6110 -32797 6286 -32763
rect 6017 -32841 6051 -32807
rect 5670 -32885 5846 -32851
rect 6667 -32635 6744 -32601
rect 6550 -32797 6726 -32763
rect 6457 -32841 6491 -32807
rect 6110 -32885 6286 -32851
rect 6550 -32885 6726 -32851
rect 7389 -32948 7677 -32913
rect 8337 -32948 8625 -32913
rect 9273 -32948 9561 -32913
rect 10204 -32948 10492 -32913
rect 11131 -32948 11419 -32913
rect 5689 -32987 5821 -32953
rect 6129 -32987 6261 -32953
rect 6569 -32987 6701 -32953
rect -12473 -34327 -12401 -33205
rect -12295 -33209 -12193 -33175
rect -11904 -33209 -11837 -33175
rect -12111 -33305 -11987 -33271
rect -12295 -33401 -12193 -33367
rect -11904 -33401 -11837 -33367
rect -12112 -33497 -11988 -33463
rect 7150 -33130 7184 -33020
rect -11413 -33241 -11358 -33176
rect -11264 -33209 -11158 -33175
rect -11584 -33350 -11516 -33343
rect -11584 -33415 -11578 -33350
rect -11578 -33415 -11523 -33350
rect -11523 -33415 -11516 -33350
rect -11584 -33423 -11516 -33415
rect -12295 -33593 -12193 -33559
rect -11897 -33593 -11837 -33559
rect -12112 -33689 -11988 -33655
rect -11585 -33657 -11532 -33543
rect -11279 -33305 -11264 -33271
rect -11264 -33305 -11245 -33271
rect -11178 -33401 -11158 -33367
rect -11158 -33401 -11144 -33367
rect -11279 -33497 -11264 -33463
rect -11264 -33497 -11245 -33463
rect -11178 -33593 -11158 -33559
rect -11158 -33593 -11144 -33559
rect -11279 -33689 -11264 -33655
rect -11264 -33689 -11245 -33655
rect -12295 -33785 -12193 -33751
rect -11880 -33785 -11837 -33751
rect -11178 -33785 -11158 -33751
rect -11158 -33785 -11144 -33751
rect -12112 -33881 -11988 -33847
rect -12296 -33977 -12194 -33943
rect -11897 -33977 -11837 -33943
rect -11278 -33881 -11264 -33847
rect -11264 -33881 -11244 -33847
rect -11178 -33977 -11158 -33943
rect -11158 -33977 -11144 -33943
rect -12112 -34073 -11988 -34039
rect -12298 -34169 -12196 -34135
rect -11903 -34169 -11837 -34135
rect -12112 -34265 -11988 -34231
rect -12298 -34361 -12196 -34327
rect -11903 -34361 -11801 -34327
rect -11279 -34073 -11264 -34039
rect -11264 -34073 -11245 -34039
rect -11577 -34263 -11524 -34130
rect -11178 -34169 -11158 -34135
rect -11158 -34169 -11144 -34135
rect -11279 -34265 -11264 -34231
rect -11264 -34265 -11245 -34231
rect -11070 -34327 -11024 -33204
rect 7245 -33315 7246 -33208
rect 7246 -33315 7280 -33208
rect 7245 -33320 7280 -33315
rect 7342 -33130 7376 -33020
rect 7534 -33130 7568 -33020
rect 7438 -33315 7472 -33208
rect 7472 -33315 7473 -33208
rect 7438 -33320 7473 -33315
rect 7726 -33130 7760 -33020
rect 7630 -33315 7664 -33208
rect 7664 -33315 7665 -33208
rect 7630 -33320 7665 -33315
rect 7918 -33130 7952 -33020
rect 7822 -33315 7856 -33208
rect 7856 -33315 7857 -33208
rect 7822 -33320 7857 -33315
rect 8098 -33130 8132 -33020
rect 8193 -33315 8194 -33208
rect 8194 -33315 8228 -33208
rect 8193 -33320 8228 -33315
rect 8290 -33130 8324 -33020
rect 8482 -33130 8516 -33020
rect 8386 -33315 8420 -33208
rect 8420 -33315 8421 -33208
rect 8386 -33320 8421 -33315
rect 8674 -33130 8708 -33020
rect 8578 -33315 8612 -33208
rect 8612 -33315 8613 -33208
rect 8578 -33320 8613 -33315
rect 8866 -33130 8900 -33020
rect 8770 -33315 8804 -33208
rect 8804 -33315 8805 -33208
rect 8770 -33320 8805 -33315
rect 9034 -33130 9068 -33020
rect 9129 -33315 9130 -33208
rect 9130 -33315 9164 -33208
rect 9129 -33320 9164 -33315
rect 9226 -33130 9260 -33020
rect 9418 -33130 9452 -33020
rect 9322 -33315 9356 -33208
rect 9356 -33315 9357 -33208
rect 9322 -33320 9357 -33315
rect 9610 -33130 9644 -33020
rect 9514 -33315 9548 -33208
rect 9548 -33315 9549 -33208
rect 9514 -33320 9549 -33315
rect 9802 -33130 9836 -33020
rect 9706 -33315 9740 -33208
rect 9740 -33315 9741 -33208
rect 9706 -33320 9741 -33315
rect 9965 -33130 9999 -33020
rect 10060 -33315 10061 -33208
rect 10061 -33315 10095 -33208
rect 10060 -33320 10095 -33315
rect 10157 -33130 10191 -33020
rect 10349 -33130 10383 -33020
rect 10253 -33315 10287 -33208
rect 10287 -33315 10288 -33208
rect 10253 -33320 10288 -33315
rect 10541 -33130 10575 -33020
rect 10445 -33315 10479 -33208
rect 10479 -33315 10480 -33208
rect 10445 -33320 10480 -33315
rect 10733 -33130 10767 -33020
rect 10637 -33315 10671 -33208
rect 10671 -33315 10672 -33208
rect 10637 -33320 10672 -33315
rect 10892 -33130 10926 -33020
rect 10987 -33315 10988 -33208
rect 10988 -33315 11022 -33208
rect 10987 -33320 11022 -33315
rect 11084 -33130 11118 -33020
rect 11276 -33130 11310 -33020
rect 11180 -33315 11214 -33208
rect 11214 -33315 11215 -33208
rect 11180 -33320 11215 -33315
rect 11468 -33130 11502 -33020
rect 11372 -33315 11406 -33208
rect 11406 -33315 11407 -33208
rect 11372 -33320 11407 -33315
rect 11660 -33130 11694 -33020
rect 11564 -33315 11598 -33208
rect 11598 -33315 11599 -33208
rect 11564 -33320 11599 -33315
rect 7198 -33408 7232 -33374
rect 7390 -33408 7424 -33374
rect 7582 -33408 7616 -33374
rect 7774 -33408 7808 -33374
rect 8146 -33408 8180 -33374
rect 8338 -33408 8372 -33374
rect 8530 -33408 8564 -33374
rect 8722 -33408 8756 -33374
rect 9082 -33408 9116 -33374
rect 9274 -33408 9308 -33374
rect 9466 -33408 9500 -33374
rect 9658 -33408 9692 -33374
rect 10013 -33408 10047 -33374
rect 10205 -33408 10239 -33374
rect 10397 -33408 10431 -33374
rect 10589 -33408 10623 -33374
rect 10940 -33408 10974 -33374
rect 11132 -33408 11166 -33374
rect 11324 -33408 11358 -33374
rect 11516 -33408 11550 -33374
rect -11264 -34361 -11158 -34327
rect 7298 -34106 7332 -33758
rect 7332 -34106 7333 -33758
rect 7298 -34158 7333 -34106
rect 7298 -34509 7332 -34158
rect 7332 -34509 7333 -34158
rect 7372 -34522 7406 -33746
rect -11553 -34533 -11510 -34528
rect -11553 -34567 -11548 -34533
rect -11548 -34567 -11514 -34533
rect -11514 -34567 -11510 -34533
rect 7756 -34522 7790 -33746
rect 8246 -34106 8280 -33758
rect 8280 -34106 8281 -33758
rect 8246 -34158 8281 -34106
rect 8246 -34509 8280 -34158
rect 8280 -34509 8281 -34158
rect 8320 -34522 8354 -33746
rect 8704 -34522 8738 -33746
rect 9182 -34106 9216 -33758
rect 9216 -34106 9217 -33758
rect 9182 -34158 9217 -34106
rect 9182 -34509 9216 -34158
rect 9216 -34509 9217 -34158
rect 9256 -34522 9290 -33746
rect 9640 -34522 9674 -33746
rect 10113 -34106 10147 -33758
rect 10147 -34106 10148 -33758
rect 10113 -34158 10148 -34106
rect 10113 -34509 10147 -34158
rect 10147 -34509 10148 -34158
rect 10187 -34522 10221 -33746
rect 10571 -34522 10605 -33746
rect 11040 -34106 11074 -33758
rect 11074 -34106 11075 -33758
rect 11040 -34158 11075 -34106
rect 11040 -34509 11074 -34158
rect 11074 -34509 11075 -34158
rect 11114 -34522 11148 -33746
rect 11498 -34522 11532 -33746
rect 11811 -34123 12168 -34072
rect 11785 -34459 11819 -34369
rect 11881 -34317 11915 -34227
rect 11977 -34459 12011 -34369
rect 12073 -34317 12107 -34227
rect 12169 -34459 12203 -34369
rect 12265 -34317 12299 -34227
rect 12361 -34459 12395 -34369
rect 12457 -34317 12491 -34227
rect 12553 -34459 12587 -34369
rect 12649 -34317 12683 -34227
rect 12986 -34293 13077 -34259
rect 12745 -34459 12779 -34369
rect 12929 -34365 12935 -34331
rect 12935 -34365 13008 -34331
rect 12170 -34555 12204 -34521
rect -11553 -34571 -11510 -34567
rect 12842 -34605 12876 -34379
rect 13052 -34461 13129 -34427
rect 12929 -34557 12935 -34523
rect 12935 -34557 13008 -34523
rect 7298 -35038 7332 -34687
rect 7332 -35038 7333 -34687
rect 7298 -35090 7333 -35038
rect 7298 -35438 7332 -35090
rect 7332 -35438 7333 -35090
rect 7372 -35450 7406 -34674
rect 7756 -35450 7790 -34674
rect 8246 -35038 8280 -34687
rect 8280 -35038 8281 -34687
rect 8246 -35090 8281 -35038
rect 8246 -35438 8280 -35090
rect 8280 -35438 8281 -35090
rect 8320 -35450 8354 -34674
rect 8704 -35450 8738 -34674
rect 9182 -35038 9216 -34687
rect 9216 -35038 9217 -34687
rect 9182 -35090 9217 -35038
rect 9182 -35438 9216 -35090
rect 9216 -35438 9217 -35090
rect 9256 -35450 9290 -34674
rect 9640 -35450 9674 -34674
rect 10113 -35037 10147 -34686
rect 10147 -35037 10148 -34686
rect 10113 -35089 10148 -35037
rect 10113 -35437 10147 -35089
rect 10147 -35437 10148 -35089
rect 10187 -35449 10221 -34673
rect 10571 -35449 10605 -34673
rect 11040 -35038 11074 -34687
rect 11074 -35038 11075 -34687
rect 11040 -35090 11075 -35038
rect 11040 -35438 11074 -35090
rect 11074 -35438 11075 -35090
rect 11114 -35450 11148 -34674
rect 12313 -34660 12347 -34626
rect 11498 -35450 11532 -34674
rect 12265 -34892 12299 -34716
rect 13052 -34653 13129 -34619
rect 12935 -34815 13111 -34781
rect 12842 -34859 12876 -34825
rect 12935 -34903 13111 -34869
rect 12183 -35036 12382 -34975
rect 12954 -35005 13086 -34971
rect 12930 -35668 12964 -35634
rect 13184 -35668 13410 -35634
rect 7198 -35822 7232 -35788
rect 7390 -35822 7424 -35788
rect 7582 -35822 7616 -35788
rect 7774 -35822 7808 -35788
rect 8146 -35822 8180 -35788
rect 8338 -35822 8372 -35788
rect 8530 -35822 8564 -35788
rect 8722 -35822 8756 -35788
rect 9082 -35822 9116 -35788
rect 9274 -35822 9308 -35788
rect 9466 -35822 9500 -35788
rect 9658 -35822 9692 -35788
rect 10013 -35821 10047 -35787
rect 10205 -35821 10239 -35787
rect 10397 -35821 10431 -35787
rect 10589 -35821 10623 -35787
rect 10940 -35822 10974 -35788
rect 11132 -35822 11166 -35788
rect 11324 -35822 11358 -35788
rect 11516 -35822 11550 -35788
rect 7245 -35881 7280 -35876
rect 7245 -35988 7246 -35881
rect 7246 -35988 7280 -35881
rect 7150 -36176 7184 -36066
rect 7342 -36176 7376 -36066
rect 7438 -35881 7473 -35876
rect 7438 -35988 7472 -35881
rect 7472 -35988 7473 -35881
rect 7534 -36176 7568 -36066
rect 7630 -35881 7665 -35876
rect 7630 -35988 7664 -35881
rect 7664 -35988 7665 -35881
rect 7726 -36176 7760 -36066
rect 7822 -35881 7857 -35876
rect 7822 -35988 7856 -35881
rect 7856 -35988 7857 -35881
rect 7918 -36176 7952 -36066
rect 8193 -35881 8228 -35876
rect 8193 -35988 8194 -35881
rect 8194 -35988 8228 -35881
rect 8098 -36176 8132 -36066
rect 8290 -36176 8324 -36066
rect 8386 -35881 8421 -35876
rect 8386 -35988 8420 -35881
rect 8420 -35988 8421 -35881
rect 8482 -36176 8516 -36066
rect 8578 -35881 8613 -35876
rect 8578 -35988 8612 -35881
rect 8612 -35988 8613 -35881
rect 8674 -36176 8708 -36066
rect 8770 -35881 8805 -35876
rect 8770 -35988 8804 -35881
rect 8804 -35988 8805 -35881
rect 8866 -36176 8900 -36066
rect 9129 -35881 9164 -35876
rect 9129 -35988 9130 -35881
rect 9130 -35988 9164 -35881
rect 9034 -36176 9068 -36066
rect 9226 -36176 9260 -36066
rect 9322 -35881 9357 -35876
rect 9322 -35988 9356 -35881
rect 9356 -35988 9357 -35881
rect 9418 -36176 9452 -36066
rect 9514 -35881 9549 -35876
rect 9514 -35988 9548 -35881
rect 9548 -35988 9549 -35881
rect 9610 -36176 9644 -36066
rect 9706 -35881 9741 -35876
rect 9706 -35988 9740 -35881
rect 9740 -35988 9741 -35881
rect 9802 -36176 9836 -36066
rect 10060 -35880 10095 -35875
rect 10060 -35987 10061 -35880
rect 10061 -35987 10095 -35880
rect 9965 -36175 9999 -36065
rect 10157 -36175 10191 -36065
rect 10253 -35880 10288 -35875
rect 10253 -35987 10287 -35880
rect 10287 -35987 10288 -35880
rect 10349 -36175 10383 -36065
rect 10445 -35880 10480 -35875
rect 10445 -35987 10479 -35880
rect 10479 -35987 10480 -35880
rect 10541 -36175 10575 -36065
rect 10637 -35880 10672 -35875
rect 10637 -35987 10671 -35880
rect 10671 -35987 10672 -35880
rect 10733 -36175 10767 -36065
rect 10987 -35881 11022 -35876
rect 10987 -35988 10988 -35881
rect 10988 -35988 11022 -35881
rect 10892 -36176 10926 -36066
rect 11084 -36176 11118 -36066
rect 11180 -35881 11215 -35876
rect 11180 -35988 11214 -35881
rect 11214 -35988 11215 -35881
rect 11276 -36176 11310 -36066
rect 11372 -35881 11407 -35876
rect 11372 -35988 11406 -35881
rect 11406 -35988 11407 -35881
rect 11468 -36176 11502 -36066
rect 11564 -35881 11599 -35876
rect 11564 -35988 11598 -35881
rect 11598 -35988 11599 -35881
rect 12784 -35878 12818 -35746
rect 12886 -35903 12920 -35727
rect 12974 -35903 13008 -35727
rect 13136 -35921 13170 -35844
rect 13232 -35727 13266 -35721
rect 13232 -35800 13266 -35727
rect 13328 -35921 13362 -35844
rect 13424 -35727 13458 -35721
rect 13424 -35800 13458 -35727
rect 13496 -35869 13530 -35778
rect 12930 -36047 12964 -36013
rect 13184 -36047 13410 -36013
rect 11660 -36176 11694 -36066
rect 7389 -36283 7677 -36248
rect 8337 -36283 8625 -36248
rect 9273 -36283 9561 -36248
rect 10204 -36282 10492 -36247
rect 11131 -36283 11419 -36248
rect 12784 -36257 12818 -36125
rect 12886 -36282 12920 -36106
rect 12974 -36282 13008 -36106
rect 13136 -36300 13170 -36223
rect 13232 -36106 13266 -36100
rect 13232 -36179 13266 -36106
rect 13328 -36300 13362 -36223
rect 13424 -36106 13458 -36100
rect 13424 -36179 13458 -36106
rect 13496 -36248 13530 -36157
<< metal1 >>
rect -27350 6877 1670 6966
rect -27525 4541 -27436 4547
rect -27350 4541 -27261 6877
rect -21822 6725 -21816 6814
rect -21727 6725 -21721 6814
rect -21816 6684 -21727 6725
rect -21821 6595 -21720 6684
rect -15130 6664 -15022 6670
rect -25114 4541 -25005 4557
rect -27436 4452 -25005 4541
rect -27525 4446 -27436 4452
rect -25114 3948 -25005 4452
rect -24042 4517 -22832 4545
rect -24042 4445 -24000 4517
rect -22878 4445 -22832 4517
rect -24042 4411 -22832 4445
rect -24042 4339 -23788 4411
rect -24042 4237 -24030 4339
rect -23996 4237 -23838 4339
rect -23804 4237 -23788 4339
rect -24042 4219 -23788 4237
rect -23662 4340 -23212 4366
rect -23662 4339 -23262 4340
rect -23662 4237 -23646 4339
rect -23612 4237 -23454 4339
rect -23420 4238 -23262 4339
rect -23228 4238 -23212 4340
rect -23420 4237 -23212 4238
rect -23662 4219 -23212 4237
rect -23086 4342 -22832 4411
rect -23086 4240 -23070 4342
rect -23036 4240 -22878 4342
rect -22844 4240 -22832 4342
rect -23086 4219 -22832 4240
rect -22656 4490 -22498 4575
rect -22656 4418 -22632 4490
rect -22560 4418 -22498 4490
rect -23950 4156 -22924 4181
rect -23950 4155 -23742 4156
rect -23950 4031 -23934 4155
rect -23900 4032 -23742 4155
rect -23708 4032 -23550 4156
rect -23516 4032 -23358 4156
rect -23324 4032 -23166 4156
rect -23132 4032 -22974 4156
rect -22940 4032 -22924 4156
rect -23900 4031 -22924 4032
rect -23950 4002 -22924 4031
rect -24042 3948 -23788 3969
rect -25120 3839 -25114 3948
rect -25005 3839 -24999 3948
rect -24042 3881 -24030 3948
rect -23996 3881 -23838 3948
rect -23804 3881 -23788 3948
rect -24042 3822 -23788 3881
rect -23662 3941 -23212 3958
rect -23662 3881 -23646 3941
rect -23612 3924 -23262 3941
rect -23612 3881 -23454 3924
rect -23420 3881 -23262 3924
rect -23228 3881 -23212 3941
rect -23662 3866 -23212 3881
rect -23086 3947 -22832 3969
rect -23086 3881 -23070 3947
rect -23036 3881 -22878 3947
rect -23086 3845 -22878 3881
rect -22844 3845 -22832 3947
rect -23086 3822 -22832 3845
rect -22656 3767 -22498 4418
rect -22431 4552 -22256 4559
rect -22431 4366 -22416 4552
rect -22230 4366 -22224 4552
rect -21815 4549 -21726 6595
rect -15022 6556 1484 6664
rect -15130 6550 -15022 6556
rect -19318 6376 -19312 6448
rect -19240 6376 -19234 6448
rect -19312 4575 -19240 6376
rect -18534 6279 -18528 6368
rect -18439 6279 -18433 6368
rect -22680 3766 -22488 3767
rect -23879 3628 -23764 3647
rect -24825 3549 -23995 3587
rect -24825 3409 -24791 3549
rect -24197 3494 -23995 3549
rect -23879 3560 -23862 3628
rect -23782 3560 -23764 3628
rect -24197 3457 -23953 3494
rect -24197 3409 -24029 3457
rect -24825 3402 -24029 3409
rect -23964 3402 -23953 3457
rect -24825 3378 -23953 3402
rect -23879 3463 -23764 3560
rect -23694 3629 -22905 3647
rect -23694 3576 -23662 3629
rect -23548 3621 -22905 3629
rect -23548 3576 -23075 3621
rect -23694 3568 -23075 3576
rect -22942 3568 -22905 3621
rect -23694 3548 -22905 3568
rect -22680 3624 -22637 3766
rect -22517 3624 -22488 3766
rect -22680 3547 -22488 3624
rect -22431 3508 -22256 4366
rect -21823 3991 -21714 4549
rect -20751 4517 -19541 4545
rect -20751 4445 -20709 4517
rect -19587 4445 -19541 4517
rect -20751 4411 -19541 4445
rect -20751 4339 -20497 4411
rect -20751 4237 -20739 4339
rect -20705 4237 -20547 4339
rect -20513 4237 -20497 4339
rect -20751 4219 -20497 4237
rect -20371 4340 -19921 4366
rect -20371 4339 -19971 4340
rect -20371 4237 -20355 4339
rect -20321 4237 -20163 4339
rect -20129 4238 -19971 4339
rect -19937 4238 -19921 4340
rect -20129 4237 -19921 4238
rect -20371 4219 -19921 4237
rect -19795 4342 -19541 4411
rect -19795 4240 -19779 4342
rect -19745 4240 -19587 4342
rect -19553 4240 -19541 4342
rect -19795 4219 -19541 4240
rect -20659 4156 -19633 4181
rect -20659 4155 -20451 4156
rect -20659 4031 -20643 4155
rect -20609 4032 -20451 4155
rect -20417 4032 -20259 4156
rect -20225 4032 -20067 4156
rect -20033 4032 -19875 4156
rect -19841 4032 -19683 4156
rect -19649 4032 -19633 4156
rect -20609 4031 -19633 4032
rect -20659 4002 -19633 4031
rect -21829 3987 -21708 3991
rect -21829 3876 -21823 3987
rect -21714 3876 -21708 3987
rect -21829 3870 -21708 3876
rect -20751 3948 -20497 3969
rect -20751 3881 -20739 3948
rect -20705 3881 -20547 3948
rect -20513 3881 -20497 3948
rect -20751 3822 -20497 3881
rect -20371 3941 -19921 3958
rect -20371 3881 -20355 3941
rect -20321 3924 -19971 3941
rect -20321 3881 -20163 3924
rect -20129 3881 -19971 3924
rect -19937 3881 -19921 3941
rect -20371 3866 -19921 3881
rect -19795 3947 -19541 3969
rect -19795 3881 -19779 3947
rect -19745 3881 -19587 3947
rect -19795 3845 -19587 3881
rect -19553 3845 -19541 3947
rect -19795 3822 -19541 3845
rect -19365 3767 -19207 4575
rect -18528 4560 -18439 6279
rect -16025 6124 -16019 6196
rect -15947 6124 -15941 6196
rect -16019 4575 -15947 6124
rect -15236 5884 -15230 5973
rect -15141 5884 -15135 5973
rect -19140 4553 -18949 4559
rect -19140 4372 -19130 4553
rect -19140 4366 -18949 4372
rect -19389 3766 -19197 3767
rect -20588 3628 -20473 3647
rect -22891 3463 -22256 3508
rect -23879 3377 -22256 3463
rect -21534 3549 -20704 3587
rect -21534 3409 -21500 3549
rect -20906 3494 -20704 3549
rect -20588 3560 -20571 3628
rect -20491 3560 -20473 3628
rect -20906 3457 -20662 3494
rect -20906 3409 -20738 3457
rect -21534 3402 -20738 3409
rect -20673 3402 -20662 3457
rect -21534 3378 -20662 3402
rect -20588 3463 -20473 3560
rect -20403 3629 -19614 3647
rect -20403 3576 -20371 3629
rect -20257 3621 -19614 3629
rect -20257 3576 -19784 3621
rect -20403 3568 -19784 3576
rect -19651 3568 -19614 3621
rect -20403 3548 -19614 3568
rect -19389 3624 -19346 3766
rect -19226 3624 -19197 3766
rect -19389 3547 -19197 3624
rect -19140 3508 -18965 4366
rect -18532 3998 -18423 4560
rect -17460 4517 -16250 4545
rect -17460 4445 -17418 4517
rect -16296 4445 -16250 4517
rect -17460 4411 -16250 4445
rect -17460 4339 -17206 4411
rect -17460 4237 -17448 4339
rect -17414 4237 -17256 4339
rect -17222 4237 -17206 4339
rect -17460 4219 -17206 4237
rect -17080 4340 -16630 4366
rect -17080 4339 -16680 4340
rect -17080 4237 -17064 4339
rect -17030 4237 -16872 4339
rect -16838 4238 -16680 4339
rect -16646 4238 -16630 4340
rect -16838 4237 -16630 4238
rect -17080 4219 -16630 4237
rect -16504 4342 -16250 4411
rect -16504 4240 -16488 4342
rect -16454 4240 -16296 4342
rect -16262 4240 -16250 4342
rect -16504 4219 -16250 4240
rect -17368 4156 -16342 4181
rect -17368 4155 -17160 4156
rect -17368 4031 -17352 4155
rect -17318 4032 -17160 4155
rect -17126 4032 -16968 4156
rect -16934 4032 -16776 4156
rect -16742 4032 -16584 4156
rect -16550 4032 -16392 4156
rect -16358 4032 -16342 4156
rect -17318 4031 -16342 4032
rect -17368 4002 -16342 4031
rect -18532 3881 -18423 3887
rect -17460 3948 -17206 3969
rect -17460 3881 -17448 3948
rect -17414 3881 -17256 3948
rect -17222 3881 -17206 3948
rect -17460 3822 -17206 3881
rect -17080 3941 -16630 3958
rect -17080 3881 -17064 3941
rect -17030 3924 -16680 3941
rect -17030 3881 -16872 3924
rect -16838 3881 -16680 3924
rect -16646 3881 -16630 3941
rect -17080 3866 -16630 3881
rect -16504 3947 -16250 3969
rect -16504 3881 -16488 3947
rect -16454 3881 -16296 3947
rect -16504 3845 -16296 3881
rect -16262 3845 -16250 3947
rect -16504 3822 -16250 3845
rect -16074 3767 -15916 4575
rect -15230 4571 -15141 5884
rect -12748 5681 -12742 5753
rect -12670 5681 -12664 5753
rect -12742 4575 -12670 5681
rect -11946 5537 -11940 5626
rect -11851 5537 -11845 5626
rect -15849 4556 -15674 4559
rect -15849 4378 -15826 4556
rect -15648 4378 -15642 4556
rect -16098 3766 -15906 3767
rect -17297 3628 -17182 3647
rect -19600 3463 -18965 3508
rect -20588 3377 -18965 3463
rect -18243 3549 -17413 3587
rect -18243 3409 -18209 3549
rect -17615 3494 -17413 3549
rect -17297 3560 -17280 3628
rect -17200 3560 -17182 3628
rect -17615 3457 -17371 3494
rect -17615 3409 -17447 3457
rect -18243 3402 -17447 3409
rect -17382 3402 -17371 3457
rect -18243 3378 -17371 3402
rect -17297 3463 -17182 3560
rect -17112 3629 -16323 3647
rect -17112 3576 -17080 3629
rect -16966 3621 -16323 3629
rect -16966 3576 -16493 3621
rect -17112 3568 -16493 3576
rect -16360 3568 -16323 3621
rect -17112 3548 -16323 3568
rect -16098 3624 -16055 3766
rect -15935 3624 -15906 3766
rect -16098 3547 -15906 3624
rect -15849 3508 -15674 4378
rect -15241 4006 -15132 4571
rect -14169 4517 -12959 4545
rect -14169 4445 -14127 4517
rect -13005 4445 -12959 4517
rect -14169 4411 -12959 4445
rect -14169 4339 -13915 4411
rect -14169 4237 -14157 4339
rect -14123 4237 -13965 4339
rect -13931 4237 -13915 4339
rect -14169 4219 -13915 4237
rect -13789 4340 -13339 4366
rect -13789 4339 -13389 4340
rect -13789 4237 -13773 4339
rect -13739 4237 -13581 4339
rect -13547 4238 -13389 4339
rect -13355 4238 -13339 4340
rect -13547 4237 -13339 4238
rect -13789 4219 -13339 4237
rect -13213 4342 -12959 4411
rect -13213 4240 -13197 4342
rect -13163 4240 -13005 4342
rect -12971 4240 -12959 4342
rect -13213 4219 -12959 4240
rect -14077 4156 -13051 4181
rect -14077 4155 -13869 4156
rect -14077 4031 -14061 4155
rect -14027 4032 -13869 4155
rect -13835 4032 -13677 4156
rect -13643 4032 -13485 4156
rect -13451 4032 -13293 4156
rect -13259 4032 -13101 4156
rect -13067 4032 -13051 4156
rect -14027 4031 -13051 4032
rect -15247 4002 -15126 4006
rect -14077 4002 -13051 4031
rect -15247 3891 -15241 4002
rect -15132 3891 -15126 4002
rect -15247 3885 -15126 3891
rect -14169 3948 -13915 3969
rect -14169 3881 -14157 3948
rect -14123 3881 -13965 3948
rect -13931 3881 -13915 3948
rect -14169 3822 -13915 3881
rect -13789 3941 -13339 3958
rect -13789 3881 -13773 3941
rect -13739 3924 -13389 3941
rect -13739 3881 -13581 3924
rect -13547 3881 -13389 3924
rect -13355 3881 -13339 3941
rect -13789 3866 -13339 3881
rect -13213 3947 -12959 3969
rect -13213 3881 -13197 3947
rect -13163 3881 -13005 3947
rect -13213 3845 -13005 3881
rect -12971 3845 -12959 3947
rect -13213 3822 -12959 3845
rect -12783 3767 -12625 4575
rect -12555 4559 -12549 4562
rect -12558 4387 -12549 4559
rect -12374 4387 -12368 4562
rect -11940 4560 -11851 5537
rect -9445 5385 -9439 5457
rect -9367 5385 -9361 5457
rect -9439 4575 -9367 5385
rect -6173 5339 -6084 5346
rect -8646 5227 -8640 5316
rect -8551 5227 -8545 5316
rect -6173 5269 -6166 5339
rect -6096 5269 -6084 5339
rect -6173 5261 -6084 5269
rect -12807 3766 -12615 3767
rect -14006 3628 -13891 3647
rect -16309 3463 -15674 3508
rect -17297 3377 -15674 3463
rect -14952 3549 -14122 3587
rect -14952 3409 -14918 3549
rect -14324 3494 -14122 3549
rect -14006 3560 -13989 3628
rect -13909 3560 -13891 3628
rect -14324 3457 -14080 3494
rect -14324 3409 -14156 3457
rect -14952 3402 -14156 3409
rect -14091 3402 -14080 3457
rect -14952 3378 -14080 3402
rect -14006 3463 -13891 3560
rect -13821 3629 -13032 3647
rect -13821 3576 -13789 3629
rect -13675 3621 -13032 3629
rect -13675 3576 -13202 3621
rect -13821 3568 -13202 3576
rect -13069 3568 -13032 3621
rect -13821 3548 -13032 3568
rect -12807 3624 -12764 3766
rect -12644 3624 -12615 3766
rect -12807 3547 -12615 3624
rect -12558 3508 -12383 4387
rect -11950 3995 -11841 4560
rect -10878 4517 -9668 4545
rect -10878 4445 -10836 4517
rect -9714 4445 -9668 4517
rect -10878 4411 -9668 4445
rect -10878 4339 -10624 4411
rect -10878 4237 -10866 4339
rect -10832 4237 -10674 4339
rect -10640 4237 -10624 4339
rect -10878 4219 -10624 4237
rect -10498 4340 -10048 4366
rect -10498 4339 -10098 4340
rect -10498 4237 -10482 4339
rect -10448 4237 -10290 4339
rect -10256 4238 -10098 4339
rect -10064 4238 -10048 4340
rect -10256 4237 -10048 4238
rect -10498 4219 -10048 4237
rect -9922 4342 -9668 4411
rect -9922 4240 -9906 4342
rect -9872 4240 -9714 4342
rect -9680 4240 -9668 4342
rect -9922 4219 -9668 4240
rect -10786 4156 -9760 4181
rect -10786 4155 -10578 4156
rect -10786 4031 -10770 4155
rect -10736 4032 -10578 4155
rect -10544 4032 -10386 4156
rect -10352 4032 -10194 4156
rect -10160 4032 -10002 4156
rect -9968 4032 -9810 4156
rect -9776 4032 -9760 4156
rect -10736 4031 -9760 4032
rect -10786 4002 -9760 4031
rect -11956 3991 -11835 3995
rect -11956 3880 -11950 3991
rect -11841 3880 -11835 3991
rect -11956 3874 -11835 3880
rect -10878 3948 -10624 3969
rect -10878 3881 -10866 3948
rect -10832 3881 -10674 3948
rect -10640 3881 -10624 3948
rect -10878 3822 -10624 3881
rect -10498 3941 -10048 3958
rect -10498 3881 -10482 3941
rect -10448 3924 -10098 3941
rect -10448 3881 -10290 3924
rect -10256 3881 -10098 3924
rect -10064 3881 -10048 3941
rect -10498 3866 -10048 3881
rect -9922 3947 -9668 3969
rect -9922 3881 -9906 3947
rect -9872 3881 -9714 3947
rect -9922 3845 -9714 3881
rect -9680 3845 -9668 3947
rect -9922 3822 -9668 3845
rect -9492 3767 -9334 4575
rect -8640 4565 -8551 5227
rect -6166 4575 -6096 5261
rect 1376 5232 1484 6556
rect 1581 6318 1670 6877
rect 1565 5925 1674 6318
rect 1795 6241 3005 6269
rect 1795 6169 1841 6241
rect 2963 6169 3005 6241
rect 1795 6135 3005 6169
rect 1795 6066 2049 6135
rect 1795 5964 1807 6066
rect 1841 5964 1999 6066
rect 2033 5964 2049 6066
rect 1795 5943 2049 5964
rect 2175 6064 2625 6090
rect 2175 5962 2191 6064
rect 2225 6063 2625 6064
rect 2225 5962 2383 6063
rect 2175 5961 2383 5962
rect 2417 5961 2575 6063
rect 2609 5961 2625 6063
rect 2175 5943 2625 5961
rect 2751 6063 3005 6135
rect 2751 5961 2767 6063
rect 2801 5961 2959 6063
rect 2993 5961 3005 6063
rect 2751 5943 3005 5961
rect 1565 5501 1674 5813
rect 1887 5880 2913 5905
rect 1887 5756 1903 5880
rect 1937 5756 2095 5880
rect 2129 5756 2287 5880
rect 2321 5756 2479 5880
rect 2513 5756 2671 5880
rect 2705 5879 2913 5880
rect 2705 5756 2863 5879
rect 1887 5755 2863 5756
rect 2897 5755 2913 5879
rect 1887 5726 2913 5755
rect 1795 5671 2049 5693
rect 1795 5569 1807 5671
rect 1841 5605 1999 5671
rect 2033 5605 2049 5671
rect 1841 5569 2049 5605
rect 2175 5665 2625 5682
rect 2175 5605 2191 5665
rect 2225 5648 2575 5665
rect 2225 5605 2383 5648
rect 2417 5605 2575 5648
rect 2609 5605 2625 5665
rect 2175 5590 2625 5605
rect 2751 5672 3005 5693
rect 2751 5605 2767 5672
rect 2801 5605 2959 5672
rect 2993 5605 3005 5672
rect 1795 5546 2049 5569
rect 2751 5546 3005 5605
rect 1552 5495 1685 5501
rect 1552 5398 1564 5495
rect 1673 5398 1685 5495
rect 3177 5474 3286 6370
rect 3401 6241 4611 6269
rect 3401 6169 3447 6241
rect 4569 6169 4611 6241
rect 3401 6135 4611 6169
rect 3401 6066 3655 6135
rect 3401 5964 3413 6066
rect 3447 5964 3605 6066
rect 3639 5964 3655 6066
rect 3401 5943 3655 5964
rect 3781 6064 4231 6090
rect 3781 5962 3797 6064
rect 3831 6063 4231 6064
rect 3831 5962 3989 6063
rect 3781 5961 3989 5962
rect 4023 5961 4181 6063
rect 4215 5961 4231 6063
rect 3781 5943 4231 5961
rect 4357 6063 4611 6135
rect 4357 5961 4373 6063
rect 4407 5961 4565 6063
rect 4599 5961 4611 6063
rect 4357 5943 4611 5961
rect 3493 5880 4519 5905
rect 3493 5756 3509 5880
rect 3543 5756 3701 5880
rect 3735 5756 3893 5880
rect 3927 5756 4085 5880
rect 4119 5756 4277 5880
rect 4311 5879 4519 5880
rect 4311 5756 4469 5879
rect 3493 5755 4469 5756
rect 4503 5755 4519 5879
rect 3493 5726 4519 5755
rect 3401 5671 3655 5693
rect 3401 5569 3413 5671
rect 3447 5605 3605 5671
rect 3639 5605 3655 5671
rect 3447 5569 3655 5605
rect 3781 5665 4231 5682
rect 3781 5605 3797 5665
rect 3831 5648 4181 5665
rect 3831 5605 3989 5648
rect 4023 5605 4181 5648
rect 4215 5605 4231 5665
rect 3781 5590 4231 5605
rect 4357 5672 4611 5693
rect 4357 5605 4373 5672
rect 4407 5605 4565 5672
rect 4599 5605 4611 5672
rect 3401 5546 3655 5569
rect 4357 5546 4611 5605
rect 4729 5541 4821 6348
rect 4861 5924 4970 6348
rect 5105 6265 6315 6267
rect 5105 6239 8026 6265
rect 5105 6167 5151 6239
rect 6273 6167 8026 6239
rect 5105 6133 8026 6167
rect 5105 6064 5359 6133
rect 5105 5962 5117 6064
rect 5151 5962 5309 6064
rect 5343 5962 5359 6064
rect 5105 5941 5359 5962
rect 5485 6062 5935 6088
rect 5485 5960 5501 6062
rect 5535 6061 5935 6062
rect 5535 5960 5693 6061
rect 5485 5959 5693 5960
rect 5727 5959 5885 6061
rect 5919 5959 5935 6061
rect 5485 5941 5935 5959
rect 6061 6061 8026 6133
rect 6061 5959 6077 6061
rect 6111 5959 6269 6061
rect 6303 5959 8026 6061
rect 6061 5944 8026 5959
rect 6061 5941 6315 5944
rect 4861 5815 4873 5924
rect 4861 5619 4970 5815
rect 5197 5878 6223 5903
rect 5197 5754 5213 5878
rect 5247 5754 5405 5878
rect 5439 5754 5597 5878
rect 5631 5754 5789 5878
rect 5823 5754 5981 5878
rect 6015 5877 6223 5878
rect 6015 5754 6173 5877
rect 5197 5753 6173 5754
rect 6207 5753 6223 5877
rect 5197 5724 6223 5753
rect 5105 5669 5359 5691
rect 1552 5392 1685 5398
rect 3165 5468 3298 5474
rect 3165 5371 3177 5468
rect 3286 5371 3298 5468
rect 4729 5472 4738 5541
rect 4807 5472 4821 5541
rect 4849 5613 4982 5619
rect 4849 5516 4861 5613
rect 4970 5516 4982 5613
rect 5105 5567 5117 5669
rect 5151 5603 5309 5669
rect 5343 5603 5359 5669
rect 5151 5567 5359 5603
rect 5485 5663 5935 5680
rect 5485 5603 5501 5663
rect 5535 5646 5885 5663
rect 5535 5603 5693 5646
rect 5727 5603 5885 5646
rect 5919 5603 5935 5663
rect 5485 5588 5935 5603
rect 6061 5670 6315 5691
rect 6061 5603 6077 5670
rect 6111 5603 6269 5670
rect 6303 5603 6315 5670
rect 5105 5544 5359 5567
rect 6061 5544 6315 5603
rect 7100 5561 8023 5944
rect 6938 5554 8023 5561
rect 4849 5510 4982 5516
rect 4729 5438 4821 5472
rect 6938 5507 6967 5554
rect 7536 5544 8023 5554
rect 7536 5507 7572 5544
rect 6938 5441 7572 5507
rect 7804 5531 8023 5544
rect 7804 5497 7872 5531
rect 7963 5497 8023 5531
rect 7804 5476 8023 5497
rect 7809 5459 8023 5476
rect 6938 5435 7573 5441
rect 1868 5353 2657 5371
rect 1868 5345 2511 5353
rect 1868 5292 1905 5345
rect 2038 5300 2511 5345
rect 2625 5300 2657 5353
rect 2038 5292 2657 5300
rect 1868 5272 2657 5292
rect 2727 5352 2842 5371
rect 3165 5365 3298 5371
rect 2727 5284 2745 5352
rect 2825 5284 2842 5352
rect 3474 5353 4263 5371
rect 3474 5345 4117 5353
rect 1358 5187 1854 5232
rect 2727 5187 2842 5284
rect 2958 5232 3129 5311
rect 3474 5292 3511 5345
rect 3644 5300 4117 5345
rect 4231 5300 4263 5353
rect 3644 5292 4263 5300
rect 3474 5272 4263 5292
rect 4333 5352 4448 5371
rect 4333 5284 4351 5352
rect 4431 5284 4448 5352
rect 5178 5351 5967 5369
rect 5178 5343 5821 5351
rect 2958 5218 3460 5232
rect 1358 5101 2842 5187
rect 2916 5187 3460 5218
rect 4333 5187 4448 5284
rect 4564 5218 4735 5311
rect 5178 5290 5215 5343
rect 5348 5298 5821 5343
rect 5935 5298 5967 5351
rect 5348 5290 5967 5298
rect 5178 5270 5967 5290
rect 6037 5350 6152 5369
rect 6037 5282 6055 5350
rect 6135 5282 6152 5350
rect 6938 5355 6951 5435
rect 6985 5355 7143 5435
rect 7177 5355 7335 5435
rect 7369 5355 7527 5435
rect 7561 5355 7573 5435
rect 6938 5349 7573 5355
rect 7709 5411 7778 5427
rect 6938 5348 7572 5349
rect 7709 5320 7728 5411
rect 7599 5319 7728 5320
rect 7031 5313 7728 5319
rect 2916 5181 4448 5187
rect 2916 5126 2927 5181
rect 2992 5126 4448 5181
rect 2916 5102 4448 5126
rect 4522 5181 4735 5218
rect 4522 5126 4533 5181
rect 4598 5159 4735 5181
rect 4598 5126 4826 5159
rect 4522 5102 4826 5126
rect 3026 5101 4448 5102
rect 1358 5089 1854 5101
rect 3026 5089 3460 5101
rect -5357 4991 -5351 5080
rect -5262 4991 -5256 5080
rect 1800 5032 1855 5048
rect -9267 4429 -9092 4559
rect -9516 3766 -9324 3767
rect -10715 3628 -10600 3647
rect -13018 3463 -12383 3508
rect -14006 3377 -12383 3463
rect -11661 3549 -10831 3587
rect -11661 3409 -11627 3549
rect -11033 3494 -10831 3549
rect -10715 3560 -10698 3628
rect -10618 3560 -10600 3628
rect -11033 3457 -10789 3494
rect -11033 3409 -10865 3457
rect -11661 3402 -10865 3409
rect -10800 3402 -10789 3457
rect -11661 3378 -10789 3402
rect -10715 3463 -10600 3560
rect -10530 3629 -9741 3647
rect -10530 3576 -10498 3629
rect -10384 3621 -9741 3629
rect -10384 3576 -9911 3621
rect -10530 3568 -9911 3576
rect -9778 3568 -9741 3621
rect -10530 3548 -9741 3568
rect -9516 3624 -9473 3766
rect -9353 3624 -9324 3766
rect -9516 3547 -9324 3624
rect -9267 3508 -9092 4252
rect -8660 4015 -8551 4565
rect -7588 4517 -6378 4545
rect -7588 4445 -7546 4517
rect -6424 4445 -6378 4517
rect -7588 4411 -6378 4445
rect -7588 4339 -7334 4411
rect -7588 4237 -7576 4339
rect -7542 4237 -7384 4339
rect -7350 4237 -7334 4339
rect -7588 4219 -7334 4237
rect -7208 4340 -6758 4366
rect -7208 4339 -6808 4340
rect -7208 4237 -7192 4339
rect -7158 4237 -7000 4339
rect -6966 4238 -6808 4339
rect -6774 4238 -6758 4340
rect -6966 4237 -6758 4238
rect -7208 4219 -6758 4237
rect -6632 4342 -6378 4411
rect -6632 4240 -6616 4342
rect -6582 4240 -6424 4342
rect -6390 4240 -6378 4342
rect -6632 4219 -6378 4240
rect -7496 4156 -6470 4181
rect -7496 4155 -7288 4156
rect -7496 4031 -7480 4155
rect -7446 4032 -7288 4155
rect -7254 4032 -7096 4156
rect -7062 4032 -6904 4156
rect -6870 4032 -6712 4156
rect -6678 4032 -6520 4156
rect -6486 4032 -6470 4156
rect -7446 4031 -6470 4032
rect -8666 4009 -8545 4015
rect -8666 3900 -8660 4009
rect -8551 3900 -8545 4009
rect -7496 4002 -6470 4031
rect -8666 3894 -8545 3900
rect -7588 3948 -7334 3969
rect -7588 3881 -7576 3948
rect -7542 3881 -7384 3948
rect -7350 3881 -7334 3948
rect -7588 3822 -7334 3881
rect -7208 3941 -6758 3958
rect -7208 3881 -7192 3941
rect -7158 3924 -6808 3941
rect -7158 3881 -7000 3924
rect -6966 3881 -6808 3924
rect -6774 3881 -6758 3941
rect -7208 3866 -6758 3881
rect -6632 3947 -6378 3969
rect -6632 3881 -6616 3947
rect -6582 3881 -6424 3947
rect -6632 3845 -6424 3881
rect -6390 3845 -6378 3947
rect -6632 3822 -6378 3845
rect -6202 3767 -6044 4575
rect -5984 4395 -5978 4570
rect -5803 4395 -5797 4570
rect -5351 4563 -5262 4991
rect 1800 4926 1807 5032
rect 1841 4926 1855 5032
rect 1887 5047 2337 5059
rect 1887 5013 1903 5047
rect 1937 5013 2095 5047
rect 2129 5046 2337 5047
rect 2129 5013 2287 5046
rect 1887 5012 2287 5013
rect 2321 5012 2337 5046
rect 1887 4991 2337 5012
rect 2463 5047 2913 5059
rect 2463 5013 2479 5047
rect 2513 5013 2671 5047
rect 2705 5013 2863 5047
rect 2897 5013 2913 5047
rect 2463 4991 2913 5013
rect 2947 5032 3002 5048
rect 1800 4860 1855 4926
rect 1985 4946 2050 4963
rect 1985 4912 1999 4946
rect 2033 4912 2050 4946
rect 1985 4860 2050 4912
rect 2178 4946 2625 4958
rect 2178 4912 2191 4946
rect 2225 4912 2383 4946
rect 2417 4912 2575 4946
rect 2609 4912 2625 4946
rect 2178 4894 2625 4912
rect 2751 4946 2816 4962
rect 2751 4912 2767 4946
rect 2801 4912 2816 4946
rect 2751 4860 2816 4912
rect 2947 4926 2959 5032
rect 2993 4926 3002 5032
rect 2947 4860 3002 4926
rect 1800 4849 3002 4860
rect 1800 4838 2301 4849
rect 2361 4838 3002 4849
rect -2881 4746 -2875 4818
rect -2803 4746 -2797 4818
rect 1800 4792 1841 4838
rect 2964 4792 3002 4838
rect 1800 4789 2301 4792
rect 2361 4789 3002 4792
rect 1800 4769 3002 4789
rect 3406 5032 3461 5048
rect 3406 4926 3413 5032
rect 3447 4926 3461 5032
rect 3493 5047 3943 5059
rect 3493 5013 3509 5047
rect 3543 5013 3701 5047
rect 3735 5046 3943 5047
rect 3735 5013 3893 5046
rect 3493 5012 3893 5013
rect 3927 5012 3943 5046
rect 3493 4991 3943 5012
rect 4069 5047 4519 5059
rect 4069 5013 4085 5047
rect 4119 5013 4277 5047
rect 4311 5013 4469 5047
rect 4503 5013 4519 5047
rect 4069 4991 4519 5013
rect 4553 5032 4608 5048
rect 3406 4860 3461 4926
rect 3591 4946 3656 4963
rect 3591 4912 3605 4946
rect 3639 4912 3656 4946
rect 3591 4860 3656 4912
rect 3784 4946 4231 4958
rect 3784 4912 3797 4946
rect 3831 4912 3989 4946
rect 4023 4912 4181 4946
rect 4215 4912 4231 4946
rect 3784 4894 4231 4912
rect 4357 4946 4422 4962
rect 4357 4912 4373 4946
rect 4407 4912 4422 4946
rect 4357 4860 4422 4912
rect 4553 4926 4565 5032
rect 4599 4926 4608 5032
rect 4553 4860 4608 4926
rect 3406 4849 4608 4860
rect 3406 4838 3907 4849
rect 3967 4838 4608 4849
rect 3406 4792 3447 4838
rect 4570 4792 4608 4838
rect 3406 4789 3907 4792
rect 3967 4789 4608 4792
rect 3406 4769 4608 4789
rect -2875 4579 -2803 4746
rect 419 4612 425 4684
rect 497 4612 503 4684
rect -2908 4575 -2758 4579
rect 425 4575 497 4612
rect 4689 4583 4826 5102
rect 4953 5087 4959 5230
rect 5028 5185 5164 5230
rect 6037 5185 6152 5282
rect 6268 5236 6439 5309
rect 6268 5216 6755 5236
rect 7031 5233 7047 5313
rect 7081 5233 7239 5313
rect 7273 5233 7431 5313
rect 7465 5233 7728 5313
rect 7031 5227 7728 5233
rect 5028 5099 6152 5185
rect 6226 5179 6755 5216
rect 6226 5124 6237 5179
rect 6302 5177 6755 5179
rect 6903 5180 7067 5198
rect 6903 5177 7017 5180
rect 6302 5145 7017 5177
rect 7051 5145 7067 5180
rect 6302 5124 7067 5145
rect 6226 5122 7067 5124
rect 6226 5100 6439 5122
rect 5028 5087 5164 5099
rect 6641 5063 7067 5122
rect 7095 5180 7355 5199
rect 7095 5145 7306 5180
rect 7340 5145 7355 5180
rect 7095 5125 7355 5145
rect 7431 5185 7728 5227
rect 7762 5185 7778 5411
rect 7809 5425 7815 5459
rect 7894 5455 8023 5459
rect 7894 5425 7900 5455
rect 7809 5267 7900 5425
rect 7809 5233 7815 5267
rect 7894 5233 7900 5267
rect 7809 5217 7900 5233
rect 7932 5363 8121 5427
rect 7932 5329 7938 5363
rect 8015 5329 8121 5363
rect 5110 5030 5165 5046
rect 5110 4924 5117 5030
rect 5151 4924 5165 5030
rect 5197 5045 5647 5057
rect 5197 5011 5213 5045
rect 5247 5011 5405 5045
rect 5439 5044 5647 5045
rect 5439 5011 5597 5044
rect 5197 5010 5597 5011
rect 5631 5010 5647 5044
rect 5197 4989 5647 5010
rect 5773 5045 6223 5057
rect 7095 5056 7145 5125
rect 7431 5097 7778 5185
rect 7932 5171 8121 5329
rect 5773 5011 5789 5045
rect 5823 5011 5981 5045
rect 6015 5011 6173 5045
rect 6207 5011 6223 5045
rect 5773 4989 6223 5011
rect 6257 5030 6312 5046
rect 7095 5034 7101 5056
rect 5110 4858 5165 4924
rect 5295 4944 5360 4961
rect 5295 4910 5309 4944
rect 5343 4910 5360 4944
rect 5295 4858 5360 4910
rect 5488 4944 5935 4956
rect 5488 4910 5501 4944
rect 5535 4910 5693 4944
rect 5727 4910 5885 4944
rect 5919 4910 5935 4944
rect 5488 4892 5935 4910
rect 6061 4944 6126 4960
rect 6061 4910 6077 4944
rect 6111 4910 6126 4944
rect 6061 4858 6126 4910
rect 6257 4924 6269 5030
rect 6303 4924 6312 5030
rect 6257 4858 6312 4924
rect 5110 4847 6312 4858
rect 5110 4836 5611 4847
rect 5671 4836 6312 4847
rect 5110 4790 5151 4836
rect 6274 4790 6312 4836
rect 5110 4787 5611 4790
rect 5671 4787 6312 4790
rect 5110 4767 6312 4787
rect 6903 5021 7101 5034
rect 7135 5021 7145 5056
rect 7173 5085 7778 5097
rect 7173 5051 7185 5085
rect 7561 5051 7778 5085
rect 7173 5046 7778 5051
rect 7173 5045 7609 5046
rect 6903 4898 7145 5021
rect 7709 4965 7778 5046
rect 7809 5137 7938 5171
rect 8015 5137 8121 5171
rect 7809 5009 8121 5137
rect 7809 4975 7821 5009
rect 7997 4975 8121 5009
rect 7809 4969 8009 4975
rect 7709 4931 7728 4965
rect 7762 4931 7778 4965
rect 7709 4914 7778 4931
rect 7809 4921 8009 4928
rect 6903 4583 7039 4898
rect 7173 4893 7573 4899
rect 7173 4859 7185 4893
rect 7561 4859 7573 4893
rect 7173 4821 7573 4859
rect 7173 4787 7200 4821
rect 7535 4787 7573 4821
rect 7173 4776 7323 4787
rect 7314 4693 7323 4776
rect 7433 4776 7573 4787
rect 7809 4887 7821 4921
rect 7997 4887 8009 4921
rect 8037 4914 8121 4975
rect 7809 4819 8009 4887
rect 7809 4802 7840 4819
rect 7809 4778 7810 4802
rect 7972 4785 8009 4819
rect 7433 4693 7441 4776
rect 7314 4684 7441 4693
rect 7919 4778 8009 4785
rect 7810 4687 7919 4693
rect -6226 3766 -6034 3767
rect -7425 3628 -7310 3647
rect -9727 3463 -9092 3508
rect -10715 3377 -9092 3463
rect -8371 3549 -7541 3587
rect -8371 3409 -8337 3549
rect -7743 3494 -7541 3549
rect -7425 3560 -7408 3628
rect -7328 3560 -7310 3628
rect -7743 3457 -7499 3494
rect -7743 3409 -7575 3457
rect -8371 3402 -7575 3409
rect -7510 3402 -7499 3457
rect -8371 3378 -7499 3402
rect -7425 3463 -7310 3560
rect -7240 3629 -6451 3647
rect -7240 3576 -7208 3629
rect -7094 3621 -6451 3629
rect -7094 3576 -6621 3621
rect -7240 3568 -6621 3576
rect -6488 3568 -6451 3621
rect -7240 3548 -6451 3568
rect -6226 3624 -6183 3766
rect -6063 3624 -6034 3766
rect -6226 3547 -6034 3624
rect -5977 3508 -5802 4395
rect -5369 4015 -5260 4563
rect -4297 4517 -3087 4545
rect -4297 4445 -4255 4517
rect -3133 4445 -3087 4517
rect -4297 4411 -3087 4445
rect -4297 4339 -4043 4411
rect -4297 4237 -4285 4339
rect -4251 4237 -4093 4339
rect -4059 4237 -4043 4339
rect -4297 4219 -4043 4237
rect -3917 4340 -3467 4366
rect -3917 4339 -3517 4340
rect -3917 4237 -3901 4339
rect -3867 4237 -3709 4339
rect -3675 4238 -3517 4339
rect -3483 4238 -3467 4340
rect -3675 4237 -3467 4238
rect -3917 4219 -3467 4237
rect -3341 4342 -3087 4411
rect -3341 4240 -3325 4342
rect -3291 4240 -3133 4342
rect -3099 4240 -3087 4342
rect -3341 4219 -3087 4240
rect -4205 4156 -3179 4181
rect -4205 4155 -3997 4156
rect -4205 4031 -4189 4155
rect -4155 4032 -3997 4155
rect -3963 4032 -3805 4156
rect -3771 4032 -3613 4156
rect -3579 4032 -3421 4156
rect -3387 4032 -3229 4156
rect -3195 4032 -3179 4156
rect -4155 4031 -3179 4032
rect -5375 4009 -5254 4015
rect -5375 3900 -5369 4009
rect -5260 3900 -5254 4009
rect -4205 4002 -3179 4031
rect -5375 3894 -5254 3900
rect -4297 3948 -4043 3969
rect -4297 3881 -4285 3948
rect -4251 3881 -4093 3948
rect -4059 3881 -4043 3948
rect -4297 3822 -4043 3881
rect -3917 3941 -3467 3958
rect -3917 3881 -3901 3941
rect -3867 3924 -3517 3941
rect -3867 3881 -3709 3924
rect -3675 3881 -3517 3924
rect -3483 3881 -3467 3941
rect -3917 3866 -3467 3881
rect -3341 3947 -3087 3969
rect -3341 3881 -3325 3947
rect -3291 3881 -3133 3947
rect -3341 3845 -3133 3881
rect -3099 3845 -3087 3947
rect -3341 3822 -3087 3845
rect -2911 3767 -2753 4575
rect -2691 4558 -2503 4564
rect -2064 4560 -2058 4562
rect -2691 4383 -2683 4558
rect -2508 4383 -2503 4558
rect -2691 4376 -2503 4383
rect -2078 4473 -2058 4560
rect -1969 4473 -1963 4562
rect -1006 4517 204 4545
rect -2935 3766 -2743 3767
rect -4134 3628 -4019 3647
rect -6437 3463 -5802 3508
rect -7425 3377 -5802 3463
rect -5080 3549 -4250 3587
rect -5080 3409 -5046 3549
rect -4452 3494 -4250 3549
rect -4134 3560 -4117 3628
rect -4037 3560 -4019 3628
rect -4452 3457 -4208 3494
rect -4452 3409 -4284 3457
rect -5080 3402 -4284 3409
rect -4219 3402 -4208 3457
rect -5080 3378 -4208 3402
rect -4134 3463 -4019 3560
rect -3949 3629 -3160 3647
rect -3949 3576 -3917 3629
rect -3803 3621 -3160 3629
rect -3803 3576 -3330 3621
rect -3949 3568 -3330 3576
rect -3197 3568 -3160 3621
rect -3949 3548 -3160 3568
rect -2935 3624 -2892 3766
rect -2772 3624 -2743 3766
rect -2935 3547 -2743 3624
rect -2686 3508 -2511 4376
rect -2078 3999 -1969 4473
rect -1006 4445 -964 4517
rect 158 4445 204 4517
rect -1006 4411 204 4445
rect -1006 4339 -752 4411
rect -1006 4237 -994 4339
rect -960 4237 -802 4339
rect -768 4237 -752 4339
rect -1006 4219 -752 4237
rect -626 4340 -176 4366
rect -626 4339 -226 4340
rect -626 4237 -610 4339
rect -576 4237 -418 4339
rect -384 4238 -226 4339
rect -192 4238 -176 4340
rect -384 4237 -176 4238
rect -626 4219 -176 4237
rect -50 4342 204 4411
rect -50 4240 -34 4342
rect 0 4240 158 4342
rect 192 4240 204 4342
rect -50 4219 204 4240
rect -914 4156 112 4181
rect -914 4155 -706 4156
rect -914 4031 -898 4155
rect -864 4032 -706 4155
rect -672 4032 -514 4156
rect -480 4032 -322 4156
rect -288 4032 -130 4156
rect -96 4032 62 4156
rect 96 4032 112 4156
rect -864 4031 112 4032
rect -914 4002 112 4031
rect -2084 3994 -1963 3999
rect -2084 3883 -2078 3994
rect -1969 3883 -1963 3994
rect -2084 3877 -1963 3883
rect -1006 3948 -752 3969
rect -1006 3881 -994 3948
rect -960 3881 -802 3948
rect -768 3881 -752 3948
rect -1006 3822 -752 3881
rect -626 3941 -176 3958
rect -626 3881 -610 3941
rect -576 3924 -226 3941
rect -576 3881 -418 3924
rect -384 3881 -226 3924
rect -192 3881 -176 3941
rect -626 3866 -176 3881
rect -50 3947 204 3969
rect -50 3881 -34 3947
rect 0 3881 158 3947
rect -50 3845 158 3881
rect 192 3845 204 3947
rect -50 3822 204 3845
rect 380 3767 538 4575
rect 605 4549 780 4559
rect 596 4377 602 4549
rect 774 4377 780 4549
rect 4689 4446 7039 4583
rect 605 4238 780 4377
rect 602 4232 780 4238
rect 596 4060 602 4232
rect 774 4060 780 4232
rect 2921 4275 2987 4281
rect 4885 4275 4951 4281
rect 2987 4209 4885 4275
rect 4951 4209 4993 4275
rect 2921 4203 2987 4209
rect 4885 4203 4951 4209
rect 602 4054 780 4060
rect 356 3766 548 3767
rect -843 3628 -728 3647
rect -3146 3463 -2511 3508
rect -4134 3377 -2511 3463
rect -1789 3549 -959 3587
rect -1789 3409 -1755 3549
rect -1161 3494 -959 3549
rect -843 3560 -826 3628
rect -746 3560 -728 3628
rect -1161 3457 -917 3494
rect -1161 3409 -993 3457
rect -1789 3402 -993 3409
rect -928 3402 -917 3457
rect -1789 3378 -917 3402
rect -843 3463 -728 3560
rect -658 3629 131 3647
rect -658 3576 -626 3629
rect -512 3621 131 3629
rect -512 3576 -39 3621
rect -658 3568 -39 3576
rect 94 3568 131 3621
rect -658 3548 131 3568
rect 356 3624 399 3766
rect 519 3624 548 3766
rect 356 3547 548 3624
rect 605 3540 780 4054
rect 5339 4083 5411 4089
rect 5339 3540 5411 4011
rect 5658 3983 7357 4027
rect 5658 3949 5721 3983
rect 5812 3949 6161 3983
rect 6252 3949 6601 3983
rect 6692 3949 7357 3983
rect 5658 3937 7357 3949
rect 5658 3911 5872 3937
rect 605 3508 5411 3540
rect 145 3463 5411 3508
rect -843 3377 5411 3463
rect -22891 3365 -22256 3377
rect -19600 3365 -18965 3377
rect -16309 3365 -15674 3377
rect -13018 3365 -12383 3377
rect -9727 3365 -9092 3377
rect -6437 3365 -5802 3377
rect -3146 3365 -2511 3377
rect 145 3365 5411 3377
rect 5558 3879 5627 3885
rect 5558 3637 5577 3810
rect 5611 3637 5627 3810
rect 5658 3877 5664 3911
rect 5743 3907 5872 3911
rect 6098 3911 6312 3937
rect 5743 3877 5749 3907
rect 5998 3879 6067 3885
rect 5658 3719 5749 3877
rect 5658 3685 5664 3719
rect 5743 3685 5749 3719
rect 5658 3669 5749 3685
rect 5781 3815 5970 3879
rect 5781 3781 5787 3815
rect 5864 3781 5970 3815
rect 5558 3535 5627 3637
rect 5781 3623 5970 3781
rect 5658 3589 5787 3623
rect 5864 3589 5970 3623
rect 5558 3417 5628 3535
rect 5658 3461 5970 3589
rect 5658 3427 5670 3461
rect 5846 3427 5970 3461
rect 5658 3421 5858 3427
rect 5558 3383 5577 3417
rect 5611 3383 5628 3417
rect 5558 3366 5628 3383
rect -24039 3308 -23984 3324
rect -24039 3202 -24030 3308
rect -23996 3202 -23984 3308
rect -23950 3323 -23500 3335
rect -23950 3289 -23934 3323
rect -23900 3289 -23742 3323
rect -23708 3289 -23550 3323
rect -23516 3289 -23500 3323
rect -23950 3267 -23500 3289
rect -23374 3323 -22924 3335
rect -23374 3322 -23166 3323
rect -23374 3288 -23358 3322
rect -23324 3289 -23166 3322
rect -23132 3289 -22974 3323
rect -22940 3289 -22924 3323
rect -23324 3288 -22924 3289
rect -23374 3267 -22924 3288
rect -22892 3308 -22837 3324
rect -24039 3136 -23984 3202
rect -23853 3222 -23788 3238
rect -23853 3188 -23838 3222
rect -23804 3188 -23788 3222
rect -23853 3136 -23788 3188
rect -23662 3222 -23215 3234
rect -23662 3188 -23646 3222
rect -23612 3188 -23454 3222
rect -23420 3188 -23262 3222
rect -23228 3188 -23215 3222
rect -23662 3170 -23215 3188
rect -23087 3222 -23022 3239
rect -23087 3188 -23070 3222
rect -23036 3188 -23022 3222
rect -23087 3136 -23022 3188
rect -22892 3202 -22878 3308
rect -22844 3202 -22837 3308
rect -22892 3136 -22837 3202
rect -24039 3125 -22837 3136
rect -24039 3114 -23398 3125
rect -23338 3114 -22837 3125
rect -24039 3068 -24001 3114
rect -22878 3068 -22837 3114
rect -24039 3065 -23398 3068
rect -23338 3065 -22837 3068
rect -24039 3045 -22837 3065
rect -20748 3308 -20693 3324
rect -20748 3202 -20739 3308
rect -20705 3202 -20693 3308
rect -20659 3323 -20209 3335
rect -20659 3289 -20643 3323
rect -20609 3289 -20451 3323
rect -20417 3289 -20259 3323
rect -20225 3289 -20209 3323
rect -20659 3267 -20209 3289
rect -20083 3323 -19633 3335
rect -20083 3322 -19875 3323
rect -20083 3288 -20067 3322
rect -20033 3289 -19875 3322
rect -19841 3289 -19683 3323
rect -19649 3289 -19633 3323
rect -20033 3288 -19633 3289
rect -20083 3267 -19633 3288
rect -19601 3308 -19546 3324
rect -20748 3136 -20693 3202
rect -20562 3222 -20497 3238
rect -20562 3188 -20547 3222
rect -20513 3188 -20497 3222
rect -20562 3136 -20497 3188
rect -20371 3222 -19924 3234
rect -20371 3188 -20355 3222
rect -20321 3188 -20163 3222
rect -20129 3188 -19971 3222
rect -19937 3188 -19924 3222
rect -20371 3170 -19924 3188
rect -19796 3222 -19731 3239
rect -19796 3188 -19779 3222
rect -19745 3188 -19731 3222
rect -19796 3136 -19731 3188
rect -19601 3202 -19587 3308
rect -19553 3202 -19546 3308
rect -19601 3136 -19546 3202
rect -20748 3125 -19546 3136
rect -20748 3114 -20107 3125
rect -20047 3114 -19546 3125
rect -20748 3068 -20710 3114
rect -19587 3068 -19546 3114
rect -20748 3065 -20107 3068
rect -20047 3065 -19546 3068
rect -20748 3045 -19546 3065
rect -17457 3308 -17402 3324
rect -17457 3202 -17448 3308
rect -17414 3202 -17402 3308
rect -17368 3323 -16918 3335
rect -17368 3289 -17352 3323
rect -17318 3289 -17160 3323
rect -17126 3289 -16968 3323
rect -16934 3289 -16918 3323
rect -17368 3267 -16918 3289
rect -16792 3323 -16342 3335
rect -16792 3322 -16584 3323
rect -16792 3288 -16776 3322
rect -16742 3289 -16584 3322
rect -16550 3289 -16392 3323
rect -16358 3289 -16342 3323
rect -16742 3288 -16342 3289
rect -16792 3267 -16342 3288
rect -16310 3308 -16255 3324
rect -17457 3136 -17402 3202
rect -17271 3222 -17206 3238
rect -17271 3188 -17256 3222
rect -17222 3188 -17206 3222
rect -17271 3136 -17206 3188
rect -17080 3222 -16633 3234
rect -17080 3188 -17064 3222
rect -17030 3188 -16872 3222
rect -16838 3188 -16680 3222
rect -16646 3188 -16633 3222
rect -17080 3170 -16633 3188
rect -16505 3222 -16440 3239
rect -16505 3188 -16488 3222
rect -16454 3188 -16440 3222
rect -16505 3136 -16440 3188
rect -16310 3202 -16296 3308
rect -16262 3202 -16255 3308
rect -16310 3136 -16255 3202
rect -17457 3125 -16255 3136
rect -17457 3114 -16816 3125
rect -16756 3114 -16255 3125
rect -17457 3068 -17419 3114
rect -16296 3068 -16255 3114
rect -17457 3065 -16816 3068
rect -16756 3065 -16255 3068
rect -17457 3045 -16255 3065
rect -14166 3308 -14111 3324
rect -14166 3202 -14157 3308
rect -14123 3202 -14111 3308
rect -14077 3323 -13627 3335
rect -14077 3289 -14061 3323
rect -14027 3289 -13869 3323
rect -13835 3289 -13677 3323
rect -13643 3289 -13627 3323
rect -14077 3267 -13627 3289
rect -13501 3323 -13051 3335
rect -13501 3322 -13293 3323
rect -13501 3288 -13485 3322
rect -13451 3289 -13293 3322
rect -13259 3289 -13101 3323
rect -13067 3289 -13051 3323
rect -13451 3288 -13051 3289
rect -13501 3267 -13051 3288
rect -13019 3308 -12964 3324
rect -14166 3136 -14111 3202
rect -13980 3222 -13915 3238
rect -13980 3188 -13965 3222
rect -13931 3188 -13915 3222
rect -13980 3136 -13915 3188
rect -13789 3222 -13342 3234
rect -13789 3188 -13773 3222
rect -13739 3188 -13581 3222
rect -13547 3188 -13389 3222
rect -13355 3188 -13342 3222
rect -13789 3170 -13342 3188
rect -13214 3222 -13149 3239
rect -13214 3188 -13197 3222
rect -13163 3188 -13149 3222
rect -13214 3136 -13149 3188
rect -13019 3202 -13005 3308
rect -12971 3202 -12964 3308
rect -13019 3136 -12964 3202
rect -14166 3125 -12964 3136
rect -14166 3114 -13525 3125
rect -13465 3114 -12964 3125
rect -14166 3068 -14128 3114
rect -13005 3068 -12964 3114
rect -14166 3065 -13525 3068
rect -13465 3065 -12964 3068
rect -14166 3045 -12964 3065
rect -10875 3308 -10820 3324
rect -10875 3202 -10866 3308
rect -10832 3202 -10820 3308
rect -10786 3323 -10336 3335
rect -10786 3289 -10770 3323
rect -10736 3289 -10578 3323
rect -10544 3289 -10386 3323
rect -10352 3289 -10336 3323
rect -10786 3267 -10336 3289
rect -10210 3323 -9760 3335
rect -10210 3322 -10002 3323
rect -10210 3288 -10194 3322
rect -10160 3289 -10002 3322
rect -9968 3289 -9810 3323
rect -9776 3289 -9760 3323
rect -10160 3288 -9760 3289
rect -10210 3267 -9760 3288
rect -9728 3308 -9673 3324
rect -10875 3136 -10820 3202
rect -10689 3222 -10624 3238
rect -10689 3188 -10674 3222
rect -10640 3188 -10624 3222
rect -10689 3136 -10624 3188
rect -10498 3222 -10051 3234
rect -10498 3188 -10482 3222
rect -10448 3188 -10290 3222
rect -10256 3188 -10098 3222
rect -10064 3188 -10051 3222
rect -10498 3170 -10051 3188
rect -9923 3222 -9858 3239
rect -9923 3188 -9906 3222
rect -9872 3188 -9858 3222
rect -9923 3136 -9858 3188
rect -9728 3202 -9714 3308
rect -9680 3202 -9673 3308
rect -9728 3136 -9673 3202
rect -10875 3125 -9673 3136
rect -10875 3114 -10234 3125
rect -10174 3114 -9673 3125
rect -10875 3068 -10837 3114
rect -9714 3068 -9673 3114
rect -10875 3065 -10234 3068
rect -10174 3065 -9673 3068
rect -10875 3045 -9673 3065
rect -7585 3308 -7530 3324
rect -7585 3202 -7576 3308
rect -7542 3202 -7530 3308
rect -7496 3323 -7046 3335
rect -7496 3289 -7480 3323
rect -7446 3289 -7288 3323
rect -7254 3289 -7096 3323
rect -7062 3289 -7046 3323
rect -7496 3267 -7046 3289
rect -6920 3323 -6470 3335
rect -6920 3322 -6712 3323
rect -6920 3288 -6904 3322
rect -6870 3289 -6712 3322
rect -6678 3289 -6520 3323
rect -6486 3289 -6470 3323
rect -6870 3288 -6470 3289
rect -6920 3267 -6470 3288
rect -6438 3308 -6383 3324
rect -7585 3136 -7530 3202
rect -7399 3222 -7334 3238
rect -7399 3188 -7384 3222
rect -7350 3188 -7334 3222
rect -7399 3136 -7334 3188
rect -7208 3222 -6761 3234
rect -7208 3188 -7192 3222
rect -7158 3188 -7000 3222
rect -6966 3188 -6808 3222
rect -6774 3188 -6761 3222
rect -7208 3170 -6761 3188
rect -6633 3222 -6568 3239
rect -6633 3188 -6616 3222
rect -6582 3188 -6568 3222
rect -6633 3136 -6568 3188
rect -6438 3202 -6424 3308
rect -6390 3202 -6383 3308
rect -6438 3136 -6383 3202
rect -7585 3125 -6383 3136
rect -7585 3114 -6944 3125
rect -6884 3114 -6383 3125
rect -7585 3068 -7547 3114
rect -6424 3068 -6383 3114
rect -7585 3065 -6944 3068
rect -6884 3065 -6383 3068
rect -7585 3045 -6383 3065
rect -4294 3308 -4239 3324
rect -4294 3202 -4285 3308
rect -4251 3202 -4239 3308
rect -4205 3323 -3755 3335
rect -4205 3289 -4189 3323
rect -4155 3289 -3997 3323
rect -3963 3289 -3805 3323
rect -3771 3289 -3755 3323
rect -4205 3267 -3755 3289
rect -3629 3323 -3179 3335
rect -3629 3322 -3421 3323
rect -3629 3288 -3613 3322
rect -3579 3289 -3421 3322
rect -3387 3289 -3229 3323
rect -3195 3289 -3179 3323
rect -3579 3288 -3179 3289
rect -3629 3267 -3179 3288
rect -3147 3308 -3092 3324
rect -4294 3136 -4239 3202
rect -4108 3222 -4043 3238
rect -4108 3188 -4093 3222
rect -4059 3188 -4043 3222
rect -4108 3136 -4043 3188
rect -3917 3222 -3470 3234
rect -3917 3188 -3901 3222
rect -3867 3188 -3709 3222
rect -3675 3188 -3517 3222
rect -3483 3188 -3470 3222
rect -3917 3170 -3470 3188
rect -3342 3222 -3277 3239
rect -3342 3188 -3325 3222
rect -3291 3188 -3277 3222
rect -3342 3136 -3277 3188
rect -3147 3202 -3133 3308
rect -3099 3202 -3092 3308
rect -3147 3136 -3092 3202
rect -4294 3125 -3092 3136
rect -4294 3114 -3653 3125
rect -3593 3114 -3092 3125
rect -4294 3068 -4256 3114
rect -3133 3068 -3092 3114
rect -4294 3065 -3653 3068
rect -3593 3065 -3092 3068
rect -4294 3045 -3092 3065
rect -1003 3308 -948 3324
rect -1003 3202 -994 3308
rect -960 3202 -948 3308
rect -914 3323 -464 3335
rect -914 3289 -898 3323
rect -864 3289 -706 3323
rect -672 3289 -514 3323
rect -480 3289 -464 3323
rect -914 3267 -464 3289
rect -338 3323 112 3335
rect -338 3322 -130 3323
rect -338 3288 -322 3322
rect -288 3289 -130 3322
rect -96 3289 62 3323
rect 96 3289 112 3323
rect -288 3288 112 3289
rect -338 3267 112 3288
rect 144 3308 199 3324
rect -1003 3136 -948 3202
rect -817 3222 -752 3238
rect -817 3188 -802 3222
rect -768 3188 -752 3222
rect -817 3136 -752 3188
rect -626 3222 -179 3234
rect -626 3188 -610 3222
rect -576 3188 -418 3222
rect -384 3188 -226 3222
rect -192 3188 -179 3222
rect -626 3170 -179 3188
rect -51 3222 14 3239
rect -51 3188 -34 3222
rect 0 3188 14 3222
rect -51 3136 14 3188
rect 144 3202 158 3308
rect 192 3202 199 3308
rect 144 3136 199 3202
rect -1003 3125 199 3136
rect -1003 3114 -362 3125
rect -302 3114 199 3125
rect -1003 3068 -965 3114
rect 158 3068 199 3114
rect -1003 3065 -362 3068
rect -302 3065 199 3068
rect -1003 3045 199 3065
rect -24716 2733 -23506 2761
rect -24716 2661 -24670 2733
rect -23548 2661 -23506 2733
rect -24716 2627 -23506 2661
rect -24716 2558 -24462 2627
rect -24716 2456 -24704 2558
rect -24670 2456 -24512 2558
rect -24478 2456 -24462 2558
rect -24716 2435 -24462 2456
rect -24336 2556 -23886 2582
rect -24336 2454 -24320 2556
rect -24286 2555 -23886 2556
rect -24286 2454 -24128 2555
rect -24336 2453 -24128 2454
rect -24094 2453 -23936 2555
rect -23902 2453 -23886 2555
rect -24336 2435 -23886 2453
rect -23760 2555 -23506 2627
rect -23760 2453 -23744 2555
rect -23710 2453 -23552 2555
rect -23518 2453 -23506 2555
rect -23760 2435 -23506 2453
rect -23157 2733 -21947 2761
rect -23157 2661 -23111 2733
rect -21989 2661 -21947 2733
rect -23157 2627 -21947 2661
rect -23157 2558 -22903 2627
rect -23157 2456 -23145 2558
rect -23111 2456 -22953 2558
rect -22919 2456 -22903 2558
rect -23157 2435 -22903 2456
rect -22777 2556 -22327 2582
rect -22777 2454 -22761 2556
rect -22727 2555 -22327 2556
rect -22727 2454 -22569 2555
rect -22777 2453 -22569 2454
rect -22535 2453 -22377 2555
rect -22343 2453 -22327 2555
rect -22777 2435 -22327 2453
rect -22201 2555 -21947 2627
rect -22201 2453 -22185 2555
rect -22151 2453 -21993 2555
rect -21959 2453 -21947 2555
rect -22201 2435 -21947 2453
rect -21425 2733 -20215 2761
rect -21425 2661 -21379 2733
rect -20257 2661 -20215 2733
rect -21425 2627 -20215 2661
rect -21425 2558 -21171 2627
rect -21425 2456 -21413 2558
rect -21379 2456 -21221 2558
rect -21187 2456 -21171 2558
rect -21425 2435 -21171 2456
rect -21045 2556 -20595 2582
rect -21045 2454 -21029 2556
rect -20995 2555 -20595 2556
rect -20995 2454 -20837 2555
rect -21045 2453 -20837 2454
rect -20803 2453 -20645 2555
rect -20611 2453 -20595 2555
rect -21045 2435 -20595 2453
rect -20469 2555 -20215 2627
rect -20469 2453 -20453 2555
rect -20419 2453 -20261 2555
rect -20227 2453 -20215 2555
rect -20469 2435 -20215 2453
rect -19866 2733 -18656 2761
rect -19866 2661 -19820 2733
rect -18698 2661 -18656 2733
rect -19866 2627 -18656 2661
rect -19866 2558 -19612 2627
rect -19866 2456 -19854 2558
rect -19820 2456 -19662 2558
rect -19628 2456 -19612 2558
rect -19866 2435 -19612 2456
rect -19486 2556 -19036 2582
rect -19486 2454 -19470 2556
rect -19436 2555 -19036 2556
rect -19436 2454 -19278 2555
rect -19486 2453 -19278 2454
rect -19244 2453 -19086 2555
rect -19052 2453 -19036 2555
rect -19486 2435 -19036 2453
rect -18910 2555 -18656 2627
rect -18910 2453 -18894 2555
rect -18860 2453 -18702 2555
rect -18668 2453 -18656 2555
rect -18910 2435 -18656 2453
rect -18134 2733 -16924 2761
rect -18134 2661 -18088 2733
rect -16966 2661 -16924 2733
rect -18134 2627 -16924 2661
rect -18134 2558 -17880 2627
rect -18134 2456 -18122 2558
rect -18088 2456 -17930 2558
rect -17896 2456 -17880 2558
rect -18134 2435 -17880 2456
rect -17754 2556 -17304 2582
rect -17754 2454 -17738 2556
rect -17704 2555 -17304 2556
rect -17704 2454 -17546 2555
rect -17754 2453 -17546 2454
rect -17512 2453 -17354 2555
rect -17320 2453 -17304 2555
rect -17754 2435 -17304 2453
rect -17178 2555 -16924 2627
rect -17178 2453 -17162 2555
rect -17128 2453 -16970 2555
rect -16936 2453 -16924 2555
rect -17178 2435 -16924 2453
rect -16575 2733 -15365 2761
rect -16575 2661 -16529 2733
rect -15407 2661 -15365 2733
rect -16575 2627 -15365 2661
rect -16575 2558 -16321 2627
rect -16575 2456 -16563 2558
rect -16529 2456 -16371 2558
rect -16337 2456 -16321 2558
rect -16575 2435 -16321 2456
rect -16195 2556 -15745 2582
rect -16195 2454 -16179 2556
rect -16145 2555 -15745 2556
rect -16145 2454 -15987 2555
rect -16195 2453 -15987 2454
rect -15953 2453 -15795 2555
rect -15761 2453 -15745 2555
rect -16195 2435 -15745 2453
rect -15619 2555 -15365 2627
rect -15619 2453 -15603 2555
rect -15569 2453 -15411 2555
rect -15377 2453 -15365 2555
rect -15619 2435 -15365 2453
rect -14843 2733 -13633 2761
rect -14843 2661 -14797 2733
rect -13675 2661 -13633 2733
rect -14843 2627 -13633 2661
rect -14843 2558 -14589 2627
rect -14843 2456 -14831 2558
rect -14797 2456 -14639 2558
rect -14605 2456 -14589 2558
rect -14843 2435 -14589 2456
rect -14463 2556 -14013 2582
rect -14463 2454 -14447 2556
rect -14413 2555 -14013 2556
rect -14413 2454 -14255 2555
rect -14463 2453 -14255 2454
rect -14221 2453 -14063 2555
rect -14029 2453 -14013 2555
rect -14463 2435 -14013 2453
rect -13887 2555 -13633 2627
rect -13887 2453 -13871 2555
rect -13837 2453 -13679 2555
rect -13645 2453 -13633 2555
rect -13887 2435 -13633 2453
rect -13284 2733 -12074 2761
rect -13284 2661 -13238 2733
rect -12116 2661 -12074 2733
rect -13284 2627 -12074 2661
rect -13284 2558 -13030 2627
rect -13284 2456 -13272 2558
rect -13238 2456 -13080 2558
rect -13046 2456 -13030 2558
rect -13284 2435 -13030 2456
rect -12904 2556 -12454 2582
rect -12904 2454 -12888 2556
rect -12854 2555 -12454 2556
rect -12854 2454 -12696 2555
rect -12904 2453 -12696 2454
rect -12662 2453 -12504 2555
rect -12470 2453 -12454 2555
rect -12904 2435 -12454 2453
rect -12328 2555 -12074 2627
rect -12328 2453 -12312 2555
rect -12278 2453 -12120 2555
rect -12086 2453 -12074 2555
rect -12328 2435 -12074 2453
rect -11552 2733 -10342 2761
rect -11552 2661 -11506 2733
rect -10384 2661 -10342 2733
rect -11552 2627 -10342 2661
rect -11552 2558 -11298 2627
rect -11552 2456 -11540 2558
rect -11506 2456 -11348 2558
rect -11314 2456 -11298 2558
rect -11552 2435 -11298 2456
rect -11172 2556 -10722 2582
rect -11172 2454 -11156 2556
rect -11122 2555 -10722 2556
rect -11122 2454 -10964 2555
rect -11172 2453 -10964 2454
rect -10930 2453 -10772 2555
rect -10738 2453 -10722 2555
rect -11172 2435 -10722 2453
rect -10596 2555 -10342 2627
rect -10596 2453 -10580 2555
rect -10546 2453 -10388 2555
rect -10354 2453 -10342 2555
rect -10596 2435 -10342 2453
rect -9993 2733 -8783 2761
rect -9993 2661 -9947 2733
rect -8825 2661 -8783 2733
rect -9993 2627 -8783 2661
rect -9993 2558 -9739 2627
rect -9993 2456 -9981 2558
rect -9947 2456 -9789 2558
rect -9755 2456 -9739 2558
rect -9993 2435 -9739 2456
rect -9613 2556 -9163 2582
rect -9613 2454 -9597 2556
rect -9563 2555 -9163 2556
rect -9563 2454 -9405 2555
rect -9613 2453 -9405 2454
rect -9371 2453 -9213 2555
rect -9179 2453 -9163 2555
rect -9613 2435 -9163 2453
rect -9037 2555 -8783 2627
rect -9037 2453 -9021 2555
rect -8987 2453 -8829 2555
rect -8795 2453 -8783 2555
rect -9037 2435 -8783 2453
rect -8262 2733 -7052 2761
rect -8262 2661 -8216 2733
rect -7094 2661 -7052 2733
rect -8262 2627 -7052 2661
rect -8262 2558 -8008 2627
rect -8262 2456 -8250 2558
rect -8216 2456 -8058 2558
rect -8024 2456 -8008 2558
rect -8262 2435 -8008 2456
rect -7882 2556 -7432 2582
rect -7882 2454 -7866 2556
rect -7832 2555 -7432 2556
rect -7832 2454 -7674 2555
rect -7882 2453 -7674 2454
rect -7640 2453 -7482 2555
rect -7448 2453 -7432 2555
rect -7882 2435 -7432 2453
rect -7306 2555 -7052 2627
rect -7306 2453 -7290 2555
rect -7256 2453 -7098 2555
rect -7064 2453 -7052 2555
rect -7306 2435 -7052 2453
rect -6703 2733 -5493 2761
rect -6703 2661 -6657 2733
rect -5535 2661 -5493 2733
rect -6703 2627 -5493 2661
rect -6703 2558 -6449 2627
rect -6703 2456 -6691 2558
rect -6657 2456 -6499 2558
rect -6465 2456 -6449 2558
rect -6703 2435 -6449 2456
rect -6323 2556 -5873 2582
rect -6323 2454 -6307 2556
rect -6273 2555 -5873 2556
rect -6273 2454 -6115 2555
rect -6323 2453 -6115 2454
rect -6081 2453 -5923 2555
rect -5889 2453 -5873 2555
rect -6323 2435 -5873 2453
rect -5747 2555 -5493 2627
rect -5747 2453 -5731 2555
rect -5697 2453 -5539 2555
rect -5505 2453 -5493 2555
rect -5747 2435 -5493 2453
rect -4971 2733 -3761 2761
rect -4971 2661 -4925 2733
rect -3803 2661 -3761 2733
rect -4971 2627 -3761 2661
rect -4971 2558 -4717 2627
rect -4971 2456 -4959 2558
rect -4925 2456 -4767 2558
rect -4733 2456 -4717 2558
rect -4971 2435 -4717 2456
rect -4591 2556 -4141 2582
rect -4591 2454 -4575 2556
rect -4541 2555 -4141 2556
rect -4541 2454 -4383 2555
rect -4591 2453 -4383 2454
rect -4349 2453 -4191 2555
rect -4157 2453 -4141 2555
rect -4591 2435 -4141 2453
rect -4015 2555 -3761 2627
rect -4015 2453 -3999 2555
rect -3965 2453 -3807 2555
rect -3773 2453 -3761 2555
rect -4015 2435 -3761 2453
rect -3412 2733 -2202 2761
rect -3412 2661 -3366 2733
rect -2244 2661 -2202 2733
rect -3412 2627 -2202 2661
rect -3412 2558 -3158 2627
rect -3412 2456 -3400 2558
rect -3366 2456 -3208 2558
rect -3174 2456 -3158 2558
rect -3412 2435 -3158 2456
rect -3032 2556 -2582 2582
rect -3032 2454 -3016 2556
rect -2982 2555 -2582 2556
rect -2982 2454 -2824 2555
rect -3032 2453 -2824 2454
rect -2790 2453 -2632 2555
rect -2598 2453 -2582 2555
rect -3032 2435 -2582 2453
rect -2456 2555 -2202 2627
rect -2456 2453 -2440 2555
rect -2406 2453 -2248 2555
rect -2214 2453 -2202 2555
rect -2456 2435 -2202 2453
rect -1680 2733 -470 2761
rect -1680 2661 -1634 2733
rect -512 2661 -470 2733
rect -1680 2627 -470 2661
rect -1680 2558 -1426 2627
rect -1680 2456 -1668 2558
rect -1634 2456 -1476 2558
rect -1442 2456 -1426 2558
rect -1680 2435 -1426 2456
rect -1300 2556 -850 2582
rect -1300 2454 -1284 2556
rect -1250 2555 -850 2556
rect -1250 2454 -1092 2555
rect -1300 2453 -1092 2454
rect -1058 2453 -900 2555
rect -866 2453 -850 2555
rect -1300 2435 -850 2453
rect -724 2555 -470 2627
rect -724 2453 -708 2555
rect -674 2453 -516 2555
rect -482 2453 -470 2555
rect -724 2435 -470 2453
rect -121 2733 1089 2761
rect -121 2661 -75 2733
rect 1047 2661 1089 2733
rect -121 2627 1089 2661
rect -121 2558 133 2627
rect -121 2456 -109 2558
rect -75 2456 83 2558
rect 117 2456 133 2558
rect -121 2435 133 2456
rect 259 2556 709 2582
rect 259 2454 275 2556
rect 309 2555 709 2556
rect 309 2454 467 2555
rect 259 2453 467 2454
rect 501 2453 659 2555
rect 693 2453 709 2555
rect 259 2435 709 2453
rect 835 2555 1089 2627
rect 835 2453 851 2555
rect 885 2453 1043 2555
rect 1077 2453 1089 2555
rect 835 2435 1089 2453
rect -24624 2372 -23598 2397
rect -24624 2248 -24608 2372
rect -24574 2248 -24416 2372
rect -24382 2248 -24224 2372
rect -24190 2248 -24032 2372
rect -23998 2248 -23840 2372
rect -23806 2371 -23598 2372
rect -23806 2248 -23648 2371
rect -24624 2247 -23648 2248
rect -23614 2247 -23598 2371
rect -24624 2218 -23598 2247
rect -23065 2372 -22039 2397
rect -23065 2248 -23049 2372
rect -23015 2248 -22857 2372
rect -22823 2248 -22665 2372
rect -22631 2248 -22473 2372
rect -22439 2248 -22281 2372
rect -22247 2371 -22039 2372
rect -22247 2248 -22089 2371
rect -23065 2247 -22089 2248
rect -22055 2247 -22039 2371
rect -23065 2218 -22039 2247
rect -21333 2372 -20307 2397
rect -21333 2248 -21317 2372
rect -21283 2248 -21125 2372
rect -21091 2248 -20933 2372
rect -20899 2248 -20741 2372
rect -20707 2248 -20549 2372
rect -20515 2371 -20307 2372
rect -20515 2248 -20357 2371
rect -21333 2247 -20357 2248
rect -20323 2247 -20307 2371
rect -21333 2218 -20307 2247
rect -19774 2372 -18748 2397
rect -19774 2248 -19758 2372
rect -19724 2248 -19566 2372
rect -19532 2248 -19374 2372
rect -19340 2248 -19182 2372
rect -19148 2248 -18990 2372
rect -18956 2371 -18748 2372
rect -18956 2248 -18798 2371
rect -19774 2247 -18798 2248
rect -18764 2247 -18748 2371
rect -19774 2218 -18748 2247
rect -18042 2372 -17016 2397
rect -18042 2248 -18026 2372
rect -17992 2248 -17834 2372
rect -17800 2248 -17642 2372
rect -17608 2248 -17450 2372
rect -17416 2248 -17258 2372
rect -17224 2371 -17016 2372
rect -17224 2248 -17066 2371
rect -18042 2247 -17066 2248
rect -17032 2247 -17016 2371
rect -18042 2218 -17016 2247
rect -16483 2372 -15457 2397
rect -16483 2248 -16467 2372
rect -16433 2248 -16275 2372
rect -16241 2248 -16083 2372
rect -16049 2248 -15891 2372
rect -15857 2248 -15699 2372
rect -15665 2371 -15457 2372
rect -15665 2248 -15507 2371
rect -16483 2247 -15507 2248
rect -15473 2247 -15457 2371
rect -16483 2218 -15457 2247
rect -14751 2372 -13725 2397
rect -14751 2248 -14735 2372
rect -14701 2248 -14543 2372
rect -14509 2248 -14351 2372
rect -14317 2248 -14159 2372
rect -14125 2248 -13967 2372
rect -13933 2371 -13725 2372
rect -13933 2248 -13775 2371
rect -14751 2247 -13775 2248
rect -13741 2247 -13725 2371
rect -14751 2218 -13725 2247
rect -13192 2372 -12166 2397
rect -13192 2248 -13176 2372
rect -13142 2248 -12984 2372
rect -12950 2248 -12792 2372
rect -12758 2248 -12600 2372
rect -12566 2248 -12408 2372
rect -12374 2371 -12166 2372
rect -12374 2248 -12216 2371
rect -13192 2247 -12216 2248
rect -12182 2247 -12166 2371
rect -13192 2218 -12166 2247
rect -11460 2372 -10434 2397
rect -11460 2248 -11444 2372
rect -11410 2248 -11252 2372
rect -11218 2248 -11060 2372
rect -11026 2248 -10868 2372
rect -10834 2248 -10676 2372
rect -10642 2371 -10434 2372
rect -10642 2248 -10484 2371
rect -11460 2247 -10484 2248
rect -10450 2247 -10434 2371
rect -11460 2218 -10434 2247
rect -9901 2372 -8875 2397
rect -9901 2248 -9885 2372
rect -9851 2248 -9693 2372
rect -9659 2248 -9501 2372
rect -9467 2248 -9309 2372
rect -9275 2248 -9117 2372
rect -9083 2371 -8875 2372
rect -9083 2248 -8925 2371
rect -9901 2247 -8925 2248
rect -8891 2247 -8875 2371
rect -9901 2218 -8875 2247
rect -8170 2372 -7144 2397
rect -8170 2248 -8154 2372
rect -8120 2248 -7962 2372
rect -7928 2248 -7770 2372
rect -7736 2248 -7578 2372
rect -7544 2248 -7386 2372
rect -7352 2371 -7144 2372
rect -7352 2248 -7194 2371
rect -8170 2247 -7194 2248
rect -7160 2247 -7144 2371
rect -8170 2218 -7144 2247
rect -6611 2372 -5585 2397
rect -6611 2248 -6595 2372
rect -6561 2248 -6403 2372
rect -6369 2248 -6211 2372
rect -6177 2248 -6019 2372
rect -5985 2248 -5827 2372
rect -5793 2371 -5585 2372
rect -5793 2248 -5635 2371
rect -6611 2247 -5635 2248
rect -5601 2247 -5585 2371
rect -6611 2218 -5585 2247
rect -4879 2372 -3853 2397
rect -4879 2248 -4863 2372
rect -4829 2248 -4671 2372
rect -4637 2248 -4479 2372
rect -4445 2248 -4287 2372
rect -4253 2248 -4095 2372
rect -4061 2371 -3853 2372
rect -4061 2248 -3903 2371
rect -4879 2247 -3903 2248
rect -3869 2247 -3853 2371
rect -4879 2218 -3853 2247
rect -3320 2372 -2294 2397
rect -3320 2248 -3304 2372
rect -3270 2248 -3112 2372
rect -3078 2248 -2920 2372
rect -2886 2248 -2728 2372
rect -2694 2248 -2536 2372
rect -2502 2371 -2294 2372
rect -2502 2248 -2344 2371
rect -3320 2247 -2344 2248
rect -2310 2247 -2294 2371
rect -3320 2218 -2294 2247
rect -1588 2372 -562 2397
rect -1588 2248 -1572 2372
rect -1538 2248 -1380 2372
rect -1346 2248 -1188 2372
rect -1154 2248 -996 2372
rect -962 2248 -804 2372
rect -770 2371 -562 2372
rect -770 2248 -612 2371
rect -1588 2247 -612 2248
rect -578 2247 -562 2371
rect -1588 2218 -562 2247
rect -29 2372 997 2397
rect -29 2248 -13 2372
rect 21 2248 179 2372
rect 213 2248 371 2372
rect 405 2248 563 2372
rect 597 2248 755 2372
rect 789 2371 997 2372
rect 789 2248 947 2371
rect -29 2247 947 2248
rect 981 2247 997 2371
rect -29 2218 997 2247
rect -24716 2163 -24462 2185
rect -24716 2061 -24704 2163
rect -24670 2097 -24512 2163
rect -24478 2097 -24462 2163
rect -24670 2061 -24462 2097
rect -24336 2157 -23886 2174
rect -24336 2097 -24320 2157
rect -24286 2140 -23936 2157
rect -24286 2097 -24128 2140
rect -24094 2097 -23936 2140
rect -23902 2097 -23886 2157
rect -24336 2082 -23886 2097
rect -23760 2164 -23506 2185
rect -23760 2097 -23744 2164
rect -23710 2097 -23552 2164
rect -23518 2097 -23506 2164
rect -24716 2038 -24462 2061
rect -23760 2038 -23506 2097
rect -23157 2163 -22903 2185
rect -23157 2061 -23145 2163
rect -23111 2097 -22953 2163
rect -22919 2097 -22903 2163
rect -23111 2061 -22903 2097
rect -22777 2157 -22327 2174
rect -22777 2097 -22761 2157
rect -22727 2140 -22377 2157
rect -22727 2097 -22569 2140
rect -22535 2097 -22377 2140
rect -22343 2097 -22327 2157
rect -22777 2082 -22327 2097
rect -22201 2164 -21947 2185
rect -22201 2097 -22185 2164
rect -22151 2097 -21993 2164
rect -21959 2097 -21947 2164
rect -23157 2038 -22903 2061
rect -22201 2038 -21947 2097
rect -21425 2163 -21171 2185
rect -21425 2061 -21413 2163
rect -21379 2097 -21221 2163
rect -21187 2097 -21171 2163
rect -21379 2061 -21171 2097
rect -21045 2157 -20595 2174
rect -21045 2097 -21029 2157
rect -20995 2140 -20645 2157
rect -20995 2097 -20837 2140
rect -20803 2097 -20645 2140
rect -20611 2097 -20595 2157
rect -21045 2082 -20595 2097
rect -20469 2164 -20215 2185
rect -20469 2097 -20453 2164
rect -20419 2097 -20261 2164
rect -20227 2097 -20215 2164
rect -21425 2038 -21171 2061
rect -20469 2038 -20215 2097
rect -19866 2163 -19612 2185
rect -19866 2061 -19854 2163
rect -19820 2097 -19662 2163
rect -19628 2097 -19612 2163
rect -19820 2061 -19612 2097
rect -19486 2157 -19036 2174
rect -19486 2097 -19470 2157
rect -19436 2140 -19086 2157
rect -19436 2097 -19278 2140
rect -19244 2097 -19086 2140
rect -19052 2097 -19036 2157
rect -19486 2082 -19036 2097
rect -18910 2164 -18656 2185
rect -18910 2097 -18894 2164
rect -18860 2097 -18702 2164
rect -18668 2097 -18656 2164
rect -19866 2038 -19612 2061
rect -18910 2038 -18656 2097
rect -18134 2163 -17880 2185
rect -18134 2061 -18122 2163
rect -18088 2097 -17930 2163
rect -17896 2097 -17880 2163
rect -18088 2061 -17880 2097
rect -17754 2157 -17304 2174
rect -17754 2097 -17738 2157
rect -17704 2140 -17354 2157
rect -17704 2097 -17546 2140
rect -17512 2097 -17354 2140
rect -17320 2097 -17304 2157
rect -17754 2082 -17304 2097
rect -17178 2164 -16924 2185
rect -17178 2097 -17162 2164
rect -17128 2097 -16970 2164
rect -16936 2097 -16924 2164
rect -18134 2038 -17880 2061
rect -17178 2038 -16924 2097
rect -16575 2163 -16321 2185
rect -16575 2061 -16563 2163
rect -16529 2097 -16371 2163
rect -16337 2097 -16321 2163
rect -16529 2061 -16321 2097
rect -16195 2157 -15745 2174
rect -16195 2097 -16179 2157
rect -16145 2140 -15795 2157
rect -16145 2097 -15987 2140
rect -15953 2097 -15795 2140
rect -15761 2097 -15745 2157
rect -16195 2082 -15745 2097
rect -15619 2164 -15365 2185
rect -15619 2097 -15603 2164
rect -15569 2097 -15411 2164
rect -15377 2097 -15365 2164
rect -16575 2038 -16321 2061
rect -15619 2038 -15365 2097
rect -14843 2163 -14589 2185
rect -14843 2061 -14831 2163
rect -14797 2097 -14639 2163
rect -14605 2097 -14589 2163
rect -14797 2061 -14589 2097
rect -14463 2157 -14013 2174
rect -14463 2097 -14447 2157
rect -14413 2140 -14063 2157
rect -14413 2097 -14255 2140
rect -14221 2097 -14063 2140
rect -14029 2097 -14013 2157
rect -14463 2082 -14013 2097
rect -13887 2164 -13633 2185
rect -13887 2097 -13871 2164
rect -13837 2097 -13679 2164
rect -13645 2097 -13633 2164
rect -14843 2038 -14589 2061
rect -13887 2038 -13633 2097
rect -13284 2163 -13030 2185
rect -13284 2061 -13272 2163
rect -13238 2097 -13080 2163
rect -13046 2097 -13030 2163
rect -13238 2061 -13030 2097
rect -12904 2157 -12454 2174
rect -12904 2097 -12888 2157
rect -12854 2140 -12504 2157
rect -12854 2097 -12696 2140
rect -12662 2097 -12504 2140
rect -12470 2097 -12454 2157
rect -12904 2082 -12454 2097
rect -12328 2164 -12074 2185
rect -12328 2097 -12312 2164
rect -12278 2097 -12120 2164
rect -12086 2097 -12074 2164
rect -13284 2038 -13030 2061
rect -12328 2038 -12074 2097
rect -11552 2163 -11298 2185
rect -11552 2061 -11540 2163
rect -11506 2097 -11348 2163
rect -11314 2097 -11298 2163
rect -11506 2061 -11298 2097
rect -11172 2157 -10722 2174
rect -11172 2097 -11156 2157
rect -11122 2140 -10772 2157
rect -11122 2097 -10964 2140
rect -10930 2097 -10772 2140
rect -10738 2097 -10722 2157
rect -11172 2082 -10722 2097
rect -10596 2164 -10342 2185
rect -10596 2097 -10580 2164
rect -10546 2097 -10388 2164
rect -10354 2097 -10342 2164
rect -11552 2038 -11298 2061
rect -10596 2038 -10342 2097
rect -9993 2163 -9739 2185
rect -9993 2061 -9981 2163
rect -9947 2097 -9789 2163
rect -9755 2097 -9739 2163
rect -9947 2061 -9739 2097
rect -9613 2157 -9163 2174
rect -9613 2097 -9597 2157
rect -9563 2140 -9213 2157
rect -9563 2097 -9405 2140
rect -9371 2097 -9213 2140
rect -9179 2097 -9163 2157
rect -9613 2082 -9163 2097
rect -9037 2164 -8783 2185
rect -9037 2097 -9021 2164
rect -8987 2097 -8829 2164
rect -8795 2097 -8783 2164
rect -9993 2038 -9739 2061
rect -9037 2038 -8783 2097
rect -8262 2163 -8008 2185
rect -8262 2061 -8250 2163
rect -8216 2097 -8058 2163
rect -8024 2097 -8008 2163
rect -8216 2061 -8008 2097
rect -7882 2157 -7432 2174
rect -7882 2097 -7866 2157
rect -7832 2140 -7482 2157
rect -7832 2097 -7674 2140
rect -7640 2097 -7482 2140
rect -7448 2097 -7432 2157
rect -7882 2082 -7432 2097
rect -7306 2164 -7052 2185
rect -7306 2097 -7290 2164
rect -7256 2097 -7098 2164
rect -7064 2097 -7052 2164
rect -8262 2038 -8008 2061
rect -7306 2038 -7052 2097
rect -6703 2163 -6449 2185
rect -6703 2061 -6691 2163
rect -6657 2097 -6499 2163
rect -6465 2097 -6449 2163
rect -6657 2061 -6449 2097
rect -6323 2157 -5873 2174
rect -6323 2097 -6307 2157
rect -6273 2140 -5923 2157
rect -6273 2097 -6115 2140
rect -6081 2097 -5923 2140
rect -5889 2097 -5873 2157
rect -6323 2082 -5873 2097
rect -5747 2164 -5493 2185
rect -5747 2097 -5731 2164
rect -5697 2097 -5539 2164
rect -5505 2097 -5493 2164
rect -6703 2038 -6449 2061
rect -5747 2038 -5493 2097
rect -4971 2163 -4717 2185
rect -4971 2061 -4959 2163
rect -4925 2097 -4767 2163
rect -4733 2097 -4717 2163
rect -4925 2061 -4717 2097
rect -4591 2157 -4141 2174
rect -4591 2097 -4575 2157
rect -4541 2140 -4191 2157
rect -4541 2097 -4383 2140
rect -4349 2097 -4191 2140
rect -4157 2097 -4141 2157
rect -4591 2082 -4141 2097
rect -4015 2164 -3761 2185
rect -4015 2097 -3999 2164
rect -3965 2097 -3807 2164
rect -3773 2097 -3761 2164
rect -4971 2038 -4717 2061
rect -4015 2038 -3761 2097
rect -3412 2163 -3158 2185
rect -3412 2061 -3400 2163
rect -3366 2097 -3208 2163
rect -3174 2097 -3158 2163
rect -3366 2061 -3158 2097
rect -3032 2157 -2582 2174
rect -3032 2097 -3016 2157
rect -2982 2140 -2632 2157
rect -2982 2097 -2824 2140
rect -2790 2097 -2632 2140
rect -2598 2097 -2582 2157
rect -3032 2082 -2582 2097
rect -2456 2164 -2202 2185
rect -2456 2097 -2440 2164
rect -2406 2097 -2248 2164
rect -2214 2097 -2202 2164
rect -3412 2038 -3158 2061
rect -2456 2038 -2202 2097
rect -1680 2163 -1426 2185
rect -1680 2061 -1668 2163
rect -1634 2097 -1476 2163
rect -1442 2097 -1426 2163
rect -1634 2061 -1426 2097
rect -1300 2157 -850 2174
rect -1300 2097 -1284 2157
rect -1250 2140 -900 2157
rect -1250 2097 -1092 2140
rect -1058 2097 -900 2140
rect -866 2097 -850 2157
rect -1300 2082 -850 2097
rect -724 2164 -470 2185
rect -724 2097 -708 2164
rect -674 2097 -516 2164
rect -482 2097 -470 2164
rect -1680 2038 -1426 2061
rect -724 2038 -470 2097
rect -121 2163 133 2185
rect -121 2061 -109 2163
rect -75 2097 83 2163
rect 117 2097 133 2163
rect -75 2061 133 2097
rect 259 2157 709 2174
rect 259 2097 275 2157
rect 309 2140 659 2157
rect 309 2097 467 2140
rect 501 2097 659 2140
rect 693 2097 709 2157
rect 259 2082 709 2097
rect 835 2164 1089 2185
rect 835 2097 851 2164
rect 885 2097 1043 2164
rect 1077 2097 1089 2164
rect -121 2038 133 2061
rect 835 2038 1089 2097
rect -24939 1938 -24804 1962
rect -24939 1828 -24921 1938
rect -24825 1830 -24804 1938
rect -21648 1938 -21513 1962
rect -23465 1903 -23274 1908
rect -23466 1893 -23274 1903
rect -23466 1886 -23364 1893
rect -23291 1886 -23274 1893
rect -24874 1828 -24804 1830
rect -24939 1808 -24804 1828
rect -24643 1845 -23854 1863
rect -24643 1837 -24000 1845
rect -24643 1784 -24606 1837
rect -24473 1792 -24000 1837
rect -23886 1792 -23854 1845
rect -24473 1784 -23854 1792
rect -24643 1764 -23854 1784
rect -23784 1844 -23669 1863
rect -23784 1776 -23766 1844
rect -23686 1776 -23669 1844
rect -23466 1803 -23439 1886
rect -24862 1705 -24657 1724
rect -24862 1597 -24818 1705
rect -24742 1679 -24657 1705
rect -23784 1679 -23669 1776
rect -23553 1789 -23439 1803
rect -23289 1789 -23274 1886
rect -23553 1773 -23274 1789
rect -23084 1845 -22295 1863
rect -23084 1837 -22441 1845
rect -23084 1784 -23047 1837
rect -22914 1792 -22441 1837
rect -22327 1792 -22295 1845
rect -22914 1784 -22295 1792
rect -23553 1710 -23382 1773
rect -23084 1764 -22295 1784
rect -22225 1844 -22110 1863
rect -22225 1776 -22207 1844
rect -22127 1776 -22110 1844
rect -21648 1828 -21630 1938
rect -21534 1830 -21513 1938
rect -18357 1938 -18222 1962
rect -20174 1903 -19983 1908
rect -20175 1893 -19983 1903
rect -20175 1886 -20073 1893
rect -20000 1886 -19983 1893
rect -21583 1828 -21513 1830
rect -21648 1808 -21513 1828
rect -21352 1845 -20563 1863
rect -21352 1837 -20709 1845
rect -24742 1597 -23669 1679
rect -24862 1593 -23669 1597
rect -23595 1673 -23382 1710
rect -23595 1618 -23584 1673
rect -23519 1618 -23382 1673
rect -23595 1594 -23382 1618
rect -23303 1698 -23098 1724
rect -23303 1601 -23263 1698
rect -23147 1679 -23098 1698
rect -22225 1679 -22110 1776
rect -21994 1710 -21714 1803
rect -21352 1784 -21315 1837
rect -21182 1792 -20709 1837
rect -20595 1792 -20563 1845
rect -21182 1784 -20563 1792
rect -21352 1764 -20563 1784
rect -20493 1844 -20378 1863
rect -20493 1776 -20475 1844
rect -20395 1776 -20378 1844
rect -20175 1803 -20148 1886
rect -23147 1601 -22110 1679
rect -23303 1593 -22110 1601
rect -22036 1673 -21714 1710
rect -22036 1618 -22025 1673
rect -21960 1618 -21714 1673
rect -22036 1594 -21714 1618
rect -24862 1581 -24657 1593
rect -23303 1581 -23098 1593
rect -24711 1524 -24656 1540
rect -24711 1418 -24704 1524
rect -24670 1418 -24656 1524
rect -24624 1539 -24174 1551
rect -24624 1505 -24608 1539
rect -24574 1505 -24416 1539
rect -24382 1538 -24174 1539
rect -24382 1505 -24224 1538
rect -24624 1504 -24224 1505
rect -24190 1504 -24174 1538
rect -24624 1483 -24174 1504
rect -24048 1539 -23598 1551
rect -24048 1505 -24032 1539
rect -23998 1505 -23840 1539
rect -23806 1505 -23648 1539
rect -23614 1505 -23598 1539
rect -24048 1483 -23598 1505
rect -23564 1524 -23509 1540
rect -24711 1352 -24656 1418
rect -24526 1438 -24461 1455
rect -24526 1404 -24512 1438
rect -24478 1404 -24461 1438
rect -24526 1352 -24461 1404
rect -24333 1438 -23886 1450
rect -24333 1404 -24320 1438
rect -24286 1404 -24128 1438
rect -24094 1404 -23936 1438
rect -23902 1404 -23886 1438
rect -24333 1386 -23886 1404
rect -23760 1438 -23695 1454
rect -23760 1404 -23744 1438
rect -23710 1404 -23695 1438
rect -23760 1352 -23695 1404
rect -23564 1418 -23552 1524
rect -23518 1418 -23509 1524
rect -23564 1352 -23509 1418
rect -24711 1341 -23509 1352
rect -24711 1330 -24210 1341
rect -24150 1330 -23509 1341
rect -24711 1284 -24670 1330
rect -23547 1284 -23509 1330
rect -24711 1281 -24210 1284
rect -24150 1281 -23509 1284
rect -24711 1261 -23509 1281
rect -23152 1524 -23097 1540
rect -23152 1418 -23145 1524
rect -23111 1418 -23097 1524
rect -23065 1539 -22615 1551
rect -23065 1505 -23049 1539
rect -23015 1505 -22857 1539
rect -22823 1538 -22615 1539
rect -22823 1505 -22665 1538
rect -23065 1504 -22665 1505
rect -22631 1504 -22615 1538
rect -23065 1483 -22615 1504
rect -22489 1539 -22039 1551
rect -22489 1505 -22473 1539
rect -22439 1505 -22281 1539
rect -22247 1505 -22089 1539
rect -22055 1505 -22039 1539
rect -22489 1483 -22039 1505
rect -22005 1524 -21950 1540
rect -23152 1352 -23097 1418
rect -22967 1438 -22902 1455
rect -22967 1404 -22953 1438
rect -22919 1404 -22902 1438
rect -22967 1352 -22902 1404
rect -22774 1438 -22327 1450
rect -22774 1404 -22761 1438
rect -22727 1404 -22569 1438
rect -22535 1404 -22377 1438
rect -22343 1404 -22327 1438
rect -22774 1386 -22327 1404
rect -22201 1438 -22136 1454
rect -22201 1404 -22185 1438
rect -22151 1404 -22136 1438
rect -22201 1352 -22136 1404
rect -22005 1418 -21993 1524
rect -21959 1418 -21950 1524
rect -22005 1352 -21950 1418
rect -23152 1341 -21950 1352
rect -23152 1330 -22651 1341
rect -22591 1330 -21950 1341
rect -23152 1284 -23111 1330
rect -21988 1284 -21950 1330
rect -21823 1407 -21714 1594
rect -21571 1705 -21366 1724
rect -21571 1597 -21527 1705
rect -21451 1679 -21366 1705
rect -20493 1679 -20378 1776
rect -20262 1789 -20148 1803
rect -19998 1789 -19983 1886
rect -20262 1773 -19983 1789
rect -19793 1845 -19004 1863
rect -19793 1837 -19150 1845
rect -19793 1784 -19756 1837
rect -19623 1792 -19150 1837
rect -19036 1792 -19004 1845
rect -19623 1784 -19004 1792
rect -20262 1710 -20091 1773
rect -19793 1764 -19004 1784
rect -18934 1844 -18819 1863
rect -18934 1776 -18916 1844
rect -18836 1776 -18819 1844
rect -18357 1828 -18339 1938
rect -18243 1830 -18222 1938
rect -15066 1938 -14931 1962
rect -16883 1903 -16692 1908
rect -16884 1893 -16692 1903
rect -16884 1886 -16782 1893
rect -16709 1886 -16692 1893
rect -18292 1828 -18222 1830
rect -18357 1808 -18222 1828
rect -18061 1845 -17272 1863
rect -18061 1837 -17418 1845
rect -21451 1597 -20378 1679
rect -21571 1593 -20378 1597
rect -20304 1673 -20091 1710
rect -20304 1618 -20293 1673
rect -20228 1618 -20091 1673
rect -20304 1594 -20091 1618
rect -20012 1698 -19807 1724
rect -20012 1601 -19972 1698
rect -19856 1679 -19807 1698
rect -18934 1679 -18819 1776
rect -18703 1710 -18423 1803
rect -18061 1784 -18024 1837
rect -17891 1792 -17418 1837
rect -17304 1792 -17272 1845
rect -17891 1784 -17272 1792
rect -18061 1764 -17272 1784
rect -17202 1844 -17087 1863
rect -17202 1776 -17184 1844
rect -17104 1776 -17087 1844
rect -16884 1803 -16857 1886
rect -19856 1601 -18819 1679
rect -20012 1593 -18819 1601
rect -18745 1673 -18423 1710
rect -18745 1618 -18734 1673
rect -18669 1618 -18423 1673
rect -18745 1594 -18423 1618
rect -21571 1581 -21366 1593
rect -20012 1581 -19807 1593
rect -21823 1321 -21814 1407
rect -21723 1321 -21714 1407
rect -21823 1309 -21714 1321
rect -21420 1524 -21365 1540
rect -21420 1418 -21413 1524
rect -21379 1418 -21365 1524
rect -21333 1539 -20883 1551
rect -21333 1505 -21317 1539
rect -21283 1505 -21125 1539
rect -21091 1538 -20883 1539
rect -21091 1505 -20933 1538
rect -21333 1504 -20933 1505
rect -20899 1504 -20883 1538
rect -21333 1483 -20883 1504
rect -20757 1539 -20307 1551
rect -20757 1505 -20741 1539
rect -20707 1505 -20549 1539
rect -20515 1505 -20357 1539
rect -20323 1505 -20307 1539
rect -20757 1483 -20307 1505
rect -20273 1524 -20218 1540
rect -21420 1352 -21365 1418
rect -21235 1438 -21170 1455
rect -21235 1404 -21221 1438
rect -21187 1404 -21170 1438
rect -21235 1352 -21170 1404
rect -21042 1438 -20595 1450
rect -21042 1404 -21029 1438
rect -20995 1404 -20837 1438
rect -20803 1404 -20645 1438
rect -20611 1404 -20595 1438
rect -21042 1386 -20595 1404
rect -20469 1438 -20404 1454
rect -20469 1404 -20453 1438
rect -20419 1404 -20404 1438
rect -20469 1352 -20404 1404
rect -20273 1418 -20261 1524
rect -20227 1418 -20218 1524
rect -20273 1352 -20218 1418
rect -21420 1341 -20218 1352
rect -21420 1330 -20919 1341
rect -20859 1330 -20218 1341
rect -23152 1281 -22651 1284
rect -22591 1281 -21950 1284
rect -23152 1261 -21950 1281
rect -21420 1284 -21379 1330
rect -20256 1284 -20218 1330
rect -21420 1281 -20919 1284
rect -20859 1281 -20218 1284
rect -21420 1261 -20218 1281
rect -19861 1524 -19806 1540
rect -19861 1418 -19854 1524
rect -19820 1418 -19806 1524
rect -19774 1539 -19324 1551
rect -19774 1505 -19758 1539
rect -19724 1505 -19566 1539
rect -19532 1538 -19324 1539
rect -19532 1505 -19374 1538
rect -19774 1504 -19374 1505
rect -19340 1504 -19324 1538
rect -19774 1483 -19324 1504
rect -19198 1539 -18748 1551
rect -19198 1505 -19182 1539
rect -19148 1505 -18990 1539
rect -18956 1505 -18798 1539
rect -18764 1505 -18748 1539
rect -19198 1483 -18748 1505
rect -18714 1524 -18659 1540
rect -19861 1352 -19806 1418
rect -19676 1438 -19611 1455
rect -19676 1404 -19662 1438
rect -19628 1404 -19611 1438
rect -19676 1352 -19611 1404
rect -19483 1438 -19036 1450
rect -19483 1404 -19470 1438
rect -19436 1404 -19278 1438
rect -19244 1404 -19086 1438
rect -19052 1404 -19036 1438
rect -19483 1386 -19036 1404
rect -18910 1438 -18845 1454
rect -18910 1404 -18894 1438
rect -18860 1404 -18845 1438
rect -18910 1352 -18845 1404
rect -18714 1418 -18702 1524
rect -18668 1418 -18659 1524
rect -18714 1352 -18659 1418
rect -19861 1341 -18659 1352
rect -19861 1330 -19360 1341
rect -19300 1330 -18659 1341
rect -19861 1284 -19820 1330
rect -18697 1284 -18659 1330
rect -18532 1407 -18423 1594
rect -18280 1705 -18075 1724
rect -18280 1597 -18236 1705
rect -18160 1679 -18075 1705
rect -17202 1679 -17087 1776
rect -16971 1789 -16857 1803
rect -16707 1789 -16692 1886
rect -16971 1773 -16692 1789
rect -16502 1845 -15713 1863
rect -16502 1837 -15859 1845
rect -16502 1784 -16465 1837
rect -16332 1792 -15859 1837
rect -15745 1792 -15713 1845
rect -16332 1784 -15713 1792
rect -16971 1710 -16800 1773
rect -16502 1764 -15713 1784
rect -15643 1844 -15528 1863
rect -15643 1776 -15625 1844
rect -15545 1776 -15528 1844
rect -15066 1828 -15048 1938
rect -14952 1830 -14931 1938
rect -11775 1938 -11640 1962
rect -13592 1903 -13401 1908
rect -13593 1893 -13401 1903
rect -13593 1886 -13491 1893
rect -13418 1886 -13401 1893
rect -15001 1828 -14931 1830
rect -15066 1808 -14931 1828
rect -14770 1845 -13981 1863
rect -14770 1837 -14127 1845
rect -18160 1597 -17087 1679
rect -18280 1593 -17087 1597
rect -17013 1673 -16800 1710
rect -17013 1618 -17002 1673
rect -16937 1618 -16800 1673
rect -17013 1594 -16800 1618
rect -16721 1698 -16516 1724
rect -16721 1601 -16681 1698
rect -16565 1679 -16516 1698
rect -15643 1679 -15528 1776
rect -15412 1710 -15132 1803
rect -14770 1784 -14733 1837
rect -14600 1792 -14127 1837
rect -14013 1792 -13981 1845
rect -14600 1784 -13981 1792
rect -14770 1764 -13981 1784
rect -13911 1844 -13796 1863
rect -13911 1776 -13893 1844
rect -13813 1776 -13796 1844
rect -13593 1803 -13566 1886
rect -16565 1601 -15528 1679
rect -16721 1593 -15528 1601
rect -15454 1673 -15132 1710
rect -15454 1618 -15443 1673
rect -15378 1618 -15132 1673
rect -15454 1594 -15132 1618
rect -18280 1581 -18075 1593
rect -16721 1581 -16516 1593
rect -18532 1321 -18523 1407
rect -18432 1321 -18423 1407
rect -18532 1309 -18423 1321
rect -18129 1524 -18074 1540
rect -18129 1418 -18122 1524
rect -18088 1418 -18074 1524
rect -18042 1539 -17592 1551
rect -18042 1505 -18026 1539
rect -17992 1505 -17834 1539
rect -17800 1538 -17592 1539
rect -17800 1505 -17642 1538
rect -18042 1504 -17642 1505
rect -17608 1504 -17592 1538
rect -18042 1483 -17592 1504
rect -17466 1539 -17016 1551
rect -17466 1505 -17450 1539
rect -17416 1505 -17258 1539
rect -17224 1505 -17066 1539
rect -17032 1505 -17016 1539
rect -17466 1483 -17016 1505
rect -16982 1524 -16927 1540
rect -18129 1352 -18074 1418
rect -17944 1438 -17879 1455
rect -17944 1404 -17930 1438
rect -17896 1404 -17879 1438
rect -17944 1352 -17879 1404
rect -17751 1438 -17304 1450
rect -17751 1404 -17738 1438
rect -17704 1404 -17546 1438
rect -17512 1404 -17354 1438
rect -17320 1404 -17304 1438
rect -17751 1386 -17304 1404
rect -17178 1438 -17113 1454
rect -17178 1404 -17162 1438
rect -17128 1404 -17113 1438
rect -17178 1352 -17113 1404
rect -16982 1418 -16970 1524
rect -16936 1418 -16927 1524
rect -16982 1352 -16927 1418
rect -18129 1341 -16927 1352
rect -18129 1330 -17628 1341
rect -17568 1330 -16927 1341
rect -19861 1281 -19360 1284
rect -19300 1281 -18659 1284
rect -19861 1261 -18659 1281
rect -18129 1284 -18088 1330
rect -16965 1284 -16927 1330
rect -18129 1281 -17628 1284
rect -17568 1281 -16927 1284
rect -18129 1261 -16927 1281
rect -16570 1524 -16515 1540
rect -16570 1418 -16563 1524
rect -16529 1418 -16515 1524
rect -16483 1539 -16033 1551
rect -16483 1505 -16467 1539
rect -16433 1505 -16275 1539
rect -16241 1538 -16033 1539
rect -16241 1505 -16083 1538
rect -16483 1504 -16083 1505
rect -16049 1504 -16033 1538
rect -16483 1483 -16033 1504
rect -15907 1539 -15457 1551
rect -15907 1505 -15891 1539
rect -15857 1505 -15699 1539
rect -15665 1505 -15507 1539
rect -15473 1505 -15457 1539
rect -15907 1483 -15457 1505
rect -15423 1524 -15368 1540
rect -16570 1352 -16515 1418
rect -16385 1438 -16320 1455
rect -16385 1404 -16371 1438
rect -16337 1404 -16320 1438
rect -16385 1352 -16320 1404
rect -16192 1438 -15745 1450
rect -16192 1404 -16179 1438
rect -16145 1404 -15987 1438
rect -15953 1404 -15795 1438
rect -15761 1404 -15745 1438
rect -16192 1386 -15745 1404
rect -15619 1438 -15554 1454
rect -15619 1404 -15603 1438
rect -15569 1404 -15554 1438
rect -15619 1352 -15554 1404
rect -15423 1418 -15411 1524
rect -15377 1418 -15368 1524
rect -15423 1352 -15368 1418
rect -16570 1341 -15368 1352
rect -16570 1330 -16069 1341
rect -16009 1330 -15368 1341
rect -16570 1284 -16529 1330
rect -15406 1284 -15368 1330
rect -15241 1407 -15132 1594
rect -14989 1705 -14784 1724
rect -14989 1597 -14945 1705
rect -14869 1679 -14784 1705
rect -13911 1679 -13796 1776
rect -13680 1789 -13566 1803
rect -13416 1789 -13401 1886
rect -13680 1773 -13401 1789
rect -13211 1845 -12422 1863
rect -13211 1837 -12568 1845
rect -13211 1784 -13174 1837
rect -13041 1792 -12568 1837
rect -12454 1792 -12422 1845
rect -13041 1784 -12422 1792
rect -13680 1710 -13509 1773
rect -13211 1764 -12422 1784
rect -12352 1844 -12237 1863
rect -12352 1776 -12334 1844
rect -12254 1776 -12237 1844
rect -11775 1828 -11757 1938
rect -11661 1830 -11640 1938
rect -8485 1938 -8350 1962
rect -10301 1903 -10110 1908
rect -10302 1893 -10110 1903
rect -10302 1886 -10200 1893
rect -10127 1886 -10110 1893
rect -11710 1828 -11640 1830
rect -11775 1808 -11640 1828
rect -11479 1845 -10690 1863
rect -11479 1837 -10836 1845
rect -14869 1597 -13796 1679
rect -14989 1593 -13796 1597
rect -13722 1673 -13509 1710
rect -13722 1618 -13711 1673
rect -13646 1618 -13509 1673
rect -13722 1594 -13509 1618
rect -13430 1698 -13225 1724
rect -13430 1601 -13390 1698
rect -13274 1679 -13225 1698
rect -12352 1679 -12237 1776
rect -12121 1710 -11841 1803
rect -11479 1784 -11442 1837
rect -11309 1792 -10836 1837
rect -10722 1792 -10690 1845
rect -11309 1784 -10690 1792
rect -11479 1764 -10690 1784
rect -10620 1844 -10505 1863
rect -10620 1776 -10602 1844
rect -10522 1776 -10505 1844
rect -10302 1803 -10275 1886
rect -13274 1601 -12237 1679
rect -13430 1593 -12237 1601
rect -12163 1673 -11841 1710
rect -12163 1618 -12152 1673
rect -12087 1618 -11841 1673
rect -12163 1594 -11841 1618
rect -14989 1581 -14784 1593
rect -13430 1581 -13225 1593
rect -15241 1321 -15232 1407
rect -15141 1321 -15132 1407
rect -15241 1309 -15132 1321
rect -14838 1524 -14783 1540
rect -14838 1418 -14831 1524
rect -14797 1418 -14783 1524
rect -14751 1539 -14301 1551
rect -14751 1505 -14735 1539
rect -14701 1505 -14543 1539
rect -14509 1538 -14301 1539
rect -14509 1505 -14351 1538
rect -14751 1504 -14351 1505
rect -14317 1504 -14301 1538
rect -14751 1483 -14301 1504
rect -14175 1539 -13725 1551
rect -14175 1505 -14159 1539
rect -14125 1505 -13967 1539
rect -13933 1505 -13775 1539
rect -13741 1505 -13725 1539
rect -14175 1483 -13725 1505
rect -13691 1524 -13636 1540
rect -14838 1352 -14783 1418
rect -14653 1438 -14588 1455
rect -14653 1404 -14639 1438
rect -14605 1404 -14588 1438
rect -14653 1352 -14588 1404
rect -14460 1438 -14013 1450
rect -14460 1404 -14447 1438
rect -14413 1404 -14255 1438
rect -14221 1404 -14063 1438
rect -14029 1404 -14013 1438
rect -14460 1386 -14013 1404
rect -13887 1438 -13822 1454
rect -13887 1404 -13871 1438
rect -13837 1404 -13822 1438
rect -13887 1352 -13822 1404
rect -13691 1418 -13679 1524
rect -13645 1418 -13636 1524
rect -13691 1352 -13636 1418
rect -14838 1341 -13636 1352
rect -14838 1330 -14337 1341
rect -14277 1330 -13636 1341
rect -16570 1281 -16069 1284
rect -16009 1281 -15368 1284
rect -16570 1261 -15368 1281
rect -14838 1284 -14797 1330
rect -13674 1284 -13636 1330
rect -14838 1281 -14337 1284
rect -14277 1281 -13636 1284
rect -14838 1261 -13636 1281
rect -13279 1524 -13224 1540
rect -13279 1418 -13272 1524
rect -13238 1418 -13224 1524
rect -13192 1539 -12742 1551
rect -13192 1505 -13176 1539
rect -13142 1505 -12984 1539
rect -12950 1538 -12742 1539
rect -12950 1505 -12792 1538
rect -13192 1504 -12792 1505
rect -12758 1504 -12742 1538
rect -13192 1483 -12742 1504
rect -12616 1539 -12166 1551
rect -12616 1505 -12600 1539
rect -12566 1505 -12408 1539
rect -12374 1505 -12216 1539
rect -12182 1505 -12166 1539
rect -12616 1483 -12166 1505
rect -12132 1524 -12077 1540
rect -13279 1352 -13224 1418
rect -13094 1438 -13029 1455
rect -13094 1404 -13080 1438
rect -13046 1404 -13029 1438
rect -13094 1352 -13029 1404
rect -12901 1438 -12454 1450
rect -12901 1404 -12888 1438
rect -12854 1404 -12696 1438
rect -12662 1404 -12504 1438
rect -12470 1404 -12454 1438
rect -12901 1386 -12454 1404
rect -12328 1438 -12263 1454
rect -12328 1404 -12312 1438
rect -12278 1404 -12263 1438
rect -12328 1352 -12263 1404
rect -12132 1418 -12120 1524
rect -12086 1418 -12077 1524
rect -12132 1352 -12077 1418
rect -13279 1341 -12077 1352
rect -13279 1330 -12778 1341
rect -12718 1330 -12077 1341
rect -13279 1284 -13238 1330
rect -12115 1284 -12077 1330
rect -11950 1407 -11841 1594
rect -11698 1705 -11493 1724
rect -11698 1597 -11654 1705
rect -11578 1679 -11493 1705
rect -10620 1679 -10505 1776
rect -10389 1789 -10275 1803
rect -10125 1789 -10110 1886
rect -10389 1773 -10110 1789
rect -9920 1845 -9131 1863
rect -9920 1837 -9277 1845
rect -9920 1784 -9883 1837
rect -9750 1792 -9277 1837
rect -9163 1792 -9131 1845
rect -9750 1784 -9131 1792
rect -10389 1710 -10218 1773
rect -9920 1764 -9131 1784
rect -9061 1844 -8946 1863
rect -9061 1776 -9043 1844
rect -8963 1776 -8946 1844
rect -8485 1828 -8467 1938
rect -8371 1830 -8350 1938
rect -5194 1938 -5059 1962
rect -7011 1903 -6820 1908
rect -7012 1893 -6820 1903
rect -7012 1886 -6910 1893
rect -6837 1886 -6820 1893
rect -8420 1828 -8350 1830
rect -8485 1808 -8350 1828
rect -8189 1845 -7400 1863
rect -8189 1837 -7546 1845
rect -11578 1597 -10505 1679
rect -11698 1593 -10505 1597
rect -10431 1673 -10218 1710
rect -10431 1618 -10420 1673
rect -10355 1618 -10218 1673
rect -10431 1594 -10218 1618
rect -10139 1698 -9934 1724
rect -10139 1601 -10099 1698
rect -9983 1679 -9934 1698
rect -9061 1679 -8946 1776
rect -8830 1710 -8550 1803
rect -8189 1784 -8152 1837
rect -8019 1792 -7546 1837
rect -7432 1792 -7400 1845
rect -8019 1784 -7400 1792
rect -8189 1764 -7400 1784
rect -7330 1844 -7215 1863
rect -7330 1776 -7312 1844
rect -7232 1776 -7215 1844
rect -7012 1803 -6985 1886
rect -9983 1601 -8946 1679
rect -10139 1593 -8946 1601
rect -8872 1673 -8550 1710
rect -8872 1618 -8861 1673
rect -8796 1618 -8550 1673
rect -8872 1594 -8550 1618
rect -11698 1581 -11493 1593
rect -10139 1581 -9934 1593
rect -11950 1321 -11941 1407
rect -11850 1321 -11841 1407
rect -11950 1309 -11841 1321
rect -11547 1524 -11492 1540
rect -11547 1418 -11540 1524
rect -11506 1418 -11492 1524
rect -11460 1539 -11010 1551
rect -11460 1505 -11444 1539
rect -11410 1505 -11252 1539
rect -11218 1538 -11010 1539
rect -11218 1505 -11060 1538
rect -11460 1504 -11060 1505
rect -11026 1504 -11010 1538
rect -11460 1483 -11010 1504
rect -10884 1539 -10434 1551
rect -10884 1505 -10868 1539
rect -10834 1505 -10676 1539
rect -10642 1505 -10484 1539
rect -10450 1505 -10434 1539
rect -10884 1483 -10434 1505
rect -10400 1524 -10345 1540
rect -11547 1352 -11492 1418
rect -11362 1438 -11297 1455
rect -11362 1404 -11348 1438
rect -11314 1404 -11297 1438
rect -11362 1352 -11297 1404
rect -11169 1438 -10722 1450
rect -11169 1404 -11156 1438
rect -11122 1404 -10964 1438
rect -10930 1404 -10772 1438
rect -10738 1404 -10722 1438
rect -11169 1386 -10722 1404
rect -10596 1438 -10531 1454
rect -10596 1404 -10580 1438
rect -10546 1404 -10531 1438
rect -10596 1352 -10531 1404
rect -10400 1418 -10388 1524
rect -10354 1418 -10345 1524
rect -10400 1352 -10345 1418
rect -11547 1341 -10345 1352
rect -11547 1330 -11046 1341
rect -10986 1330 -10345 1341
rect -13279 1281 -12778 1284
rect -12718 1281 -12077 1284
rect -13279 1261 -12077 1281
rect -11547 1284 -11506 1330
rect -10383 1284 -10345 1330
rect -11547 1281 -11046 1284
rect -10986 1281 -10345 1284
rect -11547 1261 -10345 1281
rect -9988 1524 -9933 1540
rect -9988 1418 -9981 1524
rect -9947 1418 -9933 1524
rect -9901 1539 -9451 1551
rect -9901 1505 -9885 1539
rect -9851 1505 -9693 1539
rect -9659 1538 -9451 1539
rect -9659 1505 -9501 1538
rect -9901 1504 -9501 1505
rect -9467 1504 -9451 1538
rect -9901 1483 -9451 1504
rect -9325 1539 -8875 1551
rect -9325 1505 -9309 1539
rect -9275 1505 -9117 1539
rect -9083 1505 -8925 1539
rect -8891 1505 -8875 1539
rect -9325 1483 -8875 1505
rect -8841 1524 -8786 1540
rect -9988 1352 -9933 1418
rect -9803 1438 -9738 1455
rect -9803 1404 -9789 1438
rect -9755 1404 -9738 1438
rect -9803 1352 -9738 1404
rect -9610 1438 -9163 1450
rect -9610 1404 -9597 1438
rect -9563 1404 -9405 1438
rect -9371 1404 -9213 1438
rect -9179 1404 -9163 1438
rect -9610 1386 -9163 1404
rect -9037 1438 -8972 1454
rect -9037 1404 -9021 1438
rect -8987 1404 -8972 1438
rect -9037 1352 -8972 1404
rect -8841 1418 -8829 1524
rect -8795 1418 -8786 1524
rect -8841 1352 -8786 1418
rect -9988 1341 -8786 1352
rect -9988 1330 -9487 1341
rect -9427 1330 -8786 1341
rect -9988 1284 -9947 1330
rect -8824 1284 -8786 1330
rect -8659 1407 -8550 1594
rect -8408 1705 -8203 1724
rect -8408 1597 -8364 1705
rect -8288 1679 -8203 1705
rect -7330 1679 -7215 1776
rect -7099 1789 -6985 1803
rect -6835 1789 -6820 1886
rect -7099 1773 -6820 1789
rect -6630 1845 -5841 1863
rect -6630 1837 -5987 1845
rect -6630 1784 -6593 1837
rect -6460 1792 -5987 1837
rect -5873 1792 -5841 1845
rect -6460 1784 -5841 1792
rect -7099 1710 -6928 1773
rect -6630 1764 -5841 1784
rect -5771 1844 -5656 1863
rect -5771 1776 -5753 1844
rect -5673 1776 -5656 1844
rect -5194 1828 -5176 1938
rect -5080 1830 -5059 1938
rect -1903 1938 -1768 1962
rect -3720 1903 -3529 1908
rect -3721 1893 -3529 1903
rect -3721 1886 -3619 1893
rect -3546 1886 -3529 1893
rect -5129 1828 -5059 1830
rect -5194 1808 -5059 1828
rect -4898 1845 -4109 1863
rect -4898 1837 -4255 1845
rect -8288 1597 -7215 1679
rect -8408 1593 -7215 1597
rect -7141 1673 -6928 1710
rect -7141 1618 -7130 1673
rect -7065 1618 -6928 1673
rect -7141 1594 -6928 1618
rect -6849 1698 -6644 1724
rect -6849 1601 -6809 1698
rect -6693 1679 -6644 1698
rect -5771 1679 -5656 1776
rect -5540 1710 -5260 1803
rect -4898 1784 -4861 1837
rect -4728 1792 -4255 1837
rect -4141 1792 -4109 1845
rect -4728 1784 -4109 1792
rect -4898 1764 -4109 1784
rect -4039 1844 -3924 1863
rect -4039 1776 -4021 1844
rect -3941 1776 -3924 1844
rect -3721 1803 -3694 1886
rect -6693 1601 -5656 1679
rect -6849 1593 -5656 1601
rect -5582 1673 -5260 1710
rect -5582 1618 -5571 1673
rect -5506 1618 -5260 1673
rect -5582 1594 -5260 1618
rect -8408 1581 -8203 1593
rect -6849 1581 -6644 1593
rect -8659 1321 -8650 1407
rect -8559 1321 -8550 1407
rect -8659 1309 -8550 1321
rect -8257 1524 -8202 1540
rect -8257 1418 -8250 1524
rect -8216 1418 -8202 1524
rect -8170 1539 -7720 1551
rect -8170 1505 -8154 1539
rect -8120 1505 -7962 1539
rect -7928 1538 -7720 1539
rect -7928 1505 -7770 1538
rect -8170 1504 -7770 1505
rect -7736 1504 -7720 1538
rect -8170 1483 -7720 1504
rect -7594 1539 -7144 1551
rect -7594 1505 -7578 1539
rect -7544 1505 -7386 1539
rect -7352 1505 -7194 1539
rect -7160 1505 -7144 1539
rect -7594 1483 -7144 1505
rect -7110 1524 -7055 1540
rect -8257 1352 -8202 1418
rect -8072 1438 -8007 1455
rect -8072 1404 -8058 1438
rect -8024 1404 -8007 1438
rect -8072 1352 -8007 1404
rect -7879 1438 -7432 1450
rect -7879 1404 -7866 1438
rect -7832 1404 -7674 1438
rect -7640 1404 -7482 1438
rect -7448 1404 -7432 1438
rect -7879 1386 -7432 1404
rect -7306 1438 -7241 1454
rect -7306 1404 -7290 1438
rect -7256 1404 -7241 1438
rect -7306 1352 -7241 1404
rect -7110 1418 -7098 1524
rect -7064 1418 -7055 1524
rect -7110 1352 -7055 1418
rect -8257 1341 -7055 1352
rect -8257 1330 -7756 1341
rect -7696 1330 -7055 1341
rect -9988 1281 -9487 1284
rect -9427 1281 -8786 1284
rect -9988 1261 -8786 1281
rect -8257 1284 -8216 1330
rect -7093 1284 -7055 1330
rect -8257 1281 -7756 1284
rect -7696 1281 -7055 1284
rect -8257 1261 -7055 1281
rect -6698 1524 -6643 1540
rect -6698 1418 -6691 1524
rect -6657 1418 -6643 1524
rect -6611 1539 -6161 1551
rect -6611 1505 -6595 1539
rect -6561 1505 -6403 1539
rect -6369 1538 -6161 1539
rect -6369 1505 -6211 1538
rect -6611 1504 -6211 1505
rect -6177 1504 -6161 1538
rect -6611 1483 -6161 1504
rect -6035 1539 -5585 1551
rect -6035 1505 -6019 1539
rect -5985 1505 -5827 1539
rect -5793 1505 -5635 1539
rect -5601 1505 -5585 1539
rect -6035 1483 -5585 1505
rect -5551 1524 -5496 1540
rect -6698 1352 -6643 1418
rect -6513 1438 -6448 1455
rect -6513 1404 -6499 1438
rect -6465 1404 -6448 1438
rect -6513 1352 -6448 1404
rect -6320 1438 -5873 1450
rect -6320 1404 -6307 1438
rect -6273 1404 -6115 1438
rect -6081 1404 -5923 1438
rect -5889 1404 -5873 1438
rect -6320 1386 -5873 1404
rect -5747 1438 -5682 1454
rect -5747 1404 -5731 1438
rect -5697 1404 -5682 1438
rect -5747 1352 -5682 1404
rect -5551 1418 -5539 1524
rect -5505 1418 -5496 1524
rect -5551 1352 -5496 1418
rect -6698 1341 -5496 1352
rect -6698 1330 -6197 1341
rect -6137 1330 -5496 1341
rect -6698 1284 -6657 1330
rect -5534 1284 -5496 1330
rect -5369 1407 -5260 1594
rect -5117 1705 -4912 1724
rect -5117 1597 -5073 1705
rect -4997 1679 -4912 1705
rect -4039 1679 -3924 1776
rect -3808 1789 -3694 1803
rect -3544 1789 -3529 1886
rect -3808 1773 -3529 1789
rect -3339 1845 -2550 1863
rect -3339 1837 -2696 1845
rect -3339 1784 -3302 1837
rect -3169 1792 -2696 1837
rect -2582 1792 -2550 1845
rect -3169 1784 -2550 1792
rect -3808 1710 -3637 1773
rect -3339 1764 -2550 1784
rect -2480 1844 -2365 1863
rect -2480 1776 -2462 1844
rect -2382 1776 -2365 1844
rect -1903 1828 -1885 1938
rect -1789 1830 -1768 1938
rect -429 1903 -238 1908
rect -430 1893 -238 1903
rect -430 1886 -328 1893
rect -255 1886 -238 1893
rect -1838 1828 -1768 1830
rect -1903 1808 -1768 1828
rect -1607 1845 -818 1863
rect -1607 1837 -964 1845
rect -4997 1597 -3924 1679
rect -5117 1593 -3924 1597
rect -3850 1673 -3637 1710
rect -3850 1618 -3839 1673
rect -3774 1618 -3637 1673
rect -3850 1594 -3637 1618
rect -3558 1698 -3353 1724
rect -3558 1601 -3518 1698
rect -3402 1679 -3353 1698
rect -2480 1679 -2365 1776
rect -2249 1710 -1969 1803
rect -1607 1784 -1570 1837
rect -1437 1792 -964 1837
rect -850 1792 -818 1845
rect -1437 1784 -818 1792
rect -1607 1764 -818 1784
rect -748 1844 -633 1863
rect -748 1776 -730 1844
rect -650 1776 -633 1844
rect -430 1803 -403 1886
rect -3402 1601 -2365 1679
rect -3558 1593 -2365 1601
rect -2291 1673 -1969 1710
rect -2291 1618 -2280 1673
rect -2215 1618 -1969 1673
rect -2291 1594 -1969 1618
rect -5117 1581 -4912 1593
rect -3558 1581 -3353 1593
rect -5369 1321 -5360 1407
rect -5269 1321 -5260 1407
rect -5369 1309 -5260 1321
rect -4966 1524 -4911 1540
rect -4966 1418 -4959 1524
rect -4925 1418 -4911 1524
rect -4879 1539 -4429 1551
rect -4879 1505 -4863 1539
rect -4829 1505 -4671 1539
rect -4637 1538 -4429 1539
rect -4637 1505 -4479 1538
rect -4879 1504 -4479 1505
rect -4445 1504 -4429 1538
rect -4879 1483 -4429 1504
rect -4303 1539 -3853 1551
rect -4303 1505 -4287 1539
rect -4253 1505 -4095 1539
rect -4061 1505 -3903 1539
rect -3869 1505 -3853 1539
rect -4303 1483 -3853 1505
rect -3819 1524 -3764 1540
rect -4966 1352 -4911 1418
rect -4781 1438 -4716 1455
rect -4781 1404 -4767 1438
rect -4733 1404 -4716 1438
rect -4781 1352 -4716 1404
rect -4588 1438 -4141 1450
rect -4588 1404 -4575 1438
rect -4541 1404 -4383 1438
rect -4349 1404 -4191 1438
rect -4157 1404 -4141 1438
rect -4588 1386 -4141 1404
rect -4015 1438 -3950 1454
rect -4015 1404 -3999 1438
rect -3965 1404 -3950 1438
rect -4015 1352 -3950 1404
rect -3819 1418 -3807 1524
rect -3773 1418 -3764 1524
rect -3819 1352 -3764 1418
rect -4966 1341 -3764 1352
rect -4966 1330 -4465 1341
rect -4405 1330 -3764 1341
rect -6698 1281 -6197 1284
rect -6137 1281 -5496 1284
rect -6698 1261 -5496 1281
rect -4966 1284 -4925 1330
rect -3802 1284 -3764 1330
rect -4966 1281 -4465 1284
rect -4405 1281 -3764 1284
rect -4966 1261 -3764 1281
rect -3407 1524 -3352 1540
rect -3407 1418 -3400 1524
rect -3366 1418 -3352 1524
rect -3320 1539 -2870 1551
rect -3320 1505 -3304 1539
rect -3270 1505 -3112 1539
rect -3078 1538 -2870 1539
rect -3078 1505 -2920 1538
rect -3320 1504 -2920 1505
rect -2886 1504 -2870 1538
rect -3320 1483 -2870 1504
rect -2744 1539 -2294 1551
rect -2744 1505 -2728 1539
rect -2694 1505 -2536 1539
rect -2502 1505 -2344 1539
rect -2310 1505 -2294 1539
rect -2744 1483 -2294 1505
rect -2260 1524 -2205 1540
rect -3407 1352 -3352 1418
rect -3222 1438 -3157 1455
rect -3222 1404 -3208 1438
rect -3174 1404 -3157 1438
rect -3222 1352 -3157 1404
rect -3029 1438 -2582 1450
rect -3029 1404 -3016 1438
rect -2982 1404 -2824 1438
rect -2790 1404 -2632 1438
rect -2598 1404 -2582 1438
rect -3029 1386 -2582 1404
rect -2456 1438 -2391 1454
rect -2456 1404 -2440 1438
rect -2406 1404 -2391 1438
rect -2456 1352 -2391 1404
rect -2260 1418 -2248 1524
rect -2214 1418 -2205 1524
rect -2260 1352 -2205 1418
rect -3407 1341 -2205 1352
rect -3407 1330 -2906 1341
rect -2846 1330 -2205 1341
rect -3407 1284 -3366 1330
rect -2243 1284 -2205 1330
rect -2078 1407 -1969 1594
rect -1826 1705 -1621 1724
rect -1826 1597 -1782 1705
rect -1706 1679 -1621 1705
rect -748 1679 -633 1776
rect -517 1789 -403 1803
rect -253 1789 -238 1886
rect -517 1773 -238 1789
rect -48 1845 741 1863
rect -48 1837 595 1845
rect -48 1784 -11 1837
rect 122 1792 595 1837
rect 709 1792 741 1845
rect 122 1784 741 1792
rect -517 1710 -346 1773
rect -48 1764 741 1784
rect 811 1844 926 1863
rect 811 1776 829 1844
rect 909 1776 926 1844
rect -1706 1597 -633 1679
rect -1826 1593 -633 1597
rect -559 1673 -346 1710
rect -559 1618 -548 1673
rect -483 1618 -346 1673
rect -559 1594 -346 1618
rect -267 1698 -62 1724
rect -267 1601 -227 1698
rect -111 1679 -62 1698
rect 811 1679 926 1776
rect 1042 1710 1322 1803
rect -111 1601 926 1679
rect -267 1593 926 1601
rect 1000 1673 1322 1710
rect 1000 1618 1011 1673
rect 1076 1618 1322 1673
rect 1000 1594 1322 1618
rect -1826 1581 -1621 1593
rect -267 1581 -62 1593
rect -2078 1321 -2069 1407
rect -1978 1321 -1969 1407
rect -2078 1309 -1969 1321
rect -1675 1524 -1620 1540
rect -1675 1418 -1668 1524
rect -1634 1418 -1620 1524
rect -1588 1539 -1138 1551
rect -1588 1505 -1572 1539
rect -1538 1505 -1380 1539
rect -1346 1538 -1138 1539
rect -1346 1505 -1188 1538
rect -1588 1504 -1188 1505
rect -1154 1504 -1138 1538
rect -1588 1483 -1138 1504
rect -1012 1539 -562 1551
rect -1012 1505 -996 1539
rect -962 1505 -804 1539
rect -770 1505 -612 1539
rect -578 1505 -562 1539
rect -1012 1483 -562 1505
rect -528 1524 -473 1540
rect -1675 1352 -1620 1418
rect -1490 1438 -1425 1455
rect -1490 1404 -1476 1438
rect -1442 1404 -1425 1438
rect -1490 1352 -1425 1404
rect -1297 1438 -850 1450
rect -1297 1404 -1284 1438
rect -1250 1404 -1092 1438
rect -1058 1404 -900 1438
rect -866 1404 -850 1438
rect -1297 1386 -850 1404
rect -724 1438 -659 1454
rect -724 1404 -708 1438
rect -674 1404 -659 1438
rect -724 1352 -659 1404
rect -528 1418 -516 1524
rect -482 1418 -473 1524
rect -528 1352 -473 1418
rect -1675 1341 -473 1352
rect -1675 1330 -1174 1341
rect -1114 1330 -473 1341
rect -3407 1281 -2906 1284
rect -2846 1281 -2205 1284
rect -3407 1261 -2205 1281
rect -1675 1284 -1634 1330
rect -511 1284 -473 1330
rect -1675 1281 -1174 1284
rect -1114 1281 -473 1284
rect -1675 1261 -473 1281
rect -116 1524 -61 1540
rect -116 1418 -109 1524
rect -75 1418 -61 1524
rect -29 1539 421 1551
rect -29 1505 -13 1539
rect 21 1505 179 1539
rect 213 1538 421 1539
rect 213 1505 371 1538
rect -29 1504 371 1505
rect 405 1504 421 1538
rect -29 1483 421 1504
rect 547 1539 997 1551
rect 547 1505 563 1539
rect 597 1505 755 1539
rect 789 1505 947 1539
rect 981 1505 997 1539
rect 547 1483 997 1505
rect 1031 1524 1086 1540
rect -116 1352 -61 1418
rect 69 1438 134 1455
rect 69 1404 83 1438
rect 117 1404 134 1438
rect 69 1352 134 1404
rect 262 1438 709 1450
rect 262 1404 275 1438
rect 309 1404 467 1438
rect 501 1404 659 1438
rect 693 1404 709 1438
rect 262 1386 709 1404
rect 835 1438 900 1454
rect 835 1404 851 1438
rect 885 1404 900 1438
rect 835 1352 900 1404
rect 1031 1418 1043 1524
rect 1077 1418 1086 1524
rect 1031 1352 1086 1418
rect -116 1341 1086 1352
rect -116 1330 385 1341
rect 445 1330 1086 1341
rect -116 1284 -75 1330
rect 1048 1284 1086 1330
rect 1213 1407 1322 1594
rect 1213 1321 1222 1407
rect 1313 1321 1322 1407
rect 1213 1309 1322 1321
rect -116 1281 385 1284
rect 445 1281 1086 1284
rect -116 1261 1086 1281
rect 1425 1208 1516 3365
rect 5559 3289 5628 3366
rect 5558 3230 5628 3289
rect 5658 3373 5858 3380
rect 5658 3339 5670 3373
rect 5846 3339 5858 3373
rect 5886 3366 5970 3427
rect 5658 3271 5858 3339
rect 5658 3237 5689 3271
rect 5821 3237 5858 3271
rect 5658 3230 5858 3237
rect 5901 3314 5970 3366
rect 5559 3114 5628 3230
rect 5703 3228 5823 3230
rect 5703 3176 5734 3228
rect 5786 3176 5823 3228
rect 5901 3224 5970 3245
rect 5998 3637 6017 3810
rect 6051 3637 6067 3810
rect 6098 3877 6104 3911
rect 6183 3907 6312 3911
rect 6538 3924 7357 3937
rect 6538 3911 6752 3924
rect 6183 3877 6189 3907
rect 6438 3879 6507 3885
rect 6098 3719 6189 3877
rect 6098 3685 6104 3719
rect 6183 3685 6189 3719
rect 6098 3669 6189 3685
rect 6221 3815 6410 3879
rect 6221 3781 6227 3815
rect 6304 3781 6410 3815
rect 5998 3417 6067 3637
rect 6221 3623 6410 3781
rect 6098 3589 6227 3623
rect 6304 3589 6410 3623
rect 6098 3461 6410 3589
rect 6098 3427 6110 3461
rect 6286 3427 6410 3461
rect 6098 3421 6298 3427
rect 5998 3383 6017 3417
rect 6051 3383 6067 3417
rect 5703 3145 5823 3176
rect 5559 3045 5901 3114
rect 5559 3033 5628 3045
rect -25060 1192 -23687 1208
rect -25060 1123 -23802 1192
rect -23703 1123 -23687 1192
rect -25060 1117 -23687 1123
rect -23304 1196 -20396 1208
rect -23304 1130 -23290 1196
rect -23219 1192 -20396 1196
rect -23219 1130 -20511 1192
rect -23304 1123 -20511 1130
rect -20412 1123 -20396 1192
rect -23304 1117 -20396 1123
rect -20013 1196 -17105 1208
rect -20013 1130 -19999 1196
rect -19928 1192 -17105 1196
rect -19928 1130 -17220 1192
rect -20013 1123 -17220 1130
rect -17121 1123 -17105 1192
rect -20013 1117 -17105 1123
rect -16722 1196 -13814 1208
rect -16722 1130 -16708 1196
rect -16637 1192 -13814 1196
rect -16637 1130 -13929 1192
rect -16722 1123 -13929 1130
rect -13830 1123 -13814 1192
rect -16722 1117 -13814 1123
rect -13431 1196 -10523 1208
rect -13431 1130 -13417 1196
rect -13346 1192 -10523 1196
rect -13346 1130 -10638 1192
rect -13431 1123 -10638 1130
rect -10539 1123 -10523 1192
rect -13431 1117 -10523 1123
rect -10140 1196 -7233 1208
rect -10140 1130 -10126 1196
rect -10055 1192 -7233 1196
rect -10055 1130 -7348 1192
rect -10140 1123 -7348 1130
rect -7249 1123 -7233 1192
rect -10140 1117 -7233 1123
rect -6850 1196 -3942 1208
rect -6850 1130 -6836 1196
rect -6765 1192 -3942 1196
rect -6765 1130 -4057 1192
rect -6850 1123 -4057 1130
rect -3958 1123 -3942 1192
rect -6850 1117 -3942 1123
rect -3559 1196 -651 1208
rect -3559 1130 -3545 1196
rect -3474 1192 -651 1196
rect -3474 1130 -766 1192
rect -3559 1123 -766 1130
rect -667 1123 -651 1192
rect -3559 1117 -651 1123
rect -268 1196 1516 1208
rect -268 1130 -254 1196
rect -183 1130 1516 1196
rect -268 1117 1516 1130
rect 1922 2519 2013 2538
rect 1922 2453 1934 2519
rect 2000 2453 2013 2519
rect -25060 -123 -24969 1117
rect -24421 1001 -24147 1010
rect -24421 995 -24412 1001
rect -24598 988 -24412 995
rect -24156 995 -24147 1001
rect -23132 1001 -22858 1010
rect -23132 995 -23123 1001
rect -24156 988 -23964 995
rect -24598 941 -24569 988
rect -24000 941 -23964 988
rect -24598 929 -24412 941
rect -24156 929 -23964 941
rect -24598 875 -23964 929
rect -23489 988 -23123 995
rect -22867 995 -22858 1001
rect -22415 1001 -22141 1010
rect -22415 995 -22406 1001
rect -23489 941 -23460 988
rect -23489 929 -23123 941
rect -22867 929 -22855 995
rect -23489 875 -22855 929
rect -22607 988 -22406 995
rect -22150 995 -22141 1001
rect -21130 1001 -20856 1010
rect -21130 995 -21121 1001
rect -22150 988 -21973 995
rect -22607 941 -22578 988
rect -22009 941 -21973 988
rect -22607 929 -22406 941
rect -22150 929 -21973 941
rect -22607 875 -21973 929
rect -21307 988 -21121 995
rect -20865 995 -20856 1001
rect -19841 1001 -19567 1010
rect -19841 995 -19832 1001
rect -20865 988 -20673 995
rect -21307 941 -21278 988
rect -20709 941 -20673 988
rect -21307 929 -21121 941
rect -20865 929 -20673 941
rect -21307 875 -20673 929
rect -20198 988 -19832 995
rect -19576 995 -19567 1001
rect -19124 1001 -18850 1010
rect -19124 995 -19115 1001
rect -20198 941 -20169 988
rect -20198 929 -19832 941
rect -19576 929 -19564 995
rect -20198 875 -19564 929
rect -19316 988 -19115 995
rect -18859 995 -18850 1001
rect -17839 1001 -17565 1010
rect -17839 995 -17830 1001
rect -18859 988 -18682 995
rect -19316 941 -19287 988
rect -18718 941 -18682 988
rect -19316 929 -19115 941
rect -18859 929 -18682 941
rect -19316 875 -18682 929
rect -18016 988 -17830 995
rect -17574 995 -17565 1001
rect -16550 1001 -16276 1010
rect -16550 995 -16541 1001
rect -17574 988 -17382 995
rect -18016 941 -17987 988
rect -17418 941 -17382 988
rect -18016 929 -17830 941
rect -17574 929 -17382 941
rect -18016 875 -17382 929
rect -16907 988 -16541 995
rect -16285 995 -16276 1001
rect -15833 1001 -15559 1010
rect -15833 995 -15824 1001
rect -16907 941 -16878 988
rect -16907 929 -16541 941
rect -16285 929 -16273 995
rect -16907 875 -16273 929
rect -16025 988 -15824 995
rect -15568 995 -15559 1001
rect -14548 1001 -14274 1010
rect -14548 995 -14539 1001
rect -15568 988 -15391 995
rect -16025 941 -15996 988
rect -15427 941 -15391 988
rect -16025 929 -15824 941
rect -15568 929 -15391 941
rect -16025 875 -15391 929
rect -14725 988 -14539 995
rect -14283 995 -14274 1001
rect -13259 1001 -12985 1010
rect -13259 995 -13250 1001
rect -14283 988 -14091 995
rect -14725 941 -14696 988
rect -14127 941 -14091 988
rect -14725 929 -14539 941
rect -14283 929 -14091 941
rect -14725 875 -14091 929
rect -13616 988 -13250 995
rect -12994 995 -12985 1001
rect -12542 1001 -12268 1010
rect -12542 995 -12533 1001
rect -13616 941 -13587 988
rect -13616 929 -13250 941
rect -12994 929 -12982 995
rect -13616 875 -12982 929
rect -12734 988 -12533 995
rect -12277 995 -12268 1001
rect -11257 1001 -10983 1010
rect -11257 995 -11248 1001
rect -12277 988 -12100 995
rect -12734 941 -12705 988
rect -12136 941 -12100 988
rect -12734 929 -12533 941
rect -12277 929 -12100 941
rect -12734 875 -12100 929
rect -11434 988 -11248 995
rect -10992 995 -10983 1001
rect -9968 1001 -9694 1010
rect -9968 995 -9959 1001
rect -10992 988 -10800 995
rect -11434 941 -11405 988
rect -10836 941 -10800 988
rect -11434 929 -11248 941
rect -10992 929 -10800 941
rect -11434 875 -10800 929
rect -10325 988 -9959 995
rect -9703 995 -9694 1001
rect -9251 1001 -8977 1010
rect -9251 995 -9242 1001
rect -10325 941 -10296 988
rect -10325 929 -9959 941
rect -9703 929 -9691 995
rect -10325 875 -9691 929
rect -9443 988 -9242 995
rect -8986 995 -8977 1001
rect -7967 1001 -7693 1010
rect -7967 995 -7958 1001
rect -8986 988 -8809 995
rect -9443 941 -9414 988
rect -8845 941 -8809 988
rect -9443 929 -9242 941
rect -8986 929 -8809 941
rect -9443 875 -8809 929
rect -8144 988 -7958 995
rect -7702 995 -7693 1001
rect -6678 1001 -6404 1010
rect -6678 995 -6669 1001
rect -7702 988 -7510 995
rect -8144 941 -8115 988
rect -7546 941 -7510 988
rect -8144 929 -7958 941
rect -7702 929 -7510 941
rect -8144 875 -7510 929
rect -7035 988 -6669 995
rect -6413 995 -6404 1001
rect -5961 1001 -5687 1010
rect -5961 995 -5952 1001
rect -7035 941 -7006 988
rect -7035 929 -6669 941
rect -6413 929 -6401 995
rect -7035 875 -6401 929
rect -6153 988 -5952 995
rect -5696 995 -5687 1001
rect -4676 1001 -4402 1010
rect -4676 995 -4667 1001
rect -5696 988 -5519 995
rect -6153 941 -6124 988
rect -5555 941 -5519 988
rect -6153 929 -5952 941
rect -5696 929 -5519 941
rect -6153 875 -5519 929
rect -4853 988 -4667 995
rect -4411 995 -4402 1001
rect -3387 1001 -3113 1010
rect -3387 995 -3378 1001
rect -4411 988 -4219 995
rect -4853 941 -4824 988
rect -4255 941 -4219 988
rect -4853 929 -4667 941
rect -4411 929 -4219 941
rect -4853 875 -4219 929
rect -3744 988 -3378 995
rect -3122 995 -3113 1001
rect -2670 1001 -2396 1010
rect -2670 995 -2661 1001
rect -3744 941 -3715 988
rect -3744 929 -3378 941
rect -3122 929 -3110 995
rect -3744 875 -3110 929
rect -2862 988 -2661 995
rect -2405 995 -2396 1001
rect -1385 1001 -1111 1010
rect -1385 995 -1376 1001
rect -2405 988 -2228 995
rect -2862 941 -2833 988
rect -2264 941 -2228 988
rect -2862 929 -2661 941
rect -2405 929 -2228 941
rect -2862 875 -2228 929
rect -1562 988 -1376 995
rect -1120 995 -1111 1001
rect -96 1001 178 1010
rect -96 995 -87 1001
rect -1120 988 -928 995
rect -1562 941 -1533 988
rect -964 941 -928 988
rect -1562 929 -1376 941
rect -1120 929 -928 941
rect -1562 875 -928 929
rect -453 988 -87 995
rect 169 995 178 1001
rect 621 1001 895 1010
rect 621 995 630 1001
rect -453 941 -424 988
rect -453 929 -87 941
rect 169 929 181 995
rect -453 875 181 929
rect 429 988 630 995
rect 886 995 895 1001
rect 886 988 1063 995
rect 429 941 458 988
rect 1027 941 1063 988
rect 429 929 630 941
rect 886 929 1063 941
rect 429 875 1063 929
rect -24598 869 -23963 875
rect -24598 789 -24585 869
rect -24551 789 -24393 869
rect -24359 789 -24201 869
rect -24167 789 -24009 869
rect -23975 789 -23963 869
rect -24598 783 -23963 789
rect -23489 869 -22854 875
rect -23489 789 -23476 869
rect -23442 789 -23284 869
rect -23250 789 -23092 869
rect -23058 789 -22900 869
rect -22866 789 -22854 869
rect -23489 783 -22854 789
rect -22607 869 -21972 875
rect -22607 789 -22594 869
rect -22560 789 -22402 869
rect -22368 789 -22210 869
rect -22176 789 -22018 869
rect -21984 789 -21972 869
rect -22607 783 -21972 789
rect -21307 869 -20672 875
rect -21307 789 -21294 869
rect -21260 789 -21102 869
rect -21068 789 -20910 869
rect -20876 789 -20718 869
rect -20684 789 -20672 869
rect -21307 783 -20672 789
rect -20198 869 -19563 875
rect -20198 789 -20185 869
rect -20151 789 -19993 869
rect -19959 789 -19801 869
rect -19767 789 -19609 869
rect -19575 789 -19563 869
rect -20198 783 -19563 789
rect -19316 869 -18681 875
rect -19316 789 -19303 869
rect -19269 789 -19111 869
rect -19077 789 -18919 869
rect -18885 789 -18727 869
rect -18693 789 -18681 869
rect -19316 783 -18681 789
rect -18016 869 -17381 875
rect -18016 789 -18003 869
rect -17969 789 -17811 869
rect -17777 789 -17619 869
rect -17585 789 -17427 869
rect -17393 789 -17381 869
rect -18016 783 -17381 789
rect -16907 869 -16272 875
rect -16907 789 -16894 869
rect -16860 789 -16702 869
rect -16668 789 -16510 869
rect -16476 789 -16318 869
rect -16284 789 -16272 869
rect -16907 783 -16272 789
rect -16025 869 -15390 875
rect -16025 789 -16012 869
rect -15978 789 -15820 869
rect -15786 789 -15628 869
rect -15594 789 -15436 869
rect -15402 789 -15390 869
rect -16025 783 -15390 789
rect -14725 869 -14090 875
rect -14725 789 -14712 869
rect -14678 789 -14520 869
rect -14486 789 -14328 869
rect -14294 789 -14136 869
rect -14102 789 -14090 869
rect -14725 783 -14090 789
rect -13616 869 -12981 875
rect -13616 789 -13603 869
rect -13569 789 -13411 869
rect -13377 789 -13219 869
rect -13185 789 -13027 869
rect -12993 789 -12981 869
rect -13616 783 -12981 789
rect -12734 869 -12099 875
rect -12734 789 -12721 869
rect -12687 789 -12529 869
rect -12495 789 -12337 869
rect -12303 789 -12145 869
rect -12111 789 -12099 869
rect -12734 783 -12099 789
rect -11434 869 -10799 875
rect -11434 789 -11421 869
rect -11387 789 -11229 869
rect -11195 789 -11037 869
rect -11003 789 -10845 869
rect -10811 789 -10799 869
rect -11434 783 -10799 789
rect -10325 869 -9690 875
rect -10325 789 -10312 869
rect -10278 789 -10120 869
rect -10086 789 -9928 869
rect -9894 789 -9736 869
rect -9702 789 -9690 869
rect -10325 783 -9690 789
rect -9443 869 -8808 875
rect -9443 789 -9430 869
rect -9396 789 -9238 869
rect -9204 789 -9046 869
rect -9012 789 -8854 869
rect -8820 789 -8808 869
rect -9443 783 -8808 789
rect -8144 869 -7509 875
rect -8144 789 -8131 869
rect -8097 789 -7939 869
rect -7905 789 -7747 869
rect -7713 789 -7555 869
rect -7521 789 -7509 869
rect -8144 783 -7509 789
rect -7035 869 -6400 875
rect -7035 789 -7022 869
rect -6988 789 -6830 869
rect -6796 789 -6638 869
rect -6604 789 -6446 869
rect -6412 789 -6400 869
rect -7035 783 -6400 789
rect -6153 869 -5518 875
rect -6153 789 -6140 869
rect -6106 789 -5948 869
rect -5914 789 -5756 869
rect -5722 789 -5564 869
rect -5530 789 -5518 869
rect -6153 783 -5518 789
rect -4853 869 -4218 875
rect -4853 789 -4840 869
rect -4806 789 -4648 869
rect -4614 789 -4456 869
rect -4422 789 -4264 869
rect -4230 789 -4218 869
rect -4853 783 -4218 789
rect -3744 869 -3109 875
rect -3744 789 -3731 869
rect -3697 789 -3539 869
rect -3505 789 -3347 869
rect -3313 789 -3155 869
rect -3121 789 -3109 869
rect -3744 783 -3109 789
rect -2862 869 -2227 875
rect -2862 789 -2849 869
rect -2815 789 -2657 869
rect -2623 789 -2465 869
rect -2431 789 -2273 869
rect -2239 789 -2227 869
rect -2862 783 -2227 789
rect -1562 869 -927 875
rect -1562 789 -1549 869
rect -1515 789 -1357 869
rect -1323 789 -1165 869
rect -1131 789 -973 869
rect -939 789 -927 869
rect -1562 783 -927 789
rect -453 869 182 875
rect -453 789 -440 869
rect -406 789 -248 869
rect -214 789 -56 869
rect -22 789 136 869
rect 170 789 182 869
rect -453 783 182 789
rect 429 869 1064 875
rect 429 789 442 869
rect 476 789 634 869
rect 668 789 826 869
rect 860 789 1018 869
rect 1052 789 1064 869
rect 429 783 1064 789
rect -24598 782 -23964 783
rect -23489 782 -22855 783
rect -22607 782 -21973 783
rect -21307 782 -20673 783
rect -20198 782 -19564 783
rect -19316 782 -18682 783
rect -18016 782 -17382 783
rect -16907 782 -16273 783
rect -16025 782 -15391 783
rect -14725 782 -14091 783
rect -13616 782 -12982 783
rect -12734 782 -12100 783
rect -11434 782 -10800 783
rect -10325 782 -9691 783
rect -9443 782 -8809 783
rect -8144 782 -7510 783
rect -7035 782 -6401 783
rect -6153 782 -5519 783
rect -4853 782 -4219 783
rect -3744 782 -3110 783
rect -2862 782 -2228 783
rect -1562 782 -928 783
rect -453 782 181 783
rect 429 782 1063 783
rect -24505 747 -23927 753
rect -24505 667 -24489 747
rect -24455 667 -24297 747
rect -24263 667 -24105 747
rect -24071 667 -23927 747
rect -24505 666 -23927 667
rect -24505 661 -24046 666
rect -24633 614 -24469 632
rect -24633 605 -24519 614
rect -24633 525 -24601 605
rect -24485 579 -24469 614
rect -24503 525 -24469 579
rect -24633 497 -24469 525
rect -24441 614 -24181 633
rect -24441 579 -24230 614
rect -24196 579 -24181 614
rect -24441 559 -24181 579
rect -24441 490 -24391 559
rect -24105 531 -24046 661
rect -24441 469 -24435 490
rect -24829 455 -24435 469
rect -24401 455 -24391 490
rect -24363 519 -24046 531
rect -24363 485 -24351 519
rect -23963 518 -23927 666
rect -23396 747 -22818 753
rect -23396 667 -23380 747
rect -23346 667 -23188 747
rect -23154 667 -22996 747
rect -22962 667 -22818 747
rect -23396 661 -22818 667
rect -22514 747 -21936 753
rect -22514 667 -22498 747
rect -22464 667 -22306 747
rect -22272 667 -22114 747
rect -22080 667 -21936 747
rect -22514 661 -21936 667
rect -21214 747 -20636 753
rect -21214 667 -21198 747
rect -21164 667 -21006 747
rect -20972 667 -20814 747
rect -20780 667 -20636 747
rect -21214 666 -20636 667
rect -21214 661 -20755 666
rect -23975 485 -23927 518
rect -23524 614 -23360 632
rect -23524 604 -23410 614
rect -23524 524 -23490 604
rect -23376 579 -23360 614
rect -23392 524 -23360 579
rect -23524 497 -23360 524
rect -23332 614 -23072 633
rect -23332 579 -23121 614
rect -23087 579 -23072 614
rect -23332 559 -23072 579
rect -22996 609 -22818 661
rect -22642 614 -22478 632
rect -22642 609 -22528 614
rect -22996 579 -22528 609
rect -22494 579 -22478 614
rect -24363 479 -23927 485
rect -23332 490 -23282 559
rect -22996 531 -22478 579
rect -23332 468 -23326 490
rect -24829 412 -24391 455
rect -24829 346 -24810 412
rect -24557 346 -24391 412
rect -24829 332 -24391 346
rect -23524 455 -23326 468
rect -23292 455 -23282 490
rect -23254 519 -22478 531
rect -23254 485 -23242 519
rect -22866 485 -22818 519
rect -22642 497 -22478 519
rect -22450 614 -22190 633
rect -22450 579 -22239 614
rect -22205 579 -22190 614
rect -22450 559 -22190 579
rect -22114 616 -21936 661
rect -23254 479 -22818 485
rect -22450 490 -22400 559
rect -22114 536 -22069 616
rect -21949 536 -21936 616
rect -22114 531 -21936 536
rect -22450 468 -22444 490
rect -23524 401 -23282 455
rect -23524 341 -23500 401
rect -23315 341 -23282 401
rect -24363 327 -23963 333
rect -23524 332 -23282 341
rect -22642 455 -22444 468
rect -22410 455 -22400 490
rect -22372 519 -21936 531
rect -22372 485 -22360 519
rect -21984 485 -21936 519
rect -21342 614 -21178 632
rect -21342 605 -21228 614
rect -21342 525 -21310 605
rect -21194 579 -21178 614
rect -21212 525 -21178 579
rect -21342 497 -21178 525
rect -21150 614 -20890 633
rect -21150 579 -20939 614
rect -20905 579 -20890 614
rect -21150 559 -20890 579
rect -22372 479 -21936 485
rect -21150 490 -21100 559
rect -20814 531 -20755 661
rect -21150 469 -21144 490
rect -22642 450 -22400 455
rect -22642 375 -22628 450
rect -22483 375 -22400 450
rect -24363 293 -24351 327
rect -23975 293 -23963 327
rect -24363 255 -23963 293
rect -24363 210 -24336 255
rect -24345 203 -24336 210
rect -24001 210 -23963 255
rect -23254 327 -22854 333
rect -22642 332 -22400 375
rect -21538 455 -21144 469
rect -21110 455 -21100 490
rect -21072 519 -20755 531
rect -21072 485 -21060 519
rect -20672 518 -20636 666
rect -20105 747 -19527 753
rect -20105 667 -20089 747
rect -20055 667 -19897 747
rect -19863 667 -19705 747
rect -19671 667 -19527 747
rect -20105 661 -19527 667
rect -19223 747 -18645 753
rect -19223 667 -19207 747
rect -19173 667 -19015 747
rect -18981 667 -18823 747
rect -18789 667 -18645 747
rect -19223 661 -18645 667
rect -17923 747 -17345 753
rect -17923 667 -17907 747
rect -17873 667 -17715 747
rect -17681 667 -17523 747
rect -17489 667 -17345 747
rect -17923 666 -17345 667
rect -17923 661 -17464 666
rect -20684 485 -20636 518
rect -20233 614 -20069 632
rect -20233 604 -20119 614
rect -20233 524 -20199 604
rect -20085 579 -20069 614
rect -20101 524 -20069 579
rect -20233 497 -20069 524
rect -20041 614 -19781 633
rect -20041 579 -19830 614
rect -19796 579 -19781 614
rect -20041 559 -19781 579
rect -19705 609 -19527 661
rect -19351 614 -19187 632
rect -19351 609 -19237 614
rect -19705 579 -19237 609
rect -19203 579 -19187 614
rect -21072 479 -20636 485
rect -20041 490 -19991 559
rect -19705 531 -19187 579
rect -20041 468 -20035 490
rect -21538 412 -21100 455
rect -21538 346 -21519 412
rect -21266 346 -21100 412
rect -23254 293 -23242 327
rect -22866 293 -22854 327
rect -23254 255 -22854 293
rect -23254 221 -23227 255
rect -22892 221 -22854 255
rect -23254 210 -23100 221
rect -24001 203 -23992 210
rect -24345 194 -23992 203
rect -23111 188 -23100 210
rect -23038 210 -22854 221
rect -22372 327 -21972 333
rect -21538 332 -21100 346
rect -20233 455 -20035 468
rect -20001 455 -19991 490
rect -19963 519 -19187 531
rect -19963 485 -19951 519
rect -19575 485 -19527 519
rect -19351 497 -19187 519
rect -19159 614 -18899 633
rect -19159 579 -18948 614
rect -18914 579 -18899 614
rect -19159 559 -18899 579
rect -18823 616 -18645 661
rect -19963 479 -19527 485
rect -19159 490 -19109 559
rect -18823 536 -18778 616
rect -18658 536 -18645 616
rect -18823 531 -18645 536
rect -19159 468 -19153 490
rect -20233 401 -19991 455
rect -20233 341 -20209 401
rect -20024 341 -19991 401
rect -22372 293 -22360 327
rect -21984 293 -21972 327
rect -22372 255 -21972 293
rect -21072 327 -20672 333
rect -20233 332 -19991 341
rect -19351 455 -19153 468
rect -19119 455 -19109 490
rect -19081 519 -18645 531
rect -19081 485 -19069 519
rect -18693 485 -18645 519
rect -18051 614 -17887 632
rect -18051 605 -17937 614
rect -18051 525 -18019 605
rect -17903 579 -17887 614
rect -17921 525 -17887 579
rect -18051 497 -17887 525
rect -17859 614 -17599 633
rect -17859 579 -17648 614
rect -17614 579 -17599 614
rect -17859 559 -17599 579
rect -19081 479 -18645 485
rect -17859 490 -17809 559
rect -17523 531 -17464 661
rect -17859 469 -17853 490
rect -19351 450 -19109 455
rect -19351 375 -19337 450
rect -19192 375 -19109 450
rect -21072 293 -21060 327
rect -20684 293 -20672 327
rect -22372 221 -22345 255
rect -22010 221 -21972 255
rect -22372 210 -22233 221
rect -23038 188 -23027 210
rect -23111 177 -23027 188
rect -22246 171 -22233 210
rect -22181 210 -21972 221
rect -21801 284 -21735 290
rect -22181 171 -22168 210
rect -22246 158 -22168 171
rect -25066 -214 -25060 -123
rect -24969 -214 -24963 -123
rect -21801 -492 -21735 218
rect -21072 255 -20672 293
rect -21072 210 -21045 255
rect -21054 203 -21045 210
rect -20710 210 -20672 255
rect -19963 327 -19563 333
rect -19351 332 -19109 375
rect -18247 455 -17853 469
rect -17819 455 -17809 490
rect -17781 519 -17464 531
rect -17781 485 -17769 519
rect -17381 518 -17345 666
rect -16814 747 -16236 753
rect -16814 667 -16798 747
rect -16764 667 -16606 747
rect -16572 667 -16414 747
rect -16380 667 -16236 747
rect -16814 661 -16236 667
rect -15932 747 -15354 753
rect -15932 667 -15916 747
rect -15882 667 -15724 747
rect -15690 667 -15532 747
rect -15498 667 -15354 747
rect -15932 661 -15354 667
rect -14632 747 -14054 753
rect -14632 667 -14616 747
rect -14582 667 -14424 747
rect -14390 667 -14232 747
rect -14198 667 -14054 747
rect -14632 666 -14054 667
rect -14632 661 -14173 666
rect -17393 485 -17345 518
rect -16942 614 -16778 632
rect -16942 604 -16828 614
rect -16942 524 -16908 604
rect -16794 579 -16778 614
rect -16810 524 -16778 579
rect -16942 497 -16778 524
rect -16750 614 -16490 633
rect -16750 579 -16539 614
rect -16505 579 -16490 614
rect -16750 559 -16490 579
rect -16414 609 -16236 661
rect -16060 614 -15896 632
rect -16060 609 -15946 614
rect -16414 579 -15946 609
rect -15912 579 -15896 614
rect -17781 479 -17345 485
rect -16750 490 -16700 559
rect -16414 531 -15896 579
rect -16750 468 -16744 490
rect -18247 412 -17809 455
rect -18247 346 -18228 412
rect -17975 346 -17809 412
rect -19963 293 -19951 327
rect -19575 293 -19563 327
rect -19963 255 -19563 293
rect -19963 221 -19936 255
rect -19601 221 -19563 255
rect -19963 210 -19809 221
rect -20710 203 -20701 210
rect -21054 194 -20701 203
rect -19820 188 -19809 210
rect -19747 210 -19563 221
rect -19081 327 -18681 333
rect -18247 332 -17809 346
rect -16942 455 -16744 468
rect -16710 455 -16700 490
rect -16672 519 -15896 531
rect -16672 485 -16660 519
rect -16284 485 -16236 519
rect -16060 497 -15896 519
rect -15868 614 -15608 633
rect -15868 579 -15657 614
rect -15623 579 -15608 614
rect -15868 559 -15608 579
rect -15532 616 -15354 661
rect -16672 479 -16236 485
rect -15868 490 -15818 559
rect -15532 536 -15487 616
rect -15367 536 -15354 616
rect -15532 531 -15354 536
rect -15868 468 -15862 490
rect -16942 401 -16700 455
rect -16942 341 -16918 401
rect -16733 341 -16700 401
rect -19081 293 -19069 327
rect -18693 293 -18681 327
rect -19081 255 -18681 293
rect -17781 327 -17381 333
rect -16942 332 -16700 341
rect -16060 455 -15862 468
rect -15828 455 -15818 490
rect -15790 519 -15354 531
rect -15790 485 -15778 519
rect -15402 485 -15354 519
rect -14760 614 -14596 632
rect -14760 605 -14646 614
rect -14760 525 -14728 605
rect -14612 579 -14596 614
rect -14630 525 -14596 579
rect -14760 497 -14596 525
rect -14568 614 -14308 633
rect -14568 579 -14357 614
rect -14323 579 -14308 614
rect -14568 559 -14308 579
rect -15790 479 -15354 485
rect -14568 490 -14518 559
rect -14232 531 -14173 661
rect -14568 469 -14562 490
rect -16060 450 -15818 455
rect -16060 375 -16046 450
rect -15901 375 -15818 450
rect -17781 293 -17769 327
rect -17393 293 -17381 327
rect -19081 221 -19054 255
rect -18719 221 -18681 255
rect -19081 210 -18942 221
rect -19747 188 -19736 210
rect -19820 177 -19736 188
rect -18955 171 -18942 210
rect -18890 210 -18681 221
rect -18505 283 -18439 289
rect -18890 171 -18877 210
rect -18955 158 -18877 171
rect -18505 -306 -18439 217
rect -17781 255 -17381 293
rect -17781 210 -17754 255
rect -17763 203 -17754 210
rect -17419 210 -17381 255
rect -16672 327 -16272 333
rect -16060 332 -15818 375
rect -14956 455 -14562 469
rect -14528 455 -14518 490
rect -14490 519 -14173 531
rect -14490 485 -14478 519
rect -14090 518 -14054 666
rect -13523 747 -12945 753
rect -13523 667 -13507 747
rect -13473 667 -13315 747
rect -13281 667 -13123 747
rect -13089 667 -12945 747
rect -13523 661 -12945 667
rect -12641 747 -12063 753
rect -12641 667 -12625 747
rect -12591 667 -12433 747
rect -12399 667 -12241 747
rect -12207 667 -12063 747
rect -12641 661 -12063 667
rect -11341 747 -10763 753
rect -11341 667 -11325 747
rect -11291 667 -11133 747
rect -11099 667 -10941 747
rect -10907 667 -10763 747
rect -11341 666 -10763 667
rect -11341 661 -10882 666
rect -14102 485 -14054 518
rect -13651 614 -13487 632
rect -13651 604 -13537 614
rect -13651 524 -13617 604
rect -13503 579 -13487 614
rect -13519 524 -13487 579
rect -13651 497 -13487 524
rect -13459 614 -13199 633
rect -13459 579 -13248 614
rect -13214 579 -13199 614
rect -13459 559 -13199 579
rect -13123 609 -12945 661
rect -12769 614 -12605 632
rect -12769 609 -12655 614
rect -13123 579 -12655 609
rect -12621 579 -12605 614
rect -14490 479 -14054 485
rect -13459 490 -13409 559
rect -13123 531 -12605 579
rect -13459 468 -13453 490
rect -14956 412 -14518 455
rect -14956 346 -14937 412
rect -14684 346 -14518 412
rect -16672 293 -16660 327
rect -16284 293 -16272 327
rect -16672 255 -16272 293
rect -16672 221 -16645 255
rect -16310 221 -16272 255
rect -16672 210 -16518 221
rect -17419 203 -17410 210
rect -17763 194 -17410 203
rect -16529 188 -16518 210
rect -16456 210 -16272 221
rect -15790 327 -15390 333
rect -14956 332 -14518 346
rect -13651 455 -13453 468
rect -13419 455 -13409 490
rect -13381 519 -12605 531
rect -13381 485 -13369 519
rect -12993 485 -12945 519
rect -12769 497 -12605 519
rect -12577 614 -12317 633
rect -12577 579 -12366 614
rect -12332 579 -12317 614
rect -12577 559 -12317 579
rect -12241 616 -12063 661
rect -13381 479 -12945 485
rect -12577 490 -12527 559
rect -12241 536 -12196 616
rect -12076 536 -12063 616
rect -12241 531 -12063 536
rect -12577 468 -12571 490
rect -13651 401 -13409 455
rect -13651 341 -13627 401
rect -13442 341 -13409 401
rect -15790 293 -15778 327
rect -15402 293 -15390 327
rect -14490 327 -14090 333
rect -13651 332 -13409 341
rect -12769 455 -12571 468
rect -12537 455 -12527 490
rect -12499 519 -12063 531
rect -12499 485 -12487 519
rect -12111 485 -12063 519
rect -11469 614 -11305 632
rect -11469 605 -11355 614
rect -11469 525 -11437 605
rect -11321 579 -11305 614
rect -11339 525 -11305 579
rect -11469 497 -11305 525
rect -11277 614 -11017 633
rect -11277 579 -11066 614
rect -11032 579 -11017 614
rect -11277 559 -11017 579
rect -12499 479 -12063 485
rect -11277 490 -11227 559
rect -10941 531 -10882 661
rect -11277 469 -11271 490
rect -12769 450 -12527 455
rect -12769 375 -12755 450
rect -12610 375 -12527 450
rect -15790 255 -15390 293
rect -15790 221 -15763 255
rect -15428 221 -15390 255
rect -15790 210 -15651 221
rect -16456 188 -16445 210
rect -16529 177 -16445 188
rect -15664 171 -15651 210
rect -15599 210 -15390 221
rect -15223 296 -15157 302
rect -15599 171 -15586 210
rect -15664 158 -15586 171
rect -18505 -372 -15446 -306
rect -21801 -558 -15583 -492
rect -15649 -1309 -15583 -558
rect -15512 -1138 -15446 -372
rect -15223 -948 -15157 230
rect -14490 293 -14478 327
rect -14102 293 -14090 327
rect -14490 255 -14090 293
rect -14490 210 -14463 255
rect -14472 203 -14463 210
rect -14128 210 -14090 255
rect -13381 327 -12981 333
rect -12769 332 -12527 375
rect -11665 455 -11271 469
rect -11237 455 -11227 490
rect -11199 519 -10882 531
rect -11199 485 -11187 519
rect -10799 518 -10763 666
rect -10232 747 -9654 753
rect -10232 667 -10216 747
rect -10182 667 -10024 747
rect -9990 667 -9832 747
rect -9798 667 -9654 747
rect -10232 661 -9654 667
rect -9350 747 -8772 753
rect -9350 667 -9334 747
rect -9300 667 -9142 747
rect -9108 667 -8950 747
rect -8916 667 -8772 747
rect -9350 661 -8772 667
rect -8051 747 -7473 753
rect -8051 667 -8035 747
rect -8001 667 -7843 747
rect -7809 667 -7651 747
rect -7617 667 -7473 747
rect -8051 666 -7473 667
rect -8051 661 -7592 666
rect -10811 485 -10763 518
rect -10360 614 -10196 632
rect -10360 604 -10246 614
rect -10360 524 -10326 604
rect -10212 579 -10196 614
rect -10228 524 -10196 579
rect -10360 497 -10196 524
rect -10168 614 -9908 633
rect -10168 579 -9957 614
rect -9923 579 -9908 614
rect -10168 559 -9908 579
rect -9832 609 -9654 661
rect -9478 614 -9314 632
rect -9478 609 -9364 614
rect -9832 579 -9364 609
rect -9330 579 -9314 614
rect -11199 479 -10763 485
rect -10168 490 -10118 559
rect -9832 531 -9314 579
rect -10168 468 -10162 490
rect -11665 412 -11227 455
rect -11665 346 -11646 412
rect -11393 346 -11227 412
rect -13381 293 -13369 327
rect -12993 293 -12981 327
rect -13381 255 -12981 293
rect -13381 221 -13354 255
rect -13019 221 -12981 255
rect -13381 210 -13227 221
rect -14128 203 -14119 210
rect -14472 194 -14119 203
rect -13238 188 -13227 210
rect -13165 210 -12981 221
rect -12499 327 -12099 333
rect -11665 332 -11227 346
rect -10360 455 -10162 468
rect -10128 455 -10118 490
rect -10090 519 -9314 531
rect -10090 485 -10078 519
rect -9702 485 -9654 519
rect -9478 497 -9314 519
rect -9286 614 -9026 633
rect -9286 579 -9075 614
rect -9041 579 -9026 614
rect -9286 559 -9026 579
rect -8950 616 -8772 661
rect -10090 479 -9654 485
rect -9286 490 -9236 559
rect -8950 536 -8905 616
rect -8785 536 -8772 616
rect -8950 531 -8772 536
rect -9286 468 -9280 490
rect -10360 401 -10118 455
rect -10360 341 -10336 401
rect -10151 341 -10118 401
rect -12499 293 -12487 327
rect -12111 293 -12099 327
rect -12499 255 -12099 293
rect -11199 327 -10799 333
rect -10360 332 -10118 341
rect -9478 455 -9280 468
rect -9246 455 -9236 490
rect -9208 519 -8772 531
rect -9208 485 -9196 519
rect -8820 485 -8772 519
rect -8179 614 -8015 632
rect -8179 605 -8065 614
rect -8179 525 -8147 605
rect -8031 579 -8015 614
rect -8049 525 -8015 579
rect -8179 497 -8015 525
rect -7987 614 -7727 633
rect -7987 579 -7776 614
rect -7742 579 -7727 614
rect -7987 559 -7727 579
rect -9208 479 -8772 485
rect -7987 490 -7937 559
rect -7651 531 -7592 661
rect -7987 469 -7981 490
rect -9478 450 -9236 455
rect -9478 375 -9464 450
rect -9319 375 -9236 450
rect -11199 293 -11187 327
rect -10811 293 -10799 327
rect -12499 221 -12472 255
rect -12137 221 -12099 255
rect -11969 223 -11963 289
rect -11897 223 -11891 289
rect -11199 255 -10799 293
rect -12499 210 -12360 221
rect -13165 188 -13154 210
rect -13238 177 -13154 188
rect -12373 171 -12360 210
rect -12308 210 -12099 221
rect -12308 171 -12295 210
rect -12373 158 -12295 171
rect -11963 -785 -11897 223
rect -11199 210 -11172 255
rect -11181 203 -11172 210
rect -10837 210 -10799 255
rect -10090 327 -9690 333
rect -9478 332 -9236 375
rect -8375 455 -7981 469
rect -7947 455 -7937 490
rect -7909 519 -7592 531
rect -7909 485 -7897 519
rect -7509 518 -7473 666
rect -6942 747 -6364 753
rect -6942 667 -6926 747
rect -6892 667 -6734 747
rect -6700 667 -6542 747
rect -6508 667 -6364 747
rect -6942 661 -6364 667
rect -6060 747 -5482 753
rect -6060 667 -6044 747
rect -6010 667 -5852 747
rect -5818 667 -5660 747
rect -5626 667 -5482 747
rect -6060 661 -5482 667
rect -4760 747 -4182 753
rect -4760 667 -4744 747
rect -4710 667 -4552 747
rect -4518 667 -4360 747
rect -4326 667 -4182 747
rect -4760 666 -4182 667
rect -4760 661 -4301 666
rect -7521 485 -7473 518
rect -7070 614 -6906 632
rect -7070 604 -6956 614
rect -7070 524 -7036 604
rect -6922 579 -6906 614
rect -6938 524 -6906 579
rect -7070 497 -6906 524
rect -6878 614 -6618 633
rect -6878 579 -6667 614
rect -6633 579 -6618 614
rect -6878 559 -6618 579
rect -6542 609 -6364 661
rect -6188 614 -6024 632
rect -6188 609 -6074 614
rect -6542 579 -6074 609
rect -6040 579 -6024 614
rect -7909 479 -7473 485
rect -6878 490 -6828 559
rect -6542 531 -6024 579
rect -6878 468 -6872 490
rect -8375 412 -7937 455
rect -8375 346 -8356 412
rect -8103 346 -7937 412
rect -10090 293 -10078 327
rect -9702 293 -9690 327
rect -10090 255 -9690 293
rect -10090 221 -10063 255
rect -9728 221 -9690 255
rect -10090 210 -9936 221
rect -10837 203 -10828 210
rect -11181 194 -10828 203
rect -9947 188 -9936 210
rect -9874 210 -9690 221
rect -9208 327 -8808 333
rect -8375 332 -7937 346
rect -7070 455 -6872 468
rect -6838 455 -6828 490
rect -6800 519 -6024 531
rect -6800 485 -6788 519
rect -6412 485 -6364 519
rect -6188 497 -6024 519
rect -5996 614 -5736 633
rect -5996 579 -5785 614
rect -5751 579 -5736 614
rect -5996 559 -5736 579
rect -5660 616 -5482 661
rect -6800 479 -6364 485
rect -5996 490 -5946 559
rect -5660 536 -5615 616
rect -5495 536 -5482 616
rect -5660 531 -5482 536
rect -5996 468 -5990 490
rect -7070 401 -6828 455
rect -7070 341 -7046 401
rect -6861 341 -6828 401
rect -9208 293 -9196 327
rect -8820 293 -8808 327
rect -7909 327 -7509 333
rect -7070 332 -6828 341
rect -6188 455 -5990 468
rect -5956 455 -5946 490
rect -5918 519 -5482 531
rect -5918 485 -5906 519
rect -5530 485 -5482 519
rect -4888 614 -4724 632
rect -4888 605 -4774 614
rect -4888 525 -4856 605
rect -4740 579 -4724 614
rect -4758 525 -4724 579
rect -4888 497 -4724 525
rect -4696 614 -4436 633
rect -4696 579 -4485 614
rect -4451 579 -4436 614
rect -4696 559 -4436 579
rect -5918 479 -5482 485
rect -4696 490 -4646 559
rect -4360 531 -4301 661
rect -4696 469 -4690 490
rect -6188 450 -5946 455
rect -6188 375 -6174 450
rect -6029 375 -5946 450
rect -9208 255 -8808 293
rect -9208 221 -9181 255
rect -8846 221 -8808 255
rect -9208 210 -9069 221
rect -9874 188 -9863 210
rect -9947 177 -9863 188
rect -9082 171 -9069 210
rect -9017 210 -8808 221
rect -8633 309 -8567 315
rect -9017 171 -9004 210
rect -9082 158 -9004 171
rect -8633 -618 -8567 243
rect -7909 293 -7897 327
rect -7521 293 -7509 327
rect -7909 255 -7509 293
rect -7909 210 -7882 255
rect -7891 203 -7882 210
rect -7547 210 -7509 255
rect -6800 327 -6400 333
rect -6188 332 -5946 375
rect -5084 455 -4690 469
rect -4656 455 -4646 490
rect -4618 519 -4301 531
rect -4618 485 -4606 519
rect -4218 518 -4182 666
rect -3651 747 -3073 753
rect -3651 667 -3635 747
rect -3601 667 -3443 747
rect -3409 667 -3251 747
rect -3217 667 -3073 747
rect -3651 661 -3073 667
rect -2769 747 -2191 753
rect -2769 667 -2753 747
rect -2719 667 -2561 747
rect -2527 667 -2369 747
rect -2335 667 -2191 747
rect -2769 661 -2191 667
rect -1469 747 -891 753
rect -1469 667 -1453 747
rect -1419 667 -1261 747
rect -1227 667 -1069 747
rect -1035 667 -891 747
rect -1469 666 -891 667
rect -1469 661 -1010 666
rect -4230 485 -4182 518
rect -3779 614 -3615 632
rect -3779 604 -3665 614
rect -3779 524 -3745 604
rect -3631 579 -3615 614
rect -3647 524 -3615 579
rect -3779 497 -3615 524
rect -3587 614 -3327 633
rect -3587 579 -3376 614
rect -3342 579 -3327 614
rect -3587 559 -3327 579
rect -3251 609 -3073 661
rect -2897 614 -2733 632
rect -2897 609 -2783 614
rect -3251 579 -2783 609
rect -2749 579 -2733 614
rect -4618 479 -4182 485
rect -3587 490 -3537 559
rect -3251 531 -2733 579
rect -3587 468 -3581 490
rect -5084 412 -4646 455
rect -5084 346 -5065 412
rect -4812 346 -4646 412
rect -6800 293 -6788 327
rect -6412 293 -6400 327
rect -6800 255 -6400 293
rect -6800 221 -6773 255
rect -6438 221 -6400 255
rect -6800 210 -6646 221
rect -7547 203 -7538 210
rect -7891 194 -7538 203
rect -6657 188 -6646 210
rect -6584 210 -6400 221
rect -5918 327 -5518 333
rect -5084 332 -4646 346
rect -3779 455 -3581 468
rect -3547 455 -3537 490
rect -3509 519 -2733 531
rect -3509 485 -3497 519
rect -3121 485 -3073 519
rect -2897 497 -2733 519
rect -2705 614 -2445 633
rect -2705 579 -2494 614
rect -2460 579 -2445 614
rect -2705 559 -2445 579
rect -2369 616 -2191 661
rect -3509 479 -3073 485
rect -2705 490 -2655 559
rect -2369 536 -2324 616
rect -2204 536 -2191 616
rect -2369 531 -2191 536
rect -2705 468 -2699 490
rect -3779 401 -3537 455
rect -3779 341 -3755 401
rect -3570 341 -3537 401
rect -5918 293 -5906 327
rect -5530 293 -5518 327
rect -4618 327 -4218 333
rect -3779 332 -3537 341
rect -2897 455 -2699 468
rect -2665 455 -2655 490
rect -2627 519 -2191 531
rect -2627 485 -2615 519
rect -2239 485 -2191 519
rect -1597 614 -1433 632
rect -1597 605 -1483 614
rect -1597 525 -1565 605
rect -1449 579 -1433 614
rect -1467 525 -1433 579
rect -1597 497 -1433 525
rect -1405 614 -1145 633
rect -1405 579 -1194 614
rect -1160 579 -1145 614
rect -1405 559 -1145 579
rect -2627 479 -2191 485
rect -1405 490 -1355 559
rect -1069 531 -1010 661
rect -1405 469 -1399 490
rect -2897 450 -2655 455
rect -2897 375 -2883 450
rect -2738 375 -2655 450
rect -5918 255 -5518 293
rect -5918 221 -5891 255
rect -5556 221 -5518 255
rect -5918 210 -5779 221
rect -6584 188 -6573 210
rect -6657 177 -6573 188
rect -5792 171 -5779 210
rect -5727 210 -5518 221
rect -5349 292 -5283 298
rect -5727 171 -5714 210
rect -5792 158 -5714 171
rect -5349 -421 -5283 226
rect -4618 293 -4606 327
rect -4230 293 -4218 327
rect -4618 255 -4218 293
rect -4618 210 -4591 255
rect -4600 203 -4591 210
rect -4256 210 -4218 255
rect -3509 327 -3109 333
rect -2897 332 -2655 375
rect -1793 455 -1399 469
rect -1365 455 -1355 490
rect -1327 519 -1010 531
rect -1327 485 -1315 519
rect -927 518 -891 666
rect -360 747 218 753
rect -360 667 -344 747
rect -310 667 -152 747
rect -118 667 40 747
rect 74 667 218 747
rect -360 661 218 667
rect 522 747 1100 753
rect 522 667 538 747
rect 572 667 730 747
rect 764 667 922 747
rect 956 667 1100 747
rect 522 661 1100 667
rect -939 485 -891 518
rect -488 614 -324 632
rect -488 604 -374 614
rect -488 524 -454 604
rect -340 579 -324 614
rect -356 524 -324 579
rect -488 497 -324 524
rect -296 614 -36 633
rect -296 579 -85 614
rect -51 579 -36 614
rect -296 559 -36 579
rect 40 609 218 661
rect 394 614 558 632
rect 394 609 508 614
rect 40 579 508 609
rect 542 579 558 614
rect -1327 479 -891 485
rect -296 490 -246 559
rect 40 531 558 579
rect -296 468 -290 490
rect -1793 412 -1355 455
rect -1793 346 -1774 412
rect -1521 346 -1355 412
rect -3509 293 -3497 327
rect -3121 293 -3109 327
rect -3509 255 -3109 293
rect -3509 221 -3482 255
rect -3147 221 -3109 255
rect -3509 210 -3355 221
rect -4256 203 -4247 210
rect -4600 194 -4247 203
rect -3366 188 -3355 210
rect -3293 210 -3109 221
rect -2627 327 -2227 333
rect -1793 332 -1355 346
rect -488 455 -290 468
rect -256 455 -246 490
rect -218 519 558 531
rect -218 485 -206 519
rect 170 485 218 519
rect 394 497 558 519
rect 586 614 846 633
rect 586 579 797 614
rect 831 579 846 614
rect 586 559 846 579
rect 922 616 1100 661
rect -218 479 218 485
rect 586 490 636 559
rect 922 536 967 616
rect 1087 536 1100 616
rect 922 531 1100 536
rect 586 468 592 490
rect -488 401 -246 455
rect -488 341 -464 401
rect -279 341 -246 401
rect -2627 293 -2615 327
rect -2239 293 -2227 327
rect -2627 255 -2227 293
rect -1327 327 -927 333
rect -488 332 -246 341
rect 394 455 592 468
rect 626 455 636 490
rect 664 519 1100 531
rect 664 485 676 519
rect 1052 485 1100 519
rect 664 479 1100 485
rect 394 450 636 455
rect 394 375 408 450
rect 553 375 636 450
rect -1327 293 -1315 327
rect -939 293 -927 327
rect -2627 221 -2600 255
rect -2265 221 -2227 255
rect -2627 210 -2488 221
rect -3293 188 -3282 210
rect -3366 177 -3282 188
rect -2501 171 -2488 210
rect -2436 210 -2227 221
rect -2061 261 -1995 267
rect -2436 171 -2423 210
rect -2501 158 -2423 171
rect -1327 255 -927 293
rect -1327 210 -1300 255
rect -2061 -232 -1995 195
rect -1309 203 -1300 210
rect -965 210 -927 255
rect -218 327 182 333
rect 394 332 636 375
rect -218 293 -206 327
rect 170 293 182 327
rect -218 255 182 293
rect -218 221 -191 255
rect 144 221 182 255
rect -218 210 -64 221
rect -965 203 -956 210
rect -1309 194 -956 203
rect -75 188 -64 210
rect -2 210 182 221
rect 664 327 1064 333
rect 664 293 676 327
rect 1052 293 1064 327
rect 664 255 1064 293
rect 664 221 691 255
rect 1026 221 1064 255
rect 664 210 803 221
rect -2 188 9 210
rect -75 177 9 188
rect 790 171 803 210
rect 855 210 1064 221
rect 855 171 868 210
rect 790 158 868 171
rect 248 -40 339 -34
rect 1922 -40 2013 2453
rect 5832 452 5901 3045
rect 5998 2781 6067 3383
rect 6098 3373 6298 3380
rect 6098 3339 6110 3373
rect 6286 3339 6298 3373
rect 6326 3366 6410 3427
rect 6098 3271 6298 3339
rect 6098 3237 6129 3271
rect 6261 3237 6298 3271
rect 6098 3230 6172 3237
rect 6143 3195 6172 3230
rect 6224 3230 6298 3237
rect 6341 3312 6410 3366
rect 6341 3230 6410 3243
rect 6438 3637 6457 3810
rect 6491 3637 6507 3810
rect 6538 3877 6544 3911
rect 6623 3907 6752 3911
rect 6623 3877 6629 3907
rect 6538 3719 6629 3877
rect 6538 3685 6544 3719
rect 6623 3685 6629 3719
rect 6538 3669 6629 3685
rect 6661 3815 6850 3879
rect 6661 3781 6667 3815
rect 6744 3781 6850 3815
rect 6438 3417 6507 3637
rect 6661 3623 6850 3781
rect 6538 3589 6667 3623
rect 6744 3589 6850 3623
rect 6538 3461 6850 3589
rect 6538 3427 6550 3461
rect 6726 3427 6850 3461
rect 6538 3421 6738 3427
rect 6438 3383 6457 3417
rect 6491 3383 6507 3417
rect 6224 3195 6263 3230
rect 6143 3170 6263 3195
rect 5992 2775 6073 2781
rect 5992 2706 5998 2775
rect 6067 2772 6073 2775
rect 6067 2706 6085 2772
rect 5992 2700 6073 2706
rect 5998 546 6067 2700
rect 6438 2640 6507 3383
rect 6538 3373 6738 3380
rect 6538 3339 6550 3373
rect 6726 3339 6738 3373
rect 6766 3366 6850 3427
rect 6538 3271 6738 3339
rect 6781 3321 6850 3366
rect 7254 3327 7357 3924
rect 11860 3327 12409 3328
rect 12750 3327 13092 3328
rect 6538 3237 6569 3271
rect 6701 3237 6738 3271
rect 6538 3230 6612 3237
rect 6580 3204 6612 3230
rect 6664 3230 6738 3237
rect 6780 3290 6850 3321
rect 7137 3326 7964 3327
rect 8085 3326 8912 3327
rect 9021 3326 9848 3327
rect 9952 3326 10779 3327
rect 7137 3311 10780 3326
rect 6664 3204 6700 3230
rect 6580 3161 6700 3204
rect 6438 2565 6507 2571
rect 6780 2678 6849 3290
rect 7137 3276 7389 3311
rect 7677 3276 8337 3311
rect 8625 3276 9273 3311
rect 9561 3276 10204 3311
rect 10492 3276 10780 3311
rect 7137 3215 10780 3276
rect 10879 3311 13092 3327
rect 10879 3276 11131 3311
rect 11419 3276 13092 3311
rect 10879 3215 13092 3276
rect 7138 3204 10780 3215
rect 7138 3094 7150 3204
rect 7184 3094 7342 3204
rect 7376 3094 7534 3204
rect 7568 3094 7726 3204
rect 7760 3094 7918 3204
rect 7952 3094 8098 3204
rect 8132 3094 8290 3204
rect 8324 3094 8482 3204
rect 8516 3094 8674 3204
rect 8708 3094 8866 3204
rect 8900 3094 9034 3204
rect 9068 3094 9226 3204
rect 9260 3094 9418 3204
rect 9452 3094 9610 3204
rect 9644 3094 9802 3204
rect 9836 3094 9965 3204
rect 9999 3094 10157 3204
rect 10191 3094 10349 3204
rect 10383 3094 10541 3204
rect 10575 3094 10733 3204
rect 10767 3094 10780 3204
rect 7138 3085 10780 3094
rect 10880 3204 13092 3215
rect 10880 3094 10892 3204
rect 10926 3094 11084 3204
rect 11118 3094 11276 3204
rect 11310 3094 11468 3204
rect 11502 3094 11660 3204
rect 11694 3094 13092 3204
rect 10880 3085 13092 3094
rect 7138 3016 8001 3031
rect 7138 2904 7245 3016
rect 7280 2904 7438 3016
rect 7473 2904 7630 3016
rect 7665 2904 7822 3016
rect 7857 2904 8001 3016
rect 7138 2897 8001 2904
rect 8086 3016 8949 3031
rect 8086 2904 8193 3016
rect 8228 2904 8386 3016
rect 8421 2904 8578 3016
rect 8613 2904 8770 3016
rect 8805 2904 8949 3016
rect 8086 2897 8949 2904
rect 9022 3016 9885 3031
rect 9022 2904 9129 3016
rect 9164 2904 9322 3016
rect 9357 2904 9514 3016
rect 9549 2904 9706 3016
rect 9741 2904 9885 3016
rect 9022 2897 9885 2904
rect 9953 3016 10816 3031
rect 9953 2904 10060 3016
rect 10095 2904 10253 3016
rect 10288 2904 10445 3016
rect 10480 2904 10637 3016
rect 10672 2904 10816 3016
rect 9953 2897 10816 2904
rect 10880 3016 11743 3031
rect 10880 2904 10987 3016
rect 11022 2904 11180 3016
rect 11215 2904 11372 3016
rect 11407 2904 11564 3016
rect 11599 2904 11743 3016
rect 10880 2897 11743 2904
rect 7106 2866 7158 2867
rect 7102 2861 7248 2866
rect 7102 2809 7106 2861
rect 7158 2850 7248 2861
rect 7158 2816 7198 2850
rect 7232 2816 7248 2850
rect 7158 2809 7248 2816
rect 7102 2800 7248 2809
rect 7304 2850 7441 2866
rect 7304 2816 7390 2850
rect 7424 2816 7441 2850
rect 7304 2800 7441 2816
rect 7491 2850 7632 2865
rect 7491 2816 7582 2850
rect 7616 2816 7632 2850
rect 7304 2772 7370 2800
rect 7097 2767 7370 2772
rect 7097 2715 7113 2767
rect 7165 2715 7370 2767
rect 7491 2799 7632 2816
rect 7661 2850 7825 2866
rect 7661 2816 7774 2850
rect 7808 2816 7825 2850
rect 7661 2800 7825 2816
rect 7491 2763 7557 2799
rect 7594 2798 7628 2799
rect 7097 2706 7370 2715
rect 7409 2678 7557 2763
rect 6780 2612 7327 2678
rect 7393 2612 7557 2678
rect 6780 649 6849 2612
rect 7661 2584 7727 2800
rect 7102 2518 7727 2584
rect 7106 2317 7172 2518
rect 7891 2490 8001 2897
rect 8050 2860 8196 2866
rect 8050 2808 8069 2860
rect 8122 2850 8196 2860
rect 8122 2816 8146 2850
rect 8180 2816 8196 2850
rect 8122 2808 8196 2816
rect 8050 2800 8196 2808
rect 8252 2850 8389 2866
rect 8252 2816 8338 2850
rect 8372 2816 8389 2850
rect 8252 2800 8389 2816
rect 8439 2850 8580 2865
rect 8439 2816 8530 2850
rect 8564 2816 8580 2850
rect 8252 2772 8318 2800
rect 8050 2768 8318 2772
rect 8050 2716 8057 2768
rect 8109 2716 8318 2768
rect 8439 2799 8580 2816
rect 8609 2850 8773 2866
rect 8609 2816 8722 2850
rect 8756 2816 8773 2850
rect 8609 2800 8773 2816
rect 8439 2763 8505 2799
rect 8542 2798 8576 2799
rect 8050 2706 8318 2716
rect 8357 2685 8505 2763
rect 8357 2678 8424 2685
rect 8050 2633 8424 2678
rect 8493 2633 8505 2685
rect 8050 2612 8505 2633
rect 8609 2584 8675 2800
rect 7106 2245 7172 2251
rect 7214 2478 7413 2490
rect 7214 2466 7372 2478
rect 7214 2213 7298 2466
rect 6917 2147 6966 2213
rect 7032 2147 7298 2213
rect 7214 1715 7298 2147
rect 7333 1715 7372 2466
rect 7214 1537 7227 1715
rect 7406 1702 7413 2478
rect 7405 1550 7413 1702
rect 7750 2478 8001 2490
rect 7750 1702 7756 2478
rect 7790 2475 8001 2478
rect 8050 2518 8675 2584
rect 7790 2060 8000 2475
rect 8050 2213 8116 2518
rect 8839 2490 8949 2897
rect 8986 2861 9132 2866
rect 8986 2809 9002 2861
rect 9055 2850 9132 2861
rect 9055 2816 9082 2850
rect 9116 2816 9132 2850
rect 9055 2809 9132 2816
rect 8986 2800 9132 2809
rect 9188 2850 9325 2866
rect 9188 2816 9274 2850
rect 9308 2816 9325 2850
rect 9188 2800 9325 2816
rect 9375 2850 9516 2865
rect 9375 2816 9466 2850
rect 9500 2816 9516 2850
rect 9188 2772 9254 2800
rect 8986 2763 9254 2772
rect 9375 2799 9516 2816
rect 9545 2850 9709 2866
rect 9545 2816 9658 2850
rect 9692 2816 9709 2850
rect 9545 2800 9709 2816
rect 9375 2763 9441 2799
rect 9478 2798 9512 2799
rect 8986 2711 9000 2763
rect 9052 2711 9254 2763
rect 8986 2706 9254 2711
rect 9293 2678 9441 2763
rect 8986 2672 9441 2678
rect 8986 2619 8989 2672
rect 9042 2619 9441 2672
rect 8986 2612 9441 2619
rect 9545 2584 9611 2800
rect 8050 2141 8116 2147
rect 8162 2478 8361 2490
rect 8162 2466 8320 2478
rect 7790 1994 7872 2060
rect 7938 1994 8000 2060
rect 7790 1702 8000 1994
rect 7750 1690 8000 1702
rect 8162 1715 8246 2466
rect 8281 1715 8320 2466
rect 8354 1702 8361 2478
rect 6953 1111 7019 1117
rect 7214 1111 7298 1537
rect 7019 1045 7298 1111
rect 6953 1039 7019 1045
rect 7102 891 7168 897
rect 7102 734 7168 825
rect 7214 786 7298 1045
rect 7333 786 7372 1537
rect 7214 774 7372 786
rect 7406 774 7413 1550
rect 7214 762 7413 774
rect 7750 1550 8000 1562
rect 7750 774 7756 1550
rect 7790 1267 8000 1550
rect 7790 1201 7853 1267
rect 7919 1201 8000 1267
rect 7790 777 8000 1201
rect 8340 1550 8361 1702
rect 8698 2478 8949 2490
rect 8698 1702 8704 2478
rect 8738 2475 8949 2478
rect 8986 2519 9611 2584
rect 8738 2314 8948 2475
rect 9052 2518 9611 2519
rect 9775 2562 9885 2897
rect 10706 2866 10816 2897
rect 9917 2861 10063 2866
rect 9917 2809 9933 2861
rect 9986 2850 10063 2861
rect 9986 2816 10013 2850
rect 10047 2816 10063 2850
rect 9986 2809 10063 2816
rect 9917 2800 10063 2809
rect 10119 2850 10256 2866
rect 10119 2816 10205 2850
rect 10239 2816 10256 2850
rect 10119 2800 10256 2816
rect 10306 2850 10447 2865
rect 10306 2816 10397 2850
rect 10431 2816 10447 2850
rect 10119 2772 10185 2800
rect 9917 2763 10185 2772
rect 10306 2799 10447 2816
rect 10476 2850 10640 2866
rect 10476 2816 10589 2850
rect 10623 2816 10640 2850
rect 10476 2800 10640 2816
rect 10706 2850 10990 2866
rect 10706 2816 10940 2850
rect 10974 2816 10990 2850
rect 10706 2800 10990 2816
rect 11046 2850 11183 2866
rect 11046 2816 11132 2850
rect 11166 2816 11183 2850
rect 11046 2800 11183 2816
rect 11233 2850 11374 2865
rect 11233 2816 11324 2850
rect 11358 2816 11374 2850
rect 10306 2763 10372 2799
rect 10409 2798 10443 2799
rect 9917 2711 9935 2763
rect 9987 2711 10185 2763
rect 9917 2706 10185 2711
rect 10224 2716 10372 2763
rect 10224 2678 10262 2716
rect 9917 2647 10262 2678
rect 10331 2647 10372 2716
rect 9917 2612 10372 2647
rect 10476 2584 10542 2800
rect 9775 2496 9798 2562
rect 9864 2496 9885 2562
rect 9775 2490 9885 2496
rect 8986 2435 9052 2453
rect 9098 2478 9297 2490
rect 9098 2466 9256 2478
rect 8738 2248 8818 2314
rect 8884 2248 8948 2314
rect 8738 1702 8948 2248
rect 8698 1690 8948 1702
rect 9098 1715 9182 2466
rect 9217 1715 9256 2466
rect 9290 1702 9297 2478
rect 8162 786 8246 1537
rect 8281 786 8320 1537
rect 7790 774 8001 777
rect 7750 762 8001 774
rect 7102 668 7727 734
rect 6774 580 6780 649
rect 6849 640 6855 649
rect 6849 580 7557 640
rect 6780 574 7557 580
rect 5998 482 6066 546
rect 5999 480 6066 482
rect 6132 480 7370 546
rect 7409 489 7557 574
rect 7304 452 7370 480
rect 7491 453 7557 489
rect 7594 453 7628 454
rect 5832 386 6941 452
rect 7007 436 7248 452
rect 7007 402 7198 436
rect 7232 402 7248 436
rect 7007 386 7248 402
rect 7304 436 7441 452
rect 7304 402 7390 436
rect 7424 402 7441 436
rect 7304 386 7441 402
rect 7491 436 7632 453
rect 7491 402 7582 436
rect 7616 402 7632 436
rect 7491 387 7632 402
rect 7661 452 7727 668
rect 7661 436 7825 452
rect 7661 402 7774 436
rect 7808 402 7825 436
rect 7661 386 7825 402
rect 5832 376 5901 386
rect 7891 355 8001 762
rect 8050 770 8116 776
rect 8162 774 8320 786
rect 8354 774 8361 1550
rect 8162 762 8361 774
rect 8698 1550 8948 1562
rect 8698 774 8704 1550
rect 8738 857 8948 1550
rect 9276 1550 9297 1702
rect 9634 2478 9885 2490
rect 9634 1702 9640 2478
rect 9674 2475 9885 2478
rect 9917 2518 10542 2584
rect 9674 1702 9884 2475
rect 9917 2423 9983 2518
rect 10706 2490 10816 2800
rect 11046 2772 11112 2800
rect 10844 2706 10860 2772
rect 10926 2706 11112 2772
rect 11233 2799 11374 2816
rect 11403 2850 11567 2866
rect 11403 2816 11516 2850
rect 11550 2816 11567 2850
rect 11403 2800 11567 2816
rect 11233 2763 11299 2799
rect 11336 2798 11370 2799
rect 11151 2678 11299 2763
rect 10844 2612 10858 2678
rect 10924 2612 11299 2678
rect 11403 2584 11469 2800
rect 10844 2518 10850 2584
rect 10915 2518 11469 2584
rect 11633 2490 11743 2897
rect 9917 2351 9983 2357
rect 10029 2478 10228 2490
rect 10029 2466 10187 2478
rect 9634 1690 9884 1702
rect 10029 1715 10113 2466
rect 10148 1715 10187 2466
rect 10221 1702 10228 2478
rect 8738 791 8837 857
rect 8903 791 8948 857
rect 8738 777 8948 791
rect 8989 1111 9055 1117
rect 8738 774 8949 777
rect 8698 762 8949 774
rect 8116 704 8675 734
rect 8050 668 8675 704
rect 8050 633 8505 640
rect 8050 574 8401 633
rect 8357 569 8401 574
rect 8465 569 8505 633
rect 8050 537 8318 546
rect 8050 485 8079 537
rect 8131 485 8318 537
rect 8357 489 8505 569
rect 8050 480 8318 485
rect 8252 452 8318 480
rect 8439 453 8505 489
rect 8542 453 8576 454
rect 8050 443 8196 452
rect 8050 391 8063 443
rect 8128 436 8196 443
rect 8128 402 8146 436
rect 8180 402 8196 436
rect 8128 391 8196 402
rect 8050 386 8196 391
rect 8252 436 8389 452
rect 8252 402 8338 436
rect 8372 402 8389 436
rect 8252 386 8389 402
rect 8439 436 8580 453
rect 8439 402 8530 436
rect 8564 402 8580 436
rect 8439 387 8580 402
rect 8609 452 8675 668
rect 8609 436 8773 452
rect 8609 402 8722 436
rect 8756 402 8773 436
rect 8609 386 8773 402
rect 8839 355 8949 762
rect 8989 734 9055 1045
rect 9098 786 9182 1537
rect 9217 786 9256 1537
rect 9098 774 9256 786
rect 9290 774 9297 1550
rect 9098 762 9297 774
rect 9634 1550 9884 1562
rect 9634 774 9640 1550
rect 9674 777 9884 1550
rect 10206 1551 10228 1702
rect 10565 2478 10816 2490
rect 10565 1702 10571 2478
rect 10605 2475 10816 2478
rect 10956 2478 11155 2490
rect 10605 1702 10815 2475
rect 10565 1690 10815 1702
rect 10956 2466 11114 2478
rect 10956 1715 11040 2466
rect 11075 1715 11114 2466
rect 11148 1702 11155 2478
rect 9917 989 9983 995
rect 9674 774 9885 777
rect 9634 763 9885 774
rect 9634 762 9807 763
rect 8986 668 9611 734
rect 8986 574 8993 640
rect 9059 574 9441 640
rect 8986 480 9001 546
rect 9067 480 9254 546
rect 9293 489 9441 574
rect 9188 452 9254 480
rect 9375 453 9441 489
rect 9478 453 9512 454
rect 8986 443 9132 452
rect 8986 391 8992 443
rect 9057 436 9132 443
rect 9057 402 9082 436
rect 9116 402 9132 436
rect 9057 391 9132 402
rect 8986 386 9132 391
rect 9188 436 9325 452
rect 9188 402 9274 436
rect 9308 402 9325 436
rect 9188 386 9325 402
rect 9375 436 9516 453
rect 9375 402 9466 436
rect 9500 402 9516 436
rect 9375 387 9516 402
rect 9545 452 9611 668
rect 9775 699 9807 762
rect 9873 699 9885 763
rect 9545 436 9709 452
rect 9545 402 9658 436
rect 9692 402 9709 436
rect 9545 386 9709 402
rect 9775 355 9885 699
rect 9917 735 9983 923
rect 10029 787 10113 1538
rect 10148 787 10187 1538
rect 10029 775 10187 787
rect 10221 775 10228 1551
rect 10029 763 10228 775
rect 10565 1551 10815 1563
rect 10565 775 10571 1551
rect 10605 778 10815 1551
rect 11134 1550 11155 1702
rect 11492 2478 11743 2490
rect 11492 1702 11498 2478
rect 11532 2475 11743 2478
rect 11860 2861 13092 3085
rect 11860 2658 12189 2861
rect 12410 2658 13092 2861
rect 11532 1719 11742 2475
rect 11860 2160 13092 2658
rect 11799 2152 13092 2160
rect 11799 2101 11811 2152
rect 12168 2143 13092 2152
rect 12168 2101 12180 2143
rect 11799 2094 12180 2101
rect 11860 2056 11903 2094
rect 12726 2009 13092 2143
rect 11875 1997 12689 2009
rect 12726 2002 13137 2009
rect 11875 1907 11881 1997
rect 11915 1907 12073 1997
rect 12107 1907 12265 1997
rect 12299 1907 12457 1997
rect 12491 1907 12649 1997
rect 12683 1907 12689 1997
rect 11875 1895 12689 1907
rect 12923 1965 13137 2002
rect 12923 1931 12986 1965
rect 13077 1931 13137 1965
rect 12923 1893 13137 1931
rect 11779 1855 12209 1867
rect 11779 1765 11785 1855
rect 11819 1765 11977 1855
rect 12011 1765 12169 1855
rect 12203 1765 12209 1855
rect 11779 1753 12209 1765
rect 12355 1861 12827 1867
rect 12355 1855 12892 1861
rect 12355 1765 12361 1855
rect 12395 1765 12553 1855
rect 12587 1765 12745 1855
rect 12779 1845 12892 1855
rect 12779 1765 12842 1845
rect 12355 1753 12842 1765
rect 11532 1703 12263 1719
rect 11532 1702 12170 1703
rect 11492 1690 12170 1702
rect 11737 1669 12170 1690
rect 12204 1669 12263 1703
rect 11737 1653 12263 1669
rect 12702 1619 12842 1753
rect 12876 1619 12892 1845
rect 12923 1859 12929 1893
rect 13008 1889 13137 1893
rect 13008 1859 13014 1889
rect 12923 1701 13014 1859
rect 12923 1667 12929 1701
rect 13008 1667 13014 1701
rect 12923 1651 13014 1667
rect 13046 1797 13235 1861
rect 13046 1763 13052 1797
rect 13129 1763 13235 1797
rect 11703 1598 12363 1614
rect 11703 1564 12313 1598
rect 12347 1564 12363 1598
rect 11703 1562 12363 1564
rect 10956 786 11040 1537
rect 11075 786 11114 1537
rect 10605 775 10816 778
rect 10565 763 10816 775
rect 9917 669 10542 735
rect 9917 633 10372 641
rect 9917 575 10264 633
rect 10224 573 10264 575
rect 10324 573 10372 633
rect 9917 481 9937 547
rect 10003 481 10185 547
rect 10224 490 10372 573
rect 10119 453 10185 481
rect 10306 454 10372 490
rect 10409 454 10443 455
rect 9917 443 10063 453
rect 9917 391 9951 443
rect 10016 437 10063 443
rect 10047 403 10063 437
rect 10016 391 10063 403
rect 9917 387 10063 391
rect 10119 437 10256 453
rect 10119 403 10205 437
rect 10239 403 10256 437
rect 10119 387 10256 403
rect 10306 437 10447 454
rect 10306 403 10397 437
rect 10431 403 10447 437
rect 10306 388 10447 403
rect 10476 453 10542 669
rect 10476 437 10640 453
rect 10476 403 10589 437
rect 10623 403 10640 437
rect 10476 387 10640 403
rect 10706 452 10816 763
rect 10956 774 11114 786
rect 11148 774 11155 1550
rect 10956 762 11155 774
rect 11492 1550 12363 1562
rect 11492 774 11498 1550
rect 11532 1548 12363 1550
rect 11532 1517 11815 1548
rect 11532 777 11742 1517
rect 12259 1514 12305 1520
rect 12702 1514 12892 1619
rect 13046 1605 13235 1763
rect 12259 1508 12892 1514
rect 12259 1332 12265 1508
rect 12299 1399 12892 1508
rect 12923 1571 13052 1605
rect 13129 1571 13235 1605
rect 12923 1443 13235 1571
rect 12923 1409 12935 1443
rect 13111 1409 13235 1443
rect 12923 1403 13123 1409
rect 12299 1365 12842 1399
rect 12876 1365 12892 1399
rect 12299 1348 12892 1365
rect 12923 1355 13123 1362
rect 12299 1332 12827 1348
rect 12259 1320 12827 1332
rect 12305 1316 12827 1320
rect 12923 1321 12935 1355
rect 13111 1321 13123 1355
rect 13151 1348 13235 1409
rect 12305 1315 12825 1316
rect 12305 1314 12774 1315
rect 12171 1249 12394 1256
rect 12171 1201 12183 1249
rect 12074 1188 12183 1201
rect 12382 1201 12394 1249
rect 12923 1253 13123 1321
rect 12923 1219 12954 1253
rect 13086 1219 13123 1253
rect 12921 1212 13123 1219
rect 12382 1188 12473 1201
rect 12074 1085 12233 1188
rect 12352 1085 12473 1188
rect 12921 1163 13121 1212
rect 12921 1141 12960 1163
rect 12074 1011 12473 1085
rect 12923 1044 12960 1141
rect 13079 1141 13121 1163
rect 13079 1044 13113 1141
rect 12923 986 13113 1044
rect 11532 774 11743 777
rect 11492 762 11743 774
rect 10844 668 10850 734
rect 10916 668 11469 734
rect 10844 574 10888 640
rect 10954 574 11299 640
rect 10844 480 10859 546
rect 10925 480 11112 546
rect 11151 489 11299 574
rect 11046 452 11112 480
rect 11233 453 11299 489
rect 11336 453 11370 454
rect 10706 436 10990 452
rect 10706 402 10940 436
rect 10974 402 10990 436
rect 10706 386 10990 402
rect 11046 436 11183 452
rect 11046 402 11132 436
rect 11166 402 11183 436
rect 11046 386 11183 402
rect 11233 436 11374 453
rect 11233 402 11324 436
rect 11358 402 11374 436
rect 11233 387 11374 402
rect 11403 452 11469 668
rect 11403 436 11567 452
rect 11403 402 11516 436
rect 11550 402 11567 436
rect 11403 386 11567 402
rect 10706 356 10816 386
rect 7138 348 8001 355
rect 7138 236 7245 348
rect 7280 236 7438 348
rect 7473 236 7630 348
rect 7665 236 7822 348
rect 7857 236 8001 348
rect 7138 221 8001 236
rect 8086 348 8949 355
rect 8086 236 8193 348
rect 8228 236 8386 348
rect 8421 236 8578 348
rect 8613 236 8770 348
rect 8805 236 8949 348
rect 8086 221 8949 236
rect 9022 348 9885 355
rect 9022 236 9129 348
rect 9164 236 9322 348
rect 9357 236 9514 348
rect 9549 236 9706 348
rect 9741 236 9885 348
rect 9022 221 9885 236
rect 9953 349 10816 356
rect 11633 355 11743 762
rect 9953 237 10060 349
rect 10095 237 10253 349
rect 10288 237 10445 349
rect 10480 237 10637 349
rect 10672 237 10816 349
rect 9953 222 10816 237
rect 10880 348 11743 355
rect 10880 236 10987 348
rect 11022 236 11180 348
rect 11215 236 11372 348
rect 11407 236 11564 348
rect 11599 236 11743 348
rect 10880 221 11743 236
rect 339 -131 2013 -40
rect 7137 159 10779 168
rect 11883 167 12147 178
rect 7137 158 9965 159
rect 7137 48 7150 158
rect 7184 48 7342 158
rect 7376 48 7534 158
rect 7568 48 7726 158
rect 7760 48 7918 158
rect 7952 48 8098 158
rect 8132 48 8290 158
rect 8324 48 8482 158
rect 8516 48 8674 158
rect 8708 48 8866 158
rect 8900 48 9034 158
rect 9068 48 9226 158
rect 9260 48 9418 158
rect 9452 48 9610 158
rect 9644 48 9802 158
rect 9836 49 9965 158
rect 9999 49 10157 159
rect 10191 49 10349 159
rect 10383 49 10541 159
rect 10575 49 10733 159
rect 10767 49 10779 159
rect 9836 48 10779 49
rect 7137 -23 10779 48
rect 10880 158 11894 167
rect 10880 48 10892 158
rect 10926 48 11084 158
rect 11118 48 11276 158
rect 11310 48 11468 158
rect 11502 48 11660 158
rect 11694 48 11894 158
rect 10880 37 11894 48
rect 7137 -24 10204 -23
rect 7137 -59 7389 -24
rect 7677 -59 8337 -24
rect 8625 -59 9273 -24
rect 9561 -58 10204 -24
rect 10492 -58 10779 -23
rect 9561 -59 10779 -58
rect 7137 -73 10779 -59
rect 7137 -75 7964 -73
rect 8085 -75 8912 -73
rect 9021 -75 9848 -73
rect 9952 -74 10779 -73
rect 10879 -24 11894 37
rect 10879 -59 11131 -24
rect 11419 -59 11894 -24
rect 10879 -75 11894 -59
rect 12136 -75 12147 167
rect 11883 -86 12147 -75
rect 248 -137 339 -131
rect -2061 -238 5481 -232
rect -2061 -298 5485 -238
rect -5349 -487 5327 -421
rect -8633 -684 5162 -618
rect -11963 -851 5014 -785
rect -15223 -1014 4904 -948
rect -15512 -1204 4639 -1138
rect -15649 -1375 1625 -1309
rect 1691 -1375 4493 -1309
rect 3886 -1551 3970 -1545
rect -23628 -2225 -23414 -2203
rect -24448 -2300 -23814 -2293
rect -24448 -2347 -24419 -2300
rect -23850 -2347 -23814 -2300
rect -24448 -2419 -24410 -2347
rect -23856 -2413 -23814 -2347
rect -23628 -2304 -23605 -2225
rect -23436 -2304 -23414 -2225
rect -21608 -2225 -21394 -2203
rect -23628 -2319 -23414 -2304
rect -23728 -2367 -23659 -2351
rect -23856 -2419 -23813 -2413
rect -24448 -2499 -24435 -2419
rect -24401 -2499 -24243 -2467
rect -24209 -2499 -24051 -2467
rect -24017 -2499 -23859 -2467
rect -23825 -2499 -23813 -2419
rect -24448 -2505 -23813 -2499
rect -24448 -2506 -23814 -2505
rect -23728 -2535 -23709 -2367
rect -24355 -2541 -23709 -2535
rect -24355 -2621 -24339 -2541
rect -24305 -2621 -24147 -2541
rect -24113 -2621 -23955 -2541
rect -23921 -2593 -23709 -2541
rect -23675 -2593 -23659 -2367
rect -23628 -2353 -23622 -2319
rect -23543 -2323 -23414 -2319
rect -22411 -2300 -21777 -2293
rect -23543 -2353 -23537 -2323
rect -22411 -2347 -22382 -2300
rect -21813 -2347 -21777 -2300
rect -23628 -2511 -23537 -2353
rect -23628 -2545 -23622 -2511
rect -23543 -2545 -23537 -2511
rect -23628 -2561 -23537 -2545
rect -23505 -2415 -23316 -2351
rect -23505 -2449 -23499 -2415
rect -23422 -2449 -23316 -2415
rect -23921 -2621 -23659 -2593
rect -23505 -2607 -23316 -2449
rect -22411 -2419 -22373 -2347
rect -21819 -2413 -21777 -2347
rect -21608 -2304 -21585 -2225
rect -21416 -2304 -21394 -2225
rect -19867 -2225 -19653 -2203
rect -21608 -2319 -21394 -2304
rect -21708 -2367 -21639 -2351
rect -21819 -2419 -21776 -2413
rect -22411 -2499 -22398 -2419
rect -22364 -2499 -22206 -2467
rect -22172 -2499 -22014 -2467
rect -21980 -2499 -21822 -2467
rect -21788 -2499 -21776 -2419
rect -22411 -2505 -21776 -2499
rect -22411 -2506 -21777 -2505
rect -21708 -2535 -21689 -2367
rect -24355 -2627 -23659 -2621
rect -24641 -2791 -24635 -2648
rect -24492 -2656 -24401 -2648
rect -24492 -2674 -24319 -2656
rect -24492 -2709 -24369 -2674
rect -24335 -2709 -24319 -2674
rect -24492 -2791 -24319 -2709
rect -24291 -2674 -24031 -2655
rect -24291 -2709 -24080 -2674
rect -24046 -2709 -24031 -2674
rect -24291 -2729 -24031 -2709
rect -24291 -2798 -24241 -2729
rect -23955 -2757 -23659 -2627
rect -24291 -2820 -24285 -2798
rect -24483 -2833 -24285 -2820
rect -24251 -2833 -24241 -2798
rect -24213 -2769 -23659 -2757
rect -24213 -2803 -24201 -2769
rect -23825 -2803 -23659 -2769
rect -24213 -2809 -23659 -2803
rect -23628 -2641 -23499 -2607
rect -23422 -2641 -23316 -2607
rect -22318 -2541 -21689 -2535
rect -22318 -2621 -22302 -2541
rect -22268 -2621 -22110 -2541
rect -22076 -2621 -21918 -2541
rect -21884 -2593 -21689 -2541
rect -21655 -2593 -21639 -2367
rect -21608 -2353 -21602 -2319
rect -21523 -2323 -21394 -2319
rect -20681 -2300 -20047 -2293
rect -21523 -2353 -21517 -2323
rect -20681 -2347 -20652 -2300
rect -20083 -2347 -20047 -2300
rect -21608 -2511 -21517 -2353
rect -21608 -2545 -21602 -2511
rect -21523 -2545 -21517 -2511
rect -21608 -2561 -21517 -2545
rect -21485 -2415 -21296 -2351
rect -21485 -2449 -21479 -2415
rect -21402 -2449 -21296 -2415
rect -21884 -2621 -21639 -2593
rect -21485 -2607 -21296 -2449
rect -20681 -2419 -20643 -2347
rect -20089 -2413 -20047 -2347
rect -19867 -2304 -19844 -2225
rect -19675 -2304 -19653 -2225
rect -18088 -2225 -17874 -2203
rect -19867 -2319 -19653 -2304
rect -19967 -2367 -19898 -2351
rect -20089 -2419 -20046 -2413
rect -20681 -2499 -20668 -2419
rect -20634 -2499 -20476 -2467
rect -20442 -2499 -20284 -2467
rect -20250 -2499 -20092 -2467
rect -20058 -2499 -20046 -2419
rect -20681 -2505 -20046 -2499
rect -20681 -2506 -20047 -2505
rect -19967 -2535 -19948 -2367
rect -22318 -2627 -21639 -2621
rect -23628 -2707 -23316 -2641
rect -22793 -2656 -22379 -2655
rect -22793 -2674 -22282 -2656
rect -23628 -2747 -23054 -2707
rect -23628 -2769 -23253 -2747
rect -23628 -2803 -23616 -2769
rect -23440 -2803 -23253 -2769
rect -23628 -2809 -23428 -2803
rect -24483 -2859 -24241 -2833
rect -24588 -2940 -24241 -2859
rect -23728 -2813 -23659 -2809
rect -23728 -2847 -23709 -2813
rect -23675 -2847 -23659 -2813
rect -23728 -2864 -23659 -2847
rect -23628 -2857 -23428 -2850
rect -24603 -2956 -24241 -2940
rect -23628 -2891 -23616 -2857
rect -23440 -2891 -23428 -2857
rect -23400 -2864 -23253 -2803
rect -24603 -2987 -24394 -2956
rect -24603 -3165 -24550 -2987
rect -24428 -3165 -24394 -2987
rect -24213 -2961 -23813 -2955
rect -24213 -2995 -24201 -2961
rect -23825 -2995 -23813 -2961
rect -24213 -3033 -24184 -2995
rect -24213 -3067 -24186 -3033
rect -23844 -3057 -23813 -2995
rect -23628 -2974 -23601 -2891
rect -23452 -2974 -23428 -2891
rect -23349 -2866 -23253 -2864
rect -23121 -2866 -23054 -2747
rect -22793 -2767 -22731 -2674
rect -22413 -2709 -22332 -2674
rect -22298 -2709 -22282 -2674
rect -22413 -2767 -22282 -2709
rect -22793 -2791 -22282 -2767
rect -22254 -2674 -21994 -2655
rect -22254 -2709 -22043 -2674
rect -22009 -2709 -21994 -2674
rect -22254 -2729 -21994 -2709
rect -22254 -2798 -22204 -2729
rect -21918 -2757 -21639 -2627
rect -23349 -2911 -23054 -2866
rect -22627 -2820 -22400 -2819
rect -22254 -2820 -22248 -2798
rect -22627 -2833 -22248 -2820
rect -22214 -2833 -22204 -2798
rect -22176 -2769 -21639 -2757
rect -22176 -2803 -22164 -2769
rect -21788 -2803 -21639 -2769
rect -22176 -2809 -21639 -2803
rect -21608 -2641 -21479 -2607
rect -21402 -2641 -21296 -2607
rect -20588 -2541 -19948 -2535
rect -20588 -2621 -20572 -2541
rect -20538 -2621 -20380 -2541
rect -20346 -2621 -20188 -2541
rect -20154 -2593 -19948 -2541
rect -19914 -2593 -19898 -2367
rect -19867 -2353 -19861 -2319
rect -19782 -2323 -19653 -2319
rect -18921 -2300 -18287 -2293
rect -19782 -2353 -19776 -2323
rect -18921 -2347 -18892 -2300
rect -18323 -2347 -18287 -2300
rect -19867 -2511 -19776 -2353
rect -19867 -2545 -19861 -2511
rect -19782 -2545 -19776 -2511
rect -19867 -2561 -19776 -2545
rect -19744 -2415 -19555 -2351
rect -19744 -2449 -19738 -2415
rect -19661 -2449 -19555 -2415
rect -20154 -2621 -19898 -2593
rect -19744 -2607 -19555 -2449
rect -18921 -2419 -18883 -2347
rect -18329 -2413 -18287 -2347
rect -18088 -2304 -18065 -2225
rect -17896 -2304 -17874 -2225
rect -18088 -2319 -17874 -2304
rect -18188 -2367 -18119 -2351
rect -18329 -2419 -18286 -2413
rect -18921 -2499 -18908 -2419
rect -18874 -2499 -18716 -2467
rect -18682 -2499 -18524 -2467
rect -18490 -2499 -18332 -2467
rect -18298 -2499 -18286 -2419
rect -18921 -2505 -18286 -2499
rect -18921 -2506 -18287 -2505
rect -18188 -2535 -18169 -2367
rect -20588 -2627 -19898 -2621
rect -21608 -2769 -21296 -2641
rect -21608 -2803 -21596 -2769
rect -21420 -2775 -21296 -2769
rect -20952 -2656 -20644 -2652
rect -20952 -2674 -20552 -2656
rect -20952 -2675 -20602 -2674
rect -20952 -2772 -20889 -2675
rect -20682 -2709 -20602 -2675
rect -20568 -2709 -20552 -2674
rect -20682 -2772 -20552 -2709
rect -21420 -2803 -21293 -2775
rect -21608 -2809 -21408 -2803
rect -22627 -2852 -22204 -2833
rect -23628 -2993 -23597 -2974
rect -23465 -2993 -23428 -2974
rect -23628 -3000 -23428 -2993
rect -23851 -3067 -23813 -3057
rect -24213 -3078 -23813 -3067
rect -22627 -3080 -22594 -2852
rect -22431 -2956 -22204 -2852
rect -21708 -2813 -21639 -2809
rect -21708 -2847 -21689 -2813
rect -21655 -2847 -21639 -2813
rect -21708 -2864 -21639 -2847
rect -21608 -2857 -21408 -2850
rect -21608 -2891 -21596 -2857
rect -21420 -2891 -21408 -2857
rect -21380 -2859 -21293 -2803
rect -21209 -2779 -21203 -2775
rect -21209 -2859 -21202 -2779
rect -20952 -2791 -20552 -2772
rect -20524 -2674 -20264 -2655
rect -20524 -2709 -20313 -2674
rect -20279 -2709 -20264 -2674
rect -20524 -2729 -20264 -2709
rect -20952 -2792 -20644 -2791
rect -20524 -2798 -20474 -2729
rect -20188 -2757 -19898 -2627
rect -20524 -2820 -20518 -2798
rect -21380 -2863 -21202 -2859
rect -20944 -2833 -20518 -2820
rect -20484 -2833 -20474 -2798
rect -20446 -2769 -19898 -2757
rect -20446 -2803 -20434 -2769
rect -20058 -2803 -19898 -2769
rect -20446 -2809 -19898 -2803
rect -19867 -2641 -19738 -2607
rect -19661 -2641 -19555 -2607
rect -18828 -2541 -18169 -2535
rect -18828 -2621 -18812 -2541
rect -18778 -2621 -18620 -2541
rect -18586 -2621 -18428 -2541
rect -18394 -2593 -18169 -2541
rect -18135 -2593 -18119 -2367
rect -18088 -2353 -18082 -2319
rect -18003 -2323 -17874 -2319
rect -18003 -2353 -17997 -2323
rect -18088 -2511 -17997 -2353
rect -18088 -2545 -18082 -2511
rect -18003 -2545 -17997 -2511
rect -18088 -2561 -17997 -2545
rect -17965 -2415 -17776 -2351
rect -17965 -2449 -17959 -2415
rect -17882 -2449 -17776 -2415
rect -18394 -2621 -18119 -2593
rect -17965 -2607 -17776 -2449
rect -18828 -2627 -18119 -2621
rect -19867 -2769 -19555 -2641
rect -19867 -2803 -19855 -2769
rect -19679 -2803 -19555 -2769
rect -19111 -2656 -18907 -2653
rect -19111 -2673 -18792 -2656
rect -19111 -2780 -19043 -2673
rect -18894 -2674 -18792 -2673
rect -18894 -2709 -18842 -2674
rect -18808 -2709 -18792 -2674
rect -18894 -2780 -18792 -2709
rect -19867 -2809 -19667 -2803
rect -21380 -2864 -21296 -2863
rect -22431 -3080 -22400 -2956
rect -22176 -2961 -21776 -2955
rect -22176 -2995 -22164 -2961
rect -21788 -2995 -21776 -2961
rect -22176 -3033 -22147 -2995
rect -22176 -3067 -22149 -3033
rect -21807 -3057 -21776 -2995
rect -21608 -2974 -21581 -2891
rect -21432 -2974 -21408 -2891
rect -20944 -2956 -20474 -2833
rect -19967 -2813 -19898 -2809
rect -19967 -2847 -19948 -2813
rect -19914 -2847 -19898 -2813
rect -19967 -2864 -19898 -2847
rect -19867 -2857 -19667 -2850
rect -19867 -2891 -19855 -2857
rect -19679 -2891 -19667 -2857
rect -19639 -2864 -19555 -2803
rect -19471 -2864 -19465 -2780
rect -19111 -2791 -18792 -2780
rect -18764 -2674 -18504 -2655
rect -18764 -2709 -18553 -2674
rect -18519 -2709 -18504 -2674
rect -18764 -2729 -18504 -2709
rect -19111 -2792 -18907 -2791
rect -18764 -2798 -18714 -2729
rect -18428 -2757 -18119 -2627
rect -18764 -2820 -18758 -2798
rect -19292 -2833 -18758 -2820
rect -18724 -2833 -18714 -2798
rect -18686 -2769 -18119 -2757
rect -18686 -2803 -18674 -2769
rect -18298 -2803 -18119 -2769
rect -18686 -2809 -18119 -2803
rect -18088 -2641 -17959 -2607
rect -17882 -2641 -17776 -2607
rect -18088 -2678 -17776 -2641
rect -18088 -2696 -17536 -2678
rect -18088 -2769 -17693 -2696
rect -18088 -2803 -18076 -2769
rect -17900 -2803 -17693 -2769
rect -18088 -2809 -17888 -2803
rect -20944 -2966 -20716 -2956
rect -21608 -2993 -21577 -2974
rect -21445 -2993 -21408 -2974
rect -21608 -3000 -21408 -2993
rect -21814 -3067 -21776 -3057
rect -22176 -3078 -21776 -3067
rect -20945 -3042 -20716 -2966
rect -20446 -2961 -20046 -2955
rect -20446 -2995 -20434 -2961
rect -20058 -2995 -20046 -2961
rect -20446 -3033 -20417 -2995
rect -22627 -3113 -22400 -3080
rect -24603 -3194 -24394 -3165
rect -20945 -3165 -20917 -3042
rect -20741 -3165 -20717 -3042
rect -20446 -3067 -20419 -3033
rect -20077 -3057 -20046 -2995
rect -19867 -2974 -19840 -2891
rect -19691 -2974 -19667 -2891
rect -19867 -2993 -19836 -2974
rect -19704 -2993 -19667 -2974
rect -19867 -3000 -19667 -2993
rect -19292 -2934 -18714 -2833
rect -18188 -2813 -18119 -2809
rect -18188 -2847 -18169 -2813
rect -18135 -2847 -18119 -2813
rect -18188 -2864 -18119 -2847
rect -18088 -2857 -17888 -2850
rect -20084 -3067 -20046 -3057
rect -20446 -3078 -20046 -3067
rect -19292 -3087 -19241 -2934
rect -19043 -2956 -18714 -2934
rect -18088 -2891 -18076 -2857
rect -17900 -2891 -17888 -2857
rect -17860 -2852 -17693 -2803
rect -17579 -2852 -17536 -2696
rect -17860 -2864 -17536 -2852
rect -17826 -2865 -17536 -2864
rect -19043 -3087 -18956 -2956
rect -18686 -2961 -18286 -2955
rect -18686 -2995 -18674 -2961
rect -18298 -2995 -18286 -2961
rect -18686 -3033 -18657 -2995
rect -18686 -3067 -18659 -3033
rect -18317 -3057 -18286 -2995
rect -18088 -2974 -18061 -2891
rect -17912 -2974 -17888 -2891
rect -18088 -2993 -18057 -2974
rect -17925 -2993 -17888 -2974
rect -18088 -3000 -17888 -2993
rect -18324 -3067 -18286 -3057
rect -18686 -3078 -18286 -3067
rect -19292 -3115 -18956 -3087
rect -20945 -3188 -20717 -3165
rect -23304 -3391 -11066 -3307
rect -24861 -4016 -24578 -3997
rect -24862 -4064 -24578 -4016
rect -24862 -4337 -24807 -4064
rect -24618 -4337 -24578 -4064
rect -23584 -4037 -23370 -4015
rect -24397 -4112 -23763 -4105
rect -24397 -4159 -24368 -4112
rect -23799 -4159 -23763 -4112
rect -24397 -4231 -24359 -4159
rect -23805 -4225 -23763 -4159
rect -23584 -4116 -23561 -4037
rect -23392 -4116 -23370 -4037
rect -23584 -4131 -23370 -4116
rect -23684 -4179 -23615 -4163
rect -23805 -4231 -23762 -4225
rect -24397 -4311 -24384 -4231
rect -24350 -4311 -24192 -4279
rect -24158 -4311 -24000 -4279
rect -23966 -4311 -23808 -4279
rect -23774 -4311 -23762 -4231
rect -24397 -4317 -23762 -4311
rect -24397 -4318 -23763 -4317
rect -24862 -4379 -24578 -4337
rect -23684 -4347 -23665 -4179
rect -24304 -4353 -23665 -4347
rect -24862 -4468 -24696 -4379
rect -24304 -4433 -24288 -4353
rect -24254 -4433 -24096 -4353
rect -24062 -4433 -23904 -4353
rect -23870 -4405 -23665 -4353
rect -23631 -4405 -23615 -4179
rect -23584 -4165 -23578 -4131
rect -23499 -4135 -23370 -4131
rect -23499 -4165 -23493 -4135
rect -23304 -4163 -23210 -3391
rect -23584 -4323 -23493 -4165
rect -23584 -4357 -23578 -4323
rect -23499 -4357 -23493 -4323
rect -23584 -4373 -23493 -4357
rect -23461 -4227 -23210 -4163
rect -23461 -4261 -23455 -4227
rect -23378 -4261 -23210 -4227
rect -23870 -4433 -23615 -4405
rect -23461 -4419 -23210 -4261
rect -24304 -4439 -23615 -4433
rect -24862 -4486 -24268 -4468
rect -24862 -4521 -24318 -4486
rect -24284 -4521 -24268 -4486
rect -24862 -4603 -24268 -4521
rect -24240 -4486 -23980 -4467
rect -24240 -4521 -24029 -4486
rect -23995 -4521 -23980 -4486
rect -24240 -4541 -23980 -4521
rect -24862 -7733 -24696 -4603
rect -24240 -4610 -24190 -4541
rect -23904 -4569 -23615 -4439
rect -24240 -4632 -24234 -4610
rect -24615 -4645 -24234 -4632
rect -24200 -4645 -24190 -4610
rect -24162 -4581 -23615 -4569
rect -24162 -4615 -24150 -4581
rect -23774 -4615 -23615 -4581
rect -24162 -4621 -23615 -4615
rect -23584 -4453 -23455 -4419
rect -23378 -4453 -23210 -4419
rect -23584 -4581 -23210 -4453
rect -23584 -4615 -23572 -4581
rect -23396 -4615 -23210 -4581
rect -23584 -4621 -23384 -4615
rect -23356 -4616 -23210 -4615
rect -23088 -3538 -14356 -3454
rect -24615 -4768 -24190 -4645
rect -23684 -4625 -23615 -4621
rect -23684 -4659 -23665 -4625
rect -23631 -4659 -23615 -4625
rect -23684 -4676 -23615 -4659
rect -23584 -4669 -23384 -4662
rect -23584 -4703 -23572 -4669
rect -23396 -4703 -23384 -4669
rect -23356 -4676 -23272 -4616
rect -24615 -4997 -24479 -4768
rect -24162 -4773 -23762 -4767
rect -24162 -4807 -24150 -4773
rect -23774 -4807 -23762 -4773
rect -24162 -4845 -24133 -4807
rect -24162 -4879 -24135 -4845
rect -23793 -4869 -23762 -4807
rect -23584 -4786 -23557 -4703
rect -23408 -4786 -23384 -4703
rect -23584 -4805 -23553 -4786
rect -23421 -4805 -23384 -4786
rect -23584 -4812 -23384 -4805
rect -23800 -4879 -23762 -4869
rect -24162 -4890 -23762 -4879
rect -24615 -5751 -24479 -5133
rect -23586 -5329 -23372 -5307
rect -24397 -5404 -23763 -5397
rect -24397 -5451 -24368 -5404
rect -23799 -5451 -23763 -5404
rect -24397 -5523 -24359 -5451
rect -23805 -5517 -23763 -5451
rect -23586 -5408 -23563 -5329
rect -23394 -5408 -23372 -5329
rect -23586 -5423 -23372 -5408
rect -23686 -5471 -23617 -5455
rect -23805 -5523 -23762 -5517
rect -24397 -5603 -24384 -5523
rect -24350 -5603 -24192 -5571
rect -24158 -5603 -24000 -5571
rect -23966 -5603 -23808 -5571
rect -23774 -5603 -23762 -5523
rect -24397 -5609 -23762 -5603
rect -24397 -5610 -23763 -5609
rect -23686 -5639 -23667 -5471
rect -24304 -5645 -23667 -5639
rect -24304 -5725 -24288 -5645
rect -24254 -5725 -24096 -5645
rect -24062 -5725 -23904 -5645
rect -23870 -5697 -23667 -5645
rect -23633 -5697 -23617 -5471
rect -23586 -5457 -23580 -5423
rect -23501 -5427 -23372 -5423
rect -23501 -5457 -23495 -5427
rect -23088 -5454 -22951 -3538
rect -21259 -3686 -17647 -3602
rect -21846 -4037 -21632 -4015
rect -22661 -4112 -22027 -4105
rect -22661 -4159 -22632 -4112
rect -22063 -4159 -22027 -4112
rect -22661 -4231 -22623 -4159
rect -22069 -4225 -22027 -4159
rect -21846 -4116 -21823 -4037
rect -21654 -4116 -21632 -4037
rect -21846 -4131 -21632 -4116
rect -21946 -4179 -21877 -4163
rect -22069 -4231 -22026 -4225
rect -22661 -4311 -22648 -4231
rect -22614 -4311 -22456 -4279
rect -22422 -4311 -22264 -4279
rect -22230 -4311 -22072 -4279
rect -22038 -4311 -22026 -4231
rect -22661 -4317 -22026 -4311
rect -22661 -4318 -22027 -4317
rect -21946 -4347 -21927 -4179
rect -22568 -4353 -21927 -4347
rect -22568 -4433 -22552 -4353
rect -22518 -4433 -22360 -4353
rect -22326 -4433 -22168 -4353
rect -22134 -4405 -21927 -4353
rect -21893 -4405 -21877 -4179
rect -21846 -4165 -21840 -4131
rect -21761 -4135 -21632 -4131
rect -21761 -4165 -21755 -4135
rect -21846 -4323 -21755 -4165
rect -21846 -4357 -21840 -4323
rect -21761 -4357 -21755 -4323
rect -21846 -4373 -21755 -4357
rect -21723 -4227 -21534 -4163
rect -21723 -4261 -21717 -4227
rect -21640 -4261 -21534 -4227
rect -22134 -4433 -21877 -4405
rect -21723 -4419 -21534 -4261
rect -22568 -4439 -21877 -4433
rect -22696 -4469 -22532 -4468
rect -22888 -4481 -22532 -4469
rect -22888 -4594 -22836 -4481
rect -22690 -4486 -22532 -4481
rect -22690 -4521 -22582 -4486
rect -22548 -4521 -22532 -4486
rect -22690 -4594 -22532 -4521
rect -22888 -4603 -22532 -4594
rect -22504 -4486 -22244 -4467
rect -22504 -4521 -22293 -4486
rect -22259 -4521 -22244 -4486
rect -22504 -4541 -22244 -4521
rect -22504 -4610 -22454 -4541
rect -22168 -4569 -21877 -4439
rect -22504 -4632 -22498 -4610
rect -23352 -5455 -22951 -5454
rect -23586 -5615 -23495 -5457
rect -23586 -5649 -23580 -5615
rect -23501 -5649 -23495 -5615
rect -23586 -5665 -23495 -5649
rect -23463 -5519 -22951 -5455
rect -23463 -5553 -23457 -5519
rect -23380 -5553 -22951 -5519
rect -23870 -5725 -23617 -5697
rect -23463 -5711 -22951 -5553
rect -24304 -5731 -23617 -5725
rect -24615 -5760 -24362 -5751
rect -24615 -5778 -24268 -5760
rect -24615 -5813 -24318 -5778
rect -24284 -5813 -24268 -5778
rect -24615 -5887 -24268 -5813
rect -24432 -5895 -24268 -5887
rect -24240 -5778 -23980 -5759
rect -24240 -5813 -24029 -5778
rect -23995 -5813 -23980 -5778
rect -24240 -5833 -23980 -5813
rect -24240 -5902 -24190 -5833
rect -23904 -5861 -23617 -5731
rect -24240 -5924 -24234 -5902
rect -24637 -5937 -24234 -5924
rect -24200 -5937 -24190 -5902
rect -24162 -5873 -23617 -5861
rect -24162 -5907 -24150 -5873
rect -23774 -5907 -23617 -5873
rect -24162 -5913 -23617 -5907
rect -23586 -5745 -23457 -5711
rect -23380 -5745 -22951 -5711
rect -23586 -5873 -22951 -5745
rect -23586 -5907 -23574 -5873
rect -23398 -5907 -22951 -5873
rect -22869 -4645 -22498 -4632
rect -22464 -4645 -22454 -4610
rect -22426 -4581 -21877 -4569
rect -22426 -4615 -22414 -4581
rect -22038 -4615 -21877 -4581
rect -22426 -4621 -21877 -4615
rect -21846 -4453 -21717 -4419
rect -21640 -4453 -21534 -4419
rect -21846 -4529 -21534 -4453
rect -21259 -4529 -21128 -3686
rect -17756 -3763 -17647 -3686
rect -20649 -3827 -19439 -3799
rect -20649 -3899 -20603 -3827
rect -19481 -3899 -19439 -3827
rect -20649 -3933 -19439 -3899
rect -20649 -4002 -20395 -3933
rect -20649 -4104 -20637 -4002
rect -20603 -4104 -20445 -4002
rect -20411 -4104 -20395 -4002
rect -20649 -4125 -20395 -4104
rect -20269 -4004 -19819 -3978
rect -20269 -4106 -20253 -4004
rect -20219 -4005 -19819 -4004
rect -20219 -4106 -20061 -4005
rect -20269 -4107 -20061 -4106
rect -20027 -4107 -19869 -4005
rect -19835 -4107 -19819 -4005
rect -20269 -4125 -19819 -4107
rect -19693 -4005 -19439 -3933
rect -19693 -4107 -19677 -4005
rect -19643 -4107 -19485 -4005
rect -19451 -4107 -19439 -4005
rect -19693 -4125 -19439 -4107
rect -19090 -3827 -17880 -3799
rect -19090 -3899 -19044 -3827
rect -17922 -3899 -17880 -3827
rect -17756 -3858 -17744 -3763
rect -17655 -3858 -17647 -3763
rect -14466 -3762 -14356 -3538
rect -17756 -3869 -17647 -3858
rect -17358 -3827 -16148 -3799
rect -19090 -3933 -17880 -3899
rect -19090 -4002 -18836 -3933
rect -19090 -4104 -19078 -4002
rect -19044 -4104 -18886 -4002
rect -18852 -4104 -18836 -4002
rect -19090 -4125 -18836 -4104
rect -18710 -4004 -18260 -3978
rect -18710 -4106 -18694 -4004
rect -18660 -4005 -18260 -4004
rect -18660 -4106 -18502 -4005
rect -18710 -4107 -18502 -4106
rect -18468 -4107 -18310 -4005
rect -18276 -4107 -18260 -4005
rect -18710 -4125 -18260 -4107
rect -18134 -4005 -17880 -3933
rect -18134 -4107 -18118 -4005
rect -18084 -4107 -17926 -4005
rect -17892 -4107 -17880 -4005
rect -18134 -4125 -17880 -4107
rect -17358 -3899 -17312 -3827
rect -16190 -3899 -16148 -3827
rect -17358 -3933 -16148 -3899
rect -17358 -4002 -17104 -3933
rect -17358 -4104 -17346 -4002
rect -17312 -4104 -17154 -4002
rect -17120 -4104 -17104 -4002
rect -17358 -4125 -17104 -4104
rect -16978 -4004 -16528 -3978
rect -16978 -4106 -16962 -4004
rect -16928 -4005 -16528 -4004
rect -16928 -4106 -16770 -4005
rect -16978 -4107 -16770 -4106
rect -16736 -4107 -16578 -4005
rect -16544 -4107 -16528 -4005
rect -16978 -4125 -16528 -4107
rect -16402 -4005 -16148 -3933
rect -16402 -4107 -16386 -4005
rect -16352 -4107 -16194 -4005
rect -16160 -4107 -16148 -4005
rect -16402 -4125 -16148 -4107
rect -15799 -3827 -14589 -3799
rect -15799 -3899 -15753 -3827
rect -14631 -3899 -14589 -3827
rect -15799 -3933 -14589 -3899
rect -15799 -4002 -15545 -3933
rect -15799 -4104 -15787 -4002
rect -15753 -4104 -15595 -4002
rect -15561 -4104 -15545 -4002
rect -15799 -4125 -15545 -4104
rect -15419 -4004 -14969 -3978
rect -15419 -4106 -15403 -4004
rect -15369 -4005 -14969 -4004
rect -15369 -4106 -15211 -4005
rect -15419 -4107 -15211 -4106
rect -15177 -4107 -15019 -4005
rect -14985 -4107 -14969 -4005
rect -15419 -4125 -14969 -4107
rect -14843 -4005 -14589 -3933
rect -14466 -3946 -14460 -3762
rect -14361 -3946 -14356 -3762
rect -11174 -3761 -11066 -3391
rect -14466 -3953 -14356 -3946
rect -14067 -3827 -12857 -3799
rect -14067 -3899 -14021 -3827
rect -12899 -3899 -12857 -3827
rect -14067 -3933 -12857 -3899
rect -14843 -4107 -14827 -4005
rect -14793 -4107 -14635 -4005
rect -14601 -4107 -14589 -4005
rect -14843 -4125 -14589 -4107
rect -14067 -4002 -13813 -3933
rect -14067 -4104 -14055 -4002
rect -14021 -4104 -13863 -4002
rect -13829 -4104 -13813 -4002
rect -14067 -4125 -13813 -4104
rect -13687 -4004 -13237 -3978
rect -13687 -4106 -13671 -4004
rect -13637 -4005 -13237 -4004
rect -13637 -4106 -13479 -4005
rect -13687 -4107 -13479 -4106
rect -13445 -4107 -13287 -4005
rect -13253 -4107 -13237 -4005
rect -13687 -4125 -13237 -4107
rect -13111 -4005 -12857 -3933
rect -13111 -4107 -13095 -4005
rect -13061 -4107 -12903 -4005
rect -12869 -4107 -12857 -4005
rect -13111 -4125 -12857 -4107
rect -12508 -3827 -11298 -3799
rect -12508 -3899 -12462 -3827
rect -11340 -3899 -11298 -3827
rect -12508 -3933 -11298 -3899
rect -11174 -3905 -11165 -3761
rect -11074 -3905 -11066 -3761
rect -11174 -3916 -11066 -3905
rect -10776 -3827 -9566 -3799
rect -10776 -3899 -10730 -3827
rect -9608 -3899 -9566 -3827
rect -12508 -4002 -12254 -3933
rect -12508 -4104 -12496 -4002
rect -12462 -4104 -12304 -4002
rect -12270 -4104 -12254 -4002
rect -12508 -4125 -12254 -4104
rect -12128 -4004 -11678 -3978
rect -12128 -4106 -12112 -4004
rect -12078 -4005 -11678 -4004
rect -12078 -4106 -11920 -4005
rect -12128 -4107 -11920 -4106
rect -11886 -4107 -11728 -4005
rect -11694 -4107 -11678 -4005
rect -12128 -4125 -11678 -4107
rect -11552 -4005 -11298 -3933
rect -11552 -4107 -11536 -4005
rect -11502 -4107 -11344 -4005
rect -11310 -4107 -11298 -4005
rect -11552 -4125 -11298 -4107
rect -10776 -3933 -9566 -3899
rect -10776 -4002 -10522 -3933
rect -10776 -4104 -10764 -4002
rect -10730 -4104 -10572 -4002
rect -10538 -4104 -10522 -4002
rect -10776 -4125 -10522 -4104
rect -10396 -4004 -9946 -3978
rect -10396 -4106 -10380 -4004
rect -10346 -4005 -9946 -4004
rect -10346 -4106 -10188 -4005
rect -10396 -4107 -10188 -4106
rect -10154 -4107 -9996 -4005
rect -9962 -4107 -9946 -4005
rect -10396 -4125 -9946 -4107
rect -9820 -4005 -9566 -3933
rect -9820 -4107 -9804 -4005
rect -9770 -4107 -9612 -4005
rect -9578 -4107 -9566 -4005
rect -9820 -4125 -9566 -4107
rect -9217 -3827 -8007 -3799
rect -9217 -3899 -9171 -3827
rect -8049 -3899 -8007 -3827
rect -9217 -3933 -8007 -3899
rect -9217 -4002 -8963 -3933
rect -9217 -4104 -9205 -4002
rect -9171 -4104 -9013 -4002
rect -8979 -4104 -8963 -4002
rect -9217 -4125 -8963 -4104
rect -8837 -4004 -8387 -3978
rect -8837 -4106 -8821 -4004
rect -8787 -4005 -8387 -4004
rect -8787 -4106 -8629 -4005
rect -8837 -4107 -8629 -4106
rect -8595 -4107 -8437 -4005
rect -8403 -4107 -8387 -4005
rect -8837 -4125 -8387 -4107
rect -8261 -4005 -8007 -3933
rect -8261 -4107 -8245 -4005
rect -8211 -4107 -8053 -4005
rect -8019 -4107 -8007 -4005
rect -8261 -4125 -8007 -4107
rect -20557 -4188 -19531 -4163
rect -20557 -4312 -20541 -4188
rect -20507 -4312 -20349 -4188
rect -20315 -4312 -20157 -4188
rect -20123 -4312 -19965 -4188
rect -19931 -4312 -19773 -4188
rect -19739 -4189 -19531 -4188
rect -19739 -4312 -19581 -4189
rect -20557 -4313 -19581 -4312
rect -19547 -4313 -19531 -4189
rect -20557 -4342 -19531 -4313
rect -18998 -4188 -17972 -4163
rect -18998 -4312 -18982 -4188
rect -18948 -4312 -18790 -4188
rect -18756 -4312 -18598 -4188
rect -18564 -4312 -18406 -4188
rect -18372 -4312 -18214 -4188
rect -18180 -4189 -17972 -4188
rect -18180 -4312 -18022 -4189
rect -18998 -4313 -18022 -4312
rect -17988 -4313 -17972 -4189
rect -18998 -4342 -17972 -4313
rect -17266 -4188 -16240 -4163
rect -17266 -4312 -17250 -4188
rect -17216 -4312 -17058 -4188
rect -17024 -4312 -16866 -4188
rect -16832 -4312 -16674 -4188
rect -16640 -4312 -16482 -4188
rect -16448 -4189 -16240 -4188
rect -16448 -4312 -16290 -4189
rect -17266 -4313 -16290 -4312
rect -16256 -4313 -16240 -4189
rect -17266 -4342 -16240 -4313
rect -15707 -4188 -14681 -4163
rect -15707 -4312 -15691 -4188
rect -15657 -4312 -15499 -4188
rect -15465 -4312 -15307 -4188
rect -15273 -4312 -15115 -4188
rect -15081 -4312 -14923 -4188
rect -14889 -4189 -14681 -4188
rect -14889 -4312 -14731 -4189
rect -15707 -4313 -14731 -4312
rect -14697 -4313 -14681 -4189
rect -15707 -4342 -14681 -4313
rect -13975 -4188 -12949 -4163
rect -13975 -4312 -13959 -4188
rect -13925 -4312 -13767 -4188
rect -13733 -4312 -13575 -4188
rect -13541 -4312 -13383 -4188
rect -13349 -4312 -13191 -4188
rect -13157 -4189 -12949 -4188
rect -13157 -4312 -12999 -4189
rect -13975 -4313 -12999 -4312
rect -12965 -4313 -12949 -4189
rect -13975 -4342 -12949 -4313
rect -12416 -4188 -11390 -4163
rect -12416 -4312 -12400 -4188
rect -12366 -4312 -12208 -4188
rect -12174 -4312 -12016 -4188
rect -11982 -4312 -11824 -4188
rect -11790 -4312 -11632 -4188
rect -11598 -4189 -11390 -4188
rect -11598 -4312 -11440 -4189
rect -12416 -4313 -11440 -4312
rect -11406 -4313 -11390 -4189
rect -12416 -4342 -11390 -4313
rect -10684 -4188 -9658 -4163
rect -10684 -4312 -10668 -4188
rect -10634 -4312 -10476 -4188
rect -10442 -4312 -10284 -4188
rect -10250 -4312 -10092 -4188
rect -10058 -4312 -9900 -4188
rect -9866 -4189 -9658 -4188
rect -9866 -4312 -9708 -4189
rect -10684 -4313 -9708 -4312
rect -9674 -4313 -9658 -4189
rect -10684 -4342 -9658 -4313
rect -9125 -4188 -8099 -4163
rect -9125 -4312 -9109 -4188
rect -9075 -4312 -8917 -4188
rect -8883 -4312 -8725 -4188
rect -8691 -4312 -8533 -4188
rect -8499 -4312 -8341 -4188
rect -8307 -4189 -8099 -4188
rect -8307 -4312 -8149 -4189
rect -9125 -4313 -8149 -4312
rect -8115 -4313 -8099 -4189
rect -9125 -4342 -8099 -4313
rect -20649 -4397 -20395 -4375
rect -20649 -4499 -20637 -4397
rect -20603 -4463 -20445 -4397
rect -20411 -4463 -20395 -4397
rect -20603 -4499 -20395 -4463
rect -20269 -4403 -19819 -4386
rect -20269 -4463 -20253 -4403
rect -20219 -4420 -19869 -4403
rect -20219 -4463 -20061 -4420
rect -20027 -4463 -19869 -4420
rect -19835 -4463 -19819 -4403
rect -20269 -4478 -19819 -4463
rect -19693 -4396 -19439 -4375
rect -19693 -4463 -19677 -4396
rect -19643 -4463 -19485 -4396
rect -19451 -4463 -19439 -4396
rect -20649 -4522 -20395 -4499
rect -19693 -4522 -19439 -4463
rect -19090 -4397 -18836 -4375
rect -19090 -4499 -19078 -4397
rect -19044 -4463 -18886 -4397
rect -18852 -4463 -18836 -4397
rect -19044 -4499 -18836 -4463
rect -18710 -4403 -18260 -4386
rect -18710 -4463 -18694 -4403
rect -18660 -4420 -18310 -4403
rect -18660 -4463 -18502 -4420
rect -18468 -4463 -18310 -4420
rect -18276 -4463 -18260 -4403
rect -18710 -4478 -18260 -4463
rect -18134 -4396 -17880 -4375
rect -18134 -4463 -18118 -4396
rect -18084 -4463 -17926 -4396
rect -17892 -4463 -17880 -4396
rect -19090 -4522 -18836 -4499
rect -18134 -4522 -17880 -4463
rect -17358 -4397 -17104 -4375
rect -17358 -4499 -17346 -4397
rect -17312 -4463 -17154 -4397
rect -17120 -4463 -17104 -4397
rect -17312 -4499 -17104 -4463
rect -16978 -4403 -16528 -4386
rect -16978 -4463 -16962 -4403
rect -16928 -4420 -16578 -4403
rect -16928 -4463 -16770 -4420
rect -16736 -4463 -16578 -4420
rect -16544 -4463 -16528 -4403
rect -16978 -4478 -16528 -4463
rect -16402 -4396 -16148 -4375
rect -16402 -4463 -16386 -4396
rect -16352 -4463 -16194 -4396
rect -16160 -4463 -16148 -4396
rect -17358 -4522 -17104 -4499
rect -16402 -4522 -16148 -4463
rect -15799 -4397 -15545 -4375
rect -15799 -4499 -15787 -4397
rect -15753 -4463 -15595 -4397
rect -15561 -4463 -15545 -4397
rect -15753 -4499 -15545 -4463
rect -15419 -4403 -14969 -4386
rect -15419 -4463 -15403 -4403
rect -15369 -4420 -15019 -4403
rect -15369 -4463 -15211 -4420
rect -15177 -4463 -15019 -4420
rect -14985 -4463 -14969 -4403
rect -15419 -4478 -14969 -4463
rect -14843 -4396 -14589 -4375
rect -14843 -4463 -14827 -4396
rect -14793 -4463 -14635 -4396
rect -14601 -4463 -14589 -4396
rect -15799 -4522 -15545 -4499
rect -14843 -4522 -14589 -4463
rect -14067 -4397 -13813 -4375
rect -14067 -4499 -14055 -4397
rect -14021 -4463 -13863 -4397
rect -13829 -4463 -13813 -4397
rect -14021 -4499 -13813 -4463
rect -13687 -4403 -13237 -4386
rect -13687 -4463 -13671 -4403
rect -13637 -4420 -13287 -4403
rect -13637 -4463 -13479 -4420
rect -13445 -4463 -13287 -4420
rect -13253 -4463 -13237 -4403
rect -13687 -4478 -13237 -4463
rect -13111 -4396 -12857 -4375
rect -13111 -4463 -13095 -4396
rect -13061 -4463 -12903 -4396
rect -12869 -4463 -12857 -4396
rect -14067 -4522 -13813 -4499
rect -13111 -4522 -12857 -4463
rect -12508 -4397 -12254 -4375
rect -12508 -4499 -12496 -4397
rect -12462 -4463 -12304 -4397
rect -12270 -4463 -12254 -4397
rect -12462 -4499 -12254 -4463
rect -12128 -4403 -11678 -4386
rect -12128 -4463 -12112 -4403
rect -12078 -4420 -11728 -4403
rect -12078 -4463 -11920 -4420
rect -11886 -4463 -11728 -4420
rect -11694 -4463 -11678 -4403
rect -12128 -4478 -11678 -4463
rect -11552 -4396 -11298 -4375
rect -11552 -4463 -11536 -4396
rect -11502 -4463 -11344 -4396
rect -11310 -4463 -11298 -4396
rect -12508 -4522 -12254 -4499
rect -11552 -4522 -11298 -4463
rect -10776 -4397 -10522 -4375
rect -10776 -4499 -10764 -4397
rect -10730 -4463 -10572 -4397
rect -10538 -4463 -10522 -4397
rect -10730 -4499 -10522 -4463
rect -10396 -4403 -9946 -4386
rect -10396 -4463 -10380 -4403
rect -10346 -4420 -9996 -4403
rect -10346 -4463 -10188 -4420
rect -10154 -4463 -9996 -4420
rect -9962 -4463 -9946 -4403
rect -10396 -4478 -9946 -4463
rect -9820 -4396 -9566 -4375
rect -9820 -4463 -9804 -4396
rect -9770 -4463 -9612 -4396
rect -9578 -4463 -9566 -4396
rect -10776 -4522 -10522 -4499
rect -9820 -4522 -9566 -4463
rect -9217 -4397 -8963 -4375
rect -9217 -4499 -9205 -4397
rect -9171 -4463 -9013 -4397
rect -8979 -4463 -8963 -4397
rect -9171 -4499 -8963 -4463
rect -8837 -4403 -8387 -4386
rect -8837 -4463 -8821 -4403
rect -8787 -4420 -8437 -4403
rect -8787 -4463 -8629 -4420
rect -8595 -4463 -8437 -4420
rect -8403 -4463 -8387 -4403
rect -8837 -4478 -8387 -4463
rect -8261 -4396 -8007 -4375
rect -8261 -4463 -8245 -4396
rect -8211 -4463 -8053 -4396
rect -8019 -4463 -8007 -4396
rect -9217 -4522 -8963 -4499
rect -8261 -4522 -8007 -4463
rect -21846 -4581 -21128 -4529
rect -21846 -4615 -21834 -4581
rect -21658 -4615 -21128 -4581
rect -21846 -4621 -21646 -4615
rect -22869 -4768 -22454 -4645
rect -21946 -4625 -21877 -4621
rect -21946 -4659 -21927 -4625
rect -21893 -4659 -21877 -4625
rect -21946 -4676 -21877 -4659
rect -21846 -4669 -21646 -4662
rect -21846 -4703 -21834 -4669
rect -21658 -4703 -21646 -4669
rect -21618 -4676 -21128 -4615
rect -20872 -4622 -20737 -4598
rect -22869 -4991 -22733 -4768
rect -22426 -4773 -22026 -4767
rect -22426 -4807 -22414 -4773
rect -22038 -4807 -22026 -4773
rect -22426 -4845 -22397 -4807
rect -22426 -4879 -22399 -4845
rect -22057 -4869 -22026 -4807
rect -21846 -4786 -21819 -4703
rect -21670 -4786 -21646 -4703
rect -20872 -4732 -20854 -4622
rect -20758 -4730 -20737 -4622
rect -17581 -4622 -17446 -4598
rect -19398 -4657 -19207 -4652
rect -19399 -4667 -19207 -4657
rect -19399 -4674 -19297 -4667
rect -19224 -4674 -19207 -4667
rect -20807 -4732 -20737 -4730
rect -20872 -4752 -20737 -4732
rect -20576 -4715 -19787 -4697
rect -20576 -4723 -19933 -4715
rect -21846 -4805 -21815 -4786
rect -21683 -4805 -21646 -4786
rect -20576 -4776 -20539 -4723
rect -20406 -4768 -19933 -4723
rect -19819 -4768 -19787 -4715
rect -20406 -4776 -19787 -4768
rect -20576 -4796 -19787 -4776
rect -19717 -4716 -19602 -4697
rect -19717 -4784 -19699 -4716
rect -19619 -4784 -19602 -4716
rect -19399 -4757 -19372 -4674
rect -21846 -4812 -21646 -4805
rect -22064 -4879 -22026 -4869
rect -22426 -4890 -22026 -4879
rect -20795 -4855 -20590 -4836
rect -20795 -4963 -20751 -4855
rect -20675 -4881 -20590 -4855
rect -19717 -4881 -19602 -4784
rect -19486 -4771 -19372 -4757
rect -19222 -4771 -19207 -4674
rect -19486 -4787 -19207 -4771
rect -19017 -4715 -18228 -4697
rect -19017 -4723 -18374 -4715
rect -19017 -4776 -18980 -4723
rect -18847 -4768 -18374 -4723
rect -18260 -4768 -18228 -4715
rect -18847 -4776 -18228 -4768
rect -19486 -4850 -19315 -4787
rect -19017 -4796 -18228 -4776
rect -18158 -4716 -18043 -4697
rect -18158 -4784 -18140 -4716
rect -18060 -4784 -18043 -4716
rect -17581 -4732 -17563 -4622
rect -17467 -4730 -17446 -4622
rect -14290 -4622 -14155 -4598
rect -16107 -4657 -15916 -4652
rect -16108 -4667 -15916 -4657
rect -16108 -4674 -16006 -4667
rect -15933 -4674 -15916 -4667
rect -17516 -4732 -17446 -4730
rect -17581 -4752 -17446 -4732
rect -17285 -4715 -16496 -4697
rect -17285 -4723 -16642 -4715
rect -20675 -4963 -19602 -4881
rect -20795 -4967 -19602 -4963
rect -19528 -4887 -19315 -4850
rect -19528 -4942 -19517 -4887
rect -19452 -4942 -19315 -4887
rect -19528 -4966 -19315 -4942
rect -19236 -4862 -19031 -4836
rect -19236 -4959 -19196 -4862
rect -19080 -4881 -19031 -4862
rect -18158 -4881 -18043 -4784
rect -17927 -4850 -17647 -4757
rect -17285 -4776 -17248 -4723
rect -17115 -4768 -16642 -4723
rect -16528 -4768 -16496 -4715
rect -17115 -4776 -16496 -4768
rect -17285 -4796 -16496 -4776
rect -16426 -4716 -16311 -4697
rect -16426 -4784 -16408 -4716
rect -16328 -4784 -16311 -4716
rect -16108 -4757 -16081 -4674
rect -19080 -4959 -18043 -4881
rect -19236 -4967 -18043 -4959
rect -17969 -4887 -17647 -4850
rect -17969 -4942 -17958 -4887
rect -17893 -4942 -17647 -4887
rect -17969 -4966 -17647 -4942
rect -20795 -4979 -20590 -4967
rect -19236 -4979 -19031 -4967
rect -22869 -4997 -22732 -4991
rect -22869 -5133 -22868 -4997
rect -22869 -5139 -22732 -5133
rect -20644 -5036 -20589 -5020
rect -22869 -5759 -22733 -5139
rect -20644 -5142 -20637 -5036
rect -20603 -5142 -20589 -5036
rect -20557 -5021 -20107 -5009
rect -20557 -5055 -20541 -5021
rect -20507 -5055 -20349 -5021
rect -20315 -5022 -20107 -5021
rect -20315 -5055 -20157 -5022
rect -20557 -5056 -20157 -5055
rect -20123 -5056 -20107 -5022
rect -20557 -5077 -20107 -5056
rect -19981 -5021 -19531 -5009
rect -19981 -5055 -19965 -5021
rect -19931 -5055 -19773 -5021
rect -19739 -5055 -19581 -5021
rect -19547 -5055 -19531 -5021
rect -19981 -5077 -19531 -5055
rect -19497 -5036 -19442 -5020
rect -20644 -5208 -20589 -5142
rect -20459 -5122 -20394 -5105
rect -20459 -5156 -20445 -5122
rect -20411 -5156 -20394 -5122
rect -20459 -5208 -20394 -5156
rect -20266 -5122 -19819 -5110
rect -20266 -5156 -20253 -5122
rect -20219 -5156 -20061 -5122
rect -20027 -5156 -19869 -5122
rect -19835 -5156 -19819 -5122
rect -20266 -5174 -19819 -5156
rect -19693 -5122 -19628 -5106
rect -19693 -5156 -19677 -5122
rect -19643 -5156 -19628 -5122
rect -19693 -5208 -19628 -5156
rect -19497 -5142 -19485 -5036
rect -19451 -5142 -19442 -5036
rect -19497 -5208 -19442 -5142
rect -20644 -5219 -19442 -5208
rect -20644 -5230 -20143 -5219
rect -20083 -5230 -19442 -5219
rect -20644 -5276 -20603 -5230
rect -19480 -5276 -19442 -5230
rect -20644 -5279 -20143 -5276
rect -20083 -5279 -19442 -5276
rect -20644 -5299 -19442 -5279
rect -19085 -5036 -19030 -5020
rect -19085 -5142 -19078 -5036
rect -19044 -5142 -19030 -5036
rect -18998 -5021 -18548 -5009
rect -18998 -5055 -18982 -5021
rect -18948 -5055 -18790 -5021
rect -18756 -5022 -18548 -5021
rect -18756 -5055 -18598 -5022
rect -18998 -5056 -18598 -5055
rect -18564 -5056 -18548 -5022
rect -18998 -5077 -18548 -5056
rect -18422 -5021 -17972 -5009
rect -18422 -5055 -18406 -5021
rect -18372 -5055 -18214 -5021
rect -18180 -5055 -18022 -5021
rect -17988 -5055 -17972 -5021
rect -18422 -5077 -17972 -5055
rect -17938 -5036 -17883 -5020
rect -19085 -5208 -19030 -5142
rect -18900 -5122 -18835 -5105
rect -18900 -5156 -18886 -5122
rect -18852 -5156 -18835 -5122
rect -18900 -5208 -18835 -5156
rect -18707 -5122 -18260 -5110
rect -18707 -5156 -18694 -5122
rect -18660 -5156 -18502 -5122
rect -18468 -5156 -18310 -5122
rect -18276 -5156 -18260 -5122
rect -18707 -5174 -18260 -5156
rect -18134 -5122 -18069 -5106
rect -18134 -5156 -18118 -5122
rect -18084 -5156 -18069 -5122
rect -18134 -5208 -18069 -5156
rect -17938 -5142 -17926 -5036
rect -17892 -5142 -17883 -5036
rect -17938 -5208 -17883 -5142
rect -19085 -5219 -17883 -5208
rect -19085 -5230 -18584 -5219
rect -18524 -5230 -17883 -5219
rect -19085 -5276 -19044 -5230
rect -17921 -5276 -17883 -5230
rect -17756 -5153 -17647 -4966
rect -17504 -4855 -17299 -4836
rect -17504 -4963 -17460 -4855
rect -17384 -4881 -17299 -4855
rect -16426 -4881 -16311 -4784
rect -16195 -4771 -16081 -4757
rect -15931 -4771 -15916 -4674
rect -16195 -4787 -15916 -4771
rect -15726 -4715 -14937 -4697
rect -15726 -4723 -15083 -4715
rect -15726 -4776 -15689 -4723
rect -15556 -4768 -15083 -4723
rect -14969 -4768 -14937 -4715
rect -15556 -4776 -14937 -4768
rect -16195 -4850 -16024 -4787
rect -15726 -4796 -14937 -4776
rect -14867 -4716 -14752 -4697
rect -14867 -4784 -14849 -4716
rect -14769 -4784 -14752 -4716
rect -14290 -4732 -14272 -4622
rect -14176 -4730 -14155 -4622
rect -10999 -4622 -10864 -4598
rect -12816 -4657 -12625 -4652
rect -12817 -4667 -12625 -4657
rect -12817 -4674 -12715 -4667
rect -12642 -4674 -12625 -4667
rect -14225 -4732 -14155 -4730
rect -14290 -4752 -14155 -4732
rect -13994 -4715 -13205 -4697
rect -13994 -4723 -13351 -4715
rect -17384 -4963 -16311 -4881
rect -17504 -4967 -16311 -4963
rect -16237 -4887 -16024 -4850
rect -16237 -4942 -16226 -4887
rect -16161 -4942 -16024 -4887
rect -16237 -4966 -16024 -4942
rect -15945 -4862 -15740 -4836
rect -15945 -4959 -15905 -4862
rect -15789 -4881 -15740 -4862
rect -14867 -4881 -14752 -4784
rect -14636 -4850 -14356 -4757
rect -13994 -4776 -13957 -4723
rect -13824 -4768 -13351 -4723
rect -13237 -4768 -13205 -4715
rect -13824 -4776 -13205 -4768
rect -13994 -4796 -13205 -4776
rect -13135 -4716 -13020 -4697
rect -13135 -4784 -13117 -4716
rect -13037 -4784 -13020 -4716
rect -12817 -4757 -12790 -4674
rect -15789 -4959 -14752 -4881
rect -15945 -4967 -14752 -4959
rect -14678 -4887 -14356 -4850
rect -14678 -4942 -14667 -4887
rect -14602 -4942 -14356 -4887
rect -14678 -4966 -14356 -4942
rect -17504 -4979 -17299 -4967
rect -15945 -4979 -15740 -4967
rect -17756 -5239 -17747 -5153
rect -17656 -5239 -17647 -5153
rect -17756 -5251 -17647 -5239
rect -17353 -5036 -17298 -5020
rect -17353 -5142 -17346 -5036
rect -17312 -5142 -17298 -5036
rect -17266 -5021 -16816 -5009
rect -17266 -5055 -17250 -5021
rect -17216 -5055 -17058 -5021
rect -17024 -5022 -16816 -5021
rect -17024 -5055 -16866 -5022
rect -17266 -5056 -16866 -5055
rect -16832 -5056 -16816 -5022
rect -17266 -5077 -16816 -5056
rect -16690 -5021 -16240 -5009
rect -16690 -5055 -16674 -5021
rect -16640 -5055 -16482 -5021
rect -16448 -5055 -16290 -5021
rect -16256 -5055 -16240 -5021
rect -16690 -5077 -16240 -5055
rect -16206 -5036 -16151 -5020
rect -17353 -5208 -17298 -5142
rect -17168 -5122 -17103 -5105
rect -17168 -5156 -17154 -5122
rect -17120 -5156 -17103 -5122
rect -17168 -5208 -17103 -5156
rect -16975 -5122 -16528 -5110
rect -16975 -5156 -16962 -5122
rect -16928 -5156 -16770 -5122
rect -16736 -5156 -16578 -5122
rect -16544 -5156 -16528 -5122
rect -16975 -5174 -16528 -5156
rect -16402 -5122 -16337 -5106
rect -16402 -5156 -16386 -5122
rect -16352 -5156 -16337 -5122
rect -16402 -5208 -16337 -5156
rect -16206 -5142 -16194 -5036
rect -16160 -5142 -16151 -5036
rect -16206 -5208 -16151 -5142
rect -17353 -5219 -16151 -5208
rect -17353 -5230 -16852 -5219
rect -16792 -5230 -16151 -5219
rect -19085 -5279 -18584 -5276
rect -18524 -5279 -17883 -5276
rect -19085 -5299 -17883 -5279
rect -17353 -5276 -17312 -5230
rect -16189 -5276 -16151 -5230
rect -17353 -5279 -16852 -5276
rect -16792 -5279 -16151 -5276
rect -17353 -5299 -16151 -5279
rect -15794 -5036 -15739 -5020
rect -15794 -5142 -15787 -5036
rect -15753 -5142 -15739 -5036
rect -15707 -5021 -15257 -5009
rect -15707 -5055 -15691 -5021
rect -15657 -5055 -15499 -5021
rect -15465 -5022 -15257 -5021
rect -15465 -5055 -15307 -5022
rect -15707 -5056 -15307 -5055
rect -15273 -5056 -15257 -5022
rect -15707 -5077 -15257 -5056
rect -15131 -5021 -14681 -5009
rect -15131 -5055 -15115 -5021
rect -15081 -5055 -14923 -5021
rect -14889 -5055 -14731 -5021
rect -14697 -5055 -14681 -5021
rect -15131 -5077 -14681 -5055
rect -14647 -5036 -14592 -5020
rect -15794 -5208 -15739 -5142
rect -15609 -5122 -15544 -5105
rect -15609 -5156 -15595 -5122
rect -15561 -5156 -15544 -5122
rect -15609 -5208 -15544 -5156
rect -15416 -5122 -14969 -5110
rect -15416 -5156 -15403 -5122
rect -15369 -5156 -15211 -5122
rect -15177 -5156 -15019 -5122
rect -14985 -5156 -14969 -5122
rect -15416 -5174 -14969 -5156
rect -14843 -5122 -14778 -5106
rect -14843 -5156 -14827 -5122
rect -14793 -5156 -14778 -5122
rect -14843 -5208 -14778 -5156
rect -14647 -5142 -14635 -5036
rect -14601 -5142 -14592 -5036
rect -14647 -5208 -14592 -5142
rect -15794 -5219 -14592 -5208
rect -15794 -5230 -15293 -5219
rect -15233 -5230 -14592 -5219
rect -15794 -5276 -15753 -5230
rect -14630 -5276 -14592 -5230
rect -14465 -5153 -14356 -4966
rect -14213 -4855 -14008 -4836
rect -14213 -4963 -14169 -4855
rect -14093 -4881 -14008 -4855
rect -13135 -4881 -13020 -4784
rect -12904 -4771 -12790 -4757
rect -12640 -4771 -12625 -4674
rect -12904 -4787 -12625 -4771
rect -12435 -4715 -11646 -4697
rect -12435 -4723 -11792 -4715
rect -12435 -4776 -12398 -4723
rect -12265 -4768 -11792 -4723
rect -11678 -4768 -11646 -4715
rect -12265 -4776 -11646 -4768
rect -12904 -4850 -12733 -4787
rect -12435 -4796 -11646 -4776
rect -11576 -4716 -11461 -4697
rect -11576 -4784 -11558 -4716
rect -11478 -4784 -11461 -4716
rect -10999 -4732 -10981 -4622
rect -10885 -4730 -10864 -4622
rect -9525 -4657 -9334 -4652
rect -9526 -4667 -9334 -4657
rect -9526 -4674 -9424 -4667
rect -9351 -4674 -9334 -4667
rect -10934 -4732 -10864 -4730
rect -10999 -4752 -10864 -4732
rect -10703 -4715 -9914 -4697
rect -10703 -4723 -10060 -4715
rect -14093 -4963 -13020 -4881
rect -14213 -4967 -13020 -4963
rect -12946 -4887 -12733 -4850
rect -12946 -4942 -12935 -4887
rect -12870 -4942 -12733 -4887
rect -12946 -4966 -12733 -4942
rect -12654 -4862 -12449 -4836
rect -12654 -4959 -12614 -4862
rect -12498 -4881 -12449 -4862
rect -11576 -4881 -11461 -4784
rect -11345 -4850 -11065 -4757
rect -10703 -4776 -10666 -4723
rect -10533 -4768 -10060 -4723
rect -9946 -4768 -9914 -4715
rect -10533 -4776 -9914 -4768
rect -10703 -4796 -9914 -4776
rect -9844 -4716 -9729 -4697
rect -9844 -4784 -9826 -4716
rect -9746 -4784 -9729 -4716
rect -9526 -4757 -9499 -4674
rect -12498 -4959 -11461 -4881
rect -12654 -4967 -11461 -4959
rect -11387 -4887 -11065 -4850
rect -11387 -4942 -11376 -4887
rect -11311 -4942 -11065 -4887
rect -11387 -4966 -11065 -4942
rect -14213 -4979 -14008 -4967
rect -12654 -4979 -12449 -4967
rect -14465 -5239 -14456 -5153
rect -14365 -5239 -14356 -5153
rect -14465 -5251 -14356 -5239
rect -14062 -5036 -14007 -5020
rect -14062 -5142 -14055 -5036
rect -14021 -5142 -14007 -5036
rect -13975 -5021 -13525 -5009
rect -13975 -5055 -13959 -5021
rect -13925 -5055 -13767 -5021
rect -13733 -5022 -13525 -5021
rect -13733 -5055 -13575 -5022
rect -13975 -5056 -13575 -5055
rect -13541 -5056 -13525 -5022
rect -13975 -5077 -13525 -5056
rect -13399 -5021 -12949 -5009
rect -13399 -5055 -13383 -5021
rect -13349 -5055 -13191 -5021
rect -13157 -5055 -12999 -5021
rect -12965 -5055 -12949 -5021
rect -13399 -5077 -12949 -5055
rect -12915 -5036 -12860 -5020
rect -14062 -5208 -14007 -5142
rect -13877 -5122 -13812 -5105
rect -13877 -5156 -13863 -5122
rect -13829 -5156 -13812 -5122
rect -13877 -5208 -13812 -5156
rect -13684 -5122 -13237 -5110
rect -13684 -5156 -13671 -5122
rect -13637 -5156 -13479 -5122
rect -13445 -5156 -13287 -5122
rect -13253 -5156 -13237 -5122
rect -13684 -5174 -13237 -5156
rect -13111 -5122 -13046 -5106
rect -13111 -5156 -13095 -5122
rect -13061 -5156 -13046 -5122
rect -13111 -5208 -13046 -5156
rect -12915 -5142 -12903 -5036
rect -12869 -5142 -12860 -5036
rect -12915 -5208 -12860 -5142
rect -14062 -5219 -12860 -5208
rect -14062 -5230 -13561 -5219
rect -13501 -5230 -12860 -5219
rect -15794 -5279 -15293 -5276
rect -15233 -5279 -14592 -5276
rect -15794 -5299 -14592 -5279
rect -14062 -5276 -14021 -5230
rect -12898 -5276 -12860 -5230
rect -14062 -5279 -13561 -5276
rect -13501 -5279 -12860 -5276
rect -14062 -5299 -12860 -5279
rect -12503 -5036 -12448 -5020
rect -12503 -5142 -12496 -5036
rect -12462 -5142 -12448 -5036
rect -12416 -5021 -11966 -5009
rect -12416 -5055 -12400 -5021
rect -12366 -5055 -12208 -5021
rect -12174 -5022 -11966 -5021
rect -12174 -5055 -12016 -5022
rect -12416 -5056 -12016 -5055
rect -11982 -5056 -11966 -5022
rect -12416 -5077 -11966 -5056
rect -11840 -5021 -11390 -5009
rect -11840 -5055 -11824 -5021
rect -11790 -5055 -11632 -5021
rect -11598 -5055 -11440 -5021
rect -11406 -5055 -11390 -5021
rect -11840 -5077 -11390 -5055
rect -11356 -5036 -11301 -5020
rect -12503 -5208 -12448 -5142
rect -12318 -5122 -12253 -5105
rect -12318 -5156 -12304 -5122
rect -12270 -5156 -12253 -5122
rect -12318 -5208 -12253 -5156
rect -12125 -5122 -11678 -5110
rect -12125 -5156 -12112 -5122
rect -12078 -5156 -11920 -5122
rect -11886 -5156 -11728 -5122
rect -11694 -5156 -11678 -5122
rect -12125 -5174 -11678 -5156
rect -11552 -5122 -11487 -5106
rect -11552 -5156 -11536 -5122
rect -11502 -5156 -11487 -5122
rect -11552 -5208 -11487 -5156
rect -11356 -5142 -11344 -5036
rect -11310 -5142 -11301 -5036
rect -11356 -5208 -11301 -5142
rect -12503 -5219 -11301 -5208
rect -12503 -5230 -12002 -5219
rect -11942 -5230 -11301 -5219
rect -12503 -5276 -12462 -5230
rect -11339 -5276 -11301 -5230
rect -11174 -5153 -11065 -4966
rect -10922 -4855 -10717 -4836
rect -10922 -4963 -10878 -4855
rect -10802 -4881 -10717 -4855
rect -9844 -4881 -9729 -4784
rect -9613 -4771 -9499 -4757
rect -9349 -4771 -9334 -4674
rect -9613 -4787 -9334 -4771
rect -9144 -4715 -8355 -4697
rect -9144 -4723 -8501 -4715
rect -9144 -4776 -9107 -4723
rect -8974 -4768 -8501 -4723
rect -8387 -4768 -8355 -4715
rect -8974 -4776 -8355 -4768
rect -9613 -4850 -9442 -4787
rect -9144 -4796 -8355 -4776
rect -8285 -4716 -8170 -4697
rect -8285 -4784 -8267 -4716
rect -8187 -4784 -8170 -4716
rect -10802 -4963 -9729 -4881
rect -10922 -4967 -9729 -4963
rect -9655 -4887 -9442 -4850
rect -9655 -4942 -9644 -4887
rect -9579 -4942 -9442 -4887
rect -9655 -4966 -9442 -4942
rect -9363 -4862 -9158 -4836
rect -9363 -4959 -9323 -4862
rect -9207 -4881 -9158 -4862
rect -8285 -4881 -8170 -4784
rect -8054 -4850 -7774 -4757
rect -9207 -4959 -8170 -4881
rect -9363 -4967 -8170 -4959
rect -8096 -4887 -7774 -4850
rect -8096 -4942 -8085 -4887
rect -8020 -4942 -7774 -4887
rect -8096 -4966 -7774 -4942
rect -10922 -4979 -10717 -4967
rect -9363 -4979 -9158 -4967
rect -11174 -5239 -11165 -5153
rect -11074 -5239 -11065 -5153
rect -11174 -5251 -11065 -5239
rect -10771 -5036 -10716 -5020
rect -10771 -5142 -10764 -5036
rect -10730 -5142 -10716 -5036
rect -10684 -5021 -10234 -5009
rect -10684 -5055 -10668 -5021
rect -10634 -5055 -10476 -5021
rect -10442 -5022 -10234 -5021
rect -10442 -5055 -10284 -5022
rect -10684 -5056 -10284 -5055
rect -10250 -5056 -10234 -5022
rect -10684 -5077 -10234 -5056
rect -10108 -5021 -9658 -5009
rect -10108 -5055 -10092 -5021
rect -10058 -5055 -9900 -5021
rect -9866 -5055 -9708 -5021
rect -9674 -5055 -9658 -5021
rect -10108 -5077 -9658 -5055
rect -9624 -5036 -9569 -5020
rect -10771 -5208 -10716 -5142
rect -10586 -5122 -10521 -5105
rect -10586 -5156 -10572 -5122
rect -10538 -5156 -10521 -5122
rect -10586 -5208 -10521 -5156
rect -10393 -5122 -9946 -5110
rect -10393 -5156 -10380 -5122
rect -10346 -5156 -10188 -5122
rect -10154 -5156 -9996 -5122
rect -9962 -5156 -9946 -5122
rect -10393 -5174 -9946 -5156
rect -9820 -5122 -9755 -5106
rect -9820 -5156 -9804 -5122
rect -9770 -5156 -9755 -5122
rect -9820 -5208 -9755 -5156
rect -9624 -5142 -9612 -5036
rect -9578 -5142 -9569 -5036
rect -9624 -5208 -9569 -5142
rect -10771 -5219 -9569 -5208
rect -10771 -5230 -10270 -5219
rect -10210 -5230 -9569 -5219
rect -12503 -5279 -12002 -5276
rect -11942 -5279 -11301 -5276
rect -12503 -5299 -11301 -5279
rect -10771 -5276 -10730 -5230
rect -9607 -5276 -9569 -5230
rect -10771 -5279 -10270 -5276
rect -10210 -5279 -9569 -5276
rect -10771 -5299 -9569 -5279
rect -9212 -5036 -9157 -5020
rect -9212 -5142 -9205 -5036
rect -9171 -5142 -9157 -5036
rect -9125 -5021 -8675 -5009
rect -9125 -5055 -9109 -5021
rect -9075 -5055 -8917 -5021
rect -8883 -5022 -8675 -5021
rect -8883 -5055 -8725 -5022
rect -9125 -5056 -8725 -5055
rect -8691 -5056 -8675 -5022
rect -9125 -5077 -8675 -5056
rect -8549 -5021 -8099 -5009
rect -8549 -5055 -8533 -5021
rect -8499 -5055 -8341 -5021
rect -8307 -5055 -8149 -5021
rect -8115 -5055 -8099 -5021
rect -8549 -5077 -8099 -5055
rect -8065 -5036 -8010 -5020
rect -9212 -5208 -9157 -5142
rect -9027 -5122 -8962 -5105
rect -9027 -5156 -9013 -5122
rect -8979 -5156 -8962 -5122
rect -9027 -5208 -8962 -5156
rect -8834 -5122 -8387 -5110
rect -8834 -5156 -8821 -5122
rect -8787 -5156 -8629 -5122
rect -8595 -5156 -8437 -5122
rect -8403 -5156 -8387 -5122
rect -8834 -5174 -8387 -5156
rect -8261 -5122 -8196 -5106
rect -8261 -5156 -8245 -5122
rect -8211 -5156 -8196 -5122
rect -8261 -5208 -8196 -5156
rect -8065 -5142 -8053 -5036
rect -8019 -5142 -8010 -5036
rect -8065 -5208 -8010 -5142
rect -9212 -5219 -8010 -5208
rect -9212 -5230 -8711 -5219
rect -8651 -5230 -8010 -5219
rect -9212 -5276 -9171 -5230
rect -8048 -5276 -8010 -5230
rect -7883 -5153 -7774 -4966
rect -7883 -5239 -7874 -5153
rect -7783 -5239 -7774 -5153
rect -7883 -5251 -7774 -5239
rect -9212 -5279 -8711 -5276
rect -8651 -5279 -8010 -5276
rect -9212 -5299 -8010 -5279
rect -21852 -5329 -21638 -5307
rect -22661 -5404 -22027 -5397
rect -22661 -5451 -22632 -5404
rect -22063 -5451 -22027 -5404
rect -22661 -5523 -22623 -5451
rect -22069 -5517 -22027 -5451
rect -21852 -5408 -21829 -5329
rect -21660 -5408 -21638 -5329
rect -21852 -5423 -21638 -5408
rect -21952 -5471 -21883 -5455
rect -22069 -5523 -22026 -5517
rect -22661 -5603 -22648 -5523
rect -22614 -5603 -22456 -5571
rect -22422 -5603 -22264 -5571
rect -22230 -5603 -22072 -5571
rect -22038 -5603 -22026 -5523
rect -22661 -5609 -22026 -5603
rect -22661 -5610 -22027 -5609
rect -21952 -5639 -21933 -5471
rect -22568 -5645 -21933 -5639
rect -22568 -5725 -22552 -5645
rect -22518 -5725 -22360 -5645
rect -22326 -5725 -22168 -5645
rect -22134 -5697 -21933 -5645
rect -21899 -5697 -21883 -5471
rect -21852 -5457 -21846 -5423
rect -21767 -5427 -21638 -5423
rect -21033 -5333 -20824 -5313
rect -21767 -5457 -21761 -5427
rect -21033 -5435 -21003 -5333
rect -20885 -5352 -20824 -5333
rect -8229 -5352 -8138 -5299
rect -20885 -5368 -19620 -5352
rect -20885 -5435 -19735 -5368
rect -21033 -5437 -19735 -5435
rect -19636 -5437 -19620 -5368
rect -21033 -5443 -19620 -5437
rect -19237 -5364 -16329 -5352
rect -19237 -5430 -19223 -5364
rect -19152 -5368 -16329 -5364
rect -19152 -5430 -16444 -5368
rect -19237 -5437 -16444 -5430
rect -16345 -5437 -16329 -5368
rect -19237 -5443 -16329 -5437
rect -15946 -5364 -13038 -5352
rect -15946 -5430 -15932 -5364
rect -15861 -5368 -13038 -5364
rect -15861 -5430 -13153 -5368
rect -15946 -5437 -13153 -5430
rect -13054 -5437 -13038 -5368
rect -15946 -5443 -13038 -5437
rect -12655 -5364 -9747 -5352
rect -12655 -5430 -12641 -5364
rect -12570 -5368 -9747 -5364
rect -12570 -5430 -9862 -5368
rect -12655 -5437 -9862 -5430
rect -9763 -5437 -9747 -5368
rect -12655 -5443 -9747 -5437
rect -9364 -5364 -7684 -5352
rect -9364 -5430 -9350 -5364
rect -9279 -5430 -7684 -5364
rect -9364 -5443 -7684 -5430
rect -21852 -5615 -21761 -5457
rect -21852 -5649 -21846 -5615
rect -21767 -5649 -21761 -5615
rect -21852 -5665 -21761 -5649
rect -21729 -5519 -21540 -5455
rect -21033 -5465 -20824 -5443
rect -21729 -5553 -21723 -5519
rect -21646 -5553 -21540 -5519
rect -22134 -5725 -21883 -5697
rect -21729 -5705 -21540 -5553
rect -20354 -5559 -20080 -5550
rect -20354 -5565 -20345 -5559
rect -20531 -5572 -20345 -5565
rect -20089 -5565 -20080 -5559
rect -19065 -5559 -18791 -5550
rect -19065 -5565 -19056 -5559
rect -20089 -5572 -19897 -5565
rect -20531 -5619 -20502 -5572
rect -19933 -5619 -19897 -5572
rect -20531 -5631 -20345 -5619
rect -20089 -5631 -19897 -5619
rect -20531 -5685 -19897 -5631
rect -19422 -5572 -19056 -5565
rect -18800 -5565 -18791 -5559
rect -18348 -5559 -18074 -5550
rect -18348 -5565 -18339 -5559
rect -19422 -5619 -19393 -5572
rect -19422 -5631 -19056 -5619
rect -18800 -5631 -18788 -5565
rect -19422 -5685 -18788 -5631
rect -18540 -5572 -18339 -5565
rect -18083 -5565 -18074 -5559
rect -17063 -5559 -16789 -5550
rect -17063 -5565 -17054 -5559
rect -18083 -5572 -17906 -5565
rect -18540 -5619 -18511 -5572
rect -17942 -5619 -17906 -5572
rect -18540 -5631 -18339 -5619
rect -18083 -5631 -17906 -5619
rect -18540 -5685 -17906 -5631
rect -17240 -5572 -17054 -5565
rect -16798 -5565 -16789 -5559
rect -15774 -5559 -15500 -5550
rect -15774 -5565 -15765 -5559
rect -16798 -5572 -16606 -5565
rect -17240 -5619 -17211 -5572
rect -16642 -5619 -16606 -5572
rect -17240 -5631 -17054 -5619
rect -16798 -5631 -16606 -5619
rect -17240 -5685 -16606 -5631
rect -16131 -5572 -15765 -5565
rect -15509 -5565 -15500 -5559
rect -15057 -5559 -14783 -5550
rect -15057 -5565 -15048 -5559
rect -16131 -5619 -16102 -5572
rect -16131 -5631 -15765 -5619
rect -15509 -5631 -15497 -5565
rect -16131 -5685 -15497 -5631
rect -15249 -5572 -15048 -5565
rect -14792 -5565 -14783 -5559
rect -13772 -5559 -13498 -5550
rect -13772 -5565 -13763 -5559
rect -14792 -5572 -14615 -5565
rect -15249 -5619 -15220 -5572
rect -14651 -5619 -14615 -5572
rect -15249 -5631 -15048 -5619
rect -14792 -5631 -14615 -5619
rect -15249 -5685 -14615 -5631
rect -13949 -5572 -13763 -5565
rect -13507 -5565 -13498 -5559
rect -12483 -5559 -12209 -5550
rect -12483 -5565 -12474 -5559
rect -13507 -5572 -13315 -5565
rect -13949 -5619 -13920 -5572
rect -13351 -5619 -13315 -5572
rect -13949 -5631 -13763 -5619
rect -13507 -5631 -13315 -5619
rect -13949 -5685 -13315 -5631
rect -12840 -5572 -12474 -5565
rect -12218 -5565 -12209 -5559
rect -11766 -5559 -11492 -5550
rect -11766 -5565 -11757 -5559
rect -12840 -5619 -12811 -5572
rect -12840 -5631 -12474 -5619
rect -12218 -5631 -12206 -5565
rect -12840 -5685 -12206 -5631
rect -11958 -5572 -11757 -5565
rect -11501 -5565 -11492 -5559
rect -10481 -5559 -10207 -5550
rect -10481 -5565 -10472 -5559
rect -11501 -5572 -11324 -5565
rect -11958 -5619 -11929 -5572
rect -11360 -5619 -11324 -5572
rect -11958 -5631 -11757 -5619
rect -11501 -5631 -11324 -5619
rect -11958 -5685 -11324 -5631
rect -10658 -5572 -10472 -5565
rect -10216 -5565 -10207 -5559
rect -9192 -5559 -8918 -5550
rect -9192 -5565 -9183 -5559
rect -10216 -5572 -10024 -5565
rect -10658 -5619 -10629 -5572
rect -10060 -5619 -10024 -5572
rect -10658 -5631 -10472 -5619
rect -10216 -5631 -10024 -5619
rect -10658 -5685 -10024 -5631
rect -9549 -5572 -9183 -5565
rect -8927 -5565 -8918 -5559
rect -8475 -5559 -8201 -5550
rect -8475 -5565 -8466 -5559
rect -9549 -5619 -9520 -5572
rect -9549 -5631 -9183 -5619
rect -8927 -5631 -8915 -5565
rect -9549 -5685 -8915 -5631
rect -8667 -5572 -8466 -5565
rect -8210 -5565 -8201 -5559
rect -8210 -5572 -8033 -5565
rect -8667 -5619 -8638 -5572
rect -8069 -5619 -8033 -5572
rect -8667 -5631 -8466 -5619
rect -8210 -5631 -8033 -5619
rect -8667 -5685 -8033 -5631
rect -20531 -5691 -19896 -5685
rect -21729 -5711 -21304 -5705
rect -22568 -5731 -21883 -5725
rect -22869 -5760 -22614 -5759
rect -22869 -5778 -22532 -5760
rect -22869 -5813 -22582 -5778
rect -22548 -5813 -22532 -5778
rect -22869 -5895 -22532 -5813
rect -22504 -5778 -22244 -5759
rect -22504 -5813 -22293 -5778
rect -22259 -5813 -22244 -5778
rect -22504 -5833 -22244 -5813
rect -23586 -5913 -23386 -5907
rect -24637 -6049 -24190 -5937
rect -23686 -5917 -23617 -5913
rect -23686 -5951 -23667 -5917
rect -23633 -5951 -23617 -5917
rect -23686 -5968 -23617 -5951
rect -23586 -5961 -23386 -5954
rect -24637 -6247 -24612 -6049
rect -24466 -6060 -24190 -6049
rect -23586 -5995 -23574 -5961
rect -23398 -5995 -23386 -5961
rect -23358 -5966 -22951 -5907
rect -22504 -5902 -22454 -5833
rect -22168 -5861 -21883 -5731
rect -22504 -5924 -22498 -5902
rect -22912 -5936 -22498 -5924
rect -23358 -5968 -23012 -5966
rect -24466 -6247 -24432 -6060
rect -24162 -6065 -23762 -6059
rect -24162 -6099 -24150 -6065
rect -23774 -6099 -23762 -6065
rect -24162 -6137 -24133 -6099
rect -24162 -6171 -24135 -6137
rect -23793 -6161 -23762 -6099
rect -23586 -6078 -23559 -5995
rect -23410 -6078 -23386 -5995
rect -22912 -6046 -22884 -5936
rect -22652 -5937 -22498 -5936
rect -22464 -5937 -22454 -5902
rect -22426 -5873 -21883 -5861
rect -22426 -5907 -22414 -5873
rect -22038 -5907 -21883 -5873
rect -22426 -5913 -21883 -5907
rect -21852 -5745 -21723 -5711
rect -21646 -5731 -21304 -5711
rect -21646 -5745 -21560 -5731
rect -21852 -5873 -21560 -5745
rect -21852 -5907 -21840 -5873
rect -21664 -5907 -21560 -5873
rect -21852 -5913 -21652 -5907
rect -22652 -6046 -22454 -5937
rect -21952 -5917 -21883 -5913
rect -21952 -5951 -21933 -5917
rect -21899 -5951 -21883 -5917
rect -21952 -5968 -21883 -5951
rect -21624 -5922 -21560 -5907
rect -21347 -5922 -21304 -5731
rect -20531 -5771 -20518 -5691
rect -20484 -5771 -20326 -5691
rect -20292 -5771 -20134 -5691
rect -20100 -5771 -19942 -5691
rect -19908 -5771 -19896 -5691
rect -20531 -5777 -19896 -5771
rect -19422 -5691 -18787 -5685
rect -19422 -5771 -19409 -5691
rect -19375 -5771 -19217 -5691
rect -19183 -5771 -19025 -5691
rect -18991 -5771 -18833 -5691
rect -18799 -5771 -18787 -5691
rect -19422 -5777 -18787 -5771
rect -18540 -5691 -17905 -5685
rect -18540 -5771 -18527 -5691
rect -18493 -5771 -18335 -5691
rect -18301 -5771 -18143 -5691
rect -18109 -5771 -17951 -5691
rect -17917 -5771 -17905 -5691
rect -18540 -5777 -17905 -5771
rect -17240 -5691 -16605 -5685
rect -17240 -5771 -17227 -5691
rect -17193 -5771 -17035 -5691
rect -17001 -5771 -16843 -5691
rect -16809 -5771 -16651 -5691
rect -16617 -5771 -16605 -5691
rect -17240 -5777 -16605 -5771
rect -16131 -5691 -15496 -5685
rect -16131 -5771 -16118 -5691
rect -16084 -5771 -15926 -5691
rect -15892 -5771 -15734 -5691
rect -15700 -5771 -15542 -5691
rect -15508 -5771 -15496 -5691
rect -16131 -5777 -15496 -5771
rect -15249 -5691 -14614 -5685
rect -15249 -5771 -15236 -5691
rect -15202 -5771 -15044 -5691
rect -15010 -5771 -14852 -5691
rect -14818 -5771 -14660 -5691
rect -14626 -5771 -14614 -5691
rect -15249 -5777 -14614 -5771
rect -13949 -5691 -13314 -5685
rect -13949 -5771 -13936 -5691
rect -13902 -5771 -13744 -5691
rect -13710 -5771 -13552 -5691
rect -13518 -5771 -13360 -5691
rect -13326 -5771 -13314 -5691
rect -13949 -5777 -13314 -5771
rect -12840 -5691 -12205 -5685
rect -12840 -5771 -12827 -5691
rect -12793 -5771 -12635 -5691
rect -12601 -5771 -12443 -5691
rect -12409 -5771 -12251 -5691
rect -12217 -5771 -12205 -5691
rect -12840 -5777 -12205 -5771
rect -11958 -5691 -11323 -5685
rect -11958 -5771 -11945 -5691
rect -11911 -5771 -11753 -5691
rect -11719 -5771 -11561 -5691
rect -11527 -5771 -11369 -5691
rect -11335 -5771 -11323 -5691
rect -11958 -5777 -11323 -5771
rect -10658 -5691 -10023 -5685
rect -10658 -5771 -10645 -5691
rect -10611 -5771 -10453 -5691
rect -10419 -5771 -10261 -5691
rect -10227 -5771 -10069 -5691
rect -10035 -5771 -10023 -5691
rect -10658 -5777 -10023 -5771
rect -9549 -5691 -8914 -5685
rect -9549 -5771 -9536 -5691
rect -9502 -5771 -9344 -5691
rect -9310 -5771 -9152 -5691
rect -9118 -5771 -8960 -5691
rect -8926 -5771 -8914 -5691
rect -9549 -5777 -8914 -5771
rect -8667 -5691 -8032 -5685
rect -8667 -5771 -8654 -5691
rect -8620 -5771 -8462 -5691
rect -8428 -5771 -8270 -5691
rect -8236 -5771 -8078 -5691
rect -8044 -5771 -8032 -5691
rect -8667 -5777 -8032 -5771
rect -20531 -5778 -19897 -5777
rect -19422 -5778 -18788 -5777
rect -18540 -5778 -17906 -5777
rect -17240 -5778 -16606 -5777
rect -16131 -5778 -15497 -5777
rect -15249 -5778 -14615 -5777
rect -13949 -5778 -13315 -5777
rect -12840 -5778 -12206 -5777
rect -11958 -5778 -11324 -5777
rect -10658 -5778 -10024 -5777
rect -9549 -5778 -8915 -5777
rect -8667 -5778 -8033 -5777
rect -20438 -5813 -19860 -5807
rect -20438 -5893 -20422 -5813
rect -20388 -5893 -20230 -5813
rect -20196 -5893 -20038 -5813
rect -20004 -5893 -19860 -5813
rect -20438 -5894 -19860 -5893
rect -20438 -5899 -19979 -5894
rect -21852 -5961 -21652 -5954
rect -22912 -6059 -22454 -6046
rect -21852 -5995 -21840 -5961
rect -21664 -5995 -21652 -5961
rect -21624 -5968 -21304 -5922
rect -20566 -5946 -20402 -5928
rect -20566 -5955 -20452 -5946
rect -22696 -6060 -22454 -6059
rect -23586 -6097 -23555 -6078
rect -23423 -6097 -23386 -6078
rect -23586 -6104 -23386 -6097
rect -22426 -6065 -22026 -6059
rect -22426 -6099 -22414 -6065
rect -22038 -6099 -22026 -6065
rect -23800 -6171 -23762 -6161
rect -24162 -6182 -23762 -6171
rect -22426 -6137 -22397 -6099
rect -22426 -6171 -22399 -6137
rect -22057 -6161 -22026 -6099
rect -21852 -6078 -21825 -5995
rect -21676 -6078 -21652 -5995
rect -20566 -6035 -20534 -5955
rect -20418 -5981 -20402 -5946
rect -20436 -6035 -20402 -5981
rect -20566 -6063 -20402 -6035
rect -20374 -5946 -20114 -5927
rect -20374 -5981 -20163 -5946
rect -20129 -5981 -20114 -5946
rect -20374 -6001 -20114 -5981
rect -21852 -6097 -21821 -6078
rect -21689 -6097 -21652 -6078
rect -20374 -6070 -20324 -6001
rect -20038 -6029 -19979 -5899
rect -20374 -6091 -20368 -6070
rect -21852 -6104 -21652 -6097
rect -22064 -6171 -22026 -6161
rect -22426 -6182 -22026 -6171
rect -20762 -6105 -20368 -6091
rect -20334 -6105 -20324 -6070
rect -20296 -6041 -19979 -6029
rect -20296 -6075 -20284 -6041
rect -19896 -6042 -19860 -5894
rect -19329 -5813 -18751 -5807
rect -19329 -5893 -19313 -5813
rect -19279 -5893 -19121 -5813
rect -19087 -5893 -18929 -5813
rect -18895 -5893 -18751 -5813
rect -19329 -5899 -18751 -5893
rect -18447 -5813 -17869 -5807
rect -18447 -5893 -18431 -5813
rect -18397 -5893 -18239 -5813
rect -18205 -5893 -18047 -5813
rect -18013 -5893 -17869 -5813
rect -18447 -5899 -17869 -5893
rect -17147 -5813 -16569 -5807
rect -17147 -5893 -17131 -5813
rect -17097 -5893 -16939 -5813
rect -16905 -5893 -16747 -5813
rect -16713 -5893 -16569 -5813
rect -17147 -5894 -16569 -5893
rect -17147 -5899 -16688 -5894
rect -19908 -6075 -19860 -6042
rect -19457 -5946 -19293 -5928
rect -19457 -5956 -19343 -5946
rect -19457 -6036 -19423 -5956
rect -19309 -5981 -19293 -5946
rect -19325 -6036 -19293 -5981
rect -19457 -6063 -19293 -6036
rect -19265 -5946 -19005 -5927
rect -19265 -5981 -19054 -5946
rect -19020 -5981 -19005 -5946
rect -19265 -6001 -19005 -5981
rect -18929 -5951 -18751 -5899
rect -18575 -5946 -18411 -5928
rect -18575 -5951 -18461 -5946
rect -18929 -5981 -18461 -5951
rect -18427 -5981 -18411 -5946
rect -20296 -6081 -19860 -6075
rect -19265 -6070 -19215 -6001
rect -18929 -6029 -18411 -5981
rect -19265 -6092 -19259 -6070
rect -20762 -6148 -20324 -6105
rect -20762 -6214 -20743 -6148
rect -20490 -6214 -20324 -6148
rect -20762 -6228 -20324 -6214
rect -19457 -6105 -19259 -6092
rect -19225 -6105 -19215 -6070
rect -19187 -6041 -18411 -6029
rect -19187 -6075 -19175 -6041
rect -18799 -6075 -18751 -6041
rect -18575 -6063 -18411 -6041
rect -18383 -5946 -18123 -5927
rect -18383 -5981 -18172 -5946
rect -18138 -5981 -18123 -5946
rect -18383 -6001 -18123 -5981
rect -18047 -5944 -17869 -5899
rect -19187 -6081 -18751 -6075
rect -18383 -6070 -18333 -6001
rect -18047 -6024 -18002 -5944
rect -17882 -6024 -17869 -5944
rect -18047 -6029 -17869 -6024
rect -18383 -6092 -18377 -6070
rect -19457 -6159 -19215 -6105
rect -19457 -6219 -19433 -6159
rect -19248 -6219 -19215 -6159
rect -24637 -6262 -24432 -6247
rect -20296 -6233 -19896 -6227
rect -19457 -6228 -19215 -6219
rect -18575 -6105 -18377 -6092
rect -18343 -6105 -18333 -6070
rect -18305 -6041 -17869 -6029
rect -18305 -6075 -18293 -6041
rect -17917 -6075 -17869 -6041
rect -17275 -5946 -17111 -5928
rect -17275 -5955 -17161 -5946
rect -17275 -6035 -17243 -5955
rect -17127 -5981 -17111 -5946
rect -17145 -6035 -17111 -5981
rect -17275 -6063 -17111 -6035
rect -17083 -5946 -16823 -5927
rect -17083 -5981 -16872 -5946
rect -16838 -5981 -16823 -5946
rect -17083 -6001 -16823 -5981
rect -18305 -6081 -17869 -6075
rect -17083 -6070 -17033 -6001
rect -16747 -6029 -16688 -5899
rect -17083 -6091 -17077 -6070
rect -18575 -6110 -18333 -6105
rect -18575 -6185 -18561 -6110
rect -18416 -6185 -18333 -6110
rect -20296 -6267 -20284 -6233
rect -19908 -6267 -19896 -6233
rect -20296 -6305 -19896 -6267
rect -20296 -6350 -20269 -6305
rect -20278 -6357 -20269 -6350
rect -19934 -6350 -19896 -6305
rect -19187 -6233 -18787 -6227
rect -18575 -6228 -18333 -6185
rect -17471 -6105 -17077 -6091
rect -17043 -6105 -17033 -6070
rect -17005 -6041 -16688 -6029
rect -17005 -6075 -16993 -6041
rect -16605 -6042 -16569 -5894
rect -16038 -5813 -15460 -5807
rect -16038 -5893 -16022 -5813
rect -15988 -5893 -15830 -5813
rect -15796 -5893 -15638 -5813
rect -15604 -5893 -15460 -5813
rect -16038 -5899 -15460 -5893
rect -15156 -5813 -14578 -5807
rect -15156 -5893 -15140 -5813
rect -15106 -5893 -14948 -5813
rect -14914 -5893 -14756 -5813
rect -14722 -5893 -14578 -5813
rect -15156 -5899 -14578 -5893
rect -13856 -5813 -13278 -5807
rect -13856 -5893 -13840 -5813
rect -13806 -5893 -13648 -5813
rect -13614 -5893 -13456 -5813
rect -13422 -5893 -13278 -5813
rect -13856 -5894 -13278 -5893
rect -13856 -5899 -13397 -5894
rect -16617 -6075 -16569 -6042
rect -16166 -5946 -16002 -5928
rect -16166 -5956 -16052 -5946
rect -16166 -6036 -16132 -5956
rect -16018 -5981 -16002 -5946
rect -16034 -6036 -16002 -5981
rect -16166 -6063 -16002 -6036
rect -15974 -5946 -15714 -5927
rect -15974 -5981 -15763 -5946
rect -15729 -5981 -15714 -5946
rect -15974 -6001 -15714 -5981
rect -15638 -5951 -15460 -5899
rect -15284 -5946 -15120 -5928
rect -15284 -5951 -15170 -5946
rect -15638 -5981 -15170 -5951
rect -15136 -5981 -15120 -5946
rect -17005 -6081 -16569 -6075
rect -15974 -6070 -15924 -6001
rect -15638 -6029 -15120 -5981
rect -15974 -6092 -15968 -6070
rect -17471 -6148 -17033 -6105
rect -17471 -6214 -17452 -6148
rect -17199 -6214 -17033 -6148
rect -19187 -6267 -19175 -6233
rect -18799 -6267 -18787 -6233
rect -19187 -6305 -18787 -6267
rect -19187 -6339 -19160 -6305
rect -18825 -6339 -18787 -6305
rect -19187 -6350 -19033 -6339
rect -19934 -6357 -19925 -6350
rect -20278 -6366 -19925 -6357
rect -19044 -6372 -19033 -6350
rect -18971 -6350 -18787 -6339
rect -18305 -6233 -17905 -6227
rect -17471 -6228 -17033 -6214
rect -16166 -6105 -15968 -6092
rect -15934 -6105 -15924 -6070
rect -15896 -6041 -15120 -6029
rect -15896 -6075 -15884 -6041
rect -15508 -6075 -15460 -6041
rect -15284 -6063 -15120 -6041
rect -15092 -5946 -14832 -5927
rect -15092 -5981 -14881 -5946
rect -14847 -5981 -14832 -5946
rect -15092 -6001 -14832 -5981
rect -14756 -5944 -14578 -5899
rect -15896 -6081 -15460 -6075
rect -15092 -6070 -15042 -6001
rect -14756 -6024 -14711 -5944
rect -14591 -6024 -14578 -5944
rect -14756 -6029 -14578 -6024
rect -15092 -6092 -15086 -6070
rect -16166 -6159 -15924 -6105
rect -16166 -6219 -16142 -6159
rect -15957 -6219 -15924 -6159
rect -18305 -6267 -18293 -6233
rect -17917 -6267 -17905 -6233
rect -18305 -6305 -17905 -6267
rect -18305 -6339 -18278 -6305
rect -17943 -6339 -17905 -6305
rect -18305 -6350 -18166 -6339
rect -18971 -6372 -18960 -6350
rect -19044 -6383 -18960 -6372
rect -18179 -6389 -18166 -6350
rect -18114 -6350 -17905 -6339
rect -17005 -6233 -16605 -6227
rect -16166 -6228 -15924 -6219
rect -15284 -6105 -15086 -6092
rect -15052 -6105 -15042 -6070
rect -15014 -6041 -14578 -6029
rect -15014 -6075 -15002 -6041
rect -14626 -6075 -14578 -6041
rect -13984 -5946 -13820 -5928
rect -13984 -5955 -13870 -5946
rect -13984 -6035 -13952 -5955
rect -13836 -5981 -13820 -5946
rect -13854 -6035 -13820 -5981
rect -13984 -6063 -13820 -6035
rect -13792 -5946 -13532 -5927
rect -13792 -5981 -13581 -5946
rect -13547 -5981 -13532 -5946
rect -13792 -6001 -13532 -5981
rect -15014 -6081 -14578 -6075
rect -13792 -6070 -13742 -6001
rect -13456 -6029 -13397 -5899
rect -13792 -6091 -13786 -6070
rect -15284 -6110 -15042 -6105
rect -15284 -6185 -15270 -6110
rect -15125 -6185 -15042 -6110
rect -17005 -6267 -16993 -6233
rect -16617 -6267 -16605 -6233
rect -17005 -6305 -16605 -6267
rect -17005 -6350 -16978 -6305
rect -18114 -6389 -18101 -6350
rect -16987 -6357 -16978 -6350
rect -16643 -6350 -16605 -6305
rect -15896 -6233 -15496 -6227
rect -15284 -6228 -15042 -6185
rect -14180 -6105 -13786 -6091
rect -13752 -6105 -13742 -6070
rect -13714 -6041 -13397 -6029
rect -13714 -6075 -13702 -6041
rect -13314 -6042 -13278 -5894
rect -12747 -5813 -12169 -5807
rect -12747 -5893 -12731 -5813
rect -12697 -5893 -12539 -5813
rect -12505 -5893 -12347 -5813
rect -12313 -5893 -12169 -5813
rect -12747 -5899 -12169 -5893
rect -11865 -5813 -11287 -5807
rect -11865 -5893 -11849 -5813
rect -11815 -5893 -11657 -5813
rect -11623 -5893 -11465 -5813
rect -11431 -5893 -11287 -5813
rect -11865 -5899 -11287 -5893
rect -10565 -5813 -9987 -5807
rect -10565 -5893 -10549 -5813
rect -10515 -5893 -10357 -5813
rect -10323 -5893 -10165 -5813
rect -10131 -5893 -9987 -5813
rect -10565 -5894 -9987 -5893
rect -10565 -5899 -10106 -5894
rect -13326 -6075 -13278 -6042
rect -12875 -5946 -12711 -5928
rect -12875 -5956 -12761 -5946
rect -12875 -6036 -12841 -5956
rect -12727 -5981 -12711 -5946
rect -12743 -6036 -12711 -5981
rect -12875 -6063 -12711 -6036
rect -12683 -5946 -12423 -5927
rect -12683 -5981 -12472 -5946
rect -12438 -5981 -12423 -5946
rect -12683 -6001 -12423 -5981
rect -12347 -5951 -12169 -5899
rect -11993 -5946 -11829 -5928
rect -11993 -5951 -11879 -5946
rect -12347 -5981 -11879 -5951
rect -11845 -5981 -11829 -5946
rect -13714 -6081 -13278 -6075
rect -12683 -6070 -12633 -6001
rect -12347 -6029 -11829 -5981
rect -12683 -6092 -12677 -6070
rect -14180 -6148 -13742 -6105
rect -14180 -6214 -14161 -6148
rect -13908 -6214 -13742 -6148
rect -15896 -6267 -15884 -6233
rect -15508 -6267 -15496 -6233
rect -15896 -6305 -15496 -6267
rect -15896 -6339 -15869 -6305
rect -15534 -6339 -15496 -6305
rect -15896 -6350 -15742 -6339
rect -16643 -6357 -16634 -6350
rect -16987 -6366 -16634 -6357
rect -15753 -6372 -15742 -6350
rect -15680 -6350 -15496 -6339
rect -15014 -6233 -14614 -6227
rect -14180 -6228 -13742 -6214
rect -12875 -6105 -12677 -6092
rect -12643 -6105 -12633 -6070
rect -12605 -6041 -11829 -6029
rect -12605 -6075 -12593 -6041
rect -12217 -6075 -12169 -6041
rect -11993 -6063 -11829 -6041
rect -11801 -5946 -11541 -5927
rect -11801 -5981 -11590 -5946
rect -11556 -5981 -11541 -5946
rect -11801 -6001 -11541 -5981
rect -11465 -5944 -11287 -5899
rect -12605 -6081 -12169 -6075
rect -11801 -6070 -11751 -6001
rect -11465 -6024 -11420 -5944
rect -11300 -6024 -11287 -5944
rect -11465 -6029 -11287 -6024
rect -11801 -6092 -11795 -6070
rect -12875 -6159 -12633 -6105
rect -12875 -6219 -12851 -6159
rect -12666 -6219 -12633 -6159
rect -15014 -6267 -15002 -6233
rect -14626 -6267 -14614 -6233
rect -15014 -6305 -14614 -6267
rect -15014 -6339 -14987 -6305
rect -14652 -6339 -14614 -6305
rect -15014 -6350 -14875 -6339
rect -15680 -6372 -15669 -6350
rect -15753 -6383 -15669 -6372
rect -18179 -6402 -18101 -6389
rect -14888 -6389 -14875 -6350
rect -14823 -6350 -14614 -6339
rect -13714 -6233 -13314 -6227
rect -12875 -6228 -12633 -6219
rect -11993 -6105 -11795 -6092
rect -11761 -6105 -11751 -6070
rect -11723 -6041 -11287 -6029
rect -11723 -6075 -11711 -6041
rect -11335 -6075 -11287 -6041
rect -10693 -5946 -10529 -5928
rect -10693 -5955 -10579 -5946
rect -10693 -6035 -10661 -5955
rect -10545 -5981 -10529 -5946
rect -10563 -6035 -10529 -5981
rect -10693 -6063 -10529 -6035
rect -10501 -5946 -10241 -5927
rect -10501 -5981 -10290 -5946
rect -10256 -5981 -10241 -5946
rect -10501 -6001 -10241 -5981
rect -11723 -6081 -11287 -6075
rect -10501 -6070 -10451 -6001
rect -10165 -6029 -10106 -5899
rect -10501 -6091 -10495 -6070
rect -11993 -6110 -11751 -6105
rect -11993 -6185 -11979 -6110
rect -11834 -6185 -11751 -6110
rect -13714 -6267 -13702 -6233
rect -13326 -6267 -13314 -6233
rect -13714 -6305 -13314 -6267
rect -13714 -6350 -13687 -6305
rect -14823 -6389 -14810 -6350
rect -13696 -6357 -13687 -6350
rect -13352 -6350 -13314 -6305
rect -12605 -6233 -12205 -6227
rect -11993 -6228 -11751 -6185
rect -10889 -6105 -10495 -6091
rect -10461 -6105 -10451 -6070
rect -10423 -6041 -10106 -6029
rect -10423 -6075 -10411 -6041
rect -10023 -6042 -9987 -5894
rect -9456 -5813 -8878 -5807
rect -9456 -5893 -9440 -5813
rect -9406 -5893 -9248 -5813
rect -9214 -5893 -9056 -5813
rect -9022 -5893 -8878 -5813
rect -9456 -5899 -8878 -5893
rect -8574 -5813 -7996 -5807
rect -8574 -5893 -8558 -5813
rect -8524 -5893 -8366 -5813
rect -8332 -5893 -8174 -5813
rect -8140 -5893 -7996 -5813
rect -8574 -5899 -7996 -5893
rect -10035 -6075 -9987 -6042
rect -9584 -5946 -9420 -5928
rect -9584 -5956 -9470 -5946
rect -9584 -6036 -9550 -5956
rect -9436 -5981 -9420 -5946
rect -9452 -6036 -9420 -5981
rect -9584 -6063 -9420 -6036
rect -9392 -5946 -9132 -5927
rect -9392 -5981 -9181 -5946
rect -9147 -5981 -9132 -5946
rect -9392 -6001 -9132 -5981
rect -9056 -5951 -8878 -5899
rect -8702 -5946 -8538 -5928
rect -8702 -5951 -8588 -5946
rect -9056 -5981 -8588 -5951
rect -8554 -5981 -8538 -5946
rect -10423 -6081 -9987 -6075
rect -9392 -6070 -9342 -6001
rect -9056 -6029 -8538 -5981
rect -9392 -6092 -9386 -6070
rect -10889 -6148 -10451 -6105
rect -10889 -6214 -10870 -6148
rect -10617 -6214 -10451 -6148
rect -12605 -6267 -12593 -6233
rect -12217 -6267 -12205 -6233
rect -12605 -6305 -12205 -6267
rect -12605 -6339 -12578 -6305
rect -12243 -6339 -12205 -6305
rect -12605 -6350 -12451 -6339
rect -13352 -6357 -13343 -6350
rect -13696 -6366 -13343 -6357
rect -12462 -6372 -12451 -6350
rect -12389 -6350 -12205 -6339
rect -11723 -6233 -11323 -6227
rect -10889 -6228 -10451 -6214
rect -9584 -6105 -9386 -6092
rect -9352 -6105 -9342 -6070
rect -9314 -6041 -8538 -6029
rect -9314 -6075 -9302 -6041
rect -8926 -6075 -8878 -6041
rect -8702 -6063 -8538 -6041
rect -8510 -5946 -8250 -5927
rect -8510 -5981 -8299 -5946
rect -8265 -5981 -8250 -5946
rect -8510 -6001 -8250 -5981
rect -8174 -5944 -7996 -5899
rect -9314 -6081 -8878 -6075
rect -8510 -6070 -8460 -6001
rect -8174 -6024 -8129 -5944
rect -8009 -6024 -7996 -5944
rect -8174 -6029 -7996 -6024
rect -8510 -6092 -8504 -6070
rect -9584 -6159 -9342 -6105
rect -9584 -6219 -9560 -6159
rect -9375 -6219 -9342 -6159
rect -11723 -6267 -11711 -6233
rect -11335 -6267 -11323 -6233
rect -11723 -6305 -11323 -6267
rect -11723 -6339 -11696 -6305
rect -11361 -6339 -11323 -6305
rect -11723 -6350 -11584 -6339
rect -12389 -6372 -12378 -6350
rect -12462 -6383 -12378 -6372
rect -14888 -6402 -14810 -6389
rect -11597 -6389 -11584 -6350
rect -11532 -6350 -11323 -6339
rect -10423 -6233 -10023 -6227
rect -9584 -6228 -9342 -6219
rect -8702 -6105 -8504 -6092
rect -8470 -6105 -8460 -6070
rect -8432 -6041 -7996 -6029
rect -8432 -6075 -8420 -6041
rect -8044 -6075 -7996 -6041
rect -8432 -6081 -7996 -6075
rect -8702 -6110 -8460 -6105
rect -8702 -6185 -8688 -6110
rect -8543 -6185 -8460 -6110
rect -10423 -6267 -10411 -6233
rect -10035 -6267 -10023 -6233
rect -10423 -6305 -10023 -6267
rect -10423 -6350 -10396 -6305
rect -11532 -6389 -11519 -6350
rect -10405 -6357 -10396 -6350
rect -10061 -6350 -10023 -6305
rect -9314 -6233 -8914 -6227
rect -8702 -6228 -8460 -6185
rect -9314 -6267 -9302 -6233
rect -8926 -6267 -8914 -6233
rect -9314 -6305 -8914 -6267
rect -9314 -6339 -9287 -6305
rect -8952 -6339 -8914 -6305
rect -9314 -6350 -9160 -6339
rect -10061 -6357 -10052 -6350
rect -10405 -6366 -10052 -6357
rect -9171 -6372 -9160 -6350
rect -9098 -6350 -8914 -6339
rect -8432 -6233 -8032 -6227
rect -8432 -6267 -8420 -6233
rect -8044 -6267 -8032 -6233
rect -8432 -6305 -8032 -6267
rect -7879 -6291 -7873 -6225
rect -7807 -6291 -7801 -6225
rect -8432 -6339 -8405 -6305
rect -8070 -6339 -8032 -6305
rect -8432 -6350 -8293 -6339
rect -9098 -6372 -9087 -6350
rect -9171 -6383 -9087 -6372
rect -11597 -6402 -11519 -6389
rect -8306 -6389 -8293 -6350
rect -8241 -6350 -8032 -6339
rect -8241 -6389 -8228 -6350
rect -8306 -6402 -8228 -6389
rect -7873 -6533 -7807 -6291
rect -5439 -6533 -5373 -6527
rect -23304 -6572 -23210 -6571
rect -23304 -6656 -11066 -6572
rect -7873 -6599 -5439 -6533
rect -5439 -6605 -5373 -6599
rect -23585 -7302 -23370 -7280
rect -24397 -7377 -23763 -7370
rect -24397 -7424 -24368 -7377
rect -23799 -7424 -23763 -7377
rect -23585 -7381 -23562 -7302
rect -23393 -7381 -23370 -7302
rect -23585 -7396 -23370 -7381
rect -23585 -7400 -23578 -7396
rect -24397 -7496 -24359 -7424
rect -23805 -7490 -23763 -7424
rect -23684 -7444 -23615 -7428
rect -23805 -7496 -23762 -7490
rect -24397 -7576 -24384 -7496
rect -24350 -7576 -24192 -7544
rect -24158 -7576 -24000 -7544
rect -23966 -7576 -23808 -7544
rect -23774 -7576 -23762 -7496
rect -24397 -7582 -23762 -7576
rect -24397 -7583 -23763 -7582
rect -23684 -7612 -23665 -7444
rect -24304 -7618 -23665 -7612
rect -24304 -7698 -24288 -7618
rect -24254 -7698 -24096 -7618
rect -24062 -7698 -23904 -7618
rect -23870 -7670 -23665 -7618
rect -23631 -7670 -23615 -7444
rect -23584 -7430 -23578 -7400
rect -23499 -7400 -23370 -7396
rect -23499 -7430 -23493 -7400
rect -23304 -7428 -23210 -6656
rect -23584 -7588 -23493 -7430
rect -23584 -7622 -23578 -7588
rect -23499 -7622 -23493 -7588
rect -23584 -7638 -23493 -7622
rect -23461 -7492 -23210 -7428
rect -23461 -7526 -23455 -7492
rect -23378 -7526 -23210 -7492
rect -23870 -7698 -23615 -7670
rect -23461 -7684 -23210 -7526
rect -24304 -7704 -23615 -7698
rect -24862 -7751 -24268 -7733
rect -24862 -7786 -24318 -7751
rect -24284 -7786 -24268 -7751
rect -24862 -7868 -24268 -7786
rect -24240 -7751 -23980 -7732
rect -24240 -7786 -24029 -7751
rect -23995 -7786 -23980 -7751
rect -24240 -7806 -23980 -7786
rect -24862 -10970 -24696 -7868
rect -24240 -7875 -24190 -7806
rect -23904 -7834 -23615 -7704
rect -24240 -7897 -24234 -7875
rect -24632 -7910 -24234 -7897
rect -24200 -7910 -24190 -7875
rect -24162 -7846 -23615 -7834
rect -24162 -7880 -24150 -7846
rect -23774 -7880 -23615 -7846
rect -24162 -7886 -23615 -7880
rect -23584 -7718 -23455 -7684
rect -23378 -7718 -23210 -7684
rect -23584 -7846 -23210 -7718
rect -23584 -7880 -23572 -7846
rect -23396 -7880 -23210 -7846
rect -23088 -6803 -14356 -6719
rect -23584 -7886 -23384 -7880
rect -24632 -7911 -24190 -7910
rect -24632 -8015 -24611 -7911
rect -24368 -8015 -24190 -7911
rect -23684 -7890 -23615 -7886
rect -23684 -7924 -23665 -7890
rect -23631 -7924 -23615 -7890
rect -23684 -7941 -23615 -7924
rect -23585 -7934 -23384 -7927
rect -24632 -8033 -24190 -8015
rect -23585 -7968 -23572 -7934
rect -23396 -7968 -23384 -7934
rect -23356 -7941 -23272 -7880
rect -24162 -8038 -23762 -8032
rect -24162 -8072 -24150 -8038
rect -23774 -8072 -23762 -8038
rect -24162 -8110 -24133 -8072
rect -24162 -8144 -24135 -8110
rect -23793 -8134 -23762 -8072
rect -23585 -8051 -23558 -7968
rect -23409 -8051 -23384 -7968
rect -23585 -8070 -23553 -8051
rect -23421 -8070 -23384 -8051
rect -23585 -8077 -23384 -8070
rect -23800 -8144 -23762 -8134
rect -24162 -8155 -23762 -8144
rect -23583 -8594 -23369 -8572
rect -24397 -8669 -23763 -8662
rect -24397 -8716 -24368 -8669
rect -23799 -8716 -23763 -8669
rect -24397 -8788 -24359 -8716
rect -23805 -8782 -23763 -8716
rect -23583 -8673 -23560 -8594
rect -23391 -8673 -23369 -8594
rect -23583 -8688 -23369 -8673
rect -23683 -8736 -23614 -8720
rect -23805 -8788 -23762 -8782
rect -24397 -8868 -24384 -8788
rect -24350 -8868 -24192 -8836
rect -24158 -8868 -24000 -8836
rect -23966 -8868 -23808 -8836
rect -23774 -8868 -23762 -8788
rect -24397 -8874 -23762 -8868
rect -24397 -8875 -23763 -8874
rect -23683 -8904 -23664 -8736
rect -24304 -8910 -23664 -8904
rect -24304 -8990 -24288 -8910
rect -24254 -8990 -24096 -8910
rect -24062 -8990 -23904 -8910
rect -23870 -8962 -23664 -8910
rect -23630 -8962 -23614 -8736
rect -23583 -8722 -23577 -8688
rect -23498 -8692 -23369 -8688
rect -23498 -8722 -23492 -8692
rect -23583 -8880 -23492 -8722
rect -23583 -8914 -23577 -8880
rect -23498 -8914 -23492 -8880
rect -23583 -8930 -23492 -8914
rect -23460 -8784 -23271 -8720
rect -23460 -8818 -23454 -8784
rect -23377 -8818 -23271 -8784
rect -23460 -8905 -23271 -8818
rect -23088 -8905 -22951 -6803
rect -21259 -6951 -17647 -6867
rect -21850 -7302 -21636 -7280
rect -22660 -7377 -22026 -7370
rect -22660 -7424 -22631 -7377
rect -22062 -7424 -22026 -7377
rect -22660 -7496 -22622 -7424
rect -22068 -7490 -22026 -7424
rect -21850 -7381 -21827 -7302
rect -21658 -7381 -21636 -7302
rect -21850 -7396 -21636 -7381
rect -21950 -7444 -21881 -7428
rect -22068 -7496 -22025 -7490
rect -22660 -7576 -22647 -7496
rect -22613 -7576 -22455 -7544
rect -22421 -7576 -22263 -7544
rect -22229 -7576 -22071 -7544
rect -22037 -7576 -22025 -7496
rect -22660 -7582 -22025 -7576
rect -22660 -7583 -22026 -7582
rect -21950 -7612 -21931 -7444
rect -22567 -7618 -21931 -7612
rect -22567 -7698 -22551 -7618
rect -22517 -7698 -22359 -7618
rect -22325 -7698 -22167 -7618
rect -22133 -7670 -21931 -7618
rect -21897 -7670 -21881 -7444
rect -21850 -7430 -21844 -7396
rect -21765 -7400 -21636 -7396
rect -21765 -7430 -21759 -7400
rect -21850 -7588 -21759 -7430
rect -21850 -7622 -21844 -7588
rect -21765 -7622 -21759 -7588
rect -21850 -7638 -21759 -7622
rect -21727 -7492 -21538 -7428
rect -21727 -7526 -21721 -7492
rect -21644 -7526 -21538 -7492
rect -22133 -7698 -21881 -7670
rect -21727 -7684 -21538 -7526
rect -22567 -7704 -21881 -7698
rect -22842 -7749 -22531 -7733
rect -22842 -7856 -22808 -7749
rect -22688 -7751 -22531 -7749
rect -22688 -7786 -22581 -7751
rect -22547 -7786 -22531 -7751
rect -22688 -7856 -22531 -7786
rect -22842 -7868 -22531 -7856
rect -22503 -7751 -22243 -7732
rect -22503 -7786 -22292 -7751
rect -22258 -7786 -22243 -7751
rect -22503 -7806 -22243 -7786
rect -22503 -7875 -22453 -7806
rect -22167 -7834 -21881 -7704
rect -22503 -7897 -22497 -7875
rect -22910 -7907 -22497 -7897
rect -22910 -8015 -22857 -7907
rect -22628 -7910 -22497 -7907
rect -22463 -7910 -22453 -7875
rect -22425 -7846 -21881 -7834
rect -22425 -7880 -22413 -7846
rect -22037 -7880 -21881 -7846
rect -22425 -7886 -21881 -7880
rect -21850 -7718 -21721 -7684
rect -21644 -7718 -21538 -7684
rect -21850 -7794 -21538 -7718
rect -21259 -7794 -21128 -6951
rect -17756 -7028 -17647 -6951
rect -20649 -7092 -19439 -7064
rect -20649 -7164 -20603 -7092
rect -19481 -7164 -19439 -7092
rect -20649 -7198 -19439 -7164
rect -20649 -7267 -20395 -7198
rect -20649 -7369 -20637 -7267
rect -20603 -7369 -20445 -7267
rect -20411 -7369 -20395 -7267
rect -20649 -7390 -20395 -7369
rect -20269 -7269 -19819 -7243
rect -20269 -7371 -20253 -7269
rect -20219 -7270 -19819 -7269
rect -20219 -7371 -20061 -7270
rect -20269 -7372 -20061 -7371
rect -20027 -7372 -19869 -7270
rect -19835 -7372 -19819 -7270
rect -20269 -7390 -19819 -7372
rect -19693 -7270 -19439 -7198
rect -19693 -7372 -19677 -7270
rect -19643 -7372 -19485 -7270
rect -19451 -7372 -19439 -7270
rect -19693 -7390 -19439 -7372
rect -19090 -7092 -17880 -7064
rect -19090 -7164 -19044 -7092
rect -17922 -7164 -17880 -7092
rect -17756 -7123 -17744 -7028
rect -17655 -7123 -17647 -7028
rect -14466 -7027 -14356 -6803
rect -17756 -7134 -17647 -7123
rect -17358 -7092 -16148 -7064
rect -19090 -7198 -17880 -7164
rect -19090 -7267 -18836 -7198
rect -19090 -7369 -19078 -7267
rect -19044 -7369 -18886 -7267
rect -18852 -7369 -18836 -7267
rect -19090 -7390 -18836 -7369
rect -18710 -7269 -18260 -7243
rect -18710 -7371 -18694 -7269
rect -18660 -7270 -18260 -7269
rect -18660 -7371 -18502 -7270
rect -18710 -7372 -18502 -7371
rect -18468 -7372 -18310 -7270
rect -18276 -7372 -18260 -7270
rect -18710 -7390 -18260 -7372
rect -18134 -7270 -17880 -7198
rect -18134 -7372 -18118 -7270
rect -18084 -7372 -17926 -7270
rect -17892 -7372 -17880 -7270
rect -18134 -7390 -17880 -7372
rect -17358 -7164 -17312 -7092
rect -16190 -7164 -16148 -7092
rect -17358 -7198 -16148 -7164
rect -17358 -7267 -17104 -7198
rect -17358 -7369 -17346 -7267
rect -17312 -7369 -17154 -7267
rect -17120 -7369 -17104 -7267
rect -17358 -7390 -17104 -7369
rect -16978 -7269 -16528 -7243
rect -16978 -7371 -16962 -7269
rect -16928 -7270 -16528 -7269
rect -16928 -7371 -16770 -7270
rect -16978 -7372 -16770 -7371
rect -16736 -7372 -16578 -7270
rect -16544 -7372 -16528 -7270
rect -16978 -7390 -16528 -7372
rect -16402 -7270 -16148 -7198
rect -16402 -7372 -16386 -7270
rect -16352 -7372 -16194 -7270
rect -16160 -7372 -16148 -7270
rect -16402 -7390 -16148 -7372
rect -15799 -7092 -14589 -7064
rect -15799 -7164 -15753 -7092
rect -14631 -7164 -14589 -7092
rect -15799 -7198 -14589 -7164
rect -15799 -7267 -15545 -7198
rect -15799 -7369 -15787 -7267
rect -15753 -7369 -15595 -7267
rect -15561 -7369 -15545 -7267
rect -15799 -7390 -15545 -7369
rect -15419 -7269 -14969 -7243
rect -15419 -7371 -15403 -7269
rect -15369 -7270 -14969 -7269
rect -15369 -7371 -15211 -7270
rect -15419 -7372 -15211 -7371
rect -15177 -7372 -15019 -7270
rect -14985 -7372 -14969 -7270
rect -15419 -7390 -14969 -7372
rect -14843 -7270 -14589 -7198
rect -14466 -7211 -14460 -7027
rect -14361 -7211 -14356 -7027
rect -11174 -7026 -11066 -6656
rect -14466 -7218 -14356 -7211
rect -14067 -7092 -12857 -7064
rect -14067 -7164 -14021 -7092
rect -12899 -7164 -12857 -7092
rect -14067 -7198 -12857 -7164
rect -14843 -7372 -14827 -7270
rect -14793 -7372 -14635 -7270
rect -14601 -7372 -14589 -7270
rect -14843 -7390 -14589 -7372
rect -14067 -7267 -13813 -7198
rect -14067 -7369 -14055 -7267
rect -14021 -7369 -13863 -7267
rect -13829 -7369 -13813 -7267
rect -14067 -7390 -13813 -7369
rect -13687 -7269 -13237 -7243
rect -13687 -7371 -13671 -7269
rect -13637 -7270 -13237 -7269
rect -13637 -7371 -13479 -7270
rect -13687 -7372 -13479 -7371
rect -13445 -7372 -13287 -7270
rect -13253 -7372 -13237 -7270
rect -13687 -7390 -13237 -7372
rect -13111 -7270 -12857 -7198
rect -13111 -7372 -13095 -7270
rect -13061 -7372 -12903 -7270
rect -12869 -7372 -12857 -7270
rect -13111 -7390 -12857 -7372
rect -12508 -7092 -11298 -7064
rect -12508 -7164 -12462 -7092
rect -11340 -7164 -11298 -7092
rect -12508 -7198 -11298 -7164
rect -11174 -7170 -11165 -7026
rect -11074 -7170 -11066 -7026
rect -11174 -7181 -11066 -7170
rect -10776 -7092 -9566 -7064
rect -10776 -7164 -10730 -7092
rect -9608 -7164 -9566 -7092
rect -12508 -7267 -12254 -7198
rect -12508 -7369 -12496 -7267
rect -12462 -7369 -12304 -7267
rect -12270 -7369 -12254 -7267
rect -12508 -7390 -12254 -7369
rect -12128 -7269 -11678 -7243
rect -12128 -7371 -12112 -7269
rect -12078 -7270 -11678 -7269
rect -12078 -7371 -11920 -7270
rect -12128 -7372 -11920 -7371
rect -11886 -7372 -11728 -7270
rect -11694 -7372 -11678 -7270
rect -12128 -7390 -11678 -7372
rect -11552 -7270 -11298 -7198
rect -11552 -7372 -11536 -7270
rect -11502 -7372 -11344 -7270
rect -11310 -7372 -11298 -7270
rect -11552 -7390 -11298 -7372
rect -10776 -7198 -9566 -7164
rect -10776 -7267 -10522 -7198
rect -10776 -7369 -10764 -7267
rect -10730 -7369 -10572 -7267
rect -10538 -7369 -10522 -7267
rect -10776 -7390 -10522 -7369
rect -10396 -7269 -9946 -7243
rect -10396 -7371 -10380 -7269
rect -10346 -7270 -9946 -7269
rect -10346 -7371 -10188 -7270
rect -10396 -7372 -10188 -7371
rect -10154 -7372 -9996 -7270
rect -9962 -7372 -9946 -7270
rect -10396 -7390 -9946 -7372
rect -9820 -7270 -9566 -7198
rect -9820 -7372 -9804 -7270
rect -9770 -7372 -9612 -7270
rect -9578 -7372 -9566 -7270
rect -9820 -7390 -9566 -7372
rect -9217 -7092 -8007 -7064
rect -9217 -7164 -9171 -7092
rect -8049 -7164 -8007 -7092
rect -9217 -7198 -8007 -7164
rect -9217 -7267 -8963 -7198
rect -9217 -7369 -9205 -7267
rect -9171 -7369 -9013 -7267
rect -8979 -7369 -8963 -7267
rect -9217 -7390 -8963 -7369
rect -8837 -7269 -8387 -7243
rect -8837 -7371 -8821 -7269
rect -8787 -7270 -8387 -7269
rect -8787 -7371 -8629 -7270
rect -8837 -7372 -8629 -7371
rect -8595 -7372 -8437 -7270
rect -8403 -7372 -8387 -7270
rect -8837 -7390 -8387 -7372
rect -8261 -7270 -8007 -7198
rect -8261 -7372 -8245 -7270
rect -8211 -7372 -8053 -7270
rect -8019 -7372 -8007 -7270
rect -8261 -7390 -8007 -7372
rect -20557 -7453 -19531 -7428
rect -20557 -7577 -20541 -7453
rect -20507 -7577 -20349 -7453
rect -20315 -7577 -20157 -7453
rect -20123 -7577 -19965 -7453
rect -19931 -7577 -19773 -7453
rect -19739 -7454 -19531 -7453
rect -19739 -7577 -19581 -7454
rect -20557 -7578 -19581 -7577
rect -19547 -7578 -19531 -7454
rect -20557 -7607 -19531 -7578
rect -18998 -7453 -17972 -7428
rect -18998 -7577 -18982 -7453
rect -18948 -7577 -18790 -7453
rect -18756 -7577 -18598 -7453
rect -18564 -7577 -18406 -7453
rect -18372 -7577 -18214 -7453
rect -18180 -7454 -17972 -7453
rect -18180 -7577 -18022 -7454
rect -18998 -7578 -18022 -7577
rect -17988 -7578 -17972 -7454
rect -18998 -7607 -17972 -7578
rect -17266 -7453 -16240 -7428
rect -17266 -7577 -17250 -7453
rect -17216 -7577 -17058 -7453
rect -17024 -7577 -16866 -7453
rect -16832 -7577 -16674 -7453
rect -16640 -7577 -16482 -7453
rect -16448 -7454 -16240 -7453
rect -16448 -7577 -16290 -7454
rect -17266 -7578 -16290 -7577
rect -16256 -7578 -16240 -7454
rect -17266 -7607 -16240 -7578
rect -15707 -7453 -14681 -7428
rect -15707 -7577 -15691 -7453
rect -15657 -7577 -15499 -7453
rect -15465 -7577 -15307 -7453
rect -15273 -7577 -15115 -7453
rect -15081 -7577 -14923 -7453
rect -14889 -7454 -14681 -7453
rect -14889 -7577 -14731 -7454
rect -15707 -7578 -14731 -7577
rect -14697 -7578 -14681 -7454
rect -15707 -7607 -14681 -7578
rect -13975 -7453 -12949 -7428
rect -13975 -7577 -13959 -7453
rect -13925 -7577 -13767 -7453
rect -13733 -7577 -13575 -7453
rect -13541 -7577 -13383 -7453
rect -13349 -7577 -13191 -7453
rect -13157 -7454 -12949 -7453
rect -13157 -7577 -12999 -7454
rect -13975 -7578 -12999 -7577
rect -12965 -7578 -12949 -7454
rect -13975 -7607 -12949 -7578
rect -12416 -7453 -11390 -7428
rect -12416 -7577 -12400 -7453
rect -12366 -7577 -12208 -7453
rect -12174 -7577 -12016 -7453
rect -11982 -7577 -11824 -7453
rect -11790 -7577 -11632 -7453
rect -11598 -7454 -11390 -7453
rect -11598 -7577 -11440 -7454
rect -12416 -7578 -11440 -7577
rect -11406 -7578 -11390 -7454
rect -12416 -7607 -11390 -7578
rect -10684 -7453 -9658 -7428
rect -10684 -7577 -10668 -7453
rect -10634 -7577 -10476 -7453
rect -10442 -7577 -10284 -7453
rect -10250 -7577 -10092 -7453
rect -10058 -7577 -9900 -7453
rect -9866 -7454 -9658 -7453
rect -9866 -7577 -9708 -7454
rect -10684 -7578 -9708 -7577
rect -9674 -7578 -9658 -7454
rect -10684 -7607 -9658 -7578
rect -9125 -7453 -8099 -7428
rect -9125 -7577 -9109 -7453
rect -9075 -7577 -8917 -7453
rect -8883 -7577 -8725 -7453
rect -8691 -7577 -8533 -7453
rect -8499 -7577 -8341 -7453
rect -8307 -7454 -8099 -7453
rect -8307 -7577 -8149 -7454
rect -9125 -7578 -8149 -7577
rect -8115 -7578 -8099 -7454
rect -9125 -7607 -8099 -7578
rect -20649 -7662 -20395 -7640
rect -20649 -7764 -20637 -7662
rect -20603 -7728 -20445 -7662
rect -20411 -7728 -20395 -7662
rect -20603 -7764 -20395 -7728
rect -20269 -7668 -19819 -7651
rect -20269 -7728 -20253 -7668
rect -20219 -7685 -19869 -7668
rect -20219 -7728 -20061 -7685
rect -20027 -7728 -19869 -7685
rect -19835 -7728 -19819 -7668
rect -20269 -7743 -19819 -7728
rect -19693 -7661 -19439 -7640
rect -19693 -7728 -19677 -7661
rect -19643 -7728 -19485 -7661
rect -19451 -7728 -19439 -7661
rect -20649 -7787 -20395 -7764
rect -19693 -7787 -19439 -7728
rect -19090 -7662 -18836 -7640
rect -19090 -7764 -19078 -7662
rect -19044 -7728 -18886 -7662
rect -18852 -7728 -18836 -7662
rect -19044 -7764 -18836 -7728
rect -18710 -7668 -18260 -7651
rect -18710 -7728 -18694 -7668
rect -18660 -7685 -18310 -7668
rect -18660 -7728 -18502 -7685
rect -18468 -7728 -18310 -7685
rect -18276 -7728 -18260 -7668
rect -18710 -7743 -18260 -7728
rect -18134 -7661 -17880 -7640
rect -18134 -7728 -18118 -7661
rect -18084 -7728 -17926 -7661
rect -17892 -7728 -17880 -7661
rect -19090 -7787 -18836 -7764
rect -18134 -7787 -17880 -7728
rect -17358 -7662 -17104 -7640
rect -17358 -7764 -17346 -7662
rect -17312 -7728 -17154 -7662
rect -17120 -7728 -17104 -7662
rect -17312 -7764 -17104 -7728
rect -16978 -7668 -16528 -7651
rect -16978 -7728 -16962 -7668
rect -16928 -7685 -16578 -7668
rect -16928 -7728 -16770 -7685
rect -16736 -7728 -16578 -7685
rect -16544 -7728 -16528 -7668
rect -16978 -7743 -16528 -7728
rect -16402 -7661 -16148 -7640
rect -16402 -7728 -16386 -7661
rect -16352 -7728 -16194 -7661
rect -16160 -7728 -16148 -7661
rect -17358 -7787 -17104 -7764
rect -16402 -7787 -16148 -7728
rect -15799 -7662 -15545 -7640
rect -15799 -7764 -15787 -7662
rect -15753 -7728 -15595 -7662
rect -15561 -7728 -15545 -7662
rect -15753 -7764 -15545 -7728
rect -15419 -7668 -14969 -7651
rect -15419 -7728 -15403 -7668
rect -15369 -7685 -15019 -7668
rect -15369 -7728 -15211 -7685
rect -15177 -7728 -15019 -7685
rect -14985 -7728 -14969 -7668
rect -15419 -7743 -14969 -7728
rect -14843 -7661 -14589 -7640
rect -14843 -7728 -14827 -7661
rect -14793 -7728 -14635 -7661
rect -14601 -7728 -14589 -7661
rect -15799 -7787 -15545 -7764
rect -14843 -7787 -14589 -7728
rect -14067 -7662 -13813 -7640
rect -14067 -7764 -14055 -7662
rect -14021 -7728 -13863 -7662
rect -13829 -7728 -13813 -7662
rect -14021 -7764 -13813 -7728
rect -13687 -7668 -13237 -7651
rect -13687 -7728 -13671 -7668
rect -13637 -7685 -13287 -7668
rect -13637 -7728 -13479 -7685
rect -13445 -7728 -13287 -7685
rect -13253 -7728 -13237 -7668
rect -13687 -7743 -13237 -7728
rect -13111 -7661 -12857 -7640
rect -13111 -7728 -13095 -7661
rect -13061 -7728 -12903 -7661
rect -12869 -7728 -12857 -7661
rect -14067 -7787 -13813 -7764
rect -13111 -7787 -12857 -7728
rect -12508 -7662 -12254 -7640
rect -12508 -7764 -12496 -7662
rect -12462 -7728 -12304 -7662
rect -12270 -7728 -12254 -7662
rect -12462 -7764 -12254 -7728
rect -12128 -7668 -11678 -7651
rect -12128 -7728 -12112 -7668
rect -12078 -7685 -11728 -7668
rect -12078 -7728 -11920 -7685
rect -11886 -7728 -11728 -7685
rect -11694 -7728 -11678 -7668
rect -12128 -7743 -11678 -7728
rect -11552 -7661 -11298 -7640
rect -11552 -7728 -11536 -7661
rect -11502 -7728 -11344 -7661
rect -11310 -7728 -11298 -7661
rect -12508 -7787 -12254 -7764
rect -11552 -7787 -11298 -7728
rect -10776 -7662 -10522 -7640
rect -10776 -7764 -10764 -7662
rect -10730 -7728 -10572 -7662
rect -10538 -7728 -10522 -7662
rect -10730 -7764 -10522 -7728
rect -10396 -7668 -9946 -7651
rect -10396 -7728 -10380 -7668
rect -10346 -7685 -9996 -7668
rect -10346 -7728 -10188 -7685
rect -10154 -7728 -9996 -7685
rect -9962 -7728 -9946 -7668
rect -10396 -7743 -9946 -7728
rect -9820 -7661 -9566 -7640
rect -9820 -7728 -9804 -7661
rect -9770 -7728 -9612 -7661
rect -9578 -7728 -9566 -7661
rect -10776 -7787 -10522 -7764
rect -9820 -7787 -9566 -7728
rect -9217 -7662 -8963 -7640
rect -9217 -7764 -9205 -7662
rect -9171 -7728 -9013 -7662
rect -8979 -7728 -8963 -7662
rect -9171 -7764 -8963 -7728
rect -8837 -7668 -8387 -7651
rect -8837 -7728 -8821 -7668
rect -8787 -7685 -8437 -7668
rect -8787 -7728 -8629 -7685
rect -8595 -7728 -8437 -7685
rect -8403 -7728 -8387 -7668
rect -8837 -7743 -8387 -7728
rect -8261 -7661 -8007 -7640
rect -8261 -7728 -8245 -7661
rect -8211 -7728 -8053 -7661
rect -8019 -7728 -8007 -7661
rect -9217 -7787 -8963 -7764
rect -8261 -7787 -8007 -7728
rect -21850 -7846 -21128 -7794
rect -21850 -7880 -21838 -7846
rect -21662 -7880 -21128 -7846
rect -21850 -7886 -21650 -7880
rect -22628 -8015 -22453 -7910
rect -21950 -7890 -21881 -7886
rect -21950 -7924 -21931 -7890
rect -21897 -7924 -21881 -7890
rect -21950 -7941 -21881 -7924
rect -21850 -7934 -21650 -7927
rect -22910 -8033 -22453 -8015
rect -21850 -7968 -21838 -7934
rect -21662 -7968 -21650 -7934
rect -21622 -7941 -21128 -7880
rect -20872 -7887 -20737 -7863
rect -22910 -8038 -22614 -8033
rect -22425 -8038 -22025 -8032
rect -22425 -8072 -22413 -8038
rect -22037 -8072 -22025 -8038
rect -22425 -8110 -22396 -8072
rect -22425 -8144 -22398 -8110
rect -22056 -8134 -22025 -8072
rect -21850 -8051 -21823 -7968
rect -21674 -8051 -21650 -7968
rect -20872 -7997 -20854 -7887
rect -20758 -7995 -20737 -7887
rect -17581 -7887 -17446 -7863
rect -19398 -7922 -19207 -7917
rect -19399 -7932 -19207 -7922
rect -19399 -7939 -19297 -7932
rect -19224 -7939 -19207 -7932
rect -20807 -7997 -20737 -7995
rect -20872 -8017 -20737 -7997
rect -20576 -7980 -19787 -7962
rect -20576 -7988 -19933 -7980
rect -21850 -8070 -21819 -8051
rect -21687 -8070 -21650 -8051
rect -20576 -8041 -20539 -7988
rect -20406 -8033 -19933 -7988
rect -19819 -8033 -19787 -7980
rect -20406 -8041 -19787 -8033
rect -20576 -8061 -19787 -8041
rect -19717 -7981 -19602 -7962
rect -19717 -8049 -19699 -7981
rect -19619 -8049 -19602 -7981
rect -19399 -8022 -19372 -7939
rect -21850 -8077 -21650 -8070
rect -22063 -8144 -22025 -8134
rect -22425 -8155 -22025 -8144
rect -20795 -8120 -20590 -8101
rect -20795 -8228 -20751 -8120
rect -20675 -8146 -20590 -8120
rect -19717 -8146 -19602 -8049
rect -19486 -8036 -19372 -8022
rect -19222 -8036 -19207 -7939
rect -19486 -8052 -19207 -8036
rect -19017 -7980 -18228 -7962
rect -19017 -7988 -18374 -7980
rect -19017 -8041 -18980 -7988
rect -18847 -8033 -18374 -7988
rect -18260 -8033 -18228 -7980
rect -18847 -8041 -18228 -8033
rect -19486 -8115 -19315 -8052
rect -19017 -8061 -18228 -8041
rect -18158 -7981 -18043 -7962
rect -18158 -8049 -18140 -7981
rect -18060 -8049 -18043 -7981
rect -17581 -7997 -17563 -7887
rect -17467 -7995 -17446 -7887
rect -14290 -7887 -14155 -7863
rect -16107 -7922 -15916 -7917
rect -16108 -7932 -15916 -7922
rect -16108 -7939 -16006 -7932
rect -15933 -7939 -15916 -7932
rect -17516 -7997 -17446 -7995
rect -17581 -8017 -17446 -7997
rect -17285 -7980 -16496 -7962
rect -17285 -7988 -16642 -7980
rect -20675 -8228 -19602 -8146
rect -20795 -8232 -19602 -8228
rect -19528 -8152 -19315 -8115
rect -19528 -8207 -19517 -8152
rect -19452 -8207 -19315 -8152
rect -19528 -8231 -19315 -8207
rect -19236 -8127 -19031 -8101
rect -19236 -8224 -19196 -8127
rect -19080 -8146 -19031 -8127
rect -18158 -8146 -18043 -8049
rect -17927 -8115 -17647 -8022
rect -17285 -8041 -17248 -7988
rect -17115 -8033 -16642 -7988
rect -16528 -8033 -16496 -7980
rect -17115 -8041 -16496 -8033
rect -17285 -8061 -16496 -8041
rect -16426 -7981 -16311 -7962
rect -16426 -8049 -16408 -7981
rect -16328 -8049 -16311 -7981
rect -16108 -8022 -16081 -7939
rect -19080 -8224 -18043 -8146
rect -19236 -8232 -18043 -8224
rect -17969 -8152 -17647 -8115
rect -17969 -8207 -17958 -8152
rect -17893 -8207 -17647 -8152
rect -17969 -8231 -17647 -8207
rect -20795 -8244 -20590 -8232
rect -19236 -8244 -19031 -8232
rect -20644 -8301 -20589 -8285
rect -20644 -8407 -20637 -8301
rect -20603 -8407 -20589 -8301
rect -20557 -8286 -20107 -8274
rect -20557 -8320 -20541 -8286
rect -20507 -8320 -20349 -8286
rect -20315 -8287 -20107 -8286
rect -20315 -8320 -20157 -8287
rect -20557 -8321 -20157 -8320
rect -20123 -8321 -20107 -8287
rect -20557 -8342 -20107 -8321
rect -19981 -8286 -19531 -8274
rect -19981 -8320 -19965 -8286
rect -19931 -8320 -19773 -8286
rect -19739 -8320 -19581 -8286
rect -19547 -8320 -19531 -8286
rect -19981 -8342 -19531 -8320
rect -19497 -8301 -19442 -8285
rect -20644 -8473 -20589 -8407
rect -20459 -8387 -20394 -8370
rect -20459 -8421 -20445 -8387
rect -20411 -8421 -20394 -8387
rect -20459 -8473 -20394 -8421
rect -20266 -8387 -19819 -8375
rect -20266 -8421 -20253 -8387
rect -20219 -8421 -20061 -8387
rect -20027 -8421 -19869 -8387
rect -19835 -8421 -19819 -8387
rect -20266 -8439 -19819 -8421
rect -19693 -8387 -19628 -8371
rect -19693 -8421 -19677 -8387
rect -19643 -8421 -19628 -8387
rect -19693 -8473 -19628 -8421
rect -19497 -8407 -19485 -8301
rect -19451 -8407 -19442 -8301
rect -19497 -8473 -19442 -8407
rect -20644 -8484 -19442 -8473
rect -20644 -8495 -20143 -8484
rect -20083 -8495 -19442 -8484
rect -20644 -8541 -20603 -8495
rect -19480 -8541 -19442 -8495
rect -20644 -8544 -20143 -8541
rect -20083 -8544 -19442 -8541
rect -20644 -8564 -19442 -8544
rect -19085 -8301 -19030 -8285
rect -19085 -8407 -19078 -8301
rect -19044 -8407 -19030 -8301
rect -18998 -8286 -18548 -8274
rect -18998 -8320 -18982 -8286
rect -18948 -8320 -18790 -8286
rect -18756 -8287 -18548 -8286
rect -18756 -8320 -18598 -8287
rect -18998 -8321 -18598 -8320
rect -18564 -8321 -18548 -8287
rect -18998 -8342 -18548 -8321
rect -18422 -8286 -17972 -8274
rect -18422 -8320 -18406 -8286
rect -18372 -8320 -18214 -8286
rect -18180 -8320 -18022 -8286
rect -17988 -8320 -17972 -8286
rect -18422 -8342 -17972 -8320
rect -17938 -8301 -17883 -8285
rect -19085 -8473 -19030 -8407
rect -18900 -8387 -18835 -8370
rect -18900 -8421 -18886 -8387
rect -18852 -8421 -18835 -8387
rect -18900 -8473 -18835 -8421
rect -18707 -8387 -18260 -8375
rect -18707 -8421 -18694 -8387
rect -18660 -8421 -18502 -8387
rect -18468 -8421 -18310 -8387
rect -18276 -8421 -18260 -8387
rect -18707 -8439 -18260 -8421
rect -18134 -8387 -18069 -8371
rect -18134 -8421 -18118 -8387
rect -18084 -8421 -18069 -8387
rect -18134 -8473 -18069 -8421
rect -17938 -8407 -17926 -8301
rect -17892 -8407 -17883 -8301
rect -17938 -8473 -17883 -8407
rect -19085 -8484 -17883 -8473
rect -19085 -8495 -18584 -8484
rect -18524 -8495 -17883 -8484
rect -19085 -8541 -19044 -8495
rect -17921 -8541 -17883 -8495
rect -17756 -8418 -17647 -8231
rect -17504 -8120 -17299 -8101
rect -17504 -8228 -17460 -8120
rect -17384 -8146 -17299 -8120
rect -16426 -8146 -16311 -8049
rect -16195 -8036 -16081 -8022
rect -15931 -8036 -15916 -7939
rect -16195 -8052 -15916 -8036
rect -15726 -7980 -14937 -7962
rect -15726 -7988 -15083 -7980
rect -15726 -8041 -15689 -7988
rect -15556 -8033 -15083 -7988
rect -14969 -8033 -14937 -7980
rect -15556 -8041 -14937 -8033
rect -16195 -8115 -16024 -8052
rect -15726 -8061 -14937 -8041
rect -14867 -7981 -14752 -7962
rect -14867 -8049 -14849 -7981
rect -14769 -8049 -14752 -7981
rect -14290 -7997 -14272 -7887
rect -14176 -7995 -14155 -7887
rect -10999 -7887 -10864 -7863
rect -12816 -7922 -12625 -7917
rect -12817 -7932 -12625 -7922
rect -12817 -7939 -12715 -7932
rect -12642 -7939 -12625 -7932
rect -14225 -7997 -14155 -7995
rect -14290 -8017 -14155 -7997
rect -13994 -7980 -13205 -7962
rect -13994 -7988 -13351 -7980
rect -17384 -8228 -16311 -8146
rect -17504 -8232 -16311 -8228
rect -16237 -8152 -16024 -8115
rect -16237 -8207 -16226 -8152
rect -16161 -8207 -16024 -8152
rect -16237 -8231 -16024 -8207
rect -15945 -8127 -15740 -8101
rect -15945 -8224 -15905 -8127
rect -15789 -8146 -15740 -8127
rect -14867 -8146 -14752 -8049
rect -14636 -8115 -14356 -8022
rect -13994 -8041 -13957 -7988
rect -13824 -8033 -13351 -7988
rect -13237 -8033 -13205 -7980
rect -13824 -8041 -13205 -8033
rect -13994 -8061 -13205 -8041
rect -13135 -7981 -13020 -7962
rect -13135 -8049 -13117 -7981
rect -13037 -8049 -13020 -7981
rect -12817 -8022 -12790 -7939
rect -15789 -8224 -14752 -8146
rect -15945 -8232 -14752 -8224
rect -14678 -8152 -14356 -8115
rect -14678 -8207 -14667 -8152
rect -14602 -8207 -14356 -8152
rect -14678 -8231 -14356 -8207
rect -17504 -8244 -17299 -8232
rect -15945 -8244 -15740 -8232
rect -17756 -8504 -17747 -8418
rect -17656 -8504 -17647 -8418
rect -17756 -8516 -17647 -8504
rect -17353 -8301 -17298 -8285
rect -17353 -8407 -17346 -8301
rect -17312 -8407 -17298 -8301
rect -17266 -8286 -16816 -8274
rect -17266 -8320 -17250 -8286
rect -17216 -8320 -17058 -8286
rect -17024 -8287 -16816 -8286
rect -17024 -8320 -16866 -8287
rect -17266 -8321 -16866 -8320
rect -16832 -8321 -16816 -8287
rect -17266 -8342 -16816 -8321
rect -16690 -8286 -16240 -8274
rect -16690 -8320 -16674 -8286
rect -16640 -8320 -16482 -8286
rect -16448 -8320 -16290 -8286
rect -16256 -8320 -16240 -8286
rect -16690 -8342 -16240 -8320
rect -16206 -8301 -16151 -8285
rect -17353 -8473 -17298 -8407
rect -17168 -8387 -17103 -8370
rect -17168 -8421 -17154 -8387
rect -17120 -8421 -17103 -8387
rect -17168 -8473 -17103 -8421
rect -16975 -8387 -16528 -8375
rect -16975 -8421 -16962 -8387
rect -16928 -8421 -16770 -8387
rect -16736 -8421 -16578 -8387
rect -16544 -8421 -16528 -8387
rect -16975 -8439 -16528 -8421
rect -16402 -8387 -16337 -8371
rect -16402 -8421 -16386 -8387
rect -16352 -8421 -16337 -8387
rect -16402 -8473 -16337 -8421
rect -16206 -8407 -16194 -8301
rect -16160 -8407 -16151 -8301
rect -16206 -8473 -16151 -8407
rect -17353 -8484 -16151 -8473
rect -17353 -8495 -16852 -8484
rect -16792 -8495 -16151 -8484
rect -19085 -8544 -18584 -8541
rect -18524 -8544 -17883 -8541
rect -19085 -8564 -17883 -8544
rect -17353 -8541 -17312 -8495
rect -16189 -8541 -16151 -8495
rect -17353 -8544 -16852 -8541
rect -16792 -8544 -16151 -8541
rect -17353 -8564 -16151 -8544
rect -15794 -8301 -15739 -8285
rect -15794 -8407 -15787 -8301
rect -15753 -8407 -15739 -8301
rect -15707 -8286 -15257 -8274
rect -15707 -8320 -15691 -8286
rect -15657 -8320 -15499 -8286
rect -15465 -8287 -15257 -8286
rect -15465 -8320 -15307 -8287
rect -15707 -8321 -15307 -8320
rect -15273 -8321 -15257 -8287
rect -15707 -8342 -15257 -8321
rect -15131 -8286 -14681 -8274
rect -15131 -8320 -15115 -8286
rect -15081 -8320 -14923 -8286
rect -14889 -8320 -14731 -8286
rect -14697 -8320 -14681 -8286
rect -15131 -8342 -14681 -8320
rect -14647 -8301 -14592 -8285
rect -15794 -8473 -15739 -8407
rect -15609 -8387 -15544 -8370
rect -15609 -8421 -15595 -8387
rect -15561 -8421 -15544 -8387
rect -15609 -8473 -15544 -8421
rect -15416 -8387 -14969 -8375
rect -15416 -8421 -15403 -8387
rect -15369 -8421 -15211 -8387
rect -15177 -8421 -15019 -8387
rect -14985 -8421 -14969 -8387
rect -15416 -8439 -14969 -8421
rect -14843 -8387 -14778 -8371
rect -14843 -8421 -14827 -8387
rect -14793 -8421 -14778 -8387
rect -14843 -8473 -14778 -8421
rect -14647 -8407 -14635 -8301
rect -14601 -8407 -14592 -8301
rect -14647 -8473 -14592 -8407
rect -15794 -8484 -14592 -8473
rect -15794 -8495 -15293 -8484
rect -15233 -8495 -14592 -8484
rect -15794 -8541 -15753 -8495
rect -14630 -8541 -14592 -8495
rect -14465 -8418 -14356 -8231
rect -14213 -8120 -14008 -8101
rect -14213 -8228 -14169 -8120
rect -14093 -8146 -14008 -8120
rect -13135 -8146 -13020 -8049
rect -12904 -8036 -12790 -8022
rect -12640 -8036 -12625 -7939
rect -12904 -8052 -12625 -8036
rect -12435 -7980 -11646 -7962
rect -12435 -7988 -11792 -7980
rect -12435 -8041 -12398 -7988
rect -12265 -8033 -11792 -7988
rect -11678 -8033 -11646 -7980
rect -12265 -8041 -11646 -8033
rect -12904 -8115 -12733 -8052
rect -12435 -8061 -11646 -8041
rect -11576 -7981 -11461 -7962
rect -11576 -8049 -11558 -7981
rect -11478 -8049 -11461 -7981
rect -10999 -7997 -10981 -7887
rect -10885 -7995 -10864 -7887
rect -9525 -7922 -9334 -7917
rect -9526 -7932 -9334 -7922
rect -9526 -7939 -9424 -7932
rect -9351 -7939 -9334 -7932
rect -10934 -7997 -10864 -7995
rect -10999 -8017 -10864 -7997
rect -10703 -7980 -9914 -7962
rect -10703 -7988 -10060 -7980
rect -14093 -8228 -13020 -8146
rect -14213 -8232 -13020 -8228
rect -12946 -8152 -12733 -8115
rect -12946 -8207 -12935 -8152
rect -12870 -8207 -12733 -8152
rect -12946 -8231 -12733 -8207
rect -12654 -8127 -12449 -8101
rect -12654 -8224 -12614 -8127
rect -12498 -8146 -12449 -8127
rect -11576 -8146 -11461 -8049
rect -11345 -8115 -11065 -8022
rect -10703 -8041 -10666 -7988
rect -10533 -8033 -10060 -7988
rect -9946 -8033 -9914 -7980
rect -10533 -8041 -9914 -8033
rect -10703 -8061 -9914 -8041
rect -9844 -7981 -9729 -7962
rect -9844 -8049 -9826 -7981
rect -9746 -8049 -9729 -7981
rect -9526 -8022 -9499 -7939
rect -12498 -8224 -11461 -8146
rect -12654 -8232 -11461 -8224
rect -11387 -8152 -11065 -8115
rect -11387 -8207 -11376 -8152
rect -11311 -8207 -11065 -8152
rect -11387 -8231 -11065 -8207
rect -14213 -8244 -14008 -8232
rect -12654 -8244 -12449 -8232
rect -14465 -8504 -14456 -8418
rect -14365 -8504 -14356 -8418
rect -14465 -8516 -14356 -8504
rect -14062 -8301 -14007 -8285
rect -14062 -8407 -14055 -8301
rect -14021 -8407 -14007 -8301
rect -13975 -8286 -13525 -8274
rect -13975 -8320 -13959 -8286
rect -13925 -8320 -13767 -8286
rect -13733 -8287 -13525 -8286
rect -13733 -8320 -13575 -8287
rect -13975 -8321 -13575 -8320
rect -13541 -8321 -13525 -8287
rect -13975 -8342 -13525 -8321
rect -13399 -8286 -12949 -8274
rect -13399 -8320 -13383 -8286
rect -13349 -8320 -13191 -8286
rect -13157 -8320 -12999 -8286
rect -12965 -8320 -12949 -8286
rect -13399 -8342 -12949 -8320
rect -12915 -8301 -12860 -8285
rect -14062 -8473 -14007 -8407
rect -13877 -8387 -13812 -8370
rect -13877 -8421 -13863 -8387
rect -13829 -8421 -13812 -8387
rect -13877 -8473 -13812 -8421
rect -13684 -8387 -13237 -8375
rect -13684 -8421 -13671 -8387
rect -13637 -8421 -13479 -8387
rect -13445 -8421 -13287 -8387
rect -13253 -8421 -13237 -8387
rect -13684 -8439 -13237 -8421
rect -13111 -8387 -13046 -8371
rect -13111 -8421 -13095 -8387
rect -13061 -8421 -13046 -8387
rect -13111 -8473 -13046 -8421
rect -12915 -8407 -12903 -8301
rect -12869 -8407 -12860 -8301
rect -12915 -8473 -12860 -8407
rect -14062 -8484 -12860 -8473
rect -14062 -8495 -13561 -8484
rect -13501 -8495 -12860 -8484
rect -15794 -8544 -15293 -8541
rect -15233 -8544 -14592 -8541
rect -15794 -8564 -14592 -8544
rect -14062 -8541 -14021 -8495
rect -12898 -8541 -12860 -8495
rect -14062 -8544 -13561 -8541
rect -13501 -8544 -12860 -8541
rect -14062 -8564 -12860 -8544
rect -12503 -8301 -12448 -8285
rect -12503 -8407 -12496 -8301
rect -12462 -8407 -12448 -8301
rect -12416 -8286 -11966 -8274
rect -12416 -8320 -12400 -8286
rect -12366 -8320 -12208 -8286
rect -12174 -8287 -11966 -8286
rect -12174 -8320 -12016 -8287
rect -12416 -8321 -12016 -8320
rect -11982 -8321 -11966 -8287
rect -12416 -8342 -11966 -8321
rect -11840 -8286 -11390 -8274
rect -11840 -8320 -11824 -8286
rect -11790 -8320 -11632 -8286
rect -11598 -8320 -11440 -8286
rect -11406 -8320 -11390 -8286
rect -11840 -8342 -11390 -8320
rect -11356 -8301 -11301 -8285
rect -12503 -8473 -12448 -8407
rect -12318 -8387 -12253 -8370
rect -12318 -8421 -12304 -8387
rect -12270 -8421 -12253 -8387
rect -12318 -8473 -12253 -8421
rect -12125 -8387 -11678 -8375
rect -12125 -8421 -12112 -8387
rect -12078 -8421 -11920 -8387
rect -11886 -8421 -11728 -8387
rect -11694 -8421 -11678 -8387
rect -12125 -8439 -11678 -8421
rect -11552 -8387 -11487 -8371
rect -11552 -8421 -11536 -8387
rect -11502 -8421 -11487 -8387
rect -11552 -8473 -11487 -8421
rect -11356 -8407 -11344 -8301
rect -11310 -8407 -11301 -8301
rect -11356 -8473 -11301 -8407
rect -12503 -8484 -11301 -8473
rect -12503 -8495 -12002 -8484
rect -11942 -8495 -11301 -8484
rect -12503 -8541 -12462 -8495
rect -11339 -8541 -11301 -8495
rect -11174 -8418 -11065 -8231
rect -10922 -8120 -10717 -8101
rect -10922 -8228 -10878 -8120
rect -10802 -8146 -10717 -8120
rect -9844 -8146 -9729 -8049
rect -9613 -8036 -9499 -8022
rect -9349 -8036 -9334 -7939
rect -9613 -8052 -9334 -8036
rect -9144 -7980 -8355 -7962
rect -9144 -7988 -8501 -7980
rect -9144 -8041 -9107 -7988
rect -8974 -8033 -8501 -7988
rect -8387 -8033 -8355 -7980
rect -8974 -8041 -8355 -8033
rect -9613 -8115 -9442 -8052
rect -9144 -8061 -8355 -8041
rect -8285 -7981 -8170 -7962
rect -8285 -8049 -8267 -7981
rect -8187 -8049 -8170 -7981
rect -10802 -8228 -9729 -8146
rect -10922 -8232 -9729 -8228
rect -9655 -8152 -9442 -8115
rect -9655 -8207 -9644 -8152
rect -9579 -8207 -9442 -8152
rect -9655 -8231 -9442 -8207
rect -9363 -8127 -9158 -8101
rect -9363 -8224 -9323 -8127
rect -9207 -8146 -9158 -8127
rect -8285 -8146 -8170 -8049
rect -8054 -8115 -7774 -8022
rect -9207 -8224 -8170 -8146
rect -9363 -8232 -8170 -8224
rect -8096 -8152 -7774 -8115
rect -8096 -8207 -8085 -8152
rect -8020 -8205 -7774 -8152
rect -8020 -8207 -4977 -8205
rect -8096 -8231 -4977 -8207
rect -10922 -8244 -10717 -8232
rect -9363 -8244 -9158 -8232
rect -7883 -8271 -4977 -8231
rect -11174 -8504 -11165 -8418
rect -11074 -8504 -11065 -8418
rect -11174 -8516 -11065 -8504
rect -10771 -8301 -10716 -8285
rect -10771 -8407 -10764 -8301
rect -10730 -8407 -10716 -8301
rect -10684 -8286 -10234 -8274
rect -10684 -8320 -10668 -8286
rect -10634 -8320 -10476 -8286
rect -10442 -8287 -10234 -8286
rect -10442 -8320 -10284 -8287
rect -10684 -8321 -10284 -8320
rect -10250 -8321 -10234 -8287
rect -10684 -8342 -10234 -8321
rect -10108 -8286 -9658 -8274
rect -10108 -8320 -10092 -8286
rect -10058 -8320 -9900 -8286
rect -9866 -8320 -9708 -8286
rect -9674 -8320 -9658 -8286
rect -10108 -8342 -9658 -8320
rect -9624 -8301 -9569 -8285
rect -10771 -8473 -10716 -8407
rect -10586 -8387 -10521 -8370
rect -10586 -8421 -10572 -8387
rect -10538 -8421 -10521 -8387
rect -10586 -8473 -10521 -8421
rect -10393 -8387 -9946 -8375
rect -10393 -8421 -10380 -8387
rect -10346 -8421 -10188 -8387
rect -10154 -8421 -9996 -8387
rect -9962 -8421 -9946 -8387
rect -10393 -8439 -9946 -8421
rect -9820 -8387 -9755 -8371
rect -9820 -8421 -9804 -8387
rect -9770 -8421 -9755 -8387
rect -9820 -8473 -9755 -8421
rect -9624 -8407 -9612 -8301
rect -9578 -8407 -9569 -8301
rect -9624 -8473 -9569 -8407
rect -10771 -8484 -9569 -8473
rect -10771 -8495 -10270 -8484
rect -10210 -8495 -9569 -8484
rect -12503 -8544 -12002 -8541
rect -11942 -8544 -11301 -8541
rect -12503 -8564 -11301 -8544
rect -10771 -8541 -10730 -8495
rect -9607 -8541 -9569 -8495
rect -10771 -8544 -10270 -8541
rect -10210 -8544 -9569 -8541
rect -10771 -8564 -9569 -8544
rect -9212 -8301 -9157 -8285
rect -9212 -8407 -9205 -8301
rect -9171 -8407 -9157 -8301
rect -9125 -8286 -8675 -8274
rect -9125 -8320 -9109 -8286
rect -9075 -8320 -8917 -8286
rect -8883 -8287 -8675 -8286
rect -8883 -8320 -8725 -8287
rect -9125 -8321 -8725 -8320
rect -8691 -8321 -8675 -8287
rect -9125 -8342 -8675 -8321
rect -8549 -8286 -8099 -8274
rect -8549 -8320 -8533 -8286
rect -8499 -8320 -8341 -8286
rect -8307 -8320 -8149 -8286
rect -8115 -8320 -8099 -8286
rect -8549 -8342 -8099 -8320
rect -8065 -8301 -8010 -8285
rect -9212 -8473 -9157 -8407
rect -9027 -8387 -8962 -8370
rect -9027 -8421 -9013 -8387
rect -8979 -8421 -8962 -8387
rect -9027 -8473 -8962 -8421
rect -8834 -8387 -8387 -8375
rect -8834 -8421 -8821 -8387
rect -8787 -8421 -8629 -8387
rect -8595 -8421 -8437 -8387
rect -8403 -8421 -8387 -8387
rect -8834 -8439 -8387 -8421
rect -8261 -8387 -8196 -8371
rect -8261 -8421 -8245 -8387
rect -8211 -8421 -8196 -8387
rect -8261 -8473 -8196 -8421
rect -8065 -8407 -8053 -8301
rect -8019 -8407 -8010 -8301
rect -8065 -8473 -8010 -8407
rect -9212 -8484 -8010 -8473
rect -9212 -8495 -8711 -8484
rect -8651 -8495 -8010 -8484
rect -9212 -8541 -9171 -8495
rect -8048 -8541 -8010 -8495
rect -7883 -8418 -7774 -8271
rect -7883 -8504 -7874 -8418
rect -7783 -8504 -7774 -8418
rect -7883 -8516 -7774 -8504
rect -9212 -8544 -8711 -8541
rect -8651 -8544 -8010 -8541
rect -9212 -8564 -8010 -8544
rect -21846 -8594 -21632 -8572
rect -22661 -8669 -22027 -8662
rect -22661 -8716 -22632 -8669
rect -22063 -8716 -22027 -8669
rect -22661 -8788 -22623 -8716
rect -22069 -8782 -22027 -8716
rect -21846 -8673 -21823 -8594
rect -21654 -8673 -21632 -8594
rect -21846 -8688 -21632 -8673
rect -21946 -8736 -21877 -8720
rect -22069 -8788 -22026 -8782
rect -22661 -8868 -22648 -8788
rect -22614 -8868 -22456 -8836
rect -22422 -8868 -22264 -8836
rect -22230 -8868 -22072 -8836
rect -22038 -8868 -22026 -8788
rect -22661 -8874 -22026 -8868
rect -22661 -8875 -22027 -8874
rect -21946 -8904 -21927 -8736
rect -23870 -8990 -23614 -8962
rect -23460 -8976 -22951 -8905
rect -24304 -8996 -23614 -8990
rect -24632 -9039 -24268 -9025
rect -24632 -9146 -24601 -9039
rect -24445 -9043 -24268 -9039
rect -24445 -9078 -24318 -9043
rect -24284 -9078 -24268 -9043
rect -24445 -9146 -24268 -9078
rect -24632 -9160 -24268 -9146
rect -24240 -9043 -23980 -9024
rect -24240 -9078 -24029 -9043
rect -23995 -9078 -23980 -9043
rect -24240 -9098 -23980 -9078
rect -24240 -9167 -24190 -9098
rect -23904 -9126 -23614 -8996
rect -24240 -9189 -24234 -9167
rect -24637 -9202 -24234 -9189
rect -24200 -9202 -24190 -9167
rect -24162 -9138 -23614 -9126
rect -24162 -9172 -24150 -9138
rect -23774 -9172 -23614 -9138
rect -24162 -9178 -23614 -9172
rect -23583 -9010 -23454 -8976
rect -23377 -9010 -22951 -8976
rect -22568 -8910 -21927 -8904
rect -22568 -8990 -22552 -8910
rect -22518 -8990 -22360 -8910
rect -22326 -8990 -22168 -8910
rect -22134 -8962 -21927 -8910
rect -21893 -8962 -21877 -8736
rect -21846 -8722 -21840 -8688
rect -21761 -8692 -21632 -8688
rect -21033 -8598 -20824 -8578
rect -21761 -8722 -21755 -8692
rect -21033 -8700 -21003 -8598
rect -20885 -8617 -20824 -8598
rect -8185 -8617 -8094 -8564
rect -20885 -8633 -19620 -8617
rect -20885 -8700 -19735 -8633
rect -21033 -8702 -19735 -8700
rect -19636 -8702 -19620 -8633
rect -21033 -8708 -19620 -8702
rect -19237 -8629 -16329 -8617
rect -19237 -8695 -19223 -8629
rect -19152 -8633 -16329 -8629
rect -19152 -8695 -16444 -8633
rect -19237 -8702 -16444 -8695
rect -16345 -8702 -16329 -8633
rect -19237 -8708 -16329 -8702
rect -15946 -8629 -13038 -8617
rect -15946 -8695 -15932 -8629
rect -15861 -8633 -13038 -8629
rect -15861 -8695 -13153 -8633
rect -15946 -8702 -13153 -8695
rect -13054 -8702 -13038 -8633
rect -15946 -8708 -13038 -8702
rect -12655 -8629 -9747 -8617
rect -12655 -8695 -12641 -8629
rect -12570 -8633 -9747 -8629
rect -12570 -8695 -9862 -8633
rect -12655 -8702 -9862 -8695
rect -9763 -8702 -9747 -8633
rect -12655 -8708 -9747 -8702
rect -9364 -8629 -7684 -8617
rect -9364 -8695 -9350 -8629
rect -9279 -8695 -7684 -8629
rect -9364 -8708 -7684 -8695
rect -21846 -8880 -21755 -8722
rect -21846 -8914 -21840 -8880
rect -21761 -8914 -21755 -8880
rect -21846 -8930 -21755 -8914
rect -21723 -8784 -21534 -8720
rect -21033 -8730 -20824 -8708
rect -21723 -8818 -21717 -8784
rect -21640 -8818 -21534 -8784
rect -22134 -8990 -21877 -8962
rect -21723 -8970 -21534 -8818
rect -20354 -8824 -20080 -8815
rect -20354 -8830 -20345 -8824
rect -20531 -8837 -20345 -8830
rect -20089 -8830 -20080 -8824
rect -19065 -8824 -18791 -8815
rect -19065 -8830 -19056 -8824
rect -20089 -8837 -19897 -8830
rect -20531 -8884 -20502 -8837
rect -19933 -8884 -19897 -8837
rect -20531 -8896 -20345 -8884
rect -20089 -8896 -19897 -8884
rect -20531 -8950 -19897 -8896
rect -19422 -8837 -19056 -8830
rect -18800 -8830 -18791 -8824
rect -18348 -8824 -18074 -8815
rect -18348 -8830 -18339 -8824
rect -19422 -8884 -19393 -8837
rect -19422 -8896 -19056 -8884
rect -18800 -8896 -18788 -8830
rect -19422 -8950 -18788 -8896
rect -18540 -8837 -18339 -8830
rect -18083 -8830 -18074 -8824
rect -17063 -8824 -16789 -8815
rect -17063 -8830 -17054 -8824
rect -18083 -8837 -17906 -8830
rect -18540 -8884 -18511 -8837
rect -17942 -8884 -17906 -8837
rect -18540 -8896 -18339 -8884
rect -18083 -8896 -17906 -8884
rect -18540 -8950 -17906 -8896
rect -17240 -8837 -17054 -8830
rect -16798 -8830 -16789 -8824
rect -15774 -8824 -15500 -8815
rect -15774 -8830 -15765 -8824
rect -16798 -8837 -16606 -8830
rect -17240 -8884 -17211 -8837
rect -16642 -8884 -16606 -8837
rect -17240 -8896 -17054 -8884
rect -16798 -8896 -16606 -8884
rect -17240 -8950 -16606 -8896
rect -16131 -8837 -15765 -8830
rect -15509 -8830 -15500 -8824
rect -15057 -8824 -14783 -8815
rect -15057 -8830 -15048 -8824
rect -16131 -8884 -16102 -8837
rect -16131 -8896 -15765 -8884
rect -15509 -8896 -15497 -8830
rect -16131 -8950 -15497 -8896
rect -15249 -8837 -15048 -8830
rect -14792 -8830 -14783 -8824
rect -13772 -8824 -13498 -8815
rect -13772 -8830 -13763 -8824
rect -14792 -8837 -14615 -8830
rect -15249 -8884 -15220 -8837
rect -14651 -8884 -14615 -8837
rect -15249 -8896 -15048 -8884
rect -14792 -8896 -14615 -8884
rect -15249 -8950 -14615 -8896
rect -13949 -8837 -13763 -8830
rect -13507 -8830 -13498 -8824
rect -12483 -8824 -12209 -8815
rect -12483 -8830 -12474 -8824
rect -13507 -8837 -13315 -8830
rect -13949 -8884 -13920 -8837
rect -13351 -8884 -13315 -8837
rect -13949 -8896 -13763 -8884
rect -13507 -8896 -13315 -8884
rect -13949 -8950 -13315 -8896
rect -12840 -8837 -12474 -8830
rect -12218 -8830 -12209 -8824
rect -11766 -8824 -11492 -8815
rect -11766 -8830 -11757 -8824
rect -12840 -8884 -12811 -8837
rect -12840 -8896 -12474 -8884
rect -12218 -8896 -12206 -8830
rect -12840 -8950 -12206 -8896
rect -11958 -8837 -11757 -8830
rect -11501 -8830 -11492 -8824
rect -10481 -8824 -10207 -8815
rect -10481 -8830 -10472 -8824
rect -11501 -8837 -11324 -8830
rect -11958 -8884 -11929 -8837
rect -11360 -8884 -11324 -8837
rect -11958 -8896 -11757 -8884
rect -11501 -8896 -11324 -8884
rect -11958 -8950 -11324 -8896
rect -10658 -8837 -10472 -8830
rect -10216 -8830 -10207 -8824
rect -9192 -8824 -8918 -8815
rect -9192 -8830 -9183 -8824
rect -10216 -8837 -10024 -8830
rect -10658 -8884 -10629 -8837
rect -10060 -8884 -10024 -8837
rect -10658 -8896 -10472 -8884
rect -10216 -8896 -10024 -8884
rect -10658 -8950 -10024 -8896
rect -9549 -8837 -9183 -8830
rect -8927 -8830 -8918 -8824
rect -8475 -8824 -8201 -8815
rect -8475 -8830 -8466 -8824
rect -9549 -8884 -9520 -8837
rect -9549 -8896 -9183 -8884
rect -8927 -8896 -8915 -8830
rect -9549 -8950 -8915 -8896
rect -8667 -8837 -8466 -8830
rect -8210 -8830 -8201 -8824
rect -8210 -8837 -8033 -8830
rect -8667 -8884 -8638 -8837
rect -8069 -8884 -8033 -8837
rect -8667 -8896 -8466 -8884
rect -8210 -8896 -8033 -8884
rect -8667 -8950 -8033 -8896
rect -20531 -8956 -19896 -8950
rect -21723 -8976 -21304 -8970
rect -22568 -8996 -21877 -8990
rect -23583 -9138 -22951 -9010
rect -23583 -9172 -23571 -9138
rect -23395 -9172 -22951 -9138
rect -22910 -9037 -22532 -9025
rect -22910 -9148 -22885 -9037
rect -22683 -9043 -22532 -9037
rect -22683 -9078 -22582 -9043
rect -22548 -9078 -22532 -9043
rect -22683 -9148 -22532 -9078
rect -22910 -9160 -22532 -9148
rect -22504 -9043 -22244 -9024
rect -22504 -9078 -22293 -9043
rect -22259 -9078 -22244 -9043
rect -22504 -9098 -22244 -9078
rect -23583 -9178 -23383 -9172
rect -24637 -9314 -24190 -9202
rect -23683 -9182 -23614 -9178
rect -23683 -9216 -23664 -9182
rect -23630 -9216 -23614 -9182
rect -23683 -9233 -23614 -9216
rect -23583 -9226 -23383 -9219
rect -24637 -9512 -24612 -9314
rect -24466 -9325 -24190 -9314
rect -23583 -9260 -23571 -9226
rect -23395 -9260 -23383 -9226
rect -23355 -9231 -22951 -9172
rect -22504 -9167 -22454 -9098
rect -22168 -9126 -21877 -8996
rect -22504 -9189 -22498 -9167
rect -22913 -9202 -22498 -9189
rect -22464 -9202 -22454 -9167
rect -22426 -9138 -21877 -9126
rect -22426 -9172 -22414 -9138
rect -22038 -9172 -21877 -9138
rect -22426 -9178 -21877 -9172
rect -21846 -9010 -21717 -8976
rect -21640 -9010 -21304 -8976
rect -21846 -9019 -21304 -9010
rect -21846 -9138 -21573 -9019
rect -21846 -9172 -21834 -9138
rect -21658 -9172 -21573 -9138
rect -21846 -9178 -21646 -9172
rect -22913 -9211 -22454 -9202
rect -23355 -9233 -23012 -9231
rect -24466 -9512 -24432 -9325
rect -24162 -9330 -23762 -9324
rect -24162 -9364 -24150 -9330
rect -23774 -9364 -23762 -9330
rect -24162 -9402 -24133 -9364
rect -24162 -9436 -24135 -9402
rect -23793 -9426 -23762 -9364
rect -23583 -9343 -23556 -9260
rect -23407 -9343 -23383 -9260
rect -22913 -9303 -22891 -9211
rect -22686 -9303 -22454 -9211
rect -21946 -9182 -21877 -9178
rect -21946 -9216 -21927 -9182
rect -21893 -9216 -21877 -9182
rect -21946 -9233 -21877 -9216
rect -21618 -9193 -21573 -9172
rect -21351 -9193 -21304 -9019
rect -20531 -9036 -20518 -8956
rect -20484 -9036 -20326 -8956
rect -20292 -9036 -20134 -8956
rect -20100 -9036 -19942 -8956
rect -19908 -9036 -19896 -8956
rect -20531 -9042 -19896 -9036
rect -19422 -8956 -18787 -8950
rect -19422 -9036 -19409 -8956
rect -19375 -9036 -19217 -8956
rect -19183 -9036 -19025 -8956
rect -18991 -9036 -18833 -8956
rect -18799 -9036 -18787 -8956
rect -19422 -9042 -18787 -9036
rect -18540 -8956 -17905 -8950
rect -18540 -9036 -18527 -8956
rect -18493 -9036 -18335 -8956
rect -18301 -9036 -18143 -8956
rect -18109 -9036 -17951 -8956
rect -17917 -9036 -17905 -8956
rect -18540 -9042 -17905 -9036
rect -17240 -8956 -16605 -8950
rect -17240 -9036 -17227 -8956
rect -17193 -9036 -17035 -8956
rect -17001 -9036 -16843 -8956
rect -16809 -9036 -16651 -8956
rect -16617 -9036 -16605 -8956
rect -17240 -9042 -16605 -9036
rect -16131 -8956 -15496 -8950
rect -16131 -9036 -16118 -8956
rect -16084 -9036 -15926 -8956
rect -15892 -9036 -15734 -8956
rect -15700 -9036 -15542 -8956
rect -15508 -9036 -15496 -8956
rect -16131 -9042 -15496 -9036
rect -15249 -8956 -14614 -8950
rect -15249 -9036 -15236 -8956
rect -15202 -9036 -15044 -8956
rect -15010 -9036 -14852 -8956
rect -14818 -9036 -14660 -8956
rect -14626 -9036 -14614 -8956
rect -15249 -9042 -14614 -9036
rect -13949 -8956 -13314 -8950
rect -13949 -9036 -13936 -8956
rect -13902 -9036 -13744 -8956
rect -13710 -9036 -13552 -8956
rect -13518 -9036 -13360 -8956
rect -13326 -9036 -13314 -8956
rect -13949 -9042 -13314 -9036
rect -12840 -8956 -12205 -8950
rect -12840 -9036 -12827 -8956
rect -12793 -9036 -12635 -8956
rect -12601 -9036 -12443 -8956
rect -12409 -9036 -12251 -8956
rect -12217 -9036 -12205 -8956
rect -12840 -9042 -12205 -9036
rect -11958 -8956 -11323 -8950
rect -11958 -9036 -11945 -8956
rect -11911 -9036 -11753 -8956
rect -11719 -9036 -11561 -8956
rect -11527 -9036 -11369 -8956
rect -11335 -9036 -11323 -8956
rect -11958 -9042 -11323 -9036
rect -10658 -8956 -10023 -8950
rect -10658 -9036 -10645 -8956
rect -10611 -9036 -10453 -8956
rect -10419 -9036 -10261 -8956
rect -10227 -9036 -10069 -8956
rect -10035 -9036 -10023 -8956
rect -10658 -9042 -10023 -9036
rect -9549 -8956 -8914 -8950
rect -9549 -9036 -9536 -8956
rect -9502 -9036 -9344 -8956
rect -9310 -9036 -9152 -8956
rect -9118 -9036 -8960 -8956
rect -8926 -9036 -8914 -8956
rect -9549 -9042 -8914 -9036
rect -8667 -8956 -8032 -8950
rect -8667 -9036 -8654 -8956
rect -8620 -9036 -8462 -8956
rect -8428 -9036 -8270 -8956
rect -8236 -9036 -8078 -8956
rect -8044 -9036 -8032 -8956
rect -8667 -9042 -8032 -9036
rect -20531 -9043 -19897 -9042
rect -19422 -9043 -18788 -9042
rect -18540 -9043 -17906 -9042
rect -17240 -9043 -16606 -9042
rect -16131 -9043 -15497 -9042
rect -15249 -9043 -14615 -9042
rect -13949 -9043 -13315 -9042
rect -12840 -9043 -12206 -9042
rect -11958 -9043 -11324 -9042
rect -10658 -9043 -10024 -9042
rect -9549 -9043 -8915 -9042
rect -8667 -9043 -8033 -9042
rect -20438 -9078 -19860 -9072
rect -20438 -9158 -20422 -9078
rect -20388 -9158 -20230 -9078
rect -20196 -9158 -20038 -9078
rect -20004 -9158 -19860 -9078
rect -20438 -9159 -19860 -9158
rect -20438 -9164 -19979 -9159
rect -21846 -9226 -21646 -9219
rect -22913 -9325 -22454 -9303
rect -21846 -9260 -21834 -9226
rect -21658 -9260 -21646 -9226
rect -21618 -9233 -21304 -9193
rect -20566 -9211 -20402 -9193
rect -20566 -9220 -20452 -9211
rect -23583 -9362 -23552 -9343
rect -23420 -9362 -23383 -9343
rect -23583 -9369 -23383 -9362
rect -22426 -9330 -22026 -9324
rect -22426 -9364 -22414 -9330
rect -22038 -9364 -22026 -9330
rect -23800 -9436 -23762 -9426
rect -24162 -9447 -23762 -9436
rect -22426 -9402 -22397 -9364
rect -22426 -9436 -22399 -9402
rect -22057 -9426 -22026 -9364
rect -21846 -9343 -21819 -9260
rect -21670 -9343 -21646 -9260
rect -20566 -9300 -20534 -9220
rect -20418 -9246 -20402 -9211
rect -20436 -9300 -20402 -9246
rect -20566 -9328 -20402 -9300
rect -20374 -9211 -20114 -9192
rect -20374 -9246 -20163 -9211
rect -20129 -9246 -20114 -9211
rect -20374 -9266 -20114 -9246
rect -21846 -9362 -21815 -9343
rect -21683 -9362 -21646 -9343
rect -20374 -9335 -20324 -9266
rect -20038 -9294 -19979 -9164
rect -20374 -9356 -20368 -9335
rect -21846 -9369 -21646 -9362
rect -22064 -9436 -22026 -9426
rect -22426 -9447 -22026 -9436
rect -20762 -9370 -20368 -9356
rect -20334 -9370 -20324 -9335
rect -20296 -9306 -19979 -9294
rect -20296 -9340 -20284 -9306
rect -19896 -9307 -19860 -9159
rect -19329 -9078 -18751 -9072
rect -19329 -9158 -19313 -9078
rect -19279 -9158 -19121 -9078
rect -19087 -9158 -18929 -9078
rect -18895 -9158 -18751 -9078
rect -19329 -9164 -18751 -9158
rect -18447 -9078 -17869 -9072
rect -18447 -9158 -18431 -9078
rect -18397 -9158 -18239 -9078
rect -18205 -9158 -18047 -9078
rect -18013 -9158 -17869 -9078
rect -18447 -9164 -17869 -9158
rect -17147 -9078 -16569 -9072
rect -17147 -9158 -17131 -9078
rect -17097 -9158 -16939 -9078
rect -16905 -9158 -16747 -9078
rect -16713 -9158 -16569 -9078
rect -17147 -9159 -16569 -9158
rect -17147 -9164 -16688 -9159
rect -19908 -9340 -19860 -9307
rect -19457 -9211 -19293 -9193
rect -19457 -9221 -19343 -9211
rect -19457 -9301 -19423 -9221
rect -19309 -9246 -19293 -9211
rect -19325 -9301 -19293 -9246
rect -19457 -9328 -19293 -9301
rect -19265 -9211 -19005 -9192
rect -19265 -9246 -19054 -9211
rect -19020 -9246 -19005 -9211
rect -19265 -9266 -19005 -9246
rect -18929 -9216 -18751 -9164
rect -18575 -9211 -18411 -9193
rect -18575 -9216 -18461 -9211
rect -18929 -9246 -18461 -9216
rect -18427 -9246 -18411 -9211
rect -20296 -9346 -19860 -9340
rect -19265 -9335 -19215 -9266
rect -18929 -9294 -18411 -9246
rect -19265 -9357 -19259 -9335
rect -20762 -9413 -20324 -9370
rect -20762 -9479 -20743 -9413
rect -20490 -9479 -20324 -9413
rect -20762 -9493 -20324 -9479
rect -19457 -9370 -19259 -9357
rect -19225 -9370 -19215 -9335
rect -19187 -9306 -18411 -9294
rect -19187 -9340 -19175 -9306
rect -18799 -9340 -18751 -9306
rect -18575 -9328 -18411 -9306
rect -18383 -9211 -18123 -9192
rect -18383 -9246 -18172 -9211
rect -18138 -9246 -18123 -9211
rect -18383 -9266 -18123 -9246
rect -18047 -9209 -17869 -9164
rect -19187 -9346 -18751 -9340
rect -18383 -9335 -18333 -9266
rect -18047 -9289 -18002 -9209
rect -17882 -9289 -17869 -9209
rect -18047 -9294 -17869 -9289
rect -18383 -9357 -18377 -9335
rect -19457 -9424 -19215 -9370
rect -19457 -9484 -19433 -9424
rect -19248 -9484 -19215 -9424
rect -24637 -9527 -24432 -9512
rect -20296 -9498 -19896 -9492
rect -19457 -9493 -19215 -9484
rect -18575 -9370 -18377 -9357
rect -18343 -9370 -18333 -9335
rect -18305 -9306 -17869 -9294
rect -18305 -9340 -18293 -9306
rect -17917 -9340 -17869 -9306
rect -17275 -9211 -17111 -9193
rect -17275 -9220 -17161 -9211
rect -17275 -9300 -17243 -9220
rect -17127 -9246 -17111 -9211
rect -17145 -9300 -17111 -9246
rect -17275 -9328 -17111 -9300
rect -17083 -9211 -16823 -9192
rect -17083 -9246 -16872 -9211
rect -16838 -9246 -16823 -9211
rect -17083 -9266 -16823 -9246
rect -18305 -9346 -17869 -9340
rect -17083 -9335 -17033 -9266
rect -16747 -9294 -16688 -9164
rect -17083 -9356 -17077 -9335
rect -18575 -9375 -18333 -9370
rect -18575 -9450 -18561 -9375
rect -18416 -9450 -18333 -9375
rect -20296 -9532 -20284 -9498
rect -19908 -9532 -19896 -9498
rect -20296 -9570 -19896 -9532
rect -20296 -9615 -20269 -9570
rect -20278 -9622 -20269 -9615
rect -19934 -9615 -19896 -9570
rect -19187 -9498 -18787 -9492
rect -18575 -9493 -18333 -9450
rect -17471 -9370 -17077 -9356
rect -17043 -9370 -17033 -9335
rect -17005 -9306 -16688 -9294
rect -17005 -9340 -16993 -9306
rect -16605 -9307 -16569 -9159
rect -16038 -9078 -15460 -9072
rect -16038 -9158 -16022 -9078
rect -15988 -9158 -15830 -9078
rect -15796 -9158 -15638 -9078
rect -15604 -9158 -15460 -9078
rect -16038 -9164 -15460 -9158
rect -15156 -9078 -14578 -9072
rect -15156 -9158 -15140 -9078
rect -15106 -9158 -14948 -9078
rect -14914 -9158 -14756 -9078
rect -14722 -9158 -14578 -9078
rect -15156 -9164 -14578 -9158
rect -13856 -9078 -13278 -9072
rect -13856 -9158 -13840 -9078
rect -13806 -9158 -13648 -9078
rect -13614 -9158 -13456 -9078
rect -13422 -9158 -13278 -9078
rect -13856 -9159 -13278 -9158
rect -13856 -9164 -13397 -9159
rect -16617 -9340 -16569 -9307
rect -16166 -9211 -16002 -9193
rect -16166 -9221 -16052 -9211
rect -16166 -9301 -16132 -9221
rect -16018 -9246 -16002 -9211
rect -16034 -9301 -16002 -9246
rect -16166 -9328 -16002 -9301
rect -15974 -9211 -15714 -9192
rect -15974 -9246 -15763 -9211
rect -15729 -9246 -15714 -9211
rect -15974 -9266 -15714 -9246
rect -15638 -9216 -15460 -9164
rect -15284 -9211 -15120 -9193
rect -15284 -9216 -15170 -9211
rect -15638 -9246 -15170 -9216
rect -15136 -9246 -15120 -9211
rect -17005 -9346 -16569 -9340
rect -15974 -9335 -15924 -9266
rect -15638 -9294 -15120 -9246
rect -15974 -9357 -15968 -9335
rect -17471 -9413 -17033 -9370
rect -17471 -9479 -17452 -9413
rect -17199 -9479 -17033 -9413
rect -19187 -9532 -19175 -9498
rect -18799 -9532 -18787 -9498
rect -19187 -9570 -18787 -9532
rect -19187 -9604 -19160 -9570
rect -18825 -9604 -18787 -9570
rect -19187 -9615 -19033 -9604
rect -19934 -9622 -19925 -9615
rect -20278 -9631 -19925 -9622
rect -19044 -9637 -19033 -9615
rect -18971 -9615 -18787 -9604
rect -18305 -9498 -17905 -9492
rect -17471 -9493 -17033 -9479
rect -16166 -9370 -15968 -9357
rect -15934 -9370 -15924 -9335
rect -15896 -9306 -15120 -9294
rect -15896 -9340 -15884 -9306
rect -15508 -9340 -15460 -9306
rect -15284 -9328 -15120 -9306
rect -15092 -9211 -14832 -9192
rect -15092 -9246 -14881 -9211
rect -14847 -9246 -14832 -9211
rect -15092 -9266 -14832 -9246
rect -14756 -9209 -14578 -9164
rect -15896 -9346 -15460 -9340
rect -15092 -9335 -15042 -9266
rect -14756 -9289 -14711 -9209
rect -14591 -9289 -14578 -9209
rect -14756 -9294 -14578 -9289
rect -15092 -9357 -15086 -9335
rect -16166 -9424 -15924 -9370
rect -16166 -9484 -16142 -9424
rect -15957 -9484 -15924 -9424
rect -18305 -9532 -18293 -9498
rect -17917 -9532 -17905 -9498
rect -18305 -9570 -17905 -9532
rect -18305 -9604 -18278 -9570
rect -17943 -9604 -17905 -9570
rect -18305 -9615 -18166 -9604
rect -18971 -9637 -18960 -9615
rect -19044 -9648 -18960 -9637
rect -18179 -9654 -18166 -9615
rect -18114 -9615 -17905 -9604
rect -17005 -9498 -16605 -9492
rect -16166 -9493 -15924 -9484
rect -15284 -9370 -15086 -9357
rect -15052 -9370 -15042 -9335
rect -15014 -9306 -14578 -9294
rect -15014 -9340 -15002 -9306
rect -14626 -9340 -14578 -9306
rect -13984 -9211 -13820 -9193
rect -13984 -9220 -13870 -9211
rect -13984 -9300 -13952 -9220
rect -13836 -9246 -13820 -9211
rect -13854 -9300 -13820 -9246
rect -13984 -9328 -13820 -9300
rect -13792 -9211 -13532 -9192
rect -13792 -9246 -13581 -9211
rect -13547 -9246 -13532 -9211
rect -13792 -9266 -13532 -9246
rect -15014 -9346 -14578 -9340
rect -13792 -9335 -13742 -9266
rect -13456 -9294 -13397 -9164
rect -13792 -9356 -13786 -9335
rect -15284 -9375 -15042 -9370
rect -15284 -9450 -15270 -9375
rect -15125 -9450 -15042 -9375
rect -17005 -9532 -16993 -9498
rect -16617 -9532 -16605 -9498
rect -17005 -9570 -16605 -9532
rect -17005 -9615 -16978 -9570
rect -18114 -9654 -18101 -9615
rect -16987 -9622 -16978 -9615
rect -16643 -9615 -16605 -9570
rect -15896 -9498 -15496 -9492
rect -15284 -9493 -15042 -9450
rect -14180 -9370 -13786 -9356
rect -13752 -9370 -13742 -9335
rect -13714 -9306 -13397 -9294
rect -13714 -9340 -13702 -9306
rect -13314 -9307 -13278 -9159
rect -12747 -9078 -12169 -9072
rect -12747 -9158 -12731 -9078
rect -12697 -9158 -12539 -9078
rect -12505 -9158 -12347 -9078
rect -12313 -9158 -12169 -9078
rect -12747 -9164 -12169 -9158
rect -11865 -9078 -11287 -9072
rect -11865 -9158 -11849 -9078
rect -11815 -9158 -11657 -9078
rect -11623 -9158 -11465 -9078
rect -11431 -9158 -11287 -9078
rect -11865 -9164 -11287 -9158
rect -10565 -9078 -9987 -9072
rect -10565 -9158 -10549 -9078
rect -10515 -9158 -10357 -9078
rect -10323 -9158 -10165 -9078
rect -10131 -9158 -9987 -9078
rect -10565 -9159 -9987 -9158
rect -10565 -9164 -10106 -9159
rect -13326 -9340 -13278 -9307
rect -12875 -9211 -12711 -9193
rect -12875 -9221 -12761 -9211
rect -12875 -9301 -12841 -9221
rect -12727 -9246 -12711 -9211
rect -12743 -9301 -12711 -9246
rect -12875 -9328 -12711 -9301
rect -12683 -9211 -12423 -9192
rect -12683 -9246 -12472 -9211
rect -12438 -9246 -12423 -9211
rect -12683 -9266 -12423 -9246
rect -12347 -9216 -12169 -9164
rect -11993 -9211 -11829 -9193
rect -11993 -9216 -11879 -9211
rect -12347 -9246 -11879 -9216
rect -11845 -9246 -11829 -9211
rect -13714 -9346 -13278 -9340
rect -12683 -9335 -12633 -9266
rect -12347 -9294 -11829 -9246
rect -12683 -9357 -12677 -9335
rect -14180 -9413 -13742 -9370
rect -14180 -9479 -14161 -9413
rect -13908 -9479 -13742 -9413
rect -15896 -9532 -15884 -9498
rect -15508 -9532 -15496 -9498
rect -15896 -9570 -15496 -9532
rect -15896 -9604 -15869 -9570
rect -15534 -9604 -15496 -9570
rect -15896 -9615 -15742 -9604
rect -16643 -9622 -16634 -9615
rect -16987 -9631 -16634 -9622
rect -15753 -9637 -15742 -9615
rect -15680 -9615 -15496 -9604
rect -15014 -9498 -14614 -9492
rect -14180 -9493 -13742 -9479
rect -12875 -9370 -12677 -9357
rect -12643 -9370 -12633 -9335
rect -12605 -9306 -11829 -9294
rect -12605 -9340 -12593 -9306
rect -12217 -9340 -12169 -9306
rect -11993 -9328 -11829 -9306
rect -11801 -9211 -11541 -9192
rect -11801 -9246 -11590 -9211
rect -11556 -9246 -11541 -9211
rect -11801 -9266 -11541 -9246
rect -11465 -9209 -11287 -9164
rect -12605 -9346 -12169 -9340
rect -11801 -9335 -11751 -9266
rect -11465 -9289 -11420 -9209
rect -11300 -9289 -11287 -9209
rect -11465 -9294 -11287 -9289
rect -11801 -9357 -11795 -9335
rect -12875 -9424 -12633 -9370
rect -12875 -9484 -12851 -9424
rect -12666 -9484 -12633 -9424
rect -15014 -9532 -15002 -9498
rect -14626 -9532 -14614 -9498
rect -15014 -9570 -14614 -9532
rect -15014 -9604 -14987 -9570
rect -14652 -9604 -14614 -9570
rect -15014 -9615 -14875 -9604
rect -15680 -9637 -15669 -9615
rect -15753 -9648 -15669 -9637
rect -18179 -9667 -18101 -9654
rect -14888 -9654 -14875 -9615
rect -14823 -9615 -14614 -9604
rect -13714 -9498 -13314 -9492
rect -12875 -9493 -12633 -9484
rect -11993 -9370 -11795 -9357
rect -11761 -9370 -11751 -9335
rect -11723 -9306 -11287 -9294
rect -11723 -9340 -11711 -9306
rect -11335 -9340 -11287 -9306
rect -10693 -9211 -10529 -9193
rect -10693 -9220 -10579 -9211
rect -10693 -9300 -10661 -9220
rect -10545 -9246 -10529 -9211
rect -10563 -9300 -10529 -9246
rect -10693 -9328 -10529 -9300
rect -10501 -9211 -10241 -9192
rect -10501 -9246 -10290 -9211
rect -10256 -9246 -10241 -9211
rect -10501 -9266 -10241 -9246
rect -11723 -9346 -11287 -9340
rect -10501 -9335 -10451 -9266
rect -10165 -9294 -10106 -9164
rect -10501 -9356 -10495 -9335
rect -11993 -9375 -11751 -9370
rect -11993 -9450 -11979 -9375
rect -11834 -9450 -11751 -9375
rect -13714 -9532 -13702 -9498
rect -13326 -9532 -13314 -9498
rect -13714 -9570 -13314 -9532
rect -13714 -9615 -13687 -9570
rect -14823 -9654 -14810 -9615
rect -13696 -9622 -13687 -9615
rect -13352 -9615 -13314 -9570
rect -12605 -9498 -12205 -9492
rect -11993 -9493 -11751 -9450
rect -10889 -9370 -10495 -9356
rect -10461 -9370 -10451 -9335
rect -10423 -9306 -10106 -9294
rect -10423 -9340 -10411 -9306
rect -10023 -9307 -9987 -9159
rect -9456 -9078 -8878 -9072
rect -9456 -9158 -9440 -9078
rect -9406 -9158 -9248 -9078
rect -9214 -9158 -9056 -9078
rect -9022 -9158 -8878 -9078
rect -9456 -9164 -8878 -9158
rect -8574 -9078 -7996 -9072
rect -8574 -9158 -8558 -9078
rect -8524 -9158 -8366 -9078
rect -8332 -9158 -8174 -9078
rect -8140 -9158 -7996 -9078
rect -8574 -9164 -7996 -9158
rect -10035 -9340 -9987 -9307
rect -9584 -9211 -9420 -9193
rect -9584 -9221 -9470 -9211
rect -9584 -9301 -9550 -9221
rect -9436 -9246 -9420 -9211
rect -9452 -9301 -9420 -9246
rect -9584 -9328 -9420 -9301
rect -9392 -9211 -9132 -9192
rect -9392 -9246 -9181 -9211
rect -9147 -9246 -9132 -9211
rect -9392 -9266 -9132 -9246
rect -9056 -9216 -8878 -9164
rect -8702 -9211 -8538 -9193
rect -8702 -9216 -8588 -9211
rect -9056 -9246 -8588 -9216
rect -8554 -9246 -8538 -9211
rect -10423 -9346 -9987 -9340
rect -9392 -9335 -9342 -9266
rect -9056 -9294 -8538 -9246
rect -9392 -9357 -9386 -9335
rect -10889 -9413 -10451 -9370
rect -10889 -9479 -10870 -9413
rect -10617 -9479 -10451 -9413
rect -12605 -9532 -12593 -9498
rect -12217 -9532 -12205 -9498
rect -12605 -9570 -12205 -9532
rect -12605 -9604 -12578 -9570
rect -12243 -9604 -12205 -9570
rect -12605 -9615 -12451 -9604
rect -13352 -9622 -13343 -9615
rect -13696 -9631 -13343 -9622
rect -12462 -9637 -12451 -9615
rect -12389 -9615 -12205 -9604
rect -11723 -9498 -11323 -9492
rect -10889 -9493 -10451 -9479
rect -9584 -9370 -9386 -9357
rect -9352 -9370 -9342 -9335
rect -9314 -9306 -8538 -9294
rect -9314 -9340 -9302 -9306
rect -8926 -9340 -8878 -9306
rect -8702 -9328 -8538 -9306
rect -8510 -9211 -8250 -9192
rect -8510 -9246 -8299 -9211
rect -8265 -9246 -8250 -9211
rect -8510 -9266 -8250 -9246
rect -8174 -9209 -7996 -9164
rect -9314 -9346 -8878 -9340
rect -8510 -9335 -8460 -9266
rect -8174 -9289 -8129 -9209
rect -8009 -9289 -7996 -9209
rect -8174 -9294 -7996 -9289
rect -8510 -9357 -8504 -9335
rect -9584 -9424 -9342 -9370
rect -9584 -9484 -9560 -9424
rect -9375 -9484 -9342 -9424
rect -11723 -9532 -11711 -9498
rect -11335 -9532 -11323 -9498
rect -11723 -9570 -11323 -9532
rect -11723 -9604 -11696 -9570
rect -11361 -9604 -11323 -9570
rect -11723 -9615 -11584 -9604
rect -12389 -9637 -12378 -9615
rect -12462 -9648 -12378 -9637
rect -14888 -9667 -14810 -9654
rect -11597 -9654 -11584 -9615
rect -11532 -9615 -11323 -9604
rect -10423 -9498 -10023 -9492
rect -9584 -9493 -9342 -9484
rect -8702 -9370 -8504 -9357
rect -8470 -9370 -8460 -9335
rect -8432 -9306 -7996 -9294
rect -8432 -9340 -8420 -9306
rect -8044 -9340 -7996 -9306
rect -8432 -9346 -7996 -9340
rect -8702 -9375 -8460 -9370
rect -8702 -9450 -8688 -9375
rect -8543 -9450 -8460 -9375
rect -10423 -9532 -10411 -9498
rect -10035 -9532 -10023 -9498
rect -10423 -9570 -10023 -9532
rect -10423 -9615 -10396 -9570
rect -11532 -9654 -11519 -9615
rect -10405 -9622 -10396 -9615
rect -10061 -9615 -10023 -9570
rect -9314 -9498 -8914 -9492
rect -8702 -9493 -8460 -9450
rect -9314 -9532 -9302 -9498
rect -8926 -9532 -8914 -9498
rect -9314 -9570 -8914 -9532
rect -9314 -9604 -9287 -9570
rect -8952 -9604 -8914 -9570
rect -9314 -9615 -9160 -9604
rect -10061 -9622 -10052 -9615
rect -10405 -9631 -10052 -9622
rect -9171 -9637 -9160 -9615
rect -9098 -9615 -8914 -9604
rect -8432 -9498 -8032 -9492
rect -8432 -9532 -8420 -9498
rect -8044 -9532 -8032 -9498
rect -8432 -9570 -8032 -9532
rect -8432 -9604 -8405 -9570
rect -8070 -9604 -8032 -9570
rect -8432 -9615 -8293 -9604
rect -9098 -9637 -9087 -9615
rect -9171 -9648 -9087 -9637
rect -11597 -9667 -11519 -9654
rect -8306 -9654 -8293 -9615
rect -8241 -9615 -8032 -9604
rect -8241 -9654 -8228 -9615
rect -8306 -9667 -8228 -9654
rect -23304 -9920 -11066 -9836
rect -23583 -10566 -23369 -10544
rect -24397 -10641 -23763 -10634
rect -24397 -10688 -24368 -10641
rect -23799 -10688 -23763 -10641
rect -24397 -10760 -24359 -10688
rect -23805 -10754 -23763 -10688
rect -23583 -10645 -23560 -10566
rect -23391 -10645 -23369 -10566
rect -23583 -10660 -23369 -10645
rect -23683 -10708 -23614 -10692
rect -23805 -10760 -23762 -10754
rect -24397 -10840 -24384 -10760
rect -24350 -10840 -24192 -10808
rect -24158 -10840 -24000 -10808
rect -23966 -10840 -23808 -10808
rect -23774 -10840 -23762 -10760
rect -24397 -10846 -23762 -10840
rect -24397 -10847 -23763 -10846
rect -23683 -10876 -23664 -10708
rect -24304 -10882 -23664 -10876
rect -24304 -10962 -24288 -10882
rect -24254 -10962 -24096 -10882
rect -24062 -10962 -23904 -10882
rect -23870 -10934 -23664 -10882
rect -23630 -10934 -23614 -10708
rect -23583 -10694 -23577 -10660
rect -23498 -10664 -23369 -10660
rect -23498 -10694 -23492 -10664
rect -23304 -10692 -23211 -9920
rect -23583 -10852 -23492 -10694
rect -23583 -10886 -23577 -10852
rect -23498 -10886 -23492 -10852
rect -23583 -10902 -23492 -10886
rect -23460 -10756 -23211 -10692
rect -23460 -10790 -23454 -10756
rect -23377 -10790 -23211 -10756
rect -23870 -10962 -23614 -10934
rect -23460 -10948 -23211 -10790
rect -24304 -10968 -23614 -10962
rect -24862 -11059 -24837 -10970
rect -24748 -10997 -24696 -10970
rect -24748 -11015 -24268 -10997
rect -24748 -11050 -24318 -11015
rect -24284 -11050 -24268 -11015
rect -24748 -11059 -24268 -11050
rect -24862 -11132 -24268 -11059
rect -24240 -11015 -23980 -10996
rect -24240 -11050 -24029 -11015
rect -23995 -11050 -23980 -11015
rect -24240 -11070 -23980 -11050
rect -24240 -11139 -24190 -11070
rect -23904 -11098 -23614 -10968
rect -24240 -11161 -24234 -11139
rect -24632 -11174 -24234 -11161
rect -24200 -11174 -24190 -11139
rect -24162 -11110 -23614 -11098
rect -24162 -11144 -24150 -11110
rect -23774 -11144 -23614 -11110
rect -24162 -11150 -23614 -11144
rect -23583 -10982 -23454 -10948
rect -23377 -10982 -23211 -10948
rect -23583 -11110 -23211 -10982
rect -23583 -11144 -23571 -11110
rect -23395 -11144 -23211 -11110
rect -23583 -11150 -23383 -11144
rect -24632 -11187 -24190 -11174
rect -24632 -11278 -24563 -11187
rect -24335 -11278 -24190 -11187
rect -23683 -11154 -23614 -11150
rect -23683 -11188 -23664 -11154
rect -23630 -11188 -23614 -11154
rect -23683 -11205 -23614 -11188
rect -23583 -11198 -23383 -11191
rect -24632 -11297 -24190 -11278
rect -23583 -11232 -23571 -11198
rect -23395 -11232 -23383 -11198
rect -23355 -11205 -23211 -11144
rect -23088 -10067 -14356 -9983
rect -24162 -11302 -23762 -11296
rect -24162 -11336 -24150 -11302
rect -23774 -11336 -23762 -11302
rect -24162 -11374 -24133 -11336
rect -24162 -11408 -24135 -11374
rect -23793 -11398 -23762 -11336
rect -23583 -11315 -23556 -11232
rect -23407 -11315 -23383 -11232
rect -23583 -11334 -23552 -11315
rect -23420 -11334 -23383 -11315
rect -23583 -11341 -23383 -11334
rect -23800 -11408 -23762 -11398
rect -24162 -11419 -23762 -11408
rect -23583 -11858 -23369 -11836
rect -24397 -11933 -23763 -11926
rect -24397 -11980 -24368 -11933
rect -23799 -11980 -23763 -11933
rect -24397 -12052 -24359 -11980
rect -23805 -12046 -23763 -11980
rect -23583 -11937 -23560 -11858
rect -23391 -11937 -23369 -11858
rect -23583 -11952 -23369 -11937
rect -23683 -12000 -23614 -11984
rect -23805 -12052 -23762 -12046
rect -24397 -12132 -24384 -12052
rect -24350 -12132 -24192 -12100
rect -24158 -12132 -24000 -12100
rect -23966 -12132 -23808 -12100
rect -23774 -12132 -23762 -12052
rect -24397 -12138 -23762 -12132
rect -24397 -12139 -23763 -12138
rect -23683 -12168 -23664 -12000
rect -24304 -12174 -23664 -12168
rect -24304 -12254 -24288 -12174
rect -24254 -12254 -24096 -12174
rect -24062 -12254 -23904 -12174
rect -23870 -12226 -23664 -12174
rect -23630 -12226 -23614 -12000
rect -23583 -11986 -23577 -11952
rect -23498 -11956 -23369 -11952
rect -23498 -11986 -23492 -11956
rect -23583 -12144 -23492 -11986
rect -23583 -12178 -23577 -12144
rect -23498 -12178 -23492 -12144
rect -23583 -12194 -23492 -12178
rect -23460 -12014 -23271 -11984
rect -23088 -12014 -22951 -10067
rect -21259 -10215 -17647 -10131
rect -21850 -10566 -21636 -10544
rect -22660 -10641 -22026 -10634
rect -22660 -10688 -22631 -10641
rect -22062 -10688 -22026 -10641
rect -22660 -10760 -22622 -10688
rect -22068 -10754 -22026 -10688
rect -21850 -10645 -21827 -10566
rect -21658 -10645 -21636 -10566
rect -21850 -10660 -21636 -10645
rect -21950 -10708 -21881 -10692
rect -22068 -10760 -22025 -10754
rect -22660 -10840 -22647 -10760
rect -22613 -10840 -22455 -10808
rect -22421 -10840 -22263 -10808
rect -22229 -10840 -22071 -10808
rect -22037 -10840 -22025 -10760
rect -22660 -10846 -22025 -10840
rect -22660 -10847 -22026 -10846
rect -21950 -10876 -21931 -10708
rect -22567 -10882 -21931 -10876
rect -22567 -10962 -22551 -10882
rect -22517 -10962 -22359 -10882
rect -22325 -10962 -22167 -10882
rect -22133 -10934 -21931 -10882
rect -21897 -10934 -21881 -10708
rect -21850 -10694 -21844 -10660
rect -21765 -10664 -21636 -10660
rect -21765 -10694 -21759 -10664
rect -21850 -10852 -21759 -10694
rect -21850 -10886 -21844 -10852
rect -21765 -10886 -21759 -10852
rect -21850 -10902 -21759 -10886
rect -21727 -10756 -21538 -10692
rect -21727 -10790 -21721 -10756
rect -21644 -10790 -21538 -10756
rect -22133 -10962 -21881 -10934
rect -21727 -10948 -21538 -10790
rect -22567 -10968 -21881 -10962
rect -22892 -11015 -22531 -10997
rect -22892 -11019 -22581 -11015
rect -22892 -11113 -22832 -11019
rect -22650 -11050 -22581 -11019
rect -22547 -11050 -22531 -11015
rect -22650 -11113 -22531 -11050
rect -22892 -11131 -22531 -11113
rect -22695 -11132 -22531 -11131
rect -22503 -11015 -22243 -10996
rect -22503 -11050 -22292 -11015
rect -22258 -11050 -22243 -11015
rect -22503 -11070 -22243 -11050
rect -22503 -11139 -22453 -11070
rect -22167 -11098 -21881 -10968
rect -22503 -11161 -22497 -11139
rect -22892 -11174 -22497 -11161
rect -22463 -11174 -22453 -11139
rect -22425 -11110 -21881 -11098
rect -22425 -11144 -22413 -11110
rect -22037 -11144 -21881 -11110
rect -22425 -11150 -21881 -11144
rect -21850 -10982 -21721 -10948
rect -21644 -10982 -21538 -10948
rect -21850 -11058 -21538 -10982
rect -21259 -11058 -21128 -10215
rect -17756 -10292 -17647 -10215
rect -20649 -10356 -19439 -10328
rect -20649 -10428 -20603 -10356
rect -19481 -10428 -19439 -10356
rect -20649 -10462 -19439 -10428
rect -20649 -10531 -20395 -10462
rect -20649 -10633 -20637 -10531
rect -20603 -10633 -20445 -10531
rect -20411 -10633 -20395 -10531
rect -20649 -10654 -20395 -10633
rect -20269 -10533 -19819 -10507
rect -20269 -10635 -20253 -10533
rect -20219 -10534 -19819 -10533
rect -20219 -10635 -20061 -10534
rect -20269 -10636 -20061 -10635
rect -20027 -10636 -19869 -10534
rect -19835 -10636 -19819 -10534
rect -20269 -10654 -19819 -10636
rect -19693 -10534 -19439 -10462
rect -19693 -10636 -19677 -10534
rect -19643 -10636 -19485 -10534
rect -19451 -10636 -19439 -10534
rect -19693 -10654 -19439 -10636
rect -19090 -10356 -17880 -10328
rect -19090 -10428 -19044 -10356
rect -17922 -10428 -17880 -10356
rect -17756 -10387 -17744 -10292
rect -17655 -10387 -17647 -10292
rect -14466 -10291 -14356 -10067
rect -17756 -10398 -17647 -10387
rect -17358 -10356 -16148 -10328
rect -19090 -10462 -17880 -10428
rect -19090 -10531 -18836 -10462
rect -19090 -10633 -19078 -10531
rect -19044 -10633 -18886 -10531
rect -18852 -10633 -18836 -10531
rect -19090 -10654 -18836 -10633
rect -18710 -10533 -18260 -10507
rect -18710 -10635 -18694 -10533
rect -18660 -10534 -18260 -10533
rect -18660 -10635 -18502 -10534
rect -18710 -10636 -18502 -10635
rect -18468 -10636 -18310 -10534
rect -18276 -10636 -18260 -10534
rect -18710 -10654 -18260 -10636
rect -18134 -10534 -17880 -10462
rect -18134 -10636 -18118 -10534
rect -18084 -10636 -17926 -10534
rect -17892 -10636 -17880 -10534
rect -18134 -10654 -17880 -10636
rect -17358 -10428 -17312 -10356
rect -16190 -10428 -16148 -10356
rect -17358 -10462 -16148 -10428
rect -17358 -10531 -17104 -10462
rect -17358 -10633 -17346 -10531
rect -17312 -10633 -17154 -10531
rect -17120 -10633 -17104 -10531
rect -17358 -10654 -17104 -10633
rect -16978 -10533 -16528 -10507
rect -16978 -10635 -16962 -10533
rect -16928 -10534 -16528 -10533
rect -16928 -10635 -16770 -10534
rect -16978 -10636 -16770 -10635
rect -16736 -10636 -16578 -10534
rect -16544 -10636 -16528 -10534
rect -16978 -10654 -16528 -10636
rect -16402 -10534 -16148 -10462
rect -16402 -10636 -16386 -10534
rect -16352 -10636 -16194 -10534
rect -16160 -10636 -16148 -10534
rect -16402 -10654 -16148 -10636
rect -15799 -10356 -14589 -10328
rect -15799 -10428 -15753 -10356
rect -14631 -10428 -14589 -10356
rect -15799 -10462 -14589 -10428
rect -15799 -10531 -15545 -10462
rect -15799 -10633 -15787 -10531
rect -15753 -10633 -15595 -10531
rect -15561 -10633 -15545 -10531
rect -15799 -10654 -15545 -10633
rect -15419 -10533 -14969 -10507
rect -15419 -10635 -15403 -10533
rect -15369 -10534 -14969 -10533
rect -15369 -10635 -15211 -10534
rect -15419 -10636 -15211 -10635
rect -15177 -10636 -15019 -10534
rect -14985 -10636 -14969 -10534
rect -15419 -10654 -14969 -10636
rect -14843 -10534 -14589 -10462
rect -14466 -10475 -14460 -10291
rect -14361 -10475 -14356 -10291
rect -11174 -10290 -11066 -9920
rect -14466 -10482 -14356 -10475
rect -14067 -10356 -12857 -10328
rect -14067 -10428 -14021 -10356
rect -12899 -10428 -12857 -10356
rect -14067 -10462 -12857 -10428
rect -14843 -10636 -14827 -10534
rect -14793 -10636 -14635 -10534
rect -14601 -10636 -14589 -10534
rect -14843 -10654 -14589 -10636
rect -14067 -10531 -13813 -10462
rect -14067 -10633 -14055 -10531
rect -14021 -10633 -13863 -10531
rect -13829 -10633 -13813 -10531
rect -14067 -10654 -13813 -10633
rect -13687 -10533 -13237 -10507
rect -13687 -10635 -13671 -10533
rect -13637 -10534 -13237 -10533
rect -13637 -10635 -13479 -10534
rect -13687 -10636 -13479 -10635
rect -13445 -10636 -13287 -10534
rect -13253 -10636 -13237 -10534
rect -13687 -10654 -13237 -10636
rect -13111 -10534 -12857 -10462
rect -13111 -10636 -13095 -10534
rect -13061 -10636 -12903 -10534
rect -12869 -10636 -12857 -10534
rect -13111 -10654 -12857 -10636
rect -12508 -10356 -11298 -10328
rect -12508 -10428 -12462 -10356
rect -11340 -10428 -11298 -10356
rect -12508 -10462 -11298 -10428
rect -11174 -10434 -11165 -10290
rect -11074 -10434 -11066 -10290
rect -11174 -10445 -11066 -10434
rect -10776 -10356 -9566 -10328
rect -10776 -10428 -10730 -10356
rect -9608 -10428 -9566 -10356
rect -12508 -10531 -12254 -10462
rect -12508 -10633 -12496 -10531
rect -12462 -10633 -12304 -10531
rect -12270 -10633 -12254 -10531
rect -12508 -10654 -12254 -10633
rect -12128 -10533 -11678 -10507
rect -12128 -10635 -12112 -10533
rect -12078 -10534 -11678 -10533
rect -12078 -10635 -11920 -10534
rect -12128 -10636 -11920 -10635
rect -11886 -10636 -11728 -10534
rect -11694 -10636 -11678 -10534
rect -12128 -10654 -11678 -10636
rect -11552 -10534 -11298 -10462
rect -11552 -10636 -11536 -10534
rect -11502 -10636 -11344 -10534
rect -11310 -10636 -11298 -10534
rect -11552 -10654 -11298 -10636
rect -10776 -10462 -9566 -10428
rect -10776 -10531 -10522 -10462
rect -10776 -10633 -10764 -10531
rect -10730 -10633 -10572 -10531
rect -10538 -10633 -10522 -10531
rect -10776 -10654 -10522 -10633
rect -10396 -10533 -9946 -10507
rect -10396 -10635 -10380 -10533
rect -10346 -10534 -9946 -10533
rect -10346 -10635 -10188 -10534
rect -10396 -10636 -10188 -10635
rect -10154 -10636 -9996 -10534
rect -9962 -10636 -9946 -10534
rect -10396 -10654 -9946 -10636
rect -9820 -10534 -9566 -10462
rect -9820 -10636 -9804 -10534
rect -9770 -10636 -9612 -10534
rect -9578 -10636 -9566 -10534
rect -9820 -10654 -9566 -10636
rect -9217 -10356 -8007 -10328
rect -9217 -10428 -9171 -10356
rect -8049 -10428 -8007 -10356
rect -9217 -10462 -8007 -10428
rect -9217 -10531 -8963 -10462
rect -9217 -10633 -9205 -10531
rect -9171 -10633 -9013 -10531
rect -8979 -10633 -8963 -10531
rect -9217 -10654 -8963 -10633
rect -8837 -10533 -8387 -10507
rect -8837 -10635 -8821 -10533
rect -8787 -10534 -8387 -10533
rect -8787 -10635 -8629 -10534
rect -8837 -10636 -8629 -10635
rect -8595 -10636 -8437 -10534
rect -8403 -10636 -8387 -10534
rect -8837 -10654 -8387 -10636
rect -8261 -10534 -8007 -10462
rect -8261 -10636 -8245 -10534
rect -8211 -10636 -8053 -10534
rect -8019 -10636 -8007 -10534
rect -8261 -10654 -8007 -10636
rect -20557 -10717 -19531 -10692
rect -20557 -10841 -20541 -10717
rect -20507 -10841 -20349 -10717
rect -20315 -10841 -20157 -10717
rect -20123 -10841 -19965 -10717
rect -19931 -10841 -19773 -10717
rect -19739 -10718 -19531 -10717
rect -19739 -10841 -19581 -10718
rect -20557 -10842 -19581 -10841
rect -19547 -10842 -19531 -10718
rect -20557 -10871 -19531 -10842
rect -18998 -10717 -17972 -10692
rect -18998 -10841 -18982 -10717
rect -18948 -10841 -18790 -10717
rect -18756 -10841 -18598 -10717
rect -18564 -10841 -18406 -10717
rect -18372 -10841 -18214 -10717
rect -18180 -10718 -17972 -10717
rect -18180 -10841 -18022 -10718
rect -18998 -10842 -18022 -10841
rect -17988 -10842 -17972 -10718
rect -18998 -10871 -17972 -10842
rect -17266 -10717 -16240 -10692
rect -17266 -10841 -17250 -10717
rect -17216 -10841 -17058 -10717
rect -17024 -10841 -16866 -10717
rect -16832 -10841 -16674 -10717
rect -16640 -10841 -16482 -10717
rect -16448 -10718 -16240 -10717
rect -16448 -10841 -16290 -10718
rect -17266 -10842 -16290 -10841
rect -16256 -10842 -16240 -10718
rect -17266 -10871 -16240 -10842
rect -15707 -10717 -14681 -10692
rect -15707 -10841 -15691 -10717
rect -15657 -10841 -15499 -10717
rect -15465 -10841 -15307 -10717
rect -15273 -10841 -15115 -10717
rect -15081 -10841 -14923 -10717
rect -14889 -10718 -14681 -10717
rect -14889 -10841 -14731 -10718
rect -15707 -10842 -14731 -10841
rect -14697 -10842 -14681 -10718
rect -15707 -10871 -14681 -10842
rect -13975 -10717 -12949 -10692
rect -13975 -10841 -13959 -10717
rect -13925 -10841 -13767 -10717
rect -13733 -10841 -13575 -10717
rect -13541 -10841 -13383 -10717
rect -13349 -10841 -13191 -10717
rect -13157 -10718 -12949 -10717
rect -13157 -10841 -12999 -10718
rect -13975 -10842 -12999 -10841
rect -12965 -10842 -12949 -10718
rect -13975 -10871 -12949 -10842
rect -12416 -10717 -11390 -10692
rect -12416 -10841 -12400 -10717
rect -12366 -10841 -12208 -10717
rect -12174 -10841 -12016 -10717
rect -11982 -10841 -11824 -10717
rect -11790 -10841 -11632 -10717
rect -11598 -10718 -11390 -10717
rect -11598 -10841 -11440 -10718
rect -12416 -10842 -11440 -10841
rect -11406 -10842 -11390 -10718
rect -12416 -10871 -11390 -10842
rect -10684 -10717 -9658 -10692
rect -10684 -10841 -10668 -10717
rect -10634 -10841 -10476 -10717
rect -10442 -10841 -10284 -10717
rect -10250 -10841 -10092 -10717
rect -10058 -10841 -9900 -10717
rect -9866 -10718 -9658 -10717
rect -9866 -10841 -9708 -10718
rect -10684 -10842 -9708 -10841
rect -9674 -10842 -9658 -10718
rect -10684 -10871 -9658 -10842
rect -9125 -10717 -8099 -10692
rect -9125 -10841 -9109 -10717
rect -9075 -10841 -8917 -10717
rect -8883 -10841 -8725 -10717
rect -8691 -10841 -8533 -10717
rect -8499 -10841 -8341 -10717
rect -8307 -10718 -8099 -10717
rect -8307 -10841 -8149 -10718
rect -9125 -10842 -8149 -10841
rect -8115 -10842 -8099 -10718
rect -9125 -10871 -8099 -10842
rect -20649 -10926 -20395 -10904
rect -20649 -11028 -20637 -10926
rect -20603 -10992 -20445 -10926
rect -20411 -10992 -20395 -10926
rect -20603 -11028 -20395 -10992
rect -20269 -10932 -19819 -10915
rect -20269 -10992 -20253 -10932
rect -20219 -10949 -19869 -10932
rect -20219 -10992 -20061 -10949
rect -20027 -10992 -19869 -10949
rect -19835 -10992 -19819 -10932
rect -20269 -11007 -19819 -10992
rect -19693 -10925 -19439 -10904
rect -19693 -10992 -19677 -10925
rect -19643 -10992 -19485 -10925
rect -19451 -10992 -19439 -10925
rect -20649 -11051 -20395 -11028
rect -19693 -11051 -19439 -10992
rect -19090 -10926 -18836 -10904
rect -19090 -11028 -19078 -10926
rect -19044 -10992 -18886 -10926
rect -18852 -10992 -18836 -10926
rect -19044 -11028 -18836 -10992
rect -18710 -10932 -18260 -10915
rect -18710 -10992 -18694 -10932
rect -18660 -10949 -18310 -10932
rect -18660 -10992 -18502 -10949
rect -18468 -10992 -18310 -10949
rect -18276 -10992 -18260 -10932
rect -18710 -11007 -18260 -10992
rect -18134 -10925 -17880 -10904
rect -18134 -10992 -18118 -10925
rect -18084 -10992 -17926 -10925
rect -17892 -10992 -17880 -10925
rect -19090 -11051 -18836 -11028
rect -18134 -11051 -17880 -10992
rect -17358 -10926 -17104 -10904
rect -17358 -11028 -17346 -10926
rect -17312 -10992 -17154 -10926
rect -17120 -10992 -17104 -10926
rect -17312 -11028 -17104 -10992
rect -16978 -10932 -16528 -10915
rect -16978 -10992 -16962 -10932
rect -16928 -10949 -16578 -10932
rect -16928 -10992 -16770 -10949
rect -16736 -10992 -16578 -10949
rect -16544 -10992 -16528 -10932
rect -16978 -11007 -16528 -10992
rect -16402 -10925 -16148 -10904
rect -16402 -10992 -16386 -10925
rect -16352 -10992 -16194 -10925
rect -16160 -10992 -16148 -10925
rect -17358 -11051 -17104 -11028
rect -16402 -11051 -16148 -10992
rect -15799 -10926 -15545 -10904
rect -15799 -11028 -15787 -10926
rect -15753 -10992 -15595 -10926
rect -15561 -10992 -15545 -10926
rect -15753 -11028 -15545 -10992
rect -15419 -10932 -14969 -10915
rect -15419 -10992 -15403 -10932
rect -15369 -10949 -15019 -10932
rect -15369 -10992 -15211 -10949
rect -15177 -10992 -15019 -10949
rect -14985 -10992 -14969 -10932
rect -15419 -11007 -14969 -10992
rect -14843 -10925 -14589 -10904
rect -14843 -10992 -14827 -10925
rect -14793 -10992 -14635 -10925
rect -14601 -10992 -14589 -10925
rect -15799 -11051 -15545 -11028
rect -14843 -11051 -14589 -10992
rect -14067 -10926 -13813 -10904
rect -14067 -11028 -14055 -10926
rect -14021 -10992 -13863 -10926
rect -13829 -10992 -13813 -10926
rect -14021 -11028 -13813 -10992
rect -13687 -10932 -13237 -10915
rect -13687 -10992 -13671 -10932
rect -13637 -10949 -13287 -10932
rect -13637 -10992 -13479 -10949
rect -13445 -10992 -13287 -10949
rect -13253 -10992 -13237 -10932
rect -13687 -11007 -13237 -10992
rect -13111 -10925 -12857 -10904
rect -13111 -10992 -13095 -10925
rect -13061 -10992 -12903 -10925
rect -12869 -10992 -12857 -10925
rect -14067 -11051 -13813 -11028
rect -13111 -11051 -12857 -10992
rect -12508 -10926 -12254 -10904
rect -12508 -11028 -12496 -10926
rect -12462 -10992 -12304 -10926
rect -12270 -10992 -12254 -10926
rect -12462 -11028 -12254 -10992
rect -12128 -10932 -11678 -10915
rect -12128 -10992 -12112 -10932
rect -12078 -10949 -11728 -10932
rect -12078 -10992 -11920 -10949
rect -11886 -10992 -11728 -10949
rect -11694 -10992 -11678 -10932
rect -12128 -11007 -11678 -10992
rect -11552 -10925 -11298 -10904
rect -11552 -10992 -11536 -10925
rect -11502 -10992 -11344 -10925
rect -11310 -10992 -11298 -10925
rect -12508 -11051 -12254 -11028
rect -11552 -11051 -11298 -10992
rect -10776 -10926 -10522 -10904
rect -10776 -11028 -10764 -10926
rect -10730 -10992 -10572 -10926
rect -10538 -10992 -10522 -10926
rect -10730 -11028 -10522 -10992
rect -10396 -10932 -9946 -10915
rect -10396 -10992 -10380 -10932
rect -10346 -10949 -9996 -10932
rect -10346 -10992 -10188 -10949
rect -10154 -10992 -9996 -10949
rect -9962 -10992 -9946 -10932
rect -10396 -11007 -9946 -10992
rect -9820 -10925 -9566 -10904
rect -9820 -10992 -9804 -10925
rect -9770 -10992 -9612 -10925
rect -9578 -10992 -9566 -10925
rect -10776 -11051 -10522 -11028
rect -9820 -11051 -9566 -10992
rect -9217 -10926 -8963 -10904
rect -9217 -11028 -9205 -10926
rect -9171 -10992 -9013 -10926
rect -8979 -10992 -8963 -10926
rect -9171 -11028 -8963 -10992
rect -8837 -10932 -8387 -10915
rect -8837 -10992 -8821 -10932
rect -8787 -10949 -8437 -10932
rect -8787 -10992 -8629 -10949
rect -8595 -10992 -8437 -10949
rect -8403 -10992 -8387 -10932
rect -8837 -11007 -8387 -10992
rect -8261 -10925 -8007 -10904
rect -8261 -10992 -8245 -10925
rect -8211 -10992 -8053 -10925
rect -8019 -10992 -8007 -10925
rect -9217 -11051 -8963 -11028
rect -8261 -11051 -8007 -10992
rect -21850 -11110 -21128 -11058
rect -21850 -11144 -21838 -11110
rect -21662 -11144 -21128 -11110
rect -21850 -11150 -21650 -11144
rect -22892 -11179 -22453 -11174
rect -22892 -11275 -22848 -11179
rect -22644 -11275 -22453 -11179
rect -21950 -11154 -21881 -11150
rect -21950 -11188 -21931 -11154
rect -21897 -11188 -21881 -11154
rect -21950 -11205 -21881 -11188
rect -21850 -11198 -21650 -11191
rect -22892 -11297 -22453 -11275
rect -21850 -11232 -21838 -11198
rect -21662 -11232 -21650 -11198
rect -21622 -11205 -21128 -11144
rect -20872 -11151 -20737 -11127
rect -22425 -11302 -22025 -11296
rect -22425 -11336 -22413 -11302
rect -22037 -11336 -22025 -11302
rect -22425 -11374 -22396 -11336
rect -22425 -11408 -22398 -11374
rect -22056 -11398 -22025 -11336
rect -21850 -11315 -21823 -11232
rect -21674 -11315 -21650 -11232
rect -20872 -11261 -20854 -11151
rect -20758 -11259 -20737 -11151
rect -17581 -11151 -17446 -11127
rect -19398 -11186 -19207 -11181
rect -19399 -11196 -19207 -11186
rect -19399 -11203 -19297 -11196
rect -19224 -11203 -19207 -11196
rect -20807 -11261 -20737 -11259
rect -20872 -11281 -20737 -11261
rect -20576 -11244 -19787 -11226
rect -20576 -11252 -19933 -11244
rect -21850 -11334 -21819 -11315
rect -21687 -11334 -21650 -11315
rect -20576 -11305 -20539 -11252
rect -20406 -11297 -19933 -11252
rect -19819 -11297 -19787 -11244
rect -20406 -11305 -19787 -11297
rect -20576 -11325 -19787 -11305
rect -19717 -11245 -19602 -11226
rect -19717 -11313 -19699 -11245
rect -19619 -11313 -19602 -11245
rect -19399 -11286 -19372 -11203
rect -21850 -11341 -21650 -11334
rect -22063 -11408 -22025 -11398
rect -22425 -11419 -22025 -11408
rect -20795 -11384 -20590 -11365
rect -20795 -11492 -20751 -11384
rect -20675 -11410 -20590 -11384
rect -19717 -11410 -19602 -11313
rect -19486 -11300 -19372 -11286
rect -19222 -11300 -19207 -11203
rect -19486 -11316 -19207 -11300
rect -19017 -11244 -18228 -11226
rect -19017 -11252 -18374 -11244
rect -19017 -11305 -18980 -11252
rect -18847 -11297 -18374 -11252
rect -18260 -11297 -18228 -11244
rect -18847 -11305 -18228 -11297
rect -19486 -11379 -19315 -11316
rect -19017 -11325 -18228 -11305
rect -18158 -11245 -18043 -11226
rect -18158 -11313 -18140 -11245
rect -18060 -11313 -18043 -11245
rect -17581 -11261 -17563 -11151
rect -17467 -11259 -17446 -11151
rect -14290 -11151 -14155 -11127
rect -16107 -11186 -15916 -11181
rect -16108 -11196 -15916 -11186
rect -16108 -11203 -16006 -11196
rect -15933 -11203 -15916 -11196
rect -17516 -11261 -17446 -11259
rect -17581 -11281 -17446 -11261
rect -17285 -11244 -16496 -11226
rect -17285 -11252 -16642 -11244
rect -20675 -11492 -19602 -11410
rect -20795 -11496 -19602 -11492
rect -19528 -11416 -19315 -11379
rect -19528 -11471 -19517 -11416
rect -19452 -11471 -19315 -11416
rect -19528 -11495 -19315 -11471
rect -19236 -11391 -19031 -11365
rect -19236 -11488 -19196 -11391
rect -19080 -11410 -19031 -11391
rect -18158 -11410 -18043 -11313
rect -17927 -11379 -17647 -11286
rect -17285 -11305 -17248 -11252
rect -17115 -11297 -16642 -11252
rect -16528 -11297 -16496 -11244
rect -17115 -11305 -16496 -11297
rect -17285 -11325 -16496 -11305
rect -16426 -11245 -16311 -11226
rect -16426 -11313 -16408 -11245
rect -16328 -11313 -16311 -11245
rect -16108 -11286 -16081 -11203
rect -19080 -11488 -18043 -11410
rect -19236 -11496 -18043 -11488
rect -17969 -11416 -17647 -11379
rect -17969 -11471 -17958 -11416
rect -17893 -11471 -17647 -11416
rect -17969 -11495 -17647 -11471
rect -20795 -11508 -20590 -11496
rect -19236 -11508 -19031 -11496
rect -20644 -11565 -20589 -11549
rect -20644 -11671 -20637 -11565
rect -20603 -11671 -20589 -11565
rect -20557 -11550 -20107 -11538
rect -20557 -11584 -20541 -11550
rect -20507 -11584 -20349 -11550
rect -20315 -11551 -20107 -11550
rect -20315 -11584 -20157 -11551
rect -20557 -11585 -20157 -11584
rect -20123 -11585 -20107 -11551
rect -20557 -11606 -20107 -11585
rect -19981 -11550 -19531 -11538
rect -19981 -11584 -19965 -11550
rect -19931 -11584 -19773 -11550
rect -19739 -11584 -19581 -11550
rect -19547 -11584 -19531 -11550
rect -19981 -11606 -19531 -11584
rect -19497 -11565 -19442 -11549
rect -20644 -11737 -20589 -11671
rect -20459 -11651 -20394 -11634
rect -20459 -11685 -20445 -11651
rect -20411 -11685 -20394 -11651
rect -20459 -11737 -20394 -11685
rect -20266 -11651 -19819 -11639
rect -20266 -11685 -20253 -11651
rect -20219 -11685 -20061 -11651
rect -20027 -11685 -19869 -11651
rect -19835 -11685 -19819 -11651
rect -20266 -11703 -19819 -11685
rect -19693 -11651 -19628 -11635
rect -19693 -11685 -19677 -11651
rect -19643 -11685 -19628 -11651
rect -19693 -11737 -19628 -11685
rect -19497 -11671 -19485 -11565
rect -19451 -11671 -19442 -11565
rect -19497 -11737 -19442 -11671
rect -20644 -11748 -19442 -11737
rect -20644 -11759 -20143 -11748
rect -20083 -11759 -19442 -11748
rect -20644 -11805 -20603 -11759
rect -19480 -11805 -19442 -11759
rect -20644 -11808 -20143 -11805
rect -20083 -11808 -19442 -11805
rect -20644 -11828 -19442 -11808
rect -19085 -11565 -19030 -11549
rect -19085 -11671 -19078 -11565
rect -19044 -11671 -19030 -11565
rect -18998 -11550 -18548 -11538
rect -18998 -11584 -18982 -11550
rect -18948 -11584 -18790 -11550
rect -18756 -11551 -18548 -11550
rect -18756 -11584 -18598 -11551
rect -18998 -11585 -18598 -11584
rect -18564 -11585 -18548 -11551
rect -18998 -11606 -18548 -11585
rect -18422 -11550 -17972 -11538
rect -18422 -11584 -18406 -11550
rect -18372 -11584 -18214 -11550
rect -18180 -11584 -18022 -11550
rect -17988 -11584 -17972 -11550
rect -18422 -11606 -17972 -11584
rect -17938 -11565 -17883 -11549
rect -19085 -11737 -19030 -11671
rect -18900 -11651 -18835 -11634
rect -18900 -11685 -18886 -11651
rect -18852 -11685 -18835 -11651
rect -18900 -11737 -18835 -11685
rect -18707 -11651 -18260 -11639
rect -18707 -11685 -18694 -11651
rect -18660 -11685 -18502 -11651
rect -18468 -11685 -18310 -11651
rect -18276 -11685 -18260 -11651
rect -18707 -11703 -18260 -11685
rect -18134 -11651 -18069 -11635
rect -18134 -11685 -18118 -11651
rect -18084 -11685 -18069 -11651
rect -18134 -11737 -18069 -11685
rect -17938 -11671 -17926 -11565
rect -17892 -11671 -17883 -11565
rect -17938 -11737 -17883 -11671
rect -19085 -11748 -17883 -11737
rect -19085 -11759 -18584 -11748
rect -18524 -11759 -17883 -11748
rect -19085 -11805 -19044 -11759
rect -17921 -11805 -17883 -11759
rect -17756 -11682 -17647 -11495
rect -17504 -11384 -17299 -11365
rect -17504 -11492 -17460 -11384
rect -17384 -11410 -17299 -11384
rect -16426 -11410 -16311 -11313
rect -16195 -11300 -16081 -11286
rect -15931 -11300 -15916 -11203
rect -16195 -11316 -15916 -11300
rect -15726 -11244 -14937 -11226
rect -15726 -11252 -15083 -11244
rect -15726 -11305 -15689 -11252
rect -15556 -11297 -15083 -11252
rect -14969 -11297 -14937 -11244
rect -15556 -11305 -14937 -11297
rect -16195 -11379 -16024 -11316
rect -15726 -11325 -14937 -11305
rect -14867 -11245 -14752 -11226
rect -14867 -11313 -14849 -11245
rect -14769 -11313 -14752 -11245
rect -14290 -11261 -14272 -11151
rect -14176 -11259 -14155 -11151
rect -10999 -11151 -10864 -11127
rect -12816 -11186 -12625 -11181
rect -12817 -11196 -12625 -11186
rect -12817 -11203 -12715 -11196
rect -12642 -11203 -12625 -11196
rect -14225 -11261 -14155 -11259
rect -14290 -11281 -14155 -11261
rect -13994 -11244 -13205 -11226
rect -13994 -11252 -13351 -11244
rect -17384 -11492 -16311 -11410
rect -17504 -11496 -16311 -11492
rect -16237 -11416 -16024 -11379
rect -16237 -11471 -16226 -11416
rect -16161 -11471 -16024 -11416
rect -16237 -11495 -16024 -11471
rect -15945 -11391 -15740 -11365
rect -15945 -11488 -15905 -11391
rect -15789 -11410 -15740 -11391
rect -14867 -11410 -14752 -11313
rect -14636 -11379 -14356 -11286
rect -13994 -11305 -13957 -11252
rect -13824 -11297 -13351 -11252
rect -13237 -11297 -13205 -11244
rect -13824 -11305 -13205 -11297
rect -13994 -11325 -13205 -11305
rect -13135 -11245 -13020 -11226
rect -13135 -11313 -13117 -11245
rect -13037 -11313 -13020 -11245
rect -12817 -11286 -12790 -11203
rect -15789 -11488 -14752 -11410
rect -15945 -11496 -14752 -11488
rect -14678 -11416 -14356 -11379
rect -14678 -11471 -14667 -11416
rect -14602 -11471 -14356 -11416
rect -14678 -11495 -14356 -11471
rect -17504 -11508 -17299 -11496
rect -15945 -11508 -15740 -11496
rect -17756 -11768 -17747 -11682
rect -17656 -11768 -17647 -11682
rect -17756 -11780 -17647 -11768
rect -17353 -11565 -17298 -11549
rect -17353 -11671 -17346 -11565
rect -17312 -11671 -17298 -11565
rect -17266 -11550 -16816 -11538
rect -17266 -11584 -17250 -11550
rect -17216 -11584 -17058 -11550
rect -17024 -11551 -16816 -11550
rect -17024 -11584 -16866 -11551
rect -17266 -11585 -16866 -11584
rect -16832 -11585 -16816 -11551
rect -17266 -11606 -16816 -11585
rect -16690 -11550 -16240 -11538
rect -16690 -11584 -16674 -11550
rect -16640 -11584 -16482 -11550
rect -16448 -11584 -16290 -11550
rect -16256 -11584 -16240 -11550
rect -16690 -11606 -16240 -11584
rect -16206 -11565 -16151 -11549
rect -17353 -11737 -17298 -11671
rect -17168 -11651 -17103 -11634
rect -17168 -11685 -17154 -11651
rect -17120 -11685 -17103 -11651
rect -17168 -11737 -17103 -11685
rect -16975 -11651 -16528 -11639
rect -16975 -11685 -16962 -11651
rect -16928 -11685 -16770 -11651
rect -16736 -11685 -16578 -11651
rect -16544 -11685 -16528 -11651
rect -16975 -11703 -16528 -11685
rect -16402 -11651 -16337 -11635
rect -16402 -11685 -16386 -11651
rect -16352 -11685 -16337 -11651
rect -16402 -11737 -16337 -11685
rect -16206 -11671 -16194 -11565
rect -16160 -11671 -16151 -11565
rect -16206 -11737 -16151 -11671
rect -17353 -11748 -16151 -11737
rect -17353 -11759 -16852 -11748
rect -16792 -11759 -16151 -11748
rect -19085 -11808 -18584 -11805
rect -18524 -11808 -17883 -11805
rect -19085 -11828 -17883 -11808
rect -17353 -11805 -17312 -11759
rect -16189 -11805 -16151 -11759
rect -17353 -11808 -16852 -11805
rect -16792 -11808 -16151 -11805
rect -17353 -11828 -16151 -11808
rect -15794 -11565 -15739 -11549
rect -15794 -11671 -15787 -11565
rect -15753 -11671 -15739 -11565
rect -15707 -11550 -15257 -11538
rect -15707 -11584 -15691 -11550
rect -15657 -11584 -15499 -11550
rect -15465 -11551 -15257 -11550
rect -15465 -11584 -15307 -11551
rect -15707 -11585 -15307 -11584
rect -15273 -11585 -15257 -11551
rect -15707 -11606 -15257 -11585
rect -15131 -11550 -14681 -11538
rect -15131 -11584 -15115 -11550
rect -15081 -11584 -14923 -11550
rect -14889 -11584 -14731 -11550
rect -14697 -11584 -14681 -11550
rect -15131 -11606 -14681 -11584
rect -14647 -11565 -14592 -11549
rect -15794 -11737 -15739 -11671
rect -15609 -11651 -15544 -11634
rect -15609 -11685 -15595 -11651
rect -15561 -11685 -15544 -11651
rect -15609 -11737 -15544 -11685
rect -15416 -11651 -14969 -11639
rect -15416 -11685 -15403 -11651
rect -15369 -11685 -15211 -11651
rect -15177 -11685 -15019 -11651
rect -14985 -11685 -14969 -11651
rect -15416 -11703 -14969 -11685
rect -14843 -11651 -14778 -11635
rect -14843 -11685 -14827 -11651
rect -14793 -11685 -14778 -11651
rect -14843 -11737 -14778 -11685
rect -14647 -11671 -14635 -11565
rect -14601 -11671 -14592 -11565
rect -14647 -11737 -14592 -11671
rect -15794 -11748 -14592 -11737
rect -15794 -11759 -15293 -11748
rect -15233 -11759 -14592 -11748
rect -15794 -11805 -15753 -11759
rect -14630 -11805 -14592 -11759
rect -14465 -11682 -14356 -11495
rect -14213 -11384 -14008 -11365
rect -14213 -11492 -14169 -11384
rect -14093 -11410 -14008 -11384
rect -13135 -11410 -13020 -11313
rect -12904 -11300 -12790 -11286
rect -12640 -11300 -12625 -11203
rect -12904 -11316 -12625 -11300
rect -12435 -11244 -11646 -11226
rect -12435 -11252 -11792 -11244
rect -12435 -11305 -12398 -11252
rect -12265 -11297 -11792 -11252
rect -11678 -11297 -11646 -11244
rect -12265 -11305 -11646 -11297
rect -12904 -11379 -12733 -11316
rect -12435 -11325 -11646 -11305
rect -11576 -11245 -11461 -11226
rect -11576 -11313 -11558 -11245
rect -11478 -11313 -11461 -11245
rect -10999 -11261 -10981 -11151
rect -10885 -11259 -10864 -11151
rect -5043 -11161 -4977 -8271
rect -9525 -11186 -9334 -11181
rect -9526 -11196 -9334 -11186
rect -9526 -11203 -9424 -11196
rect -9351 -11203 -9334 -11196
rect -10934 -11261 -10864 -11259
rect -10999 -11281 -10864 -11261
rect -10703 -11244 -9914 -11226
rect -10703 -11252 -10060 -11244
rect -14093 -11492 -13020 -11410
rect -14213 -11496 -13020 -11492
rect -12946 -11416 -12733 -11379
rect -12946 -11471 -12935 -11416
rect -12870 -11471 -12733 -11416
rect -12946 -11495 -12733 -11471
rect -12654 -11391 -12449 -11365
rect -12654 -11488 -12614 -11391
rect -12498 -11410 -12449 -11391
rect -11576 -11410 -11461 -11313
rect -11345 -11379 -11065 -11286
rect -10703 -11305 -10666 -11252
rect -10533 -11297 -10060 -11252
rect -9946 -11297 -9914 -11244
rect -10533 -11305 -9914 -11297
rect -10703 -11325 -9914 -11305
rect -9844 -11245 -9729 -11226
rect -9844 -11313 -9826 -11245
rect -9746 -11313 -9729 -11245
rect -9526 -11286 -9499 -11203
rect -12498 -11488 -11461 -11410
rect -12654 -11496 -11461 -11488
rect -11387 -11416 -11065 -11379
rect -11387 -11471 -11376 -11416
rect -11311 -11471 -11065 -11416
rect -11387 -11495 -11065 -11471
rect -14213 -11508 -14008 -11496
rect -12654 -11508 -12449 -11496
rect -14465 -11768 -14456 -11682
rect -14365 -11768 -14356 -11682
rect -14465 -11780 -14356 -11768
rect -14062 -11565 -14007 -11549
rect -14062 -11671 -14055 -11565
rect -14021 -11671 -14007 -11565
rect -13975 -11550 -13525 -11538
rect -13975 -11584 -13959 -11550
rect -13925 -11584 -13767 -11550
rect -13733 -11551 -13525 -11550
rect -13733 -11584 -13575 -11551
rect -13975 -11585 -13575 -11584
rect -13541 -11585 -13525 -11551
rect -13975 -11606 -13525 -11585
rect -13399 -11550 -12949 -11538
rect -13399 -11584 -13383 -11550
rect -13349 -11584 -13191 -11550
rect -13157 -11584 -12999 -11550
rect -12965 -11584 -12949 -11550
rect -13399 -11606 -12949 -11584
rect -12915 -11565 -12860 -11549
rect -14062 -11737 -14007 -11671
rect -13877 -11651 -13812 -11634
rect -13877 -11685 -13863 -11651
rect -13829 -11685 -13812 -11651
rect -13877 -11737 -13812 -11685
rect -13684 -11651 -13237 -11639
rect -13684 -11685 -13671 -11651
rect -13637 -11685 -13479 -11651
rect -13445 -11685 -13287 -11651
rect -13253 -11685 -13237 -11651
rect -13684 -11703 -13237 -11685
rect -13111 -11651 -13046 -11635
rect -13111 -11685 -13095 -11651
rect -13061 -11685 -13046 -11651
rect -13111 -11737 -13046 -11685
rect -12915 -11671 -12903 -11565
rect -12869 -11671 -12860 -11565
rect -12915 -11737 -12860 -11671
rect -14062 -11748 -12860 -11737
rect -14062 -11759 -13561 -11748
rect -13501 -11759 -12860 -11748
rect -15794 -11808 -15293 -11805
rect -15233 -11808 -14592 -11805
rect -15794 -11828 -14592 -11808
rect -14062 -11805 -14021 -11759
rect -12898 -11805 -12860 -11759
rect -14062 -11808 -13561 -11805
rect -13501 -11808 -12860 -11805
rect -14062 -11828 -12860 -11808
rect -12503 -11565 -12448 -11549
rect -12503 -11671 -12496 -11565
rect -12462 -11671 -12448 -11565
rect -12416 -11550 -11966 -11538
rect -12416 -11584 -12400 -11550
rect -12366 -11584 -12208 -11550
rect -12174 -11551 -11966 -11550
rect -12174 -11584 -12016 -11551
rect -12416 -11585 -12016 -11584
rect -11982 -11585 -11966 -11551
rect -12416 -11606 -11966 -11585
rect -11840 -11550 -11390 -11538
rect -11840 -11584 -11824 -11550
rect -11790 -11584 -11632 -11550
rect -11598 -11584 -11440 -11550
rect -11406 -11584 -11390 -11550
rect -11840 -11606 -11390 -11584
rect -11356 -11565 -11301 -11549
rect -12503 -11737 -12448 -11671
rect -12318 -11651 -12253 -11634
rect -12318 -11685 -12304 -11651
rect -12270 -11685 -12253 -11651
rect -12318 -11737 -12253 -11685
rect -12125 -11651 -11678 -11639
rect -12125 -11685 -12112 -11651
rect -12078 -11685 -11920 -11651
rect -11886 -11685 -11728 -11651
rect -11694 -11685 -11678 -11651
rect -12125 -11703 -11678 -11685
rect -11552 -11651 -11487 -11635
rect -11552 -11685 -11536 -11651
rect -11502 -11685 -11487 -11651
rect -11552 -11737 -11487 -11685
rect -11356 -11671 -11344 -11565
rect -11310 -11671 -11301 -11565
rect -11356 -11737 -11301 -11671
rect -12503 -11748 -11301 -11737
rect -12503 -11759 -12002 -11748
rect -11942 -11759 -11301 -11748
rect -12503 -11805 -12462 -11759
rect -11339 -11805 -11301 -11759
rect -11174 -11682 -11065 -11495
rect -10922 -11384 -10717 -11365
rect -10922 -11492 -10878 -11384
rect -10802 -11410 -10717 -11384
rect -9844 -11410 -9729 -11313
rect -9613 -11300 -9499 -11286
rect -9349 -11300 -9334 -11203
rect -9613 -11316 -9334 -11300
rect -9144 -11244 -8355 -11226
rect -9144 -11252 -8501 -11244
rect -9144 -11305 -9107 -11252
rect -8974 -11297 -8501 -11252
rect -8387 -11297 -8355 -11244
rect -8974 -11305 -8355 -11297
rect -9613 -11379 -9442 -11316
rect -9144 -11325 -8355 -11305
rect -8285 -11245 -8170 -11226
rect -5043 -11233 -4977 -11227
rect -8285 -11313 -8267 -11245
rect -8187 -11313 -8170 -11245
rect -10802 -11492 -9729 -11410
rect -10922 -11496 -9729 -11492
rect -9655 -11416 -9442 -11379
rect -9655 -11471 -9644 -11416
rect -9579 -11471 -9442 -11416
rect -9655 -11495 -9442 -11471
rect -9363 -11391 -9158 -11365
rect -9363 -11488 -9323 -11391
rect -9207 -11410 -9158 -11391
rect -8285 -11410 -8170 -11313
rect -8054 -11379 -7774 -11286
rect -9207 -11488 -8170 -11410
rect -9363 -11496 -8170 -11488
rect -8096 -11416 -7774 -11379
rect -8096 -11471 -8085 -11416
rect -8020 -11471 -7774 -11416
rect -8096 -11495 -7774 -11471
rect -10922 -11508 -10717 -11496
rect -9363 -11508 -9158 -11496
rect -11174 -11768 -11165 -11682
rect -11074 -11768 -11065 -11682
rect -11174 -11780 -11065 -11768
rect -10771 -11565 -10716 -11549
rect -10771 -11671 -10764 -11565
rect -10730 -11671 -10716 -11565
rect -10684 -11550 -10234 -11538
rect -10684 -11584 -10668 -11550
rect -10634 -11584 -10476 -11550
rect -10442 -11551 -10234 -11550
rect -10442 -11584 -10284 -11551
rect -10684 -11585 -10284 -11584
rect -10250 -11585 -10234 -11551
rect -10684 -11606 -10234 -11585
rect -10108 -11550 -9658 -11538
rect -10108 -11584 -10092 -11550
rect -10058 -11584 -9900 -11550
rect -9866 -11584 -9708 -11550
rect -9674 -11584 -9658 -11550
rect -10108 -11606 -9658 -11584
rect -9624 -11565 -9569 -11549
rect -10771 -11737 -10716 -11671
rect -10586 -11651 -10521 -11634
rect -10586 -11685 -10572 -11651
rect -10538 -11685 -10521 -11651
rect -10586 -11737 -10521 -11685
rect -10393 -11651 -9946 -11639
rect -10393 -11685 -10380 -11651
rect -10346 -11685 -10188 -11651
rect -10154 -11685 -9996 -11651
rect -9962 -11685 -9946 -11651
rect -10393 -11703 -9946 -11685
rect -9820 -11651 -9755 -11635
rect -9820 -11685 -9804 -11651
rect -9770 -11685 -9755 -11651
rect -9820 -11737 -9755 -11685
rect -9624 -11671 -9612 -11565
rect -9578 -11671 -9569 -11565
rect -9624 -11737 -9569 -11671
rect -10771 -11748 -9569 -11737
rect -10771 -11759 -10270 -11748
rect -10210 -11759 -9569 -11748
rect -12503 -11808 -12002 -11805
rect -11942 -11808 -11301 -11805
rect -12503 -11828 -11301 -11808
rect -10771 -11805 -10730 -11759
rect -9607 -11805 -9569 -11759
rect -10771 -11808 -10270 -11805
rect -10210 -11808 -9569 -11805
rect -10771 -11828 -9569 -11808
rect -9212 -11565 -9157 -11549
rect -9212 -11671 -9205 -11565
rect -9171 -11671 -9157 -11565
rect -9125 -11550 -8675 -11538
rect -9125 -11584 -9109 -11550
rect -9075 -11584 -8917 -11550
rect -8883 -11551 -8675 -11550
rect -8883 -11584 -8725 -11551
rect -9125 -11585 -8725 -11584
rect -8691 -11585 -8675 -11551
rect -9125 -11606 -8675 -11585
rect -8549 -11550 -8099 -11538
rect -8549 -11584 -8533 -11550
rect -8499 -11584 -8341 -11550
rect -8307 -11584 -8149 -11550
rect -8115 -11584 -8099 -11550
rect -8549 -11606 -8099 -11584
rect -8065 -11565 -8010 -11549
rect -9212 -11737 -9157 -11671
rect -9027 -11651 -8962 -11634
rect -9027 -11685 -9013 -11651
rect -8979 -11685 -8962 -11651
rect -9027 -11737 -8962 -11685
rect -8834 -11651 -8387 -11639
rect -8834 -11685 -8821 -11651
rect -8787 -11685 -8629 -11651
rect -8595 -11685 -8437 -11651
rect -8403 -11685 -8387 -11651
rect -8834 -11703 -8387 -11685
rect -8261 -11651 -8196 -11635
rect -8261 -11685 -8245 -11651
rect -8211 -11685 -8196 -11651
rect -8261 -11736 -8196 -11685
rect -8065 -11671 -8053 -11565
rect -8019 -11671 -8010 -11565
rect -8261 -11737 -8114 -11736
rect -8065 -11737 -8010 -11671
rect -9212 -11748 -8010 -11737
rect -9212 -11759 -8711 -11748
rect -8651 -11759 -8010 -11748
rect -9212 -11805 -9171 -11759
rect -8048 -11805 -8010 -11759
rect -7883 -11682 -7774 -11495
rect -7883 -11768 -7874 -11682
rect -7783 -11723 -7774 -11682
rect -7783 -11768 473 -11723
rect -7883 -11780 473 -11768
rect -7881 -11789 473 -11780
rect -9212 -11808 -8711 -11805
rect -8651 -11808 -8010 -11805
rect -9212 -11828 -8010 -11808
rect -21854 -11858 -21640 -11836
rect -23460 -12048 -22951 -12014
rect -23460 -12082 -23454 -12048
rect -23377 -12082 -22951 -12048
rect -23870 -12254 -23614 -12226
rect -23460 -12240 -22951 -12082
rect -22660 -11933 -22026 -11926
rect -22660 -11980 -22631 -11933
rect -22062 -11980 -22026 -11933
rect -22660 -12052 -22622 -11980
rect -22068 -12046 -22026 -11980
rect -21854 -11937 -21831 -11858
rect -21662 -11937 -21640 -11858
rect -21854 -11952 -21640 -11937
rect -21954 -12000 -21885 -11984
rect -22068 -12052 -22025 -12046
rect -22660 -12132 -22647 -12052
rect -22613 -12132 -22455 -12100
rect -22421 -12132 -22263 -12100
rect -22229 -12132 -22071 -12100
rect -22037 -12132 -22025 -12052
rect -22660 -12138 -22025 -12132
rect -22660 -12139 -22026 -12138
rect -21954 -12168 -21935 -12000
rect -24304 -12260 -23614 -12254
rect -24632 -12307 -24268 -12289
rect -24632 -12313 -24318 -12307
rect -24632 -12400 -24570 -12313
rect -24353 -12342 -24318 -12313
rect -24284 -12342 -24268 -12307
rect -24353 -12400 -24268 -12342
rect -24632 -12424 -24268 -12400
rect -24240 -12307 -23980 -12288
rect -24240 -12342 -24029 -12307
rect -23995 -12342 -23980 -12307
rect -24240 -12362 -23980 -12342
rect -24240 -12431 -24190 -12362
rect -23904 -12390 -23614 -12260
rect -24240 -12453 -24234 -12431
rect -24637 -12466 -24234 -12453
rect -24200 -12466 -24190 -12431
rect -24162 -12402 -23614 -12390
rect -24162 -12436 -24150 -12402
rect -23774 -12436 -23614 -12402
rect -24162 -12442 -23614 -12436
rect -23583 -12274 -23454 -12240
rect -23377 -12274 -22951 -12240
rect -22567 -12174 -21935 -12168
rect -22567 -12254 -22551 -12174
rect -22517 -12254 -22359 -12174
rect -22325 -12254 -22167 -12174
rect -22133 -12226 -21935 -12174
rect -21901 -12226 -21885 -12000
rect -21854 -11986 -21848 -11952
rect -21769 -11956 -21640 -11952
rect -21033 -11862 -20824 -11842
rect -21769 -11986 -21763 -11956
rect -21033 -11964 -21003 -11862
rect -20885 -11881 -20824 -11862
rect -8205 -11881 -8114 -11828
rect -20885 -11897 -19620 -11881
rect -20885 -11964 -19735 -11897
rect -21033 -11966 -19735 -11964
rect -19636 -11966 -19620 -11897
rect -21033 -11972 -19620 -11966
rect -19237 -11893 -16329 -11881
rect -19237 -11959 -19223 -11893
rect -19152 -11897 -16329 -11893
rect -19152 -11959 -16444 -11897
rect -19237 -11966 -16444 -11959
rect -16345 -11966 -16329 -11897
rect -19237 -11972 -16329 -11966
rect -15946 -11893 -13038 -11881
rect -15946 -11959 -15932 -11893
rect -15861 -11897 -13038 -11893
rect -15861 -11959 -13153 -11897
rect -15946 -11966 -13153 -11959
rect -13054 -11966 -13038 -11897
rect -15946 -11972 -13038 -11966
rect -12655 -11893 -9747 -11881
rect -12655 -11959 -12641 -11893
rect -12570 -11897 -9747 -11893
rect -12570 -11959 -9862 -11897
rect -12655 -11966 -9862 -11959
rect -9763 -11966 -9747 -11897
rect -12655 -11972 -9747 -11966
rect -9364 -11893 -7684 -11881
rect -9364 -11959 -9350 -11893
rect -9279 -11959 -7684 -11893
rect -9364 -11972 -7684 -11959
rect -21854 -12144 -21763 -11986
rect -21854 -12178 -21848 -12144
rect -21769 -12178 -21763 -12144
rect -21854 -12194 -21763 -12178
rect -21731 -12048 -21542 -11984
rect -21033 -11994 -20824 -11972
rect -21731 -12082 -21725 -12048
rect -21648 -12082 -21542 -12048
rect -22133 -12254 -21885 -12226
rect -21731 -12234 -21542 -12082
rect -20354 -12088 -20080 -12079
rect -20354 -12094 -20345 -12088
rect -20531 -12101 -20345 -12094
rect -20089 -12094 -20080 -12088
rect -19065 -12088 -18791 -12079
rect -19065 -12094 -19056 -12088
rect -20089 -12101 -19897 -12094
rect -20531 -12148 -20502 -12101
rect -19933 -12148 -19897 -12101
rect -20531 -12160 -20345 -12148
rect -20089 -12160 -19897 -12148
rect -20531 -12214 -19897 -12160
rect -19422 -12101 -19056 -12094
rect -18800 -12094 -18791 -12088
rect -18348 -12088 -18074 -12079
rect -18348 -12094 -18339 -12088
rect -19422 -12148 -19393 -12101
rect -19422 -12160 -19056 -12148
rect -18800 -12160 -18788 -12094
rect -19422 -12214 -18788 -12160
rect -18540 -12101 -18339 -12094
rect -18083 -12094 -18074 -12088
rect -17063 -12088 -16789 -12079
rect -17063 -12094 -17054 -12088
rect -18083 -12101 -17906 -12094
rect -18540 -12148 -18511 -12101
rect -17942 -12148 -17906 -12101
rect -18540 -12160 -18339 -12148
rect -18083 -12160 -17906 -12148
rect -18540 -12214 -17906 -12160
rect -17240 -12101 -17054 -12094
rect -16798 -12094 -16789 -12088
rect -15774 -12088 -15500 -12079
rect -15774 -12094 -15765 -12088
rect -16798 -12101 -16606 -12094
rect -17240 -12148 -17211 -12101
rect -16642 -12148 -16606 -12101
rect -17240 -12160 -17054 -12148
rect -16798 -12160 -16606 -12148
rect -17240 -12214 -16606 -12160
rect -16131 -12101 -15765 -12094
rect -15509 -12094 -15500 -12088
rect -15057 -12088 -14783 -12079
rect -15057 -12094 -15048 -12088
rect -16131 -12148 -16102 -12101
rect -16131 -12160 -15765 -12148
rect -15509 -12160 -15497 -12094
rect -16131 -12214 -15497 -12160
rect -15249 -12101 -15048 -12094
rect -14792 -12094 -14783 -12088
rect -13772 -12088 -13498 -12079
rect -13772 -12094 -13763 -12088
rect -14792 -12101 -14615 -12094
rect -15249 -12148 -15220 -12101
rect -14651 -12148 -14615 -12101
rect -15249 -12160 -15048 -12148
rect -14792 -12160 -14615 -12148
rect -15249 -12214 -14615 -12160
rect -13949 -12101 -13763 -12094
rect -13507 -12094 -13498 -12088
rect -12483 -12088 -12209 -12079
rect -12483 -12094 -12474 -12088
rect -13507 -12101 -13315 -12094
rect -13949 -12148 -13920 -12101
rect -13351 -12148 -13315 -12101
rect -13949 -12160 -13763 -12148
rect -13507 -12160 -13315 -12148
rect -13949 -12214 -13315 -12160
rect -12840 -12101 -12474 -12094
rect -12218 -12094 -12209 -12088
rect -11766 -12088 -11492 -12079
rect -11766 -12094 -11757 -12088
rect -12840 -12148 -12811 -12101
rect -12840 -12160 -12474 -12148
rect -12218 -12160 -12206 -12094
rect -12840 -12214 -12206 -12160
rect -11958 -12101 -11757 -12094
rect -11501 -12094 -11492 -12088
rect -10481 -12088 -10207 -12079
rect -10481 -12094 -10472 -12088
rect -11501 -12101 -11324 -12094
rect -11958 -12148 -11929 -12101
rect -11360 -12148 -11324 -12101
rect -11958 -12160 -11757 -12148
rect -11501 -12160 -11324 -12148
rect -11958 -12214 -11324 -12160
rect -10658 -12101 -10472 -12094
rect -10216 -12094 -10207 -12088
rect -9192 -12088 -8918 -12079
rect -9192 -12094 -9183 -12088
rect -10216 -12101 -10024 -12094
rect -10658 -12148 -10629 -12101
rect -10060 -12148 -10024 -12101
rect -10658 -12160 -10472 -12148
rect -10216 -12160 -10024 -12148
rect -10658 -12214 -10024 -12160
rect -9549 -12101 -9183 -12094
rect -8927 -12094 -8918 -12088
rect -8475 -12088 -8201 -12079
rect -8475 -12094 -8466 -12088
rect -9549 -12148 -9520 -12101
rect -9549 -12160 -9183 -12148
rect -8927 -12160 -8915 -12094
rect -9549 -12214 -8915 -12160
rect -8667 -12101 -8466 -12094
rect -8210 -12094 -8201 -12088
rect -8210 -12101 -8033 -12094
rect -8667 -12148 -8638 -12101
rect -8069 -12148 -8033 -12101
rect -8667 -12160 -8466 -12148
rect -8210 -12160 -8033 -12148
rect -8667 -12214 -8033 -12160
rect -20531 -12220 -19896 -12214
rect -21731 -12240 -21304 -12234
rect -22567 -12260 -21885 -12254
rect -23583 -12402 -22951 -12274
rect -23583 -12436 -23571 -12402
rect -23395 -12436 -22951 -12402
rect -22910 -12307 -22531 -12289
rect -22910 -12316 -22581 -12307
rect -22910 -12408 -22868 -12316
rect -22670 -12342 -22581 -12316
rect -22547 -12342 -22531 -12307
rect -22670 -12408 -22531 -12342
rect -22910 -12424 -22531 -12408
rect -22503 -12307 -22243 -12288
rect -22503 -12342 -22292 -12307
rect -22258 -12342 -22243 -12307
rect -22503 -12362 -22243 -12342
rect -23583 -12442 -23383 -12436
rect -24637 -12578 -24190 -12466
rect -23683 -12446 -23614 -12442
rect -23683 -12480 -23664 -12446
rect -23630 -12480 -23614 -12446
rect -23683 -12497 -23614 -12480
rect -23583 -12490 -23383 -12483
rect -24637 -12776 -24612 -12578
rect -24466 -12589 -24190 -12578
rect -23583 -12524 -23571 -12490
rect -23395 -12524 -23383 -12490
rect -23355 -12495 -22951 -12436
rect -22503 -12431 -22453 -12362
rect -22167 -12390 -21885 -12260
rect -22503 -12453 -22497 -12431
rect -22695 -12454 -22497 -12453
rect -22773 -12466 -22497 -12454
rect -22463 -12466 -22453 -12431
rect -22425 -12402 -21885 -12390
rect -22425 -12436 -22413 -12402
rect -22037 -12436 -21885 -12402
rect -22425 -12442 -21885 -12436
rect -21854 -12274 -21725 -12240
rect -21648 -12274 -21304 -12240
rect -21854 -12276 -21304 -12274
rect -21854 -12402 -21554 -12276
rect -21854 -12436 -21842 -12402
rect -21666 -12436 -21554 -12402
rect -21854 -12442 -21654 -12436
rect -22773 -12472 -22453 -12466
rect -23355 -12497 -23012 -12495
rect -24466 -12776 -24432 -12589
rect -24162 -12594 -23762 -12588
rect -24162 -12628 -24150 -12594
rect -23774 -12628 -23762 -12594
rect -24162 -12666 -24133 -12628
rect -24162 -12700 -24135 -12666
rect -23793 -12690 -23762 -12628
rect -23583 -12607 -23556 -12524
rect -23407 -12607 -23383 -12524
rect -22773 -12560 -22730 -12472
rect -22611 -12560 -22453 -12472
rect -21954 -12446 -21885 -12442
rect -21954 -12480 -21935 -12446
rect -21901 -12480 -21885 -12446
rect -21954 -12497 -21885 -12480
rect -21626 -12462 -21554 -12436
rect -21355 -12462 -21304 -12276
rect -20531 -12300 -20518 -12220
rect -20484 -12300 -20326 -12220
rect -20292 -12300 -20134 -12220
rect -20100 -12300 -19942 -12220
rect -19908 -12300 -19896 -12220
rect -20531 -12306 -19896 -12300
rect -19422 -12220 -18787 -12214
rect -19422 -12300 -19409 -12220
rect -19375 -12300 -19217 -12220
rect -19183 -12300 -19025 -12220
rect -18991 -12300 -18833 -12220
rect -18799 -12300 -18787 -12220
rect -19422 -12306 -18787 -12300
rect -18540 -12220 -17905 -12214
rect -18540 -12300 -18527 -12220
rect -18493 -12300 -18335 -12220
rect -18301 -12300 -18143 -12220
rect -18109 -12300 -17951 -12220
rect -17917 -12300 -17905 -12220
rect -18540 -12306 -17905 -12300
rect -17240 -12220 -16605 -12214
rect -17240 -12300 -17227 -12220
rect -17193 -12300 -17035 -12220
rect -17001 -12300 -16843 -12220
rect -16809 -12300 -16651 -12220
rect -16617 -12300 -16605 -12220
rect -17240 -12306 -16605 -12300
rect -16131 -12220 -15496 -12214
rect -16131 -12300 -16118 -12220
rect -16084 -12300 -15926 -12220
rect -15892 -12300 -15734 -12220
rect -15700 -12300 -15542 -12220
rect -15508 -12300 -15496 -12220
rect -16131 -12306 -15496 -12300
rect -15249 -12220 -14614 -12214
rect -15249 -12300 -15236 -12220
rect -15202 -12300 -15044 -12220
rect -15010 -12300 -14852 -12220
rect -14818 -12300 -14660 -12220
rect -14626 -12300 -14614 -12220
rect -15249 -12306 -14614 -12300
rect -13949 -12220 -13314 -12214
rect -13949 -12300 -13936 -12220
rect -13902 -12300 -13744 -12220
rect -13710 -12300 -13552 -12220
rect -13518 -12300 -13360 -12220
rect -13326 -12300 -13314 -12220
rect -13949 -12306 -13314 -12300
rect -12840 -12220 -12205 -12214
rect -12840 -12300 -12827 -12220
rect -12793 -12300 -12635 -12220
rect -12601 -12300 -12443 -12220
rect -12409 -12300 -12251 -12220
rect -12217 -12300 -12205 -12220
rect -12840 -12306 -12205 -12300
rect -11958 -12220 -11323 -12214
rect -11958 -12300 -11945 -12220
rect -11911 -12300 -11753 -12220
rect -11719 -12300 -11561 -12220
rect -11527 -12300 -11369 -12220
rect -11335 -12300 -11323 -12220
rect -11958 -12306 -11323 -12300
rect -10658 -12220 -10023 -12214
rect -10658 -12300 -10645 -12220
rect -10611 -12300 -10453 -12220
rect -10419 -12300 -10261 -12220
rect -10227 -12300 -10069 -12220
rect -10035 -12300 -10023 -12220
rect -10658 -12306 -10023 -12300
rect -9549 -12220 -8914 -12214
rect -9549 -12300 -9536 -12220
rect -9502 -12300 -9344 -12220
rect -9310 -12300 -9152 -12220
rect -9118 -12300 -8960 -12220
rect -8926 -12300 -8914 -12220
rect -9549 -12306 -8914 -12300
rect -8667 -12220 -8032 -12214
rect -8667 -12300 -8654 -12220
rect -8620 -12300 -8462 -12220
rect -8428 -12300 -8270 -12220
rect -8236 -12300 -8078 -12220
rect -8044 -12300 -8032 -12220
rect -8667 -12306 -8032 -12300
rect -20531 -12307 -19897 -12306
rect -19422 -12307 -18788 -12306
rect -18540 -12307 -17906 -12306
rect -17240 -12307 -16606 -12306
rect -16131 -12307 -15497 -12306
rect -15249 -12307 -14615 -12306
rect -13949 -12307 -13315 -12306
rect -12840 -12307 -12206 -12306
rect -11958 -12307 -11324 -12306
rect -10658 -12307 -10024 -12306
rect -9549 -12307 -8915 -12306
rect -8667 -12307 -8033 -12306
rect -20438 -12342 -19860 -12336
rect -20438 -12422 -20422 -12342
rect -20388 -12422 -20230 -12342
rect -20196 -12422 -20038 -12342
rect -20004 -12422 -19860 -12342
rect -20438 -12423 -19860 -12422
rect -20438 -12428 -19979 -12423
rect -21854 -12490 -21654 -12483
rect -22773 -12589 -22453 -12560
rect -21854 -12524 -21842 -12490
rect -21666 -12524 -21654 -12490
rect -21626 -12497 -21304 -12462
rect -20566 -12475 -20402 -12457
rect -20566 -12484 -20452 -12475
rect -23583 -12626 -23552 -12607
rect -23420 -12626 -23383 -12607
rect -23583 -12633 -23383 -12626
rect -22425 -12594 -22025 -12588
rect -22425 -12628 -22413 -12594
rect -22037 -12628 -22025 -12594
rect -23800 -12700 -23762 -12690
rect -24162 -12711 -23762 -12700
rect -22425 -12666 -22396 -12628
rect -22425 -12700 -22398 -12666
rect -22056 -12690 -22025 -12628
rect -21854 -12607 -21827 -12524
rect -21678 -12607 -21654 -12524
rect -20566 -12564 -20534 -12484
rect -20418 -12510 -20402 -12475
rect -20436 -12564 -20402 -12510
rect -20566 -12592 -20402 -12564
rect -20374 -12475 -20114 -12456
rect -20374 -12510 -20163 -12475
rect -20129 -12510 -20114 -12475
rect -20374 -12530 -20114 -12510
rect -21854 -12626 -21823 -12607
rect -21691 -12626 -21654 -12607
rect -20374 -12599 -20324 -12530
rect -20038 -12558 -19979 -12428
rect -20374 -12620 -20368 -12599
rect -21854 -12633 -21654 -12626
rect -22063 -12700 -22025 -12690
rect -22425 -12711 -22025 -12700
rect -20762 -12634 -20368 -12620
rect -20334 -12634 -20324 -12599
rect -20296 -12570 -19979 -12558
rect -20296 -12604 -20284 -12570
rect -19896 -12571 -19860 -12423
rect -19329 -12342 -18751 -12336
rect -19329 -12422 -19313 -12342
rect -19279 -12422 -19121 -12342
rect -19087 -12422 -18929 -12342
rect -18895 -12422 -18751 -12342
rect -19329 -12428 -18751 -12422
rect -18447 -12342 -17869 -12336
rect -18447 -12422 -18431 -12342
rect -18397 -12422 -18239 -12342
rect -18205 -12422 -18047 -12342
rect -18013 -12422 -17869 -12342
rect -18447 -12428 -17869 -12422
rect -17147 -12342 -16569 -12336
rect -17147 -12422 -17131 -12342
rect -17097 -12422 -16939 -12342
rect -16905 -12422 -16747 -12342
rect -16713 -12422 -16569 -12342
rect -17147 -12423 -16569 -12422
rect -17147 -12428 -16688 -12423
rect -19908 -12604 -19860 -12571
rect -19457 -12475 -19293 -12457
rect -19457 -12485 -19343 -12475
rect -19457 -12565 -19423 -12485
rect -19309 -12510 -19293 -12475
rect -19325 -12565 -19293 -12510
rect -19457 -12592 -19293 -12565
rect -19265 -12475 -19005 -12456
rect -19265 -12510 -19054 -12475
rect -19020 -12510 -19005 -12475
rect -19265 -12530 -19005 -12510
rect -18929 -12480 -18751 -12428
rect -18575 -12475 -18411 -12457
rect -18575 -12480 -18461 -12475
rect -18929 -12510 -18461 -12480
rect -18427 -12510 -18411 -12475
rect -20296 -12610 -19860 -12604
rect -19265 -12599 -19215 -12530
rect -18929 -12558 -18411 -12510
rect -19265 -12621 -19259 -12599
rect -20762 -12677 -20324 -12634
rect -20762 -12743 -20743 -12677
rect -20490 -12743 -20324 -12677
rect -20762 -12757 -20324 -12743
rect -19457 -12634 -19259 -12621
rect -19225 -12634 -19215 -12599
rect -19187 -12570 -18411 -12558
rect -19187 -12604 -19175 -12570
rect -18799 -12604 -18751 -12570
rect -18575 -12592 -18411 -12570
rect -18383 -12475 -18123 -12456
rect -18383 -12510 -18172 -12475
rect -18138 -12510 -18123 -12475
rect -18383 -12530 -18123 -12510
rect -18047 -12473 -17869 -12428
rect -19187 -12610 -18751 -12604
rect -18383 -12599 -18333 -12530
rect -18047 -12553 -18002 -12473
rect -17882 -12553 -17869 -12473
rect -18047 -12558 -17869 -12553
rect -18383 -12621 -18377 -12599
rect -19457 -12688 -19215 -12634
rect -19457 -12748 -19433 -12688
rect -19248 -12748 -19215 -12688
rect -24637 -12791 -24432 -12776
rect -20296 -12762 -19896 -12756
rect -19457 -12757 -19215 -12748
rect -18575 -12634 -18377 -12621
rect -18343 -12634 -18333 -12599
rect -18305 -12570 -17869 -12558
rect -18305 -12604 -18293 -12570
rect -17917 -12604 -17869 -12570
rect -17275 -12475 -17111 -12457
rect -17275 -12484 -17161 -12475
rect -17275 -12564 -17243 -12484
rect -17127 -12510 -17111 -12475
rect -17145 -12564 -17111 -12510
rect -17275 -12592 -17111 -12564
rect -17083 -12475 -16823 -12456
rect -17083 -12510 -16872 -12475
rect -16838 -12510 -16823 -12475
rect -17083 -12530 -16823 -12510
rect -18305 -12610 -17869 -12604
rect -17083 -12599 -17033 -12530
rect -16747 -12558 -16688 -12428
rect -17083 -12620 -17077 -12599
rect -18575 -12639 -18333 -12634
rect -18575 -12714 -18561 -12639
rect -18416 -12714 -18333 -12639
rect -20296 -12796 -20284 -12762
rect -19908 -12796 -19896 -12762
rect -20296 -12834 -19896 -12796
rect -20296 -12879 -20269 -12834
rect -20278 -12886 -20269 -12879
rect -19934 -12879 -19896 -12834
rect -19187 -12762 -18787 -12756
rect -18575 -12757 -18333 -12714
rect -17471 -12634 -17077 -12620
rect -17043 -12634 -17033 -12599
rect -17005 -12570 -16688 -12558
rect -17005 -12604 -16993 -12570
rect -16605 -12571 -16569 -12423
rect -16038 -12342 -15460 -12336
rect -16038 -12422 -16022 -12342
rect -15988 -12422 -15830 -12342
rect -15796 -12422 -15638 -12342
rect -15604 -12422 -15460 -12342
rect -16038 -12428 -15460 -12422
rect -15156 -12342 -14578 -12336
rect -15156 -12422 -15140 -12342
rect -15106 -12422 -14948 -12342
rect -14914 -12422 -14756 -12342
rect -14722 -12422 -14578 -12342
rect -15156 -12428 -14578 -12422
rect -13856 -12342 -13278 -12336
rect -13856 -12422 -13840 -12342
rect -13806 -12422 -13648 -12342
rect -13614 -12422 -13456 -12342
rect -13422 -12422 -13278 -12342
rect -13856 -12423 -13278 -12422
rect -13856 -12428 -13397 -12423
rect -16617 -12604 -16569 -12571
rect -16166 -12475 -16002 -12457
rect -16166 -12485 -16052 -12475
rect -16166 -12565 -16132 -12485
rect -16018 -12510 -16002 -12475
rect -16034 -12565 -16002 -12510
rect -16166 -12592 -16002 -12565
rect -15974 -12475 -15714 -12456
rect -15974 -12510 -15763 -12475
rect -15729 -12510 -15714 -12475
rect -15974 -12530 -15714 -12510
rect -15638 -12480 -15460 -12428
rect -15284 -12475 -15120 -12457
rect -15284 -12480 -15170 -12475
rect -15638 -12510 -15170 -12480
rect -15136 -12510 -15120 -12475
rect -17005 -12610 -16569 -12604
rect -15974 -12599 -15924 -12530
rect -15638 -12558 -15120 -12510
rect -15974 -12621 -15968 -12599
rect -17471 -12677 -17033 -12634
rect -17471 -12743 -17452 -12677
rect -17199 -12743 -17033 -12677
rect -19187 -12796 -19175 -12762
rect -18799 -12796 -18787 -12762
rect -19187 -12834 -18787 -12796
rect -19187 -12868 -19160 -12834
rect -18825 -12868 -18787 -12834
rect -19187 -12879 -19033 -12868
rect -19934 -12886 -19925 -12879
rect -20278 -12895 -19925 -12886
rect -19044 -12901 -19033 -12879
rect -18971 -12879 -18787 -12868
rect -18305 -12762 -17905 -12756
rect -17471 -12757 -17033 -12743
rect -16166 -12634 -15968 -12621
rect -15934 -12634 -15924 -12599
rect -15896 -12570 -15120 -12558
rect -15896 -12604 -15884 -12570
rect -15508 -12604 -15460 -12570
rect -15284 -12592 -15120 -12570
rect -15092 -12475 -14832 -12456
rect -15092 -12510 -14881 -12475
rect -14847 -12510 -14832 -12475
rect -15092 -12530 -14832 -12510
rect -14756 -12473 -14578 -12428
rect -15896 -12610 -15460 -12604
rect -15092 -12599 -15042 -12530
rect -14756 -12553 -14711 -12473
rect -14591 -12553 -14578 -12473
rect -14756 -12558 -14578 -12553
rect -15092 -12621 -15086 -12599
rect -16166 -12688 -15924 -12634
rect -16166 -12748 -16142 -12688
rect -15957 -12748 -15924 -12688
rect -18305 -12796 -18293 -12762
rect -17917 -12796 -17905 -12762
rect -18305 -12834 -17905 -12796
rect -18305 -12868 -18278 -12834
rect -17943 -12868 -17905 -12834
rect -18305 -12879 -18166 -12868
rect -18971 -12901 -18960 -12879
rect -19044 -12912 -18960 -12901
rect -18179 -12918 -18166 -12879
rect -18114 -12879 -17905 -12868
rect -17005 -12762 -16605 -12756
rect -16166 -12757 -15924 -12748
rect -15284 -12634 -15086 -12621
rect -15052 -12634 -15042 -12599
rect -15014 -12570 -14578 -12558
rect -15014 -12604 -15002 -12570
rect -14626 -12604 -14578 -12570
rect -13984 -12475 -13820 -12457
rect -13984 -12484 -13870 -12475
rect -13984 -12564 -13952 -12484
rect -13836 -12510 -13820 -12475
rect -13854 -12564 -13820 -12510
rect -13984 -12592 -13820 -12564
rect -13792 -12475 -13532 -12456
rect -13792 -12510 -13581 -12475
rect -13547 -12510 -13532 -12475
rect -13792 -12530 -13532 -12510
rect -15014 -12610 -14578 -12604
rect -13792 -12599 -13742 -12530
rect -13456 -12558 -13397 -12428
rect -13792 -12620 -13786 -12599
rect -15284 -12639 -15042 -12634
rect -15284 -12714 -15270 -12639
rect -15125 -12714 -15042 -12639
rect -17005 -12796 -16993 -12762
rect -16617 -12796 -16605 -12762
rect -17005 -12834 -16605 -12796
rect -17005 -12879 -16978 -12834
rect -18114 -12918 -18101 -12879
rect -16987 -12886 -16978 -12879
rect -16643 -12879 -16605 -12834
rect -15896 -12762 -15496 -12756
rect -15284 -12757 -15042 -12714
rect -14180 -12634 -13786 -12620
rect -13752 -12634 -13742 -12599
rect -13714 -12570 -13397 -12558
rect -13714 -12604 -13702 -12570
rect -13314 -12571 -13278 -12423
rect -12747 -12342 -12169 -12336
rect -12747 -12422 -12731 -12342
rect -12697 -12422 -12539 -12342
rect -12505 -12422 -12347 -12342
rect -12313 -12422 -12169 -12342
rect -12747 -12428 -12169 -12422
rect -11865 -12342 -11287 -12336
rect -11865 -12422 -11849 -12342
rect -11815 -12422 -11657 -12342
rect -11623 -12422 -11465 -12342
rect -11431 -12422 -11287 -12342
rect -11865 -12428 -11287 -12422
rect -10565 -12342 -9987 -12336
rect -10565 -12422 -10549 -12342
rect -10515 -12422 -10357 -12342
rect -10323 -12422 -10165 -12342
rect -10131 -12422 -9987 -12342
rect -10565 -12423 -9987 -12422
rect -10565 -12428 -10106 -12423
rect -13326 -12604 -13278 -12571
rect -12875 -12475 -12711 -12457
rect -12875 -12485 -12761 -12475
rect -12875 -12565 -12841 -12485
rect -12727 -12510 -12711 -12475
rect -12743 -12565 -12711 -12510
rect -12875 -12592 -12711 -12565
rect -12683 -12475 -12423 -12456
rect -12683 -12510 -12472 -12475
rect -12438 -12510 -12423 -12475
rect -12683 -12530 -12423 -12510
rect -12347 -12480 -12169 -12428
rect -11993 -12475 -11829 -12457
rect -11993 -12480 -11879 -12475
rect -12347 -12510 -11879 -12480
rect -11845 -12510 -11829 -12475
rect -13714 -12610 -13278 -12604
rect -12683 -12599 -12633 -12530
rect -12347 -12558 -11829 -12510
rect -12683 -12621 -12677 -12599
rect -14180 -12677 -13742 -12634
rect -14180 -12743 -14161 -12677
rect -13908 -12743 -13742 -12677
rect -15896 -12796 -15884 -12762
rect -15508 -12796 -15496 -12762
rect -15896 -12834 -15496 -12796
rect -15896 -12868 -15869 -12834
rect -15534 -12868 -15496 -12834
rect -15896 -12879 -15742 -12868
rect -16643 -12886 -16634 -12879
rect -16987 -12895 -16634 -12886
rect -15753 -12901 -15742 -12879
rect -15680 -12879 -15496 -12868
rect -15014 -12762 -14614 -12756
rect -14180 -12757 -13742 -12743
rect -12875 -12634 -12677 -12621
rect -12643 -12634 -12633 -12599
rect -12605 -12570 -11829 -12558
rect -12605 -12604 -12593 -12570
rect -12217 -12604 -12169 -12570
rect -11993 -12592 -11829 -12570
rect -11801 -12475 -11541 -12456
rect -11801 -12510 -11590 -12475
rect -11556 -12510 -11541 -12475
rect -11801 -12530 -11541 -12510
rect -11465 -12473 -11287 -12428
rect -12605 -12610 -12169 -12604
rect -11801 -12599 -11751 -12530
rect -11465 -12553 -11420 -12473
rect -11300 -12553 -11287 -12473
rect -11465 -12558 -11287 -12553
rect -11801 -12621 -11795 -12599
rect -12875 -12688 -12633 -12634
rect -12875 -12748 -12851 -12688
rect -12666 -12748 -12633 -12688
rect -15014 -12796 -15002 -12762
rect -14626 -12796 -14614 -12762
rect -15014 -12834 -14614 -12796
rect -15014 -12868 -14987 -12834
rect -14652 -12868 -14614 -12834
rect -15014 -12879 -14875 -12868
rect -15680 -12901 -15669 -12879
rect -15753 -12912 -15669 -12901
rect -18179 -12931 -18101 -12918
rect -14888 -12918 -14875 -12879
rect -14823 -12879 -14614 -12868
rect -13714 -12762 -13314 -12756
rect -12875 -12757 -12633 -12748
rect -11993 -12634 -11795 -12621
rect -11761 -12634 -11751 -12599
rect -11723 -12570 -11287 -12558
rect -11723 -12604 -11711 -12570
rect -11335 -12604 -11287 -12570
rect -10693 -12475 -10529 -12457
rect -10693 -12484 -10579 -12475
rect -10693 -12564 -10661 -12484
rect -10545 -12510 -10529 -12475
rect -10563 -12564 -10529 -12510
rect -10693 -12592 -10529 -12564
rect -10501 -12475 -10241 -12456
rect -10501 -12510 -10290 -12475
rect -10256 -12510 -10241 -12475
rect -10501 -12530 -10241 -12510
rect -11723 -12610 -11287 -12604
rect -10501 -12599 -10451 -12530
rect -10165 -12558 -10106 -12428
rect -10501 -12620 -10495 -12599
rect -11993 -12639 -11751 -12634
rect -11993 -12714 -11979 -12639
rect -11834 -12714 -11751 -12639
rect -13714 -12796 -13702 -12762
rect -13326 -12796 -13314 -12762
rect -13714 -12834 -13314 -12796
rect -13714 -12879 -13687 -12834
rect -14823 -12918 -14810 -12879
rect -13696 -12886 -13687 -12879
rect -13352 -12879 -13314 -12834
rect -12605 -12762 -12205 -12756
rect -11993 -12757 -11751 -12714
rect -10889 -12634 -10495 -12620
rect -10461 -12634 -10451 -12599
rect -10423 -12570 -10106 -12558
rect -10423 -12604 -10411 -12570
rect -10023 -12571 -9987 -12423
rect -9456 -12342 -8878 -12336
rect -9456 -12422 -9440 -12342
rect -9406 -12422 -9248 -12342
rect -9214 -12422 -9056 -12342
rect -9022 -12422 -8878 -12342
rect -9456 -12428 -8878 -12422
rect -8574 -12342 -7996 -12336
rect -8574 -12422 -8558 -12342
rect -8524 -12422 -8366 -12342
rect -8332 -12422 -8174 -12342
rect -8140 -12422 -7996 -12342
rect -8574 -12428 -7996 -12422
rect -10035 -12604 -9987 -12571
rect -9584 -12475 -9420 -12457
rect -9584 -12485 -9470 -12475
rect -9584 -12565 -9550 -12485
rect -9436 -12510 -9420 -12475
rect -9452 -12565 -9420 -12510
rect -9584 -12592 -9420 -12565
rect -9392 -12475 -9132 -12456
rect -9392 -12510 -9181 -12475
rect -9147 -12510 -9132 -12475
rect -9392 -12530 -9132 -12510
rect -9056 -12480 -8878 -12428
rect -8702 -12475 -8538 -12457
rect -8702 -12480 -8588 -12475
rect -9056 -12510 -8588 -12480
rect -8554 -12510 -8538 -12475
rect -10423 -12610 -9987 -12604
rect -9392 -12599 -9342 -12530
rect -9056 -12558 -8538 -12510
rect -9392 -12621 -9386 -12599
rect -10889 -12677 -10451 -12634
rect -10889 -12743 -10870 -12677
rect -10617 -12743 -10451 -12677
rect -12605 -12796 -12593 -12762
rect -12217 -12796 -12205 -12762
rect -12605 -12834 -12205 -12796
rect -12605 -12868 -12578 -12834
rect -12243 -12868 -12205 -12834
rect -12605 -12879 -12451 -12868
rect -13352 -12886 -13343 -12879
rect -13696 -12895 -13343 -12886
rect -12462 -12901 -12451 -12879
rect -12389 -12879 -12205 -12868
rect -11723 -12762 -11323 -12756
rect -10889 -12757 -10451 -12743
rect -9584 -12634 -9386 -12621
rect -9352 -12634 -9342 -12599
rect -9314 -12570 -8538 -12558
rect -9314 -12604 -9302 -12570
rect -8926 -12604 -8878 -12570
rect -8702 -12592 -8538 -12570
rect -8510 -12475 -8250 -12456
rect -8510 -12510 -8299 -12475
rect -8265 -12510 -8250 -12475
rect -8510 -12530 -8250 -12510
rect -8174 -12473 -7996 -12428
rect -9314 -12610 -8878 -12604
rect -8510 -12599 -8460 -12530
rect -8174 -12553 -8129 -12473
rect -8009 -12553 -7996 -12473
rect -8174 -12558 -7996 -12553
rect -8510 -12621 -8504 -12599
rect -9584 -12688 -9342 -12634
rect -9584 -12748 -9560 -12688
rect -9375 -12748 -9342 -12688
rect -11723 -12796 -11711 -12762
rect -11335 -12796 -11323 -12762
rect -11723 -12834 -11323 -12796
rect -11723 -12868 -11696 -12834
rect -11361 -12868 -11323 -12834
rect -11723 -12879 -11584 -12868
rect -12389 -12901 -12378 -12879
rect -12462 -12912 -12378 -12901
rect -14888 -12931 -14810 -12918
rect -11597 -12918 -11584 -12879
rect -11532 -12879 -11323 -12868
rect -10423 -12762 -10023 -12756
rect -9584 -12757 -9342 -12748
rect -8702 -12634 -8504 -12621
rect -8470 -12634 -8460 -12599
rect -8432 -12570 -7996 -12558
rect -8432 -12604 -8420 -12570
rect -8044 -12604 -7996 -12570
rect -8432 -12610 -7996 -12604
rect -1325 -12387 295 -12321
rect -8702 -12639 -8460 -12634
rect -8702 -12714 -8688 -12639
rect -8543 -12714 -8460 -12639
rect -10423 -12796 -10411 -12762
rect -10035 -12796 -10023 -12762
rect -10423 -12834 -10023 -12796
rect -10423 -12879 -10396 -12834
rect -11532 -12918 -11519 -12879
rect -10405 -12886 -10396 -12879
rect -10061 -12879 -10023 -12834
rect -9314 -12762 -8914 -12756
rect -8702 -12757 -8460 -12714
rect -9314 -12796 -9302 -12762
rect -8926 -12796 -8914 -12762
rect -9314 -12834 -8914 -12796
rect -9314 -12868 -9287 -12834
rect -8952 -12868 -8914 -12834
rect -9314 -12879 -9160 -12868
rect -10061 -12886 -10052 -12879
rect -10405 -12895 -10052 -12886
rect -9171 -12901 -9160 -12879
rect -9098 -12879 -8914 -12868
rect -8432 -12762 -8032 -12756
rect -8432 -12796 -8420 -12762
rect -8044 -12796 -8032 -12762
rect -8432 -12834 -8032 -12796
rect -8432 -12868 -8405 -12834
rect -8070 -12868 -8032 -12834
rect -8432 -12879 -8293 -12868
rect -9098 -12901 -9087 -12879
rect -9171 -12912 -9087 -12901
rect -11597 -12931 -11519 -12918
rect -8306 -12918 -8293 -12879
rect -8241 -12879 -8032 -12868
rect -7799 -12798 -7688 -12792
rect -1325 -12797 -1259 -12387
rect -8241 -12918 -8228 -12879
rect -7799 -12915 -7688 -12909
rect -6359 -12863 -1259 -12797
rect -1209 -12549 125 -12483
rect -8306 -12931 -8228 -12918
rect -6359 -13379 -6293 -12863
rect -1209 -12927 -1143 -12549
rect -11157 -13445 -11151 -13379
rect -11085 -13445 -6293 -13379
rect -6213 -12993 -1143 -12927
rect -1076 -12682 -57 -12623
rect -6213 -13577 -6147 -12993
rect -1076 -13069 -1017 -12682
rect -768 -12818 -684 -12812
rect -684 -12902 -676 -12834
rect -768 -12932 -676 -12902
rect -14449 -13643 -14443 -13577
rect -14377 -13643 -6147 -13577
rect -6088 -13128 -1017 -13069
rect -760 -13066 -676 -12932
rect -6088 -13700 -6029 -13128
rect -760 -13150 -374 -13066
rect -768 -13259 -684 -13258
rect -5292 -13312 -5286 -13259
rect -5233 -13312 -682 -13259
rect -5814 -13408 -5730 -13402
rect -5730 -13492 -850 -13408
rect -5814 -13498 -5730 -13492
rect -17736 -13759 -17730 -13700
rect -17671 -13759 -6029 -13700
rect -1242 -13666 -1058 -13623
rect -1242 -13720 -1201 -13666
rect -4632 -13818 -4626 -13734
rect -4542 -13818 -3436 -13734
rect -2068 -13750 -1201 -13720
rect -1117 -13750 -1058 -13666
rect -2068 -13804 -1058 -13750
rect -14814 -13976 -14808 -13924
rect -14756 -13976 -14750 -13924
rect -11441 -13973 -10779 -13897
rect -5376 -13928 -5370 -13876
rect -5318 -13880 -5312 -13876
rect -5174 -13880 -3570 -13860
rect -5318 -13924 -3570 -13880
rect -5318 -13928 -5312 -13924
rect -5174 -13944 -3570 -13924
rect -17535 -14465 -16984 -14463
rect -21025 -14475 -20959 -14469
rect -20959 -14541 -19311 -14475
rect -21025 -14547 -20959 -14541
rect -24197 -14835 -22338 -14766
rect -24197 -14844 -23005 -14835
rect -24197 -14880 -24115 -14844
rect -24449 -14917 -24357 -14916
rect -24569 -14928 -24356 -14917
rect -24569 -14953 -24443 -14928
rect -24847 -15194 -24735 -15186
rect -24569 -15194 -24562 -14953
rect -24847 -15290 -24839 -15194
rect -24743 -15290 -24562 -15194
rect -24847 -15298 -24735 -15290
rect -24569 -15522 -24562 -15290
rect -24515 -14962 -24443 -14953
rect -24363 -14962 -24356 -14928
rect -24515 -15120 -24356 -14962
rect -24515 -15154 -24443 -15120
rect -24363 -15154 -24356 -15120
rect -24515 -15312 -24356 -15154
rect -24515 -15346 -24443 -15312
rect -24363 -15346 -24356 -15312
rect -24515 -15504 -24356 -15346
rect -24327 -14928 -24053 -14880
rect -24327 -15024 -24093 -14928
rect -24327 -15058 -24321 -15024
rect -24241 -15058 -24093 -15024
rect -24327 -15216 -24235 -15058
rect -24327 -15250 -24321 -15216
rect -24241 -15250 -24235 -15216
rect -24327 -15408 -24235 -15250
rect -24207 -15149 -24133 -15134
rect -24207 -15183 -24188 -15149
rect -24153 -15183 -24133 -15149
rect -24207 -15344 -24133 -15183
rect -24105 -15304 -24093 -15058
rect -24059 -15304 -24053 -14928
rect -24105 -15316 -24053 -15304
rect -23907 -14928 -23784 -14916
rect -23907 -15304 -23901 -14928
rect -23867 -14954 -23784 -14928
rect -23867 -15289 -23829 -14954
rect -23795 -15075 -23784 -14954
rect -23795 -15176 -23421 -15075
rect -23320 -15176 -23314 -15075
rect -23795 -15289 -23784 -15176
rect -23867 -15304 -23784 -15289
rect -23907 -15316 -23784 -15304
rect -24207 -15354 -23906 -15344
rect -24207 -15388 -24064 -15354
rect -24029 -15388 -23906 -15354
rect -24207 -15394 -23906 -15388
rect -24327 -15442 -24321 -15408
rect -24241 -15442 -24235 -15408
rect -24327 -15458 -24235 -15442
rect -24206 -15438 -24071 -15422
rect -24515 -15522 -24443 -15504
rect -24569 -15538 -24443 -15522
rect -24363 -15538 -24356 -15504
rect -24569 -15551 -24356 -15538
rect -24206 -15472 -24188 -15438
rect -24153 -15472 -24071 -15438
rect -24206 -15586 -24071 -15472
rect -24936 -15658 -24916 -15586
rect -24844 -15658 -24071 -15586
rect -24042 -15739 -23906 -15394
rect -24936 -15828 -24903 -15739
rect -24812 -15828 -23906 -15739
rect -24189 -15968 -23005 -15959
rect -24189 -16037 -22526 -15968
rect -24189 -16065 -24107 -16037
rect -24448 -16102 -24356 -16101
rect -24568 -16113 -24355 -16102
rect -24568 -16138 -24442 -16113
rect -24843 -16368 -24731 -16360
rect -24568 -16368 -24561 -16138
rect -24843 -16464 -24835 -16368
rect -24739 -16464 -24561 -16368
rect -24843 -16472 -24731 -16464
rect -24568 -16707 -24561 -16464
rect -24514 -16147 -24442 -16138
rect -24362 -16147 -24355 -16113
rect -24514 -16305 -24355 -16147
rect -24514 -16339 -24442 -16305
rect -24362 -16339 -24355 -16305
rect -24514 -16497 -24355 -16339
rect -24514 -16531 -24442 -16497
rect -24362 -16531 -24355 -16497
rect -24514 -16689 -24355 -16531
rect -24326 -16113 -24052 -16065
rect -24326 -16209 -24092 -16113
rect -24326 -16243 -24320 -16209
rect -24240 -16243 -24092 -16209
rect -24326 -16401 -24234 -16243
rect -24326 -16435 -24320 -16401
rect -24240 -16435 -24234 -16401
rect -24326 -16593 -24234 -16435
rect -24206 -16334 -24132 -16319
rect -24206 -16368 -24187 -16334
rect -24152 -16368 -24132 -16334
rect -24206 -16529 -24132 -16368
rect -24104 -16489 -24092 -16243
rect -24058 -16489 -24052 -16113
rect -24104 -16501 -24052 -16489
rect -23906 -16113 -23783 -16101
rect -23906 -16489 -23900 -16113
rect -23866 -16139 -23783 -16113
rect -23866 -16474 -23828 -16139
rect -23794 -16271 -23783 -16139
rect -23794 -16372 -23378 -16271
rect -23277 -16372 -23271 -16271
rect -23794 -16474 -23783 -16372
rect -23866 -16489 -23783 -16474
rect -23906 -16501 -23783 -16489
rect -24206 -16539 -23905 -16529
rect -24206 -16573 -24063 -16539
rect -24028 -16573 -23905 -16539
rect -24206 -16579 -23905 -16573
rect -24326 -16627 -24320 -16593
rect -24240 -16627 -24234 -16593
rect -24326 -16643 -24234 -16627
rect -24205 -16623 -24070 -16607
rect -24514 -16707 -24442 -16689
rect -24568 -16723 -24442 -16707
rect -24362 -16723 -24355 -16689
rect -24568 -16736 -24355 -16723
rect -24205 -16657 -24187 -16623
rect -24152 -16657 -24070 -16623
rect -24205 -16770 -24070 -16657
rect -24936 -16842 -24908 -16770
rect -24836 -16842 -24070 -16770
rect -24041 -16923 -23905 -16579
rect -24936 -17012 -24925 -16923
rect -24836 -17012 -23905 -16923
rect -24181 -17233 -22632 -17164
rect -24181 -17242 -23005 -17233
rect -24181 -17278 -24099 -17242
rect -24443 -17315 -24351 -17314
rect -24563 -17326 -24350 -17315
rect -24563 -17351 -24437 -17326
rect -24837 -17600 -24725 -17592
rect -24563 -17600 -24556 -17351
rect -24837 -17696 -24829 -17600
rect -24733 -17696 -24556 -17600
rect -24837 -17704 -24725 -17696
rect -24563 -17920 -24556 -17696
rect -24509 -17360 -24437 -17351
rect -24357 -17360 -24350 -17326
rect -24509 -17518 -24350 -17360
rect -24509 -17552 -24437 -17518
rect -24357 -17552 -24350 -17518
rect -24509 -17710 -24350 -17552
rect -24509 -17744 -24437 -17710
rect -24357 -17744 -24350 -17710
rect -24509 -17902 -24350 -17744
rect -24321 -17326 -24047 -17278
rect -24321 -17422 -24087 -17326
rect -24321 -17456 -24315 -17422
rect -24235 -17456 -24087 -17422
rect -24321 -17614 -24229 -17456
rect -24321 -17648 -24315 -17614
rect -24235 -17648 -24229 -17614
rect -24321 -17806 -24229 -17648
rect -24201 -17547 -24127 -17532
rect -24201 -17581 -24182 -17547
rect -24147 -17581 -24127 -17547
rect -24201 -17742 -24127 -17581
rect -24099 -17702 -24087 -17456
rect -24053 -17702 -24047 -17326
rect -24099 -17714 -24047 -17702
rect -23901 -17326 -23778 -17314
rect -23901 -17702 -23895 -17326
rect -23861 -17352 -23778 -17326
rect -23861 -17687 -23823 -17352
rect -23789 -17483 -23778 -17352
rect -23789 -17584 -23369 -17483
rect -23268 -17584 -23262 -17483
rect -23789 -17687 -23778 -17584
rect -23861 -17702 -23778 -17687
rect -23901 -17714 -23778 -17702
rect -24201 -17752 -23900 -17742
rect -24201 -17786 -24058 -17752
rect -24023 -17786 -23900 -17752
rect -24201 -17792 -23900 -17786
rect -24321 -17840 -24315 -17806
rect -24235 -17840 -24229 -17806
rect -24321 -17856 -24229 -17840
rect -24200 -17836 -24065 -17820
rect -24509 -17920 -24437 -17902
rect -24563 -17936 -24437 -17920
rect -24357 -17936 -24350 -17902
rect -24563 -17949 -24350 -17936
rect -24200 -17870 -24182 -17836
rect -24147 -17870 -24065 -17836
rect -24200 -17984 -24065 -17870
rect -24936 -18054 -24921 -17984
rect -24851 -18054 -24065 -17984
rect -24036 -18128 -23900 -17792
rect -24936 -18217 -24917 -18128
rect -24824 -18217 -23900 -18128
rect -24197 -18276 -23005 -18266
rect -24197 -18344 -22744 -18276
rect -24197 -18397 -24115 -18344
rect -23061 -18345 -22744 -18344
rect -24428 -18434 -24336 -18433
rect -24548 -18445 -24335 -18434
rect -24548 -18470 -24422 -18445
rect -24823 -18714 -24711 -18706
rect -24548 -18714 -24541 -18470
rect -24823 -18810 -24815 -18714
rect -24719 -18810 -24541 -18714
rect -24823 -18818 -24711 -18810
rect -24548 -19039 -24541 -18810
rect -24494 -18479 -24422 -18470
rect -24342 -18479 -24335 -18445
rect -24494 -18637 -24335 -18479
rect -24494 -18671 -24422 -18637
rect -24342 -18671 -24335 -18637
rect -24494 -18829 -24335 -18671
rect -24494 -18863 -24422 -18829
rect -24342 -18863 -24335 -18829
rect -24494 -19021 -24335 -18863
rect -24306 -18445 -24032 -18397
rect -24306 -18541 -24072 -18445
rect -24306 -18575 -24300 -18541
rect -24220 -18575 -24072 -18541
rect -24306 -18733 -24214 -18575
rect -24306 -18767 -24300 -18733
rect -24220 -18767 -24214 -18733
rect -24306 -18925 -24214 -18767
rect -24186 -18666 -24112 -18651
rect -24186 -18700 -24167 -18666
rect -24132 -18700 -24112 -18666
rect -24186 -18861 -24112 -18700
rect -24084 -18821 -24072 -18575
rect -24038 -18821 -24032 -18445
rect -24084 -18833 -24032 -18821
rect -23886 -18445 -23763 -18433
rect -23886 -18821 -23880 -18445
rect -23846 -18471 -23763 -18445
rect -23846 -18806 -23808 -18471
rect -23774 -18624 -23763 -18471
rect -23774 -18725 -23361 -18624
rect -23260 -18725 -23254 -18624
rect -23774 -18806 -23763 -18725
rect -23846 -18821 -23763 -18806
rect -23886 -18833 -23763 -18821
rect -24186 -18871 -23885 -18861
rect -24186 -18905 -24043 -18871
rect -24008 -18905 -23885 -18871
rect -24186 -18911 -23885 -18905
rect -24306 -18959 -24300 -18925
rect -24220 -18959 -24214 -18925
rect -24306 -18975 -24214 -18959
rect -24185 -18955 -24050 -18939
rect -24494 -19039 -24422 -19021
rect -24548 -19055 -24422 -19039
rect -24342 -19055 -24335 -19021
rect -24548 -19068 -24335 -19055
rect -24185 -18989 -24167 -18955
rect -24132 -18989 -24050 -18955
rect -24185 -19103 -24050 -18989
rect -24936 -19175 -24870 -19103
rect -24798 -19175 -24050 -19103
rect -24021 -19256 -23885 -18911
rect -24936 -19345 -24889 -19256
rect -24796 -19345 -23885 -19256
rect -24144 -19460 -23005 -19455
rect -24144 -19529 -22872 -19460
rect -24144 -19533 -23005 -19529
rect -24144 -19591 -24062 -19533
rect -24426 -19628 -24334 -19627
rect -24546 -19639 -24333 -19628
rect -24546 -19664 -24420 -19639
rect -24823 -19908 -24711 -19900
rect -24546 -19908 -24539 -19664
rect -24823 -20004 -24815 -19908
rect -24719 -20004 -24539 -19908
rect -24823 -20012 -24711 -20004
rect -24546 -20233 -24539 -20004
rect -24492 -19673 -24420 -19664
rect -24340 -19673 -24333 -19639
rect -24492 -19831 -24333 -19673
rect -24492 -19865 -24420 -19831
rect -24340 -19865 -24333 -19831
rect -24492 -20023 -24333 -19865
rect -24492 -20057 -24420 -20023
rect -24340 -20057 -24333 -20023
rect -24492 -20215 -24333 -20057
rect -24304 -19639 -24030 -19591
rect -24304 -19735 -24070 -19639
rect -24304 -19769 -24298 -19735
rect -24218 -19769 -24070 -19735
rect -24304 -19927 -24212 -19769
rect -24304 -19961 -24298 -19927
rect -24218 -19961 -24212 -19927
rect -24304 -20119 -24212 -19961
rect -24184 -19860 -24110 -19845
rect -24184 -19894 -24165 -19860
rect -24130 -19894 -24110 -19860
rect -24184 -20055 -24110 -19894
rect -24082 -20015 -24070 -19769
rect -24036 -20015 -24030 -19639
rect -24082 -20027 -24030 -20015
rect -23884 -19639 -23761 -19627
rect -23884 -20015 -23878 -19639
rect -23844 -19665 -23761 -19639
rect -23844 -20000 -23806 -19665
rect -23772 -19796 -23761 -19665
rect -23772 -19897 -23338 -19796
rect -23237 -19897 -23231 -19796
rect -23772 -20000 -23761 -19897
rect -23844 -20015 -23761 -20000
rect -23884 -20027 -23761 -20015
rect -24184 -20065 -23883 -20055
rect -24184 -20099 -24041 -20065
rect -24006 -20099 -23883 -20065
rect -24184 -20105 -23883 -20099
rect -24304 -20153 -24298 -20119
rect -24218 -20153 -24212 -20119
rect -24304 -20169 -24212 -20153
rect -24183 -20149 -24048 -20133
rect -24492 -20233 -24420 -20215
rect -24546 -20249 -24420 -20233
rect -24340 -20249 -24333 -20215
rect -24546 -20262 -24333 -20249
rect -24183 -20183 -24165 -20149
rect -24130 -20183 -24048 -20149
rect -24956 -20291 -24844 -20290
rect -24183 -20291 -24048 -20183
rect -24956 -20363 -24936 -20291
rect -24864 -20363 -24048 -20291
rect -24956 -20364 -24844 -20363
rect -24940 -20444 -24792 -20436
rect -24019 -20444 -23883 -20105
rect -22941 -20239 -22872 -19529
rect -22813 -19759 -22744 -18345
rect -22701 -19259 -22632 -17233
rect -22595 -18779 -22526 -16037
rect -22407 -18279 -22338 -14835
rect -20405 -17936 -20399 -17934
rect -21574 -17984 -20399 -17936
rect -21574 -18020 -21061 -17984
rect -20405 -17986 -20399 -17984
rect -20347 -17986 -20341 -17934
rect -21722 -18094 -21602 -18034
rect -21722 -18117 -21678 -18094
rect -21935 -18169 -21929 -18117
rect -21877 -18169 -21678 -18117
rect -21722 -18185 -21678 -18169
rect -21644 -18157 -21602 -18094
rect -21574 -18042 -21122 -18020
rect -21574 -18119 -21510 -18042
rect -21476 -18119 -21318 -18042
rect -21284 -18048 -21122 -18042
rect -21284 -18060 -21116 -18048
rect -21284 -18119 -21156 -18060
rect -21574 -18125 -21156 -18119
rect -21644 -18163 -21364 -18157
rect -21644 -18185 -21606 -18163
rect -21722 -18242 -21606 -18185
rect -21572 -18242 -21414 -18163
rect -21380 -18242 -21364 -18163
rect -21722 -18248 -21364 -18242
rect -21318 -18236 -21156 -18125
rect -21122 -18236 -21116 -18060
rect -21318 -18248 -21116 -18236
rect -21075 -18060 -20925 -18048
rect -21075 -18236 -21068 -18060
rect -21034 -18085 -20925 -18060
rect -21034 -18217 -20966 -18085
rect -20932 -18174 -20643 -18085
rect -20554 -18174 -20548 -18085
rect -20932 -18217 -20925 -18174
rect -21034 -18236 -20925 -18217
rect -21075 -18248 -20925 -18236
rect -22407 -18295 -21061 -18279
rect -22407 -18329 -21558 -18295
rect -21332 -18329 -21112 -18295
rect -21078 -18329 -21061 -18295
rect -22407 -18348 -21061 -18329
rect -20414 -18434 -20362 -18428
rect -21573 -18484 -20414 -18436
rect -21573 -18520 -21060 -18484
rect -20356 -18436 -20350 -18434
rect -20356 -18484 -20349 -18436
rect -20356 -18486 -20350 -18484
rect -20414 -18492 -20362 -18486
rect -21721 -18594 -21601 -18534
rect -21721 -18626 -21677 -18594
rect -21941 -18678 -21935 -18626
rect -21883 -18678 -21677 -18626
rect -21721 -18685 -21677 -18678
rect -21643 -18657 -21601 -18594
rect -21573 -18542 -21121 -18520
rect -21573 -18619 -21509 -18542
rect -21475 -18619 -21317 -18542
rect -21283 -18548 -21121 -18542
rect -21283 -18560 -21115 -18548
rect -21283 -18619 -21155 -18560
rect -21573 -18625 -21155 -18619
rect -21643 -18663 -21363 -18657
rect -21643 -18685 -21605 -18663
rect -21721 -18742 -21605 -18685
rect -21571 -18742 -21413 -18663
rect -21379 -18742 -21363 -18663
rect -21721 -18748 -21363 -18742
rect -21317 -18736 -21155 -18625
rect -21121 -18736 -21115 -18560
rect -21317 -18748 -21115 -18736
rect -21074 -18560 -20924 -18548
rect -21074 -18736 -21067 -18560
rect -21033 -18578 -20924 -18560
rect -21033 -18585 -20650 -18578
rect -21033 -18717 -20965 -18585
rect -20931 -18667 -20650 -18585
rect -20561 -18667 -20555 -18578
rect -20931 -18717 -20924 -18667
rect -19377 -18705 -19311 -14541
rect -17535 -14511 -16983 -14465
rect -17535 -14545 -17523 -14511
rect -17433 -14516 -16983 -14511
rect -17433 -14545 -16982 -14516
rect -17535 -14579 -16982 -14545
rect -17535 -14588 -16423 -14579
rect -17677 -14607 -17563 -14601
rect -17677 -14641 -17665 -14607
rect -17575 -14641 -17563 -14607
rect -17677 -14799 -17563 -14641
rect -17677 -14833 -17665 -14799
rect -17575 -14833 -17563 -14799
rect -17677 -14991 -17563 -14833
rect -17535 -14703 -17421 -14588
rect -17535 -14737 -17523 -14703
rect -17433 -14737 -17421 -14703
rect -17535 -14895 -17421 -14737
rect -17535 -14929 -17523 -14895
rect -17433 -14929 -17421 -14895
rect -17182 -14648 -16423 -14588
rect -17535 -14935 -17421 -14929
rect -17677 -15025 -17665 -14991
rect -17575 -15025 -17563 -14991
rect -17828 -15122 -17762 -15110
rect -18084 -15281 -17986 -15269
rect -17828 -15281 -17820 -15122
rect -18084 -15355 -18072 -15281
rect -17998 -15355 -17820 -15281
rect -18084 -15367 -17986 -15355
rect -17828 -15479 -17820 -15355
rect -17769 -15479 -17762 -15122
rect -17677 -15183 -17563 -15025
rect -17282 -14943 -17216 -14927
rect -17282 -14977 -17266 -14943
rect -17232 -14977 -17216 -14943
rect -17677 -15217 -17665 -15183
rect -17575 -15217 -17563 -15183
rect -17677 -15375 -17563 -15217
rect -17677 -15409 -17665 -15375
rect -17575 -15409 -17563 -15375
rect -17677 -15415 -17563 -15409
rect -17535 -15087 -17421 -15081
rect -17535 -15121 -17523 -15087
rect -17433 -15121 -17421 -15087
rect -17535 -15279 -17421 -15121
rect -17535 -15313 -17523 -15279
rect -17433 -15313 -17421 -15279
rect -17828 -15491 -17762 -15479
rect -17535 -15471 -17421 -15313
rect -17535 -15505 -17523 -15471
rect -17433 -15505 -17421 -15471
rect -17535 -15511 -17421 -15505
rect -17387 -15086 -17321 -15027
rect -17387 -15120 -17371 -15086
rect -17337 -15120 -17321 -15086
rect -17978 -15586 -17880 -15576
rect -17978 -15658 -17966 -15586
rect -17894 -15590 -17880 -15586
rect -17387 -15590 -17321 -15120
rect -17894 -15656 -17321 -15590
rect -17894 -15658 -17880 -15656
rect -17978 -15666 -17880 -15658
rect -17282 -15724 -17216 -14977
rect -17182 -14985 -16982 -14648
rect -16924 -14908 -16850 -14896
rect -17188 -14991 -16988 -14985
rect -17188 -15025 -17176 -14991
rect -17000 -15025 -16988 -14991
rect -17188 -15031 -16988 -15025
rect -16924 -15107 -16917 -14908
rect -16856 -15107 -16850 -14908
rect -16924 -15119 -16850 -15107
rect -16902 -15311 -16856 -15119
rect -16924 -15330 -16836 -15311
rect -16924 -15382 -16905 -15330
rect -16853 -15382 -16836 -15330
rect -16924 -15401 -16836 -15382
rect -18133 -15738 -17216 -15724
rect -18133 -15827 -18123 -15738
rect -18034 -15790 -17216 -15738
rect -18034 -15827 -18005 -15790
rect -18133 -15847 -18005 -15827
rect -17535 -15865 -16984 -15863
rect -17535 -15899 -16983 -15865
rect -17535 -15911 -16583 -15899
rect -17535 -15945 -17523 -15911
rect -17433 -15945 -16583 -15911
rect -17535 -15968 -16583 -15945
rect -17535 -15988 -16982 -15968
rect -17677 -16007 -17563 -16001
rect -17677 -16041 -17665 -16007
rect -17575 -16041 -17563 -16007
rect -17677 -16199 -17563 -16041
rect -17677 -16233 -17665 -16199
rect -17575 -16233 -17563 -16199
rect -17677 -16391 -17563 -16233
rect -17535 -16103 -17421 -15988
rect -17535 -16137 -17523 -16103
rect -17433 -16137 -17421 -16103
rect -17535 -16295 -17421 -16137
rect -17535 -16329 -17523 -16295
rect -17433 -16329 -17421 -16295
rect -17535 -16335 -17421 -16329
rect -17677 -16425 -17665 -16391
rect -17575 -16425 -17563 -16391
rect -17828 -16522 -17762 -16510
rect -18096 -16683 -17998 -16671
rect -17828 -16683 -17820 -16522
rect -18096 -16757 -18084 -16683
rect -18010 -16757 -17820 -16683
rect -18096 -16769 -17998 -16757
rect -17828 -16879 -17820 -16757
rect -17769 -16879 -17762 -16522
rect -17677 -16583 -17563 -16425
rect -17282 -16343 -17216 -16327
rect -17282 -16377 -17266 -16343
rect -17232 -16377 -17216 -16343
rect -17677 -16617 -17665 -16583
rect -17575 -16617 -17563 -16583
rect -17677 -16775 -17563 -16617
rect -17677 -16809 -17665 -16775
rect -17575 -16809 -17563 -16775
rect -17677 -16815 -17563 -16809
rect -17535 -16487 -17421 -16481
rect -17535 -16521 -17523 -16487
rect -17433 -16521 -17421 -16487
rect -17535 -16679 -17421 -16521
rect -17535 -16713 -17523 -16679
rect -17433 -16713 -17421 -16679
rect -17828 -16891 -17762 -16879
rect -17535 -16871 -17421 -16713
rect -17535 -16905 -17523 -16871
rect -17433 -16905 -17421 -16871
rect -17535 -16911 -17421 -16905
rect -17387 -16486 -17321 -16427
rect -17387 -16520 -17371 -16486
rect -17337 -16520 -17321 -16486
rect -18082 -16980 -18010 -16974
rect -18010 -16988 -17892 -16980
rect -17387 -16988 -17321 -16520
rect -18010 -17052 -17321 -16988
rect -18082 -17058 -18010 -17052
rect -17964 -17054 -17321 -17052
rect -18096 -17113 -17992 -17102
rect -17282 -17112 -17216 -16377
rect -17182 -16385 -16982 -15988
rect -16924 -16308 -16850 -16296
rect -17188 -16391 -16988 -16385
rect -17188 -16425 -17176 -16391
rect -17000 -16425 -16988 -16391
rect -17188 -16431 -16988 -16425
rect -16924 -16507 -16917 -16308
rect -16856 -16507 -16850 -16308
rect -16924 -16519 -16850 -16507
rect -16906 -16717 -16852 -16519
rect -16924 -16735 -16834 -16717
rect -16924 -16789 -16906 -16735
rect -16852 -16789 -16834 -16735
rect -16924 -16807 -16834 -16789
rect -17964 -17113 -17216 -17112
rect -18096 -17202 -18089 -17113
rect -18000 -17178 -17216 -17113
rect -18000 -17202 -17830 -17178
rect -18096 -17208 -17992 -17202
rect -17535 -17265 -16984 -17263
rect -17535 -17311 -16983 -17265
rect -17535 -17345 -17523 -17311
rect -17433 -17316 -16983 -17311
rect -17433 -17319 -16982 -17316
rect -17433 -17345 -16703 -17319
rect -17535 -17388 -16703 -17345
rect -17677 -17407 -17563 -17401
rect -17677 -17441 -17665 -17407
rect -17575 -17441 -17563 -17407
rect -17677 -17599 -17563 -17441
rect -17677 -17633 -17665 -17599
rect -17575 -17633 -17563 -17599
rect -17677 -17791 -17563 -17633
rect -17535 -17503 -17421 -17388
rect -17535 -17537 -17523 -17503
rect -17433 -17537 -17421 -17503
rect -17535 -17695 -17421 -17537
rect -17535 -17729 -17523 -17695
rect -17433 -17729 -17421 -17695
rect -17535 -17735 -17421 -17729
rect -17677 -17825 -17665 -17791
rect -17575 -17825 -17563 -17791
rect -17828 -17922 -17762 -17910
rect -18100 -18069 -18002 -18057
rect -17828 -18069 -17820 -17922
rect -18100 -18143 -18088 -18069
rect -18014 -18143 -17820 -18069
rect -18100 -18155 -18002 -18143
rect -17828 -18279 -17820 -18143
rect -17769 -18279 -17762 -17922
rect -17677 -17983 -17563 -17825
rect -17282 -17743 -17216 -17727
rect -17282 -17777 -17266 -17743
rect -17232 -17777 -17216 -17743
rect -17677 -18017 -17665 -17983
rect -17575 -18017 -17563 -17983
rect -17677 -18175 -17563 -18017
rect -17677 -18209 -17665 -18175
rect -17575 -18209 -17563 -18175
rect -17677 -18215 -17563 -18209
rect -17535 -17887 -17421 -17881
rect -17535 -17921 -17523 -17887
rect -17433 -17921 -17421 -17887
rect -17535 -18079 -17421 -17921
rect -17535 -18113 -17523 -18079
rect -17433 -18113 -17421 -18079
rect -17828 -18291 -17762 -18279
rect -17535 -18271 -17421 -18113
rect -17535 -18305 -17523 -18271
rect -17433 -18305 -17421 -18271
rect -17535 -18311 -17421 -18305
rect -17387 -17886 -17321 -17827
rect -17387 -17920 -17371 -17886
rect -17337 -17920 -17321 -17886
rect -18065 -18385 -17995 -18379
rect -17995 -18396 -17893 -18385
rect -17387 -18396 -17321 -17920
rect -17995 -18455 -17321 -18396
rect -18065 -18461 -17995 -18455
rect -17964 -18462 -17321 -18455
rect -18099 -18515 -18010 -18509
rect -17282 -18514 -17216 -17777
rect -17182 -17785 -16982 -17388
rect -16924 -17708 -16850 -17696
rect -17188 -17791 -16988 -17785
rect -17188 -17825 -17176 -17791
rect -17000 -17825 -16988 -17791
rect -17188 -17831 -16988 -17825
rect -16924 -17907 -16917 -17708
rect -16856 -17907 -16850 -17708
rect -16924 -17919 -16850 -17907
rect -17054 -18167 -16968 -18151
rect -17054 -18219 -17036 -18167
rect -16984 -18175 -16968 -18167
rect -16916 -18175 -16872 -17919
rect -16984 -18211 -16872 -18175
rect -16984 -18219 -16968 -18211
rect -17054 -18237 -16968 -18219
rect -17964 -18515 -17216 -18514
rect -18010 -18580 -17216 -18515
rect -18010 -18604 -17834 -18580
rect -18099 -18610 -18010 -18604
rect -17535 -18665 -16984 -18663
rect -21033 -18736 -20924 -18717
rect -21074 -18748 -20924 -18736
rect -19383 -18771 -19377 -18705
rect -19311 -18771 -19305 -18705
rect -17535 -18711 -16983 -18665
rect -17535 -18745 -17523 -18711
rect -17433 -18716 -16983 -18711
rect -17433 -18745 -16982 -18716
rect -22595 -18795 -21060 -18779
rect -22595 -18829 -21557 -18795
rect -21331 -18829 -21111 -18795
rect -21077 -18829 -21060 -18795
rect -17535 -18788 -16982 -18745
rect -22595 -18848 -21060 -18829
rect -17677 -18807 -17563 -18801
rect -17677 -18841 -17665 -18807
rect -17575 -18841 -17563 -18807
rect -20406 -18914 -20340 -18908
rect -20406 -18916 -20399 -18914
rect -21574 -18964 -20399 -18916
rect -21574 -19000 -21061 -18964
rect -20406 -18966 -20399 -18964
rect -20347 -18966 -20340 -18914
rect -20406 -18972 -20340 -18966
rect -17677 -18999 -17563 -18841
rect -21722 -19074 -21602 -19014
rect -21722 -19109 -21678 -19074
rect -21941 -19161 -21935 -19109
rect -21883 -19161 -21678 -19109
rect -21722 -19165 -21678 -19161
rect -21644 -19137 -21602 -19074
rect -21574 -19022 -21122 -19000
rect -21574 -19099 -21510 -19022
rect -21476 -19099 -21318 -19022
rect -21284 -19028 -21122 -19022
rect -21284 -19040 -21116 -19028
rect -21284 -19099 -21156 -19040
rect -21574 -19105 -21156 -19099
rect -21644 -19143 -21364 -19137
rect -21644 -19165 -21606 -19143
rect -21722 -19222 -21606 -19165
rect -21572 -19222 -21414 -19143
rect -21380 -19222 -21364 -19143
rect -21722 -19228 -21364 -19222
rect -21318 -19216 -21156 -19105
rect -21122 -19216 -21116 -19040
rect -21318 -19228 -21116 -19216
rect -21075 -19040 -20925 -19028
rect -21075 -19216 -21068 -19040
rect -21034 -19064 -20925 -19040
rect -17677 -19033 -17665 -18999
rect -17575 -19033 -17563 -18999
rect -21034 -19065 -20651 -19064
rect -21034 -19197 -20966 -19065
rect -20932 -19153 -20651 -19065
rect -20562 -19153 -20556 -19064
rect -20932 -19197 -20925 -19153
rect -21034 -19216 -20925 -19197
rect -21075 -19228 -20925 -19216
rect -17677 -19191 -17563 -19033
rect -17535 -18903 -17421 -18788
rect -17535 -18937 -17523 -18903
rect -17433 -18937 -17421 -18903
rect -17535 -19095 -17421 -18937
rect -17535 -19129 -17523 -19095
rect -17433 -19129 -17421 -19095
rect -17182 -18959 -16982 -18788
rect -16772 -18812 -16703 -17388
rect -16652 -18650 -16583 -15968
rect -16492 -18150 -16423 -14648
rect -14806 -17799 -14758 -13976
rect -11441 -14057 -11365 -13973
rect -10855 -14032 -10779 -13973
rect -14708 -14088 -14656 -14082
rect -14708 -14146 -14656 -14140
rect -14808 -17807 -14756 -17799
rect -15983 -17855 -14756 -17807
rect -15983 -17891 -15470 -17855
rect -14808 -17863 -14756 -17855
rect -16131 -17965 -16011 -17905
rect -16131 -17988 -16087 -17965
rect -16344 -18040 -16338 -17988
rect -16286 -18040 -16087 -17988
rect -16131 -18056 -16087 -18040
rect -16053 -18028 -16011 -17965
rect -15983 -17913 -15531 -17891
rect -15983 -17990 -15919 -17913
rect -15885 -17990 -15727 -17913
rect -15693 -17919 -15531 -17913
rect -15693 -17931 -15525 -17919
rect -15693 -17990 -15565 -17931
rect -15983 -17996 -15565 -17990
rect -16053 -18034 -15773 -18028
rect -16053 -18056 -16015 -18034
rect -16131 -18113 -16015 -18056
rect -15981 -18113 -15823 -18034
rect -15789 -18113 -15773 -18034
rect -16131 -18119 -15773 -18113
rect -15727 -18107 -15565 -17996
rect -15531 -18107 -15525 -17931
rect -15727 -18119 -15525 -18107
rect -15484 -17931 -15334 -17919
rect -15484 -18107 -15477 -17931
rect -15443 -17956 -15334 -17931
rect -15443 -18088 -15375 -17956
rect -15341 -18045 -15052 -17956
rect -14963 -18045 -14957 -17956
rect -15341 -18088 -15334 -18045
rect -15443 -18107 -15334 -18088
rect -15484 -18119 -15334 -18107
rect -16492 -18166 -15470 -18150
rect -16492 -18200 -15967 -18166
rect -15741 -18200 -15521 -18166
rect -15487 -18200 -15470 -18166
rect -16492 -18219 -15470 -18200
rect -14706 -18307 -14658 -14146
rect -12501 -14193 -12175 -14181
rect -12501 -14223 -12295 -14193
rect -12501 -15345 -12473 -14223
rect -12401 -14227 -12295 -14223
rect -12193 -14227 -12175 -14193
rect -12401 -14385 -12175 -14227
rect -11925 -14193 -11778 -14181
rect -11925 -14227 -11904 -14193
rect -11837 -14227 -11778 -14193
rect -12401 -14419 -12295 -14385
rect -12193 -14419 -12175 -14385
rect -12401 -14435 -12175 -14419
rect -12137 -14289 -11958 -14273
rect -12137 -14323 -12111 -14289
rect -11987 -14323 -11958 -14289
rect -12401 -15137 -12367 -14435
rect -12137 -14481 -11958 -14323
rect -11925 -14385 -11778 -14227
rect -11543 -14194 -11334 -14057
rect -5969 -14065 -5963 -13983
rect -5881 -14065 -3716 -13983
rect -10855 -14114 -10779 -14108
rect -4932 -14122 -4271 -14103
rect -6954 -14142 -6902 -14136
rect -11543 -14228 -11413 -14194
rect -11450 -14259 -11413 -14228
rect -11358 -14259 -11334 -14194
rect -11280 -14193 -11001 -14184
rect -11280 -14227 -11264 -14193
rect -11158 -14222 -11001 -14193
rect -11158 -14227 -11070 -14222
rect -11280 -14239 -11070 -14227
rect -11450 -14270 -11334 -14259
rect -11291 -14289 -11223 -14273
rect -11291 -14323 -11279 -14289
rect -11245 -14323 -11223 -14289
rect -11925 -14419 -11904 -14385
rect -11837 -14419 -11778 -14385
rect -11925 -14435 -11778 -14419
rect -11603 -14361 -11333 -14344
rect -11603 -14441 -11584 -14361
rect -11516 -14441 -11333 -14361
rect -11603 -14459 -11333 -14441
rect -12137 -14515 -12112 -14481
rect -11988 -14515 -11958 -14481
rect -12322 -14577 -12175 -14561
rect -12322 -14611 -12295 -14577
rect -12193 -14611 -12175 -14577
rect -12322 -14769 -12175 -14611
rect -12322 -14803 -12295 -14769
rect -12193 -14803 -12175 -14769
rect -12322 -14961 -12175 -14803
rect -12322 -14995 -12296 -14961
rect -12194 -14995 -12175 -14961
rect -12322 -15011 -12175 -14995
rect -12137 -14673 -11958 -14515
rect -11603 -14561 -11504 -14529
rect -12137 -14707 -12112 -14673
rect -11988 -14707 -11958 -14673
rect -12137 -14865 -11958 -14707
rect -12137 -14899 -12112 -14865
rect -11988 -14899 -11958 -14865
rect -12137 -15057 -11958 -14899
rect -11914 -14577 -11822 -14561
rect -11914 -14611 -11897 -14577
rect -11837 -14611 -11822 -14577
rect -11914 -14769 -11822 -14611
rect -11914 -14803 -11880 -14769
rect -11837 -14803 -11822 -14769
rect -11914 -14961 -11822 -14803
rect -11914 -14995 -11897 -14961
rect -11837 -14995 -11822 -14961
rect -11914 -15011 -11822 -14995
rect -11603 -14675 -11585 -14561
rect -11532 -14675 -11504 -14561
rect -12137 -15091 -12112 -15057
rect -11988 -15091 -11958 -15057
rect -12401 -15153 -12175 -15137
rect -12401 -15187 -12298 -15153
rect -12196 -15187 -12175 -15153
rect -12401 -15345 -12175 -15187
rect -12137 -15249 -11958 -15091
rect -12137 -15283 -12112 -15249
rect -11988 -15283 -11958 -15249
rect -12137 -15299 -11958 -15283
rect -11925 -15153 -11778 -15137
rect -11925 -15187 -11903 -15153
rect -11837 -15187 -11778 -15153
rect -12501 -15379 -12298 -15345
rect -12196 -15379 -12175 -15345
rect -12501 -15391 -12175 -15379
rect -11925 -15345 -11778 -15187
rect -11603 -15148 -11504 -14675
rect -11603 -15281 -11577 -15148
rect -11524 -15281 -11504 -15148
rect -11603 -15318 -11504 -15281
rect -11419 -15332 -11333 -14459
rect -11291 -14481 -11223 -14323
rect -11092 -14370 -11070 -14239
rect -11194 -14385 -11070 -14370
rect -11194 -14419 -11178 -14385
rect -11144 -14419 -11070 -14385
rect -11194 -14435 -11070 -14419
rect -11291 -14515 -11279 -14481
rect -11245 -14515 -11223 -14481
rect -11291 -14673 -11223 -14515
rect -11291 -14707 -11279 -14673
rect -11245 -14707 -11223 -14673
rect -11291 -14723 -11223 -14707
rect -11190 -14577 -11126 -14561
rect -11190 -14611 -11178 -14577
rect -11144 -14611 -11126 -14577
rect -11190 -14769 -11126 -14611
rect -11190 -14803 -11178 -14769
rect -11144 -14803 -11126 -14769
rect -11291 -14865 -11223 -14849
rect -11291 -14899 -11278 -14865
rect -11244 -14899 -11223 -14865
rect -11291 -15057 -11223 -14899
rect -11190 -14961 -11126 -14803
rect -11190 -14995 -11178 -14961
rect -11144 -14995 -11126 -14961
rect -11190 -15008 -11126 -14995
rect -11092 -14825 -11070 -14435
rect -11024 -14825 -11001 -14222
rect -11092 -14885 -11081 -14825
rect -11021 -14885 -11001 -14825
rect -11291 -15091 -11279 -15057
rect -11245 -15091 -11223 -15057
rect -11291 -15249 -11223 -15091
rect -11092 -15136 -11070 -14885
rect -11195 -15153 -11070 -15136
rect -11195 -15187 -11178 -15153
rect -11144 -15187 -11070 -15153
rect -11195 -15201 -11070 -15187
rect -11291 -15283 -11279 -15249
rect -11245 -15283 -11223 -15249
rect -11291 -15299 -11223 -15283
rect -11092 -15331 -11070 -15201
rect -11925 -15379 -11903 -15345
rect -11801 -15379 -11778 -15345
rect -11925 -15391 -11778 -15379
rect -11464 -15537 -11321 -15332
rect -11280 -15345 -11070 -15331
rect -11024 -15345 -11001 -14885
rect -11280 -15379 -11264 -15345
rect -11158 -15379 -11001 -15345
rect -11280 -15386 -11001 -15379
rect -10850 -14331 -10795 -14325
rect -12730 -15586 -12656 -15570
rect -12612 -15586 -11481 -15582
rect -12730 -15658 -12724 -15586
rect -12652 -15594 -11481 -15586
rect -12652 -15658 -11567 -15594
rect -12730 -15666 -12656 -15658
rect -12612 -15668 -11567 -15658
rect -11493 -15668 -11481 -15594
rect -12612 -15674 -11481 -15668
rect -12566 -15738 -12440 -15728
rect -11442 -15738 -11343 -15537
rect -12612 -15837 -12555 -15738
rect -12456 -15837 -11343 -15738
rect -12566 -15848 -12440 -15837
rect -14618 -16016 -14612 -15964
rect -14560 -16016 -14554 -15964
rect -15982 -18355 -14658 -18307
rect -15982 -18391 -15469 -18355
rect -16130 -18465 -16010 -18405
rect -16130 -18497 -16086 -18465
rect -16350 -18549 -16344 -18497
rect -16292 -18549 -16086 -18497
rect -16130 -18556 -16086 -18549
rect -16052 -18528 -16010 -18465
rect -15982 -18413 -15530 -18391
rect -15982 -18490 -15918 -18413
rect -15884 -18490 -15726 -18413
rect -15692 -18419 -15530 -18413
rect -15692 -18431 -15524 -18419
rect -15692 -18490 -15564 -18431
rect -15982 -18496 -15564 -18490
rect -16052 -18534 -15772 -18528
rect -16052 -18556 -16014 -18534
rect -16130 -18613 -16014 -18556
rect -15980 -18613 -15822 -18534
rect -15788 -18613 -15772 -18534
rect -16130 -18619 -15772 -18613
rect -15726 -18607 -15564 -18496
rect -15530 -18607 -15524 -18431
rect -15726 -18619 -15524 -18607
rect -15483 -18431 -15333 -18419
rect -15483 -18607 -15476 -18431
rect -15442 -18449 -15333 -18431
rect -15442 -18456 -15059 -18449
rect -15442 -18588 -15374 -18456
rect -15340 -18538 -15059 -18456
rect -14970 -18538 -14964 -18449
rect -15340 -18588 -15333 -18538
rect -15442 -18607 -15333 -18588
rect -15483 -18619 -15333 -18607
rect -16652 -18666 -15469 -18650
rect -16652 -18700 -15966 -18666
rect -15740 -18700 -15520 -18666
rect -15486 -18700 -15469 -18666
rect -16652 -18719 -15469 -18700
rect -14610 -18787 -14562 -16016
rect -14496 -16186 -14444 -16180
rect -14496 -16244 -14444 -16238
rect -16772 -18881 -16502 -18812
rect -17182 -19028 -16712 -18959
rect -17535 -19135 -17421 -19129
rect -17677 -19225 -17665 -19191
rect -17575 -19225 -17563 -19191
rect -22701 -19275 -21061 -19259
rect -22701 -19309 -21558 -19275
rect -21332 -19309 -21112 -19275
rect -21078 -19309 -21061 -19275
rect -22701 -19328 -21061 -19309
rect -17828 -19322 -17762 -19310
rect -20410 -19416 -20404 -19414
rect -21574 -19464 -20404 -19416
rect -21574 -19500 -21061 -19464
rect -20410 -19466 -20404 -19464
rect -20352 -19466 -20346 -19414
rect -18098 -19475 -18000 -19463
rect -17828 -19475 -17820 -19322
rect -21722 -19574 -21602 -19514
rect -21722 -19631 -21678 -19574
rect -21941 -19683 -21935 -19631
rect -21883 -19665 -21678 -19631
rect -21644 -19637 -21602 -19574
rect -21574 -19522 -21122 -19500
rect -21574 -19599 -21510 -19522
rect -21476 -19599 -21318 -19522
rect -21284 -19528 -21122 -19522
rect -21284 -19540 -21116 -19528
rect -21284 -19599 -21156 -19540
rect -21574 -19605 -21156 -19599
rect -21644 -19643 -21364 -19637
rect -21644 -19665 -21606 -19643
rect -21883 -19683 -21606 -19665
rect -21722 -19722 -21606 -19683
rect -21572 -19722 -21414 -19643
rect -21380 -19722 -21364 -19643
rect -21722 -19728 -21364 -19722
rect -21318 -19716 -21156 -19605
rect -21122 -19716 -21116 -19540
rect -21318 -19728 -21116 -19716
rect -21075 -19540 -20925 -19528
rect -21075 -19716 -21068 -19540
rect -21034 -19565 -20925 -19540
rect -18098 -19549 -18086 -19475
rect -18012 -19549 -17820 -19475
rect -18098 -19561 -18000 -19549
rect -21034 -19697 -20966 -19565
rect -20932 -19571 -20925 -19565
rect -20932 -19660 -20655 -19571
rect -20566 -19660 -20560 -19571
rect -18024 -19622 -17942 -19614
rect -20932 -19697 -20925 -19660
rect -18024 -19685 -18016 -19622
rect -17953 -19685 -17942 -19622
rect -18024 -19692 -17942 -19685
rect -17828 -19679 -17820 -19549
rect -17769 -19679 -17762 -19322
rect -17677 -19383 -17563 -19225
rect -17282 -19143 -17216 -19127
rect -17282 -19177 -17266 -19143
rect -17232 -19177 -17216 -19143
rect -17677 -19417 -17665 -19383
rect -17575 -19417 -17563 -19383
rect -17677 -19575 -17563 -19417
rect -17677 -19609 -17665 -19575
rect -17575 -19609 -17563 -19575
rect -17677 -19615 -17563 -19609
rect -17535 -19287 -17421 -19281
rect -17535 -19321 -17523 -19287
rect -17433 -19321 -17421 -19287
rect -17535 -19479 -17421 -19321
rect -17535 -19513 -17523 -19479
rect -17433 -19513 -17421 -19479
rect -17828 -19691 -17762 -19679
rect -17535 -19671 -17421 -19513
rect -21034 -19716 -20925 -19697
rect -21075 -19728 -20925 -19716
rect -22813 -19775 -21061 -19759
rect -22813 -19809 -21558 -19775
rect -21332 -19809 -21112 -19775
rect -21078 -19809 -21061 -19775
rect -22813 -19828 -21061 -19809
rect -18016 -19780 -17953 -19692
rect -17535 -19705 -17523 -19671
rect -17433 -19705 -17421 -19671
rect -17535 -19711 -17421 -19705
rect -17387 -19286 -17321 -19227
rect -17387 -19320 -17371 -19286
rect -17337 -19320 -17321 -19286
rect -17387 -19780 -17321 -19320
rect -18016 -19846 -17321 -19780
rect -18016 -19847 -17953 -19846
rect -20324 -19894 -20272 -19888
rect -21574 -19944 -20324 -19896
rect -21574 -19980 -21061 -19944
rect -17282 -19898 -17216 -19177
rect -17182 -19185 -16982 -19028
rect -16924 -19108 -16850 -19096
rect -17188 -19191 -16988 -19185
rect -17188 -19225 -17176 -19191
rect -17000 -19225 -16988 -19191
rect -17188 -19231 -16988 -19225
rect -16924 -19307 -16917 -19108
rect -16856 -19307 -16850 -19108
rect -16924 -19319 -16850 -19307
rect -16918 -19609 -16872 -19319
rect -16934 -19622 -16854 -19609
rect -16934 -19674 -16921 -19622
rect -16869 -19674 -16854 -19622
rect -16934 -19689 -16854 -19674
rect -16781 -19628 -16712 -19028
rect -16571 -19128 -16502 -18881
rect -15983 -18835 -14562 -18787
rect -15983 -18871 -15470 -18835
rect -16131 -18945 -16011 -18885
rect -16131 -18980 -16087 -18945
rect -16350 -19032 -16344 -18980
rect -16292 -19032 -16087 -18980
rect -16131 -19036 -16087 -19032
rect -16053 -19008 -16011 -18945
rect -15983 -18893 -15531 -18871
rect -15983 -18970 -15919 -18893
rect -15885 -18970 -15727 -18893
rect -15693 -18899 -15531 -18893
rect -15693 -18911 -15525 -18899
rect -15693 -18970 -15565 -18911
rect -15983 -18976 -15565 -18970
rect -16053 -19014 -15773 -19008
rect -16053 -19036 -16015 -19014
rect -16131 -19093 -16015 -19036
rect -15981 -19093 -15823 -19014
rect -15789 -19093 -15773 -19014
rect -16131 -19099 -15773 -19093
rect -15727 -19087 -15565 -18976
rect -15531 -19087 -15525 -18911
rect -15727 -19099 -15525 -19087
rect -15484 -18911 -15334 -18899
rect -15484 -19087 -15477 -18911
rect -15443 -18935 -15334 -18911
rect -15443 -18936 -15060 -18935
rect -15443 -19068 -15375 -18936
rect -15341 -19024 -15060 -18936
rect -14971 -19024 -14965 -18935
rect -15341 -19068 -15334 -19024
rect -15443 -19087 -15334 -19068
rect -15484 -19099 -15334 -19087
rect -16571 -19130 -16288 -19128
rect -16571 -19146 -15470 -19130
rect -16571 -19180 -15967 -19146
rect -15741 -19180 -15521 -19146
rect -15487 -19180 -15470 -19146
rect -16571 -19197 -15470 -19180
rect -16402 -19199 -15470 -19197
rect -14494 -19287 -14446 -16244
rect -10850 -16457 -10795 -14386
rect -10307 -14771 -10252 -14765
rect -10849 -16681 -10797 -16457
rect -11453 -16770 -10779 -16681
rect -11453 -16873 -11364 -16770
rect -10307 -16774 -10252 -14826
rect -6954 -15246 -6902 -14194
rect -4932 -14156 -4768 -14122
rect -4542 -14156 -4322 -14122
rect -4288 -14156 -4271 -14122
rect -4932 -14172 -4271 -14156
rect -4932 -14203 -4869 -14172
rect -4932 -14209 -4574 -14203
rect -4932 -14248 -4816 -14209
rect -5026 -14254 -4816 -14248
rect -4910 -14266 -4816 -14254
rect -4910 -14357 -4888 -14266
rect -4854 -14288 -4816 -14266
rect -4782 -14288 -4624 -14209
rect -4590 -14288 -4574 -14209
rect -4854 -14294 -4574 -14288
rect -4528 -14215 -4326 -14203
rect -4854 -14357 -4812 -14294
rect -4528 -14326 -4366 -14215
rect -4910 -14370 -4812 -14357
rect -5026 -14376 -4812 -14370
rect -4932 -14417 -4812 -14376
rect -4784 -14332 -4366 -14326
rect -4784 -14409 -4720 -14332
rect -4686 -14409 -4528 -14332
rect -4494 -14391 -4366 -14332
rect -4332 -14391 -4326 -14215
rect -4494 -14403 -4326 -14391
rect -4285 -14215 -4135 -14203
rect -4285 -14391 -4278 -14215
rect -4244 -14234 -4135 -14215
rect -4244 -14366 -4176 -14234
rect -4142 -14250 -4135 -14234
rect -4142 -14347 -4004 -14250
rect -3907 -14347 -3901 -14250
rect -4142 -14366 -4135 -14347
rect -4244 -14391 -4135 -14366
rect -4285 -14403 -4135 -14391
rect -4494 -14409 -4332 -14403
rect -4784 -14431 -4332 -14409
rect -3798 -14431 -3716 -14065
rect -6966 -15248 -6902 -15246
rect -8135 -15296 -6902 -15248
rect -8135 -15332 -7622 -15296
rect -6966 -15298 -6902 -15296
rect -6834 -14490 -6782 -14484
rect -8283 -15406 -8163 -15346
rect -8283 -15429 -8239 -15406
rect -8496 -15481 -8490 -15429
rect -8438 -15481 -8239 -15429
rect -8690 -15496 -8594 -15486
rect -8690 -15568 -8676 -15496
rect -8604 -15568 -8594 -15496
rect -8283 -15497 -8239 -15481
rect -8205 -15469 -8163 -15406
rect -8135 -15354 -7683 -15332
rect -8135 -15431 -8071 -15354
rect -8037 -15431 -7879 -15354
rect -7845 -15360 -7683 -15354
rect -7845 -15372 -7677 -15360
rect -7845 -15431 -7717 -15372
rect -8135 -15437 -7717 -15431
rect -8205 -15475 -7925 -15469
rect -8205 -15497 -8167 -15475
rect -8283 -15554 -8167 -15497
rect -8133 -15554 -7975 -15475
rect -7941 -15554 -7925 -15475
rect -8283 -15560 -7925 -15554
rect -7879 -15548 -7717 -15437
rect -7683 -15548 -7677 -15372
rect -7879 -15560 -7677 -15548
rect -7636 -15372 -7486 -15360
rect -7636 -15548 -7629 -15372
rect -7595 -15397 -7486 -15372
rect -7595 -15529 -7527 -15397
rect -7493 -15486 -7204 -15397
rect -7115 -15486 -7109 -15397
rect -7493 -15529 -7486 -15486
rect -7595 -15548 -7486 -15529
rect -7636 -15560 -7486 -15548
rect -8690 -15586 -8594 -15568
rect -8690 -15588 -8476 -15586
rect -8676 -15591 -8476 -15588
rect -8676 -15607 -7622 -15591
rect -8676 -15641 -8119 -15607
rect -7893 -15641 -7673 -15607
rect -7639 -15641 -7622 -15607
rect -8676 -15658 -7622 -15641
rect -8554 -15660 -7622 -15658
rect -6834 -15746 -6782 -14542
rect -5048 -14494 -4864 -14446
rect -5048 -14566 -5008 -14494
rect -4936 -14543 -4864 -14494
rect -4784 -14491 -3716 -14431
rect -4784 -14515 -3899 -14491
rect -4936 -14562 -4271 -14543
rect -4936 -14566 -4768 -14562
rect -5048 -14596 -4768 -14566
rect -4542 -14596 -4322 -14562
rect -4288 -14596 -4271 -14562
rect -5048 -14612 -4271 -14596
rect -3958 -14557 -3899 -14515
rect -3833 -14556 -3716 -14491
rect -3833 -14557 -3774 -14556
rect -3958 -14612 -3774 -14557
rect -4932 -14649 -4574 -14643
rect -4932 -14706 -4816 -14649
rect -4932 -14797 -4888 -14706
rect -4854 -14728 -4816 -14706
rect -4782 -14728 -4624 -14649
rect -4590 -14728 -4574 -14649
rect -4854 -14734 -4574 -14728
rect -4528 -14655 -4326 -14643
rect -4854 -14797 -4812 -14734
rect -4528 -14766 -4366 -14655
rect -6662 -14860 -6614 -14850
rect -4932 -14853 -4812 -14797
rect -6674 -14870 -6600 -14860
rect -6674 -14922 -6664 -14870
rect -6612 -14922 -6600 -14870
rect -6674 -14930 -6600 -14922
rect -5048 -14887 -4812 -14853
rect -6970 -15748 -6782 -15746
rect -8134 -15796 -6782 -15748
rect -8134 -15832 -7621 -15796
rect -6970 -15798 -6782 -15796
rect -8282 -15906 -8162 -15846
rect -8282 -15938 -8238 -15906
rect -8502 -15990 -8496 -15938
rect -8444 -15990 -8238 -15938
rect -8282 -15997 -8238 -15990
rect -8204 -15969 -8162 -15906
rect -8134 -15854 -7682 -15832
rect -8134 -15931 -8070 -15854
rect -8036 -15931 -7878 -15854
rect -7844 -15860 -7682 -15854
rect -7844 -15872 -7676 -15860
rect -7844 -15931 -7716 -15872
rect -8134 -15937 -7716 -15931
rect -8204 -15975 -7924 -15969
rect -8204 -15997 -8166 -15975
rect -8282 -16054 -8166 -15997
rect -8132 -16054 -7974 -15975
rect -7940 -16054 -7924 -15975
rect -8282 -16060 -7924 -16054
rect -7878 -16048 -7716 -15937
rect -7682 -16048 -7676 -15872
rect -7878 -16060 -7676 -16048
rect -7635 -15872 -7485 -15860
rect -7635 -16048 -7628 -15872
rect -7594 -15890 -7485 -15872
rect -7594 -15897 -7211 -15890
rect -7594 -16029 -7526 -15897
rect -7492 -15979 -7211 -15897
rect -7122 -15979 -7116 -15890
rect -7492 -16029 -7485 -15979
rect -7594 -16048 -7485 -16029
rect -7635 -16060 -7485 -16048
rect -8554 -16091 -8482 -16087
rect -8554 -16107 -7621 -16091
rect -8554 -16140 -8118 -16107
rect -8570 -16141 -8118 -16140
rect -7892 -16141 -7672 -16107
rect -7638 -16141 -7621 -16107
rect -8570 -16152 -7621 -16141
rect -8570 -16224 -8554 -16152
rect -8482 -16160 -7621 -16152
rect -8482 -16224 -8470 -16160
rect -8570 -16236 -8470 -16224
rect -6662 -16228 -6614 -14930
rect -5048 -14991 -5020 -14887
rect -4916 -14991 -4812 -14887
rect -4784 -14772 -4366 -14766
rect -4784 -14849 -4720 -14772
rect -4686 -14849 -4528 -14772
rect -4494 -14831 -4366 -14772
rect -4332 -14831 -4326 -14655
rect -4494 -14843 -4326 -14831
rect -4285 -14655 -4135 -14643
rect -4285 -14831 -4278 -14655
rect -4244 -14674 -4135 -14655
rect -4244 -14806 -4176 -14674
rect -4142 -14806 -4135 -14674
rect -4244 -14831 -4135 -14806
rect -4285 -14843 -4135 -14831
rect -4494 -14849 -4332 -14843
rect -4784 -14871 -4332 -14849
rect -4784 -14941 -4271 -14871
rect -4784 -14975 -4768 -14941
rect -4542 -14975 -4322 -14941
rect -4288 -14975 -4271 -14941
rect -4784 -14991 -4271 -14975
rect -4232 -14883 -4135 -14843
rect -4232 -14980 -4004 -14883
rect -3907 -14980 -3901 -14883
rect -5048 -15022 -4812 -14991
rect -4232 -15022 -4135 -14980
rect -5048 -15023 -4574 -15022
rect -4932 -15028 -4574 -15023
rect -4932 -15085 -4816 -15028
rect -4932 -15176 -4888 -15085
rect -4854 -15107 -4816 -15085
rect -4782 -15107 -4624 -15028
rect -4590 -15107 -4574 -15028
rect -4854 -15113 -4574 -15107
rect -4528 -15034 -4326 -15022
rect -4854 -15176 -4812 -15113
rect -4528 -15145 -4366 -15034
rect -4932 -15236 -4812 -15176
rect -4784 -15151 -4366 -15145
rect -4784 -15228 -4720 -15151
rect -4686 -15228 -4528 -15151
rect -4494 -15210 -4366 -15151
rect -4332 -15210 -4326 -15034
rect -4494 -15222 -4326 -15210
rect -4285 -15034 -4135 -15022
rect -4285 -15210 -4278 -15034
rect -4244 -15053 -4135 -15034
rect -4244 -15185 -4176 -15053
rect -4142 -15185 -4135 -15053
rect -3654 -15182 -3570 -13944
rect -4244 -15210 -4135 -15185
rect -4285 -15222 -4135 -15210
rect -4494 -15228 -4332 -15222
rect -4784 -15250 -4332 -15228
rect -4044 -15250 -3570 -15182
rect -5048 -15306 -4864 -15265
rect -5048 -15378 -4966 -15306
rect -4894 -15362 -4864 -15306
rect -4784 -15266 -3570 -15250
rect -4784 -15334 -3774 -15266
rect -4894 -15378 -4271 -15362
rect -5048 -15381 -4271 -15378
rect -5048 -15415 -4768 -15381
rect -4542 -15415 -4322 -15381
rect -4288 -15415 -4271 -15381
rect -5048 -15431 -4271 -15415
rect -3958 -15431 -3774 -15334
rect -4932 -15468 -4574 -15462
rect -4932 -15525 -4816 -15468
rect -4932 -15616 -4888 -15525
rect -4854 -15547 -4816 -15525
rect -4782 -15547 -4624 -15468
rect -4590 -15547 -4574 -15468
rect -4854 -15553 -4574 -15547
rect -4528 -15474 -4326 -15462
rect -4854 -15616 -4812 -15553
rect -4528 -15585 -4366 -15474
rect -4932 -15672 -4812 -15616
rect -5048 -15706 -4812 -15672
rect -5048 -15810 -5020 -15706
rect -4916 -15810 -4812 -15706
rect -4784 -15591 -4366 -15585
rect -4784 -15668 -4720 -15591
rect -4686 -15668 -4528 -15591
rect -4494 -15650 -4366 -15591
rect -4332 -15650 -4326 -15474
rect -4494 -15662 -4326 -15650
rect -4285 -15474 -4135 -15462
rect -4285 -15650 -4278 -15474
rect -4244 -15493 -4135 -15474
rect -4244 -15625 -4176 -15493
rect -4142 -15625 -4135 -15493
rect -4244 -15650 -4135 -15625
rect -4285 -15662 -4135 -15650
rect -4494 -15668 -4332 -15662
rect -4784 -15690 -4332 -15668
rect -4784 -15760 -4271 -15690
rect -4784 -15794 -4768 -15760
rect -4542 -15794 -4322 -15760
rect -4288 -15794 -4271 -15760
rect -4784 -15810 -4271 -15794
rect -4232 -15702 -4135 -15662
rect -4232 -15799 -4004 -15702
rect -3907 -15799 -3901 -15702
rect -5048 -15841 -4812 -15810
rect -4232 -15841 -4135 -15799
rect -5048 -15842 -4574 -15841
rect -4932 -15847 -4574 -15842
rect -4932 -15904 -4816 -15847
rect -4932 -15995 -4888 -15904
rect -4854 -15926 -4816 -15904
rect -4782 -15926 -4624 -15847
rect -4590 -15926 -4574 -15847
rect -4854 -15932 -4574 -15926
rect -4528 -15853 -4326 -15841
rect -4854 -15995 -4812 -15932
rect -4528 -15964 -4366 -15853
rect -4932 -16055 -4812 -15995
rect -4784 -15970 -4366 -15964
rect -4784 -16047 -4720 -15970
rect -4686 -16047 -4528 -15970
rect -4494 -16029 -4366 -15970
rect -4332 -16029 -4326 -15853
rect -4494 -16041 -4326 -16029
rect -4285 -15853 -4135 -15841
rect -4285 -16029 -4278 -15853
rect -4244 -15872 -4135 -15853
rect -4244 -16004 -4176 -15872
rect -4142 -16004 -4135 -15872
rect -4244 -16029 -4135 -16004
rect -4285 -16041 -4135 -16029
rect -4494 -16047 -4332 -16041
rect -4784 -16069 -4332 -16047
rect -3520 -16069 -3436 -13818
rect -2216 -13878 -2096 -13818
rect -2216 -13969 -2172 -13878
rect -2138 -13941 -2096 -13878
rect -2068 -13826 -1616 -13804
rect -2068 -13903 -2004 -13826
rect -1970 -13903 -1812 -13826
rect -1778 -13832 -1616 -13826
rect -1778 -13844 -1610 -13832
rect -1778 -13903 -1650 -13844
rect -2068 -13909 -1650 -13903
rect -2138 -13947 -1858 -13941
rect -2138 -13969 -2100 -13947
rect -2216 -14026 -2100 -13969
rect -2066 -14026 -1908 -13947
rect -1874 -14026 -1858 -13947
rect -2216 -14031 -1858 -14026
rect -2332 -14032 -1858 -14031
rect -1812 -14020 -1650 -13909
rect -1616 -14020 -1610 -13844
rect -1812 -14032 -1610 -14020
rect -1569 -13844 -1419 -13832
rect -1569 -14020 -1562 -13844
rect -1528 -13869 -1419 -13844
rect -1528 -14001 -1460 -13869
rect -1426 -14001 -1419 -13869
rect -1528 -14020 -1419 -14001
rect -1569 -14032 -1419 -14020
rect -2332 -14063 -2096 -14032
rect -2332 -14167 -2304 -14063
rect -2200 -14167 -2096 -14063
rect -2332 -14201 -2096 -14167
rect -2216 -14257 -2096 -14201
rect -2216 -14348 -2172 -14257
rect -2138 -14320 -2096 -14257
rect -2068 -14079 -1555 -14063
rect -2068 -14113 -2052 -14079
rect -1826 -14113 -1606 -14079
rect -1572 -14113 -1555 -14079
rect -2068 -14183 -1555 -14113
rect -1516 -14074 -1419 -14032
rect -1516 -14171 -1288 -14074
rect -1191 -14171 -1185 -14074
rect -2068 -14205 -1616 -14183
rect -2068 -14282 -2004 -14205
rect -1970 -14282 -1812 -14205
rect -1778 -14211 -1616 -14205
rect -1516 -14211 -1419 -14171
rect -1778 -14223 -1610 -14211
rect -1778 -14282 -1650 -14223
rect -2068 -14288 -1650 -14282
rect -2138 -14326 -1858 -14320
rect -2138 -14348 -2100 -14326
rect -2216 -14405 -2100 -14348
rect -2066 -14405 -1908 -14326
rect -1874 -14405 -1858 -14326
rect -2216 -14411 -1858 -14405
rect -1812 -14399 -1650 -14288
rect -1616 -14399 -1610 -14223
rect -1812 -14411 -1610 -14399
rect -1569 -14223 -1419 -14211
rect -1569 -14399 -1562 -14223
rect -1528 -14248 -1419 -14223
rect -1528 -14380 -1460 -14248
rect -1426 -14380 -1419 -14248
rect -1528 -14399 -1419 -14380
rect -1569 -14411 -1419 -14399
rect -2332 -14458 -1555 -14442
rect -2332 -14492 -2052 -14458
rect -1826 -14492 -1606 -14458
rect -1572 -14492 -1555 -14458
rect -2332 -14494 -1555 -14492
rect -2332 -14566 -2288 -14494
rect -2216 -14511 -1555 -14494
rect -2216 -14566 -2148 -14511
rect -1242 -14539 -1058 -14442
rect -934 -14539 -850 -13492
rect -2332 -14608 -2148 -14566
rect -2068 -14623 -850 -14539
rect -2216 -14697 -2096 -14637
rect -2216 -14788 -2172 -14697
rect -2138 -14760 -2096 -14697
rect -2068 -14645 -1616 -14623
rect -2068 -14722 -2004 -14645
rect -1970 -14722 -1812 -14645
rect -1778 -14651 -1616 -14645
rect -1778 -14663 -1610 -14651
rect -1778 -14722 -1650 -14663
rect -2068 -14728 -1650 -14722
rect -2138 -14766 -1858 -14760
rect -2138 -14788 -2100 -14766
rect -2216 -14845 -2100 -14788
rect -2066 -14845 -1908 -14766
rect -1874 -14845 -1858 -14766
rect -2216 -14850 -1858 -14845
rect -2332 -14851 -1858 -14850
rect -1812 -14839 -1650 -14728
rect -1616 -14839 -1610 -14663
rect -1812 -14851 -1610 -14839
rect -1569 -14663 -1419 -14651
rect -1569 -14839 -1562 -14663
rect -1528 -14688 -1419 -14663
rect -1528 -14820 -1460 -14688
rect -1426 -14820 -1419 -14688
rect -1528 -14839 -1419 -14820
rect -1569 -14851 -1419 -14839
rect -2332 -14882 -2096 -14851
rect -2332 -14986 -2304 -14882
rect -2200 -14986 -2096 -14882
rect -2332 -15020 -2096 -14986
rect -2216 -15076 -2096 -15020
rect -2216 -15167 -2172 -15076
rect -2138 -15139 -2096 -15076
rect -2068 -14898 -1555 -14882
rect -2068 -14932 -2052 -14898
rect -1826 -14932 -1606 -14898
rect -1572 -14932 -1555 -14898
rect -2068 -15002 -1555 -14932
rect -1516 -14893 -1419 -14851
rect -1516 -14990 -1288 -14893
rect -1191 -14990 -1185 -14893
rect -2068 -15024 -1616 -15002
rect -2068 -15101 -2004 -15024
rect -1970 -15101 -1812 -15024
rect -1778 -15030 -1616 -15024
rect -1516 -15030 -1419 -14990
rect -1778 -15042 -1610 -15030
rect -1778 -15101 -1650 -15042
rect -2068 -15107 -1650 -15101
rect -2138 -15145 -1858 -15139
rect -2138 -15167 -2100 -15145
rect -2216 -15224 -2100 -15167
rect -2066 -15224 -1908 -15145
rect -1874 -15224 -1858 -15145
rect -2216 -15230 -1858 -15224
rect -1812 -15218 -1650 -15107
rect -1616 -15218 -1610 -15042
rect -1812 -15230 -1610 -15218
rect -1569 -15042 -1419 -15030
rect -1569 -15218 -1562 -15042
rect -1528 -15067 -1419 -15042
rect -1528 -15199 -1460 -15067
rect -1426 -15199 -1419 -15067
rect -1528 -15218 -1419 -15199
rect -1569 -15230 -1419 -15218
rect -2332 -15277 -1555 -15261
rect -2332 -15306 -2052 -15277
rect -2332 -15378 -2264 -15306
rect -2192 -15311 -2052 -15306
rect -1826 -15311 -1606 -15277
rect -1572 -15311 -1555 -15277
rect -2192 -15330 -1555 -15311
rect -2192 -15378 -2148 -15330
rect -1242 -15358 -1058 -15261
rect -768 -15358 -684 -13312
rect -2332 -15427 -2148 -15378
rect -2068 -15442 -684 -15358
rect -2216 -15516 -2096 -15456
rect -2216 -15607 -2172 -15516
rect -2138 -15579 -2096 -15516
rect -2068 -15464 -1616 -15442
rect -2068 -15541 -2004 -15464
rect -1970 -15541 -1812 -15464
rect -1778 -15470 -1616 -15464
rect -1778 -15482 -1610 -15470
rect -1778 -15541 -1650 -15482
rect -2068 -15547 -1650 -15541
rect -2138 -15585 -1858 -15579
rect -2138 -15607 -2100 -15585
rect -2216 -15664 -2100 -15607
rect -2066 -15664 -1908 -15585
rect -1874 -15664 -1858 -15585
rect -2216 -15669 -1858 -15664
rect -2332 -15670 -1858 -15669
rect -1812 -15658 -1650 -15547
rect -1616 -15658 -1610 -15482
rect -1812 -15670 -1610 -15658
rect -1569 -15482 -1419 -15470
rect -1569 -15658 -1562 -15482
rect -1528 -15507 -1419 -15482
rect -1528 -15639 -1460 -15507
rect -1426 -15639 -1419 -15507
rect -1528 -15658 -1419 -15639
rect -1569 -15670 -1419 -15658
rect -2332 -15701 -2096 -15670
rect -2332 -15805 -2304 -15701
rect -2200 -15805 -2096 -15701
rect -2332 -15839 -2096 -15805
rect -2216 -15895 -2096 -15839
rect -2216 -15986 -2172 -15895
rect -2138 -15958 -2096 -15895
rect -2068 -15717 -1555 -15701
rect -2068 -15751 -2052 -15717
rect -1826 -15751 -1606 -15717
rect -1572 -15751 -1555 -15717
rect -2068 -15821 -1555 -15751
rect -1516 -15712 -1419 -15670
rect -1516 -15809 -1288 -15712
rect -1191 -15809 -1185 -15712
rect -2068 -15843 -1616 -15821
rect -2068 -15920 -2004 -15843
rect -1970 -15920 -1812 -15843
rect -1778 -15849 -1616 -15843
rect -1516 -15849 -1419 -15809
rect -1778 -15861 -1610 -15849
rect -1778 -15920 -1650 -15861
rect -2068 -15926 -1650 -15920
rect -2138 -15964 -1858 -15958
rect -2138 -15986 -2100 -15964
rect -2216 -16043 -2100 -15986
rect -2066 -16043 -1908 -15964
rect -1874 -16043 -1858 -15964
rect -2216 -16049 -1858 -16043
rect -1812 -16037 -1650 -15926
rect -1616 -16037 -1610 -15861
rect -1812 -16049 -1610 -16037
rect -1569 -15861 -1419 -15849
rect -1569 -16037 -1562 -15861
rect -1528 -15886 -1419 -15861
rect -1528 -16018 -1460 -15886
rect -1426 -16018 -1419 -15886
rect -1528 -16037 -1419 -16018
rect -1569 -16049 -1419 -16037
rect -8135 -16276 -6614 -16228
rect -5048 -16125 -4864 -16084
rect -5048 -16195 -4995 -16125
rect -4925 -16181 -4864 -16125
rect -4784 -16153 -3436 -16069
rect -2332 -16096 -1555 -16080
rect -2332 -16125 -2052 -16096
rect -4925 -16195 -4271 -16181
rect -5048 -16200 -4271 -16195
rect -5048 -16234 -4768 -16200
rect -4542 -16234 -4322 -16200
rect -4288 -16234 -4271 -16200
rect -5048 -16250 -4271 -16234
rect -3958 -16250 -3774 -16153
rect -2332 -16195 -2285 -16125
rect -2215 -16130 -2052 -16125
rect -1826 -16130 -1606 -16096
rect -1572 -16130 -1555 -16096
rect -2215 -16149 -1555 -16130
rect -2215 -16195 -2148 -16149
rect -1242 -16177 -1058 -16080
rect -458 -16177 -374 -13150
rect -2332 -16246 -2148 -16195
rect -2068 -16261 -368 -16177
rect -8135 -16312 -7622 -16276
rect -4932 -16287 -4574 -16281
rect -8283 -16386 -8163 -16326
rect -8283 -16421 -8239 -16386
rect -8502 -16473 -8496 -16421
rect -8444 -16473 -8239 -16421
rect -8283 -16477 -8239 -16473
rect -8205 -16449 -8163 -16386
rect -8135 -16334 -7683 -16312
rect -8135 -16411 -8071 -16334
rect -8037 -16411 -7879 -16334
rect -7845 -16340 -7683 -16334
rect -7845 -16352 -7677 -16340
rect -7845 -16411 -7717 -16352
rect -8135 -16417 -7717 -16411
rect -8205 -16455 -7925 -16449
rect -8205 -16477 -8167 -16455
rect -8283 -16534 -8167 -16477
rect -8133 -16534 -7975 -16455
rect -7941 -16534 -7925 -16455
rect -8283 -16540 -7925 -16534
rect -7879 -16528 -7717 -16417
rect -7683 -16528 -7677 -16352
rect -7879 -16540 -7677 -16528
rect -7636 -16352 -7486 -16340
rect -7636 -16528 -7629 -16352
rect -7595 -16376 -7486 -16352
rect -4932 -16344 -4816 -16287
rect -7595 -16377 -7212 -16376
rect -7595 -16509 -7527 -16377
rect -7493 -16465 -7212 -16377
rect -7123 -16465 -7117 -16376
rect -4932 -16435 -4888 -16344
rect -4854 -16366 -4816 -16344
rect -4782 -16366 -4624 -16287
rect -4590 -16366 -4574 -16287
rect -4854 -16372 -4574 -16366
rect -4528 -16293 -4326 -16281
rect -4854 -16435 -4812 -16372
rect -4528 -16404 -4366 -16293
rect -7493 -16509 -7486 -16465
rect -4932 -16491 -4812 -16435
rect -7595 -16528 -7486 -16509
rect -7636 -16540 -7486 -16528
rect -5048 -16525 -4812 -16491
rect -8554 -16587 -7622 -16571
rect -8554 -16621 -8119 -16587
rect -7893 -16621 -7673 -16587
rect -7639 -16621 -7622 -16587
rect -8554 -16640 -7622 -16621
rect -5048 -16629 -5020 -16525
rect -4916 -16629 -4812 -16525
rect -4784 -16410 -4366 -16404
rect -4784 -16487 -4720 -16410
rect -4686 -16487 -4528 -16410
rect -4494 -16469 -4366 -16410
rect -4332 -16469 -4326 -16293
rect -4494 -16481 -4326 -16469
rect -4285 -16293 -4135 -16281
rect -4285 -16469 -4278 -16293
rect -4244 -16312 -4135 -16293
rect -4244 -16444 -4176 -16312
rect -4142 -16444 -4135 -16312
rect -4244 -16469 -4135 -16444
rect -4285 -16481 -4135 -16469
rect -4494 -16487 -4332 -16481
rect -4784 -16509 -4332 -16487
rect -4784 -16579 -4271 -16509
rect -4784 -16613 -4768 -16579
rect -4542 -16613 -4322 -16579
rect -4288 -16613 -4271 -16579
rect -4784 -16629 -4271 -16613
rect -4232 -16521 -4135 -16481
rect -2216 -16335 -2096 -16275
rect -2216 -16426 -2172 -16335
rect -2138 -16398 -2096 -16335
rect -2068 -16283 -1616 -16261
rect -2068 -16360 -2004 -16283
rect -1970 -16360 -1812 -16283
rect -1778 -16289 -1616 -16283
rect -1778 -16301 -1610 -16289
rect -1778 -16360 -1650 -16301
rect -2068 -16366 -1650 -16360
rect -2138 -16404 -1858 -16398
rect -2138 -16426 -2100 -16404
rect -2216 -16483 -2100 -16426
rect -2066 -16483 -1908 -16404
rect -1874 -16483 -1858 -16404
rect -2216 -16488 -1858 -16483
rect -2332 -16489 -1858 -16488
rect -1812 -16477 -1650 -16366
rect -1616 -16477 -1610 -16301
rect -1812 -16489 -1610 -16477
rect -1569 -16301 -1419 -16289
rect -1569 -16477 -1562 -16301
rect -1528 -16326 -1419 -16301
rect -1528 -16458 -1460 -16326
rect -1426 -16458 -1419 -16326
rect -1528 -16477 -1419 -16458
rect -1569 -16489 -1419 -16477
rect -2332 -16520 -2096 -16489
rect -4232 -16618 -4004 -16521
rect -3907 -16618 -3901 -16521
rect -8551 -16685 -8482 -16640
rect -5048 -16660 -4812 -16629
rect -4232 -16660 -4135 -16618
rect -2332 -16624 -2304 -16520
rect -2200 -16624 -2096 -16520
rect -2332 -16658 -2096 -16624
rect -5048 -16661 -4574 -16660
rect -4932 -16666 -4574 -16661
rect -4932 -16723 -4816 -16666
rect -8551 -16760 -8482 -16754
rect -12499 -17009 -12173 -16997
rect -12499 -17039 -12293 -17009
rect -12499 -18161 -12471 -17039
rect -12399 -17043 -12293 -17039
rect -12191 -17043 -12173 -17009
rect -12399 -17201 -12173 -17043
rect -11923 -17009 -11776 -16997
rect -11923 -17043 -11902 -17009
rect -11835 -17043 -11776 -17009
rect -12399 -17235 -12293 -17201
rect -12191 -17235 -12173 -17201
rect -12399 -17251 -12173 -17235
rect -12135 -17105 -11956 -17089
rect -12135 -17139 -12109 -17105
rect -11985 -17139 -11956 -17105
rect -12399 -17953 -12365 -17251
rect -12135 -17297 -11956 -17139
rect -11923 -17201 -11776 -17043
rect -11541 -17010 -11332 -16873
rect -11541 -17044 -11411 -17010
rect -11448 -17075 -11411 -17044
rect -11356 -17075 -11332 -17010
rect -11278 -17009 -10999 -17000
rect -11278 -17043 -11262 -17009
rect -11156 -17038 -10999 -17009
rect -11156 -17043 -11068 -17038
rect -11278 -17055 -11068 -17043
rect -11448 -17086 -11332 -17075
rect -11289 -17105 -11221 -17089
rect -11289 -17139 -11277 -17105
rect -11243 -17139 -11221 -17105
rect -11923 -17235 -11902 -17201
rect -11835 -17235 -11776 -17201
rect -11923 -17251 -11776 -17235
rect -11601 -17177 -11331 -17160
rect -11601 -17257 -11582 -17177
rect -11514 -17257 -11331 -17177
rect -11601 -17275 -11331 -17257
rect -12135 -17331 -12110 -17297
rect -11986 -17331 -11956 -17297
rect -12320 -17393 -12173 -17377
rect -12320 -17427 -12293 -17393
rect -12191 -17427 -12173 -17393
rect -12320 -17585 -12173 -17427
rect -12320 -17619 -12293 -17585
rect -12191 -17619 -12173 -17585
rect -12320 -17777 -12173 -17619
rect -12320 -17811 -12294 -17777
rect -12192 -17811 -12173 -17777
rect -12320 -17827 -12173 -17811
rect -12135 -17489 -11956 -17331
rect -11601 -17377 -11502 -17345
rect -12135 -17523 -12110 -17489
rect -11986 -17523 -11956 -17489
rect -12135 -17681 -11956 -17523
rect -12135 -17715 -12110 -17681
rect -11986 -17715 -11956 -17681
rect -12135 -17873 -11956 -17715
rect -11912 -17393 -11820 -17377
rect -11912 -17427 -11895 -17393
rect -11835 -17427 -11820 -17393
rect -11912 -17585 -11820 -17427
rect -11912 -17619 -11878 -17585
rect -11835 -17619 -11820 -17585
rect -11912 -17777 -11820 -17619
rect -11912 -17811 -11895 -17777
rect -11835 -17811 -11820 -17777
rect -11912 -17827 -11820 -17811
rect -11601 -17491 -11583 -17377
rect -11530 -17491 -11502 -17377
rect -12135 -17907 -12110 -17873
rect -11986 -17907 -11956 -17873
rect -12399 -17969 -12173 -17953
rect -12399 -18003 -12296 -17969
rect -12194 -18003 -12173 -17969
rect -12399 -18161 -12173 -18003
rect -12135 -18065 -11956 -17907
rect -12135 -18099 -12110 -18065
rect -11986 -18099 -11956 -18065
rect -12135 -18115 -11956 -18099
rect -11923 -17969 -11776 -17953
rect -11923 -18003 -11901 -17969
rect -11835 -18003 -11776 -17969
rect -12499 -18195 -12296 -18161
rect -12194 -18195 -12173 -18161
rect -12499 -18207 -12173 -18195
rect -11923 -18161 -11776 -18003
rect -11601 -17964 -11502 -17491
rect -11601 -18097 -11575 -17964
rect -11522 -18097 -11502 -17964
rect -11601 -18134 -11502 -18097
rect -11417 -18148 -11331 -17275
rect -11289 -17297 -11221 -17139
rect -11090 -17186 -11068 -17055
rect -11192 -17201 -11068 -17186
rect -11192 -17235 -11176 -17201
rect -11142 -17235 -11068 -17201
rect -11192 -17251 -11068 -17235
rect -11289 -17331 -11277 -17297
rect -11243 -17331 -11221 -17297
rect -11289 -17489 -11221 -17331
rect -11289 -17523 -11277 -17489
rect -11243 -17523 -11221 -17489
rect -11289 -17539 -11221 -17523
rect -11188 -17393 -11124 -17377
rect -11188 -17427 -11176 -17393
rect -11142 -17427 -11124 -17393
rect -11188 -17585 -11124 -17427
rect -11188 -17619 -11176 -17585
rect -11142 -17619 -11124 -17585
rect -11289 -17681 -11221 -17665
rect -11289 -17715 -11276 -17681
rect -11242 -17715 -11221 -17681
rect -11289 -17873 -11221 -17715
rect -11188 -17777 -11124 -17619
rect -11188 -17811 -11176 -17777
rect -11142 -17811 -11124 -17777
rect -11188 -17824 -11124 -17811
rect -11090 -17641 -11068 -17251
rect -11022 -17641 -10999 -17038
rect -11090 -17701 -11079 -17641
rect -11019 -17701 -10999 -17641
rect -11289 -17907 -11277 -17873
rect -11243 -17907 -11221 -17873
rect -11289 -18065 -11221 -17907
rect -11090 -17952 -11068 -17701
rect -11193 -17969 -11068 -17952
rect -11193 -18003 -11176 -17969
rect -11142 -18003 -11068 -17969
rect -11193 -18017 -11068 -18003
rect -11289 -18099 -11277 -18065
rect -11243 -18099 -11221 -18065
rect -11289 -18115 -11221 -18099
rect -11090 -18147 -11068 -18017
rect -11923 -18195 -11901 -18161
rect -11799 -18195 -11776 -18161
rect -11923 -18207 -11776 -18195
rect -11462 -18353 -11319 -18148
rect -11278 -18161 -11068 -18147
rect -11022 -18161 -10999 -17701
rect -11278 -18195 -11262 -18161
rect -11156 -18195 -10999 -18161
rect -11278 -18202 -10999 -18195
rect -12666 -18391 -12594 -18390
rect -12666 -18396 -11479 -18391
rect -12594 -18403 -11479 -18396
rect -12594 -18468 -11565 -18403
rect -12666 -18474 -11565 -18468
rect -12612 -18477 -11565 -18474
rect -11491 -18477 -11479 -18403
rect -12612 -18483 -11479 -18477
rect -11436 -18559 -11345 -18353
rect -12612 -18567 -11345 -18559
rect -12633 -18573 -11345 -18567
rect -12544 -18650 -11345 -18573
rect -12544 -18662 -12494 -18650
rect -12633 -18668 -12544 -18662
rect -15983 -19335 -14446 -19287
rect -15983 -19371 -15470 -19335
rect -16131 -19445 -16011 -19385
rect -16131 -19502 -16087 -19445
rect -16350 -19554 -16344 -19502
rect -16292 -19536 -16087 -19502
rect -16053 -19508 -16011 -19445
rect -15983 -19393 -15531 -19371
rect -15983 -19470 -15919 -19393
rect -15885 -19470 -15727 -19393
rect -15693 -19399 -15531 -19393
rect -15693 -19411 -15525 -19399
rect -15693 -19470 -15565 -19411
rect -15983 -19476 -15565 -19470
rect -16053 -19514 -15773 -19508
rect -16053 -19536 -16015 -19514
rect -16292 -19554 -16015 -19536
rect -16131 -19593 -16015 -19554
rect -15981 -19593 -15823 -19514
rect -15789 -19593 -15773 -19514
rect -16131 -19599 -15773 -19593
rect -15727 -19587 -15565 -19476
rect -15531 -19587 -15525 -19411
rect -15727 -19599 -15525 -19587
rect -15484 -19411 -15334 -19399
rect -15484 -19587 -15477 -19411
rect -15443 -19436 -15334 -19411
rect -15443 -19568 -15375 -19436
rect -15341 -19442 -15334 -19436
rect -15341 -19531 -15064 -19442
rect -14975 -19531 -14969 -19442
rect -15341 -19568 -15334 -19531
rect -15443 -19587 -15334 -19568
rect -15484 -19599 -15334 -19587
rect -10328 -19622 -10233 -16774
rect -8135 -16776 -5186 -16728
rect -8135 -16812 -7622 -16776
rect -8283 -16886 -8163 -16826
rect -8283 -16943 -8239 -16886
rect -8502 -16995 -8496 -16943
rect -8444 -16977 -8239 -16943
rect -8205 -16949 -8163 -16886
rect -8135 -16834 -7683 -16812
rect -8135 -16911 -8071 -16834
rect -8037 -16911 -7879 -16834
rect -7845 -16840 -7683 -16834
rect -7845 -16852 -7677 -16840
rect -7845 -16911 -7717 -16852
rect -8135 -16917 -7717 -16911
rect -8205 -16955 -7925 -16949
rect -8205 -16977 -8167 -16955
rect -8444 -16995 -8167 -16977
rect -8283 -17034 -8167 -16995
rect -8133 -17034 -7975 -16955
rect -7941 -17034 -7925 -16955
rect -8283 -17040 -7925 -17034
rect -7879 -17028 -7717 -16917
rect -7683 -17028 -7677 -16852
rect -7879 -17040 -7677 -17028
rect -7636 -16852 -7486 -16840
rect -7636 -17028 -7629 -16852
rect -7595 -16877 -7486 -16852
rect -7595 -17009 -7527 -16877
rect -7493 -16883 -7486 -16877
rect -7493 -16972 -7216 -16883
rect -7127 -16972 -7121 -16883
rect -7493 -17009 -7486 -16972
rect -7595 -17028 -7486 -17009
rect -7636 -17040 -7486 -17028
rect -8554 -17087 -7622 -17071
rect -8554 -17121 -8119 -17087
rect -7893 -17121 -7673 -17087
rect -7639 -17121 -7622 -17087
rect -8554 -17140 -7622 -17121
rect -8549 -17188 -8480 -17140
rect -5397 -17149 -5307 -17148
rect -5407 -17154 -5288 -17149
rect -8560 -17205 -8464 -17188
rect -8560 -17274 -8549 -17205
rect -8480 -17274 -8464 -17205
rect -8560 -17286 -8464 -17274
rect -8135 -17256 -5536 -17208
rect -5407 -17243 -5397 -17154
rect -5307 -17243 -5288 -17154
rect -5407 -17252 -5288 -17243
rect -8135 -17292 -7622 -17256
rect -8283 -17366 -8163 -17306
rect -8283 -17412 -8239 -17366
rect -8499 -17464 -8493 -17412
rect -8441 -17457 -8239 -17412
rect -8205 -17429 -8163 -17366
rect -8135 -17314 -7683 -17292
rect -8135 -17391 -8071 -17314
rect -8037 -17391 -7879 -17314
rect -7845 -17320 -7683 -17314
rect -7845 -17332 -7677 -17320
rect -7845 -17391 -7717 -17332
rect -8135 -17397 -7717 -17391
rect -8205 -17435 -7925 -17429
rect -8205 -17457 -8167 -17435
rect -8441 -17464 -8167 -17457
rect -8283 -17514 -8167 -17464
rect -8133 -17514 -7975 -17435
rect -7941 -17514 -7925 -17435
rect -8283 -17520 -7925 -17514
rect -7879 -17508 -7717 -17397
rect -7683 -17508 -7677 -17332
rect -7879 -17520 -7677 -17508
rect -7636 -17332 -7486 -17320
rect -7636 -17508 -7629 -17332
rect -7595 -17357 -7486 -17332
rect -7595 -17489 -7527 -17357
rect -7493 -17358 -7486 -17357
rect -7493 -17447 -7215 -17358
rect -7126 -17447 -7120 -17358
rect -7493 -17489 -7486 -17447
rect -7595 -17508 -7486 -17489
rect -7636 -17520 -7486 -17508
rect -8554 -17567 -7622 -17551
rect -8554 -17601 -8119 -17567
rect -7893 -17601 -7673 -17567
rect -7639 -17601 -7622 -17567
rect -8554 -17615 -7622 -17601
rect -8485 -17620 -7622 -17615
rect -8554 -17690 -8485 -17684
rect -8135 -17716 -5652 -17668
rect -8135 -17752 -7622 -17716
rect -8283 -17826 -8163 -17766
rect -8283 -17869 -8239 -17826
rect -8497 -17921 -8491 -17869
rect -8439 -17917 -8239 -17869
rect -8205 -17889 -8163 -17826
rect -8135 -17774 -7683 -17752
rect -8135 -17851 -8071 -17774
rect -8037 -17851 -7879 -17774
rect -7845 -17780 -7683 -17774
rect -7845 -17792 -7677 -17780
rect -7845 -17851 -7717 -17792
rect -8135 -17857 -7717 -17851
rect -8205 -17895 -7925 -17889
rect -8205 -17917 -8167 -17895
rect -8439 -17921 -8167 -17917
rect -8283 -17974 -8167 -17921
rect -8133 -17974 -7975 -17895
rect -7941 -17974 -7925 -17895
rect -8283 -17980 -7925 -17974
rect -7879 -17968 -7717 -17857
rect -7683 -17968 -7677 -17792
rect -7879 -17980 -7677 -17968
rect -7636 -17792 -7486 -17780
rect -7636 -17968 -7629 -17792
rect -7595 -17810 -7486 -17792
rect -7595 -17817 -7210 -17810
rect -7595 -17949 -7527 -17817
rect -7493 -17899 -7210 -17817
rect -7121 -17899 -7115 -17810
rect -7493 -17949 -7486 -17899
rect -7595 -17968 -7486 -17949
rect -7636 -17980 -7486 -17968
rect -8554 -18027 -7622 -18011
rect -8554 -18061 -8119 -18027
rect -7893 -18061 -7673 -18027
rect -7639 -18061 -7622 -18027
rect -8554 -18080 -7622 -18061
rect -8554 -18097 -8485 -18080
rect -8554 -18172 -8485 -18166
rect -8149 -18176 -5804 -18128
rect -8149 -18212 -7636 -18176
rect -8297 -18286 -8177 -18226
rect -8297 -18334 -8253 -18286
rect -8495 -18386 -8489 -18334
rect -8437 -18377 -8253 -18334
rect -8219 -18349 -8177 -18286
rect -8149 -18234 -7697 -18212
rect -8149 -18311 -8085 -18234
rect -8051 -18311 -7893 -18234
rect -7859 -18240 -7697 -18234
rect -7859 -18252 -7691 -18240
rect -7859 -18311 -7731 -18252
rect -8149 -18317 -7731 -18311
rect -8219 -18355 -7939 -18349
rect -8219 -18377 -8181 -18355
rect -8437 -18386 -8181 -18377
rect -8297 -18434 -8181 -18386
rect -8147 -18434 -7989 -18355
rect -7955 -18434 -7939 -18355
rect -8297 -18440 -7939 -18434
rect -7893 -18428 -7731 -18317
rect -7697 -18428 -7691 -18252
rect -7893 -18440 -7691 -18428
rect -7650 -18252 -7500 -18240
rect -7650 -18428 -7643 -18252
rect -7609 -18277 -7210 -18252
rect -7609 -18409 -7541 -18277
rect -7507 -18341 -7210 -18277
rect -7121 -18341 -7115 -18252
rect -7507 -18409 -7500 -18341
rect -7609 -18428 -7500 -18409
rect -7650 -18440 -7500 -18428
rect -8554 -18487 -7636 -18471
rect -8554 -18521 -8133 -18487
rect -7907 -18521 -7687 -18487
rect -7653 -18521 -7636 -18487
rect -8554 -18540 -7636 -18521
rect -8554 -18567 -8485 -18540
rect -8554 -18642 -8485 -18636
rect -8147 -18656 -5982 -18608
rect -8147 -18692 -7634 -18656
rect -8295 -18766 -8175 -18706
rect -8295 -18815 -8251 -18766
rect -8491 -18867 -8485 -18815
rect -8433 -18857 -8251 -18815
rect -8217 -18829 -8175 -18766
rect -8147 -18714 -7695 -18692
rect -8147 -18791 -8083 -18714
rect -8049 -18791 -7891 -18714
rect -7857 -18720 -7695 -18714
rect -7857 -18732 -7689 -18720
rect -7857 -18791 -7729 -18732
rect -8147 -18797 -7729 -18791
rect -8217 -18835 -7937 -18829
rect -8217 -18857 -8179 -18835
rect -8433 -18867 -8179 -18857
rect -8295 -18914 -8179 -18867
rect -8145 -18914 -7987 -18835
rect -7953 -18914 -7937 -18835
rect -8295 -18920 -7937 -18914
rect -7891 -18908 -7729 -18797
rect -7695 -18908 -7689 -18732
rect -7891 -18920 -7689 -18908
rect -7648 -18732 -7498 -18720
rect -7648 -18908 -7641 -18732
rect -7607 -18733 -7498 -18732
rect -7607 -18757 -7216 -18733
rect -7607 -18889 -7539 -18757
rect -7505 -18822 -7216 -18757
rect -7127 -18822 -7121 -18733
rect -7505 -18889 -7498 -18822
rect -7607 -18908 -7498 -18889
rect -7648 -18920 -7498 -18908
rect -8584 -18951 -8512 -18948
rect -8584 -18967 -7634 -18951
rect -8584 -19001 -8131 -18967
rect -7905 -19001 -7685 -18967
rect -7651 -19001 -7634 -18967
rect -8584 -19020 -7634 -19001
rect -8584 -19098 -8512 -19020
rect -8590 -19170 -8584 -19098
rect -8512 -19170 -8506 -19098
rect -16781 -19630 -16370 -19628
rect -16781 -19646 -15470 -19630
rect -16781 -19680 -15967 -19646
rect -15741 -19680 -15521 -19646
rect -15487 -19680 -15470 -19646
rect -16781 -19697 -15470 -19680
rect -16430 -19699 -15470 -19697
rect -11456 -19717 -10233 -19622
rect -15983 -19815 -14758 -19767
rect -15983 -19851 -15470 -19815
rect -20324 -19952 -20272 -19946
rect -17994 -19907 -17216 -19898
rect -17994 -19978 -17986 -19907
rect -17915 -19964 -17216 -19907
rect -16131 -19925 -16011 -19865
rect -17915 -19978 -17906 -19964
rect -16131 -19971 -16087 -19925
rect -21722 -20054 -21602 -19994
rect -21722 -20100 -21678 -20054
rect -21938 -20152 -21932 -20100
rect -21880 -20145 -21678 -20100
rect -21644 -20117 -21602 -20054
rect -21574 -20002 -21122 -19980
rect -17994 -19986 -17906 -19978
rect -21574 -20079 -21510 -20002
rect -21476 -20079 -21318 -20002
rect -21284 -20008 -21122 -20002
rect -21284 -20020 -21116 -20008
rect -21284 -20079 -21156 -20020
rect -21574 -20085 -21156 -20079
rect -21644 -20123 -21364 -20117
rect -21644 -20145 -21606 -20123
rect -21880 -20152 -21606 -20145
rect -21722 -20202 -21606 -20152
rect -21572 -20202 -21414 -20123
rect -21380 -20202 -21364 -20123
rect -21722 -20208 -21364 -20202
rect -21318 -20196 -21156 -20085
rect -21122 -20196 -21116 -20020
rect -21318 -20208 -21116 -20196
rect -21075 -20020 -20925 -20008
rect -21075 -20196 -21068 -20020
rect -21034 -20045 -20925 -20020
rect -16347 -20023 -16341 -19971
rect -16289 -20016 -16087 -19971
rect -16053 -19988 -16011 -19925
rect -15983 -19873 -15531 -19851
rect -14808 -19866 -14760 -19815
rect -11456 -19830 -11361 -19717
rect -15983 -19950 -15919 -19873
rect -15885 -19950 -15727 -19873
rect -15693 -19879 -15531 -19873
rect -15693 -19891 -15525 -19879
rect -15693 -19950 -15565 -19891
rect -15983 -19956 -15565 -19950
rect -16053 -19994 -15773 -19988
rect -16053 -20016 -16015 -19994
rect -16289 -20023 -16015 -20016
rect -21034 -20177 -20966 -20045
rect -20932 -20046 -20925 -20045
rect -20932 -20135 -20654 -20046
rect -20565 -20135 -20559 -20046
rect -17535 -20065 -16984 -20063
rect -17535 -20111 -16983 -20065
rect -16131 -20073 -16015 -20023
rect -15981 -20073 -15823 -19994
rect -15789 -20073 -15773 -19994
rect -16131 -20079 -15773 -20073
rect -15727 -20067 -15565 -19956
rect -15531 -20067 -15525 -19891
rect -15727 -20079 -15525 -20067
rect -15484 -19891 -15334 -19879
rect -15484 -20067 -15477 -19891
rect -15443 -19916 -15334 -19891
rect -15443 -20048 -15375 -19916
rect -15341 -19917 -15334 -19916
rect -15341 -20006 -15063 -19917
rect -14974 -20006 -14968 -19917
rect -14814 -19918 -14808 -19866
rect -14756 -19918 -14750 -19866
rect -12499 -19966 -12173 -19954
rect -12499 -19996 -12293 -19966
rect -15341 -20048 -15334 -20006
rect -15443 -20067 -15334 -20048
rect -15484 -20079 -15334 -20067
rect -20932 -20177 -20925 -20135
rect -21034 -20196 -20925 -20177
rect -21075 -20208 -20925 -20196
rect -17535 -20145 -17523 -20111
rect -17433 -20116 -16983 -20111
rect -16430 -20113 -15470 -20110
rect -17433 -20145 -16982 -20116
rect -17535 -20188 -16982 -20145
rect -17677 -20207 -17563 -20201
rect -22941 -20255 -21061 -20239
rect -22941 -20289 -21558 -20255
rect -21332 -20289 -21112 -20255
rect -21078 -20289 -21061 -20255
rect -22941 -20308 -21061 -20289
rect -17677 -20241 -17665 -20207
rect -17575 -20241 -17563 -20207
rect -20405 -20356 -20399 -20354
rect -24940 -20533 -24902 -20444
rect -24811 -20533 -23883 -20444
rect -21574 -20404 -20399 -20356
rect -21574 -20440 -21061 -20404
rect -20405 -20406 -20399 -20404
rect -20347 -20406 -20341 -20354
rect -17677 -20399 -17563 -20241
rect -17677 -20433 -17665 -20399
rect -17575 -20433 -17563 -20399
rect -21722 -20514 -21602 -20454
rect -24940 -20534 -24792 -20533
rect -21722 -20557 -21678 -20514
rect -21936 -20609 -21930 -20557
rect -21878 -20605 -21678 -20557
rect -21644 -20577 -21602 -20514
rect -21574 -20462 -21122 -20440
rect -21574 -20539 -21510 -20462
rect -21476 -20539 -21318 -20462
rect -21284 -20468 -21122 -20462
rect -21284 -20480 -21116 -20468
rect -21284 -20539 -21156 -20480
rect -21574 -20545 -21156 -20539
rect -21644 -20583 -21364 -20577
rect -21644 -20605 -21606 -20583
rect -21878 -20609 -21606 -20605
rect -24128 -20656 -23005 -20655
rect -24128 -20699 -22824 -20656
rect -21722 -20662 -21606 -20609
rect -21572 -20662 -21414 -20583
rect -21380 -20662 -21364 -20583
rect -21722 -20668 -21364 -20662
rect -21318 -20656 -21156 -20545
rect -21122 -20656 -21116 -20480
rect -21318 -20668 -21116 -20656
rect -21075 -20480 -20925 -20468
rect -21075 -20656 -21068 -20480
rect -21034 -20498 -20925 -20480
rect -21034 -20505 -20649 -20498
rect -21034 -20637 -20966 -20505
rect -20932 -20587 -20649 -20505
rect -20560 -20587 -20554 -20498
rect -20932 -20637 -20925 -20587
rect -21034 -20656 -20925 -20637
rect -21075 -20668 -20925 -20656
rect -17677 -20591 -17563 -20433
rect -17535 -20303 -17421 -20188
rect -17535 -20337 -17523 -20303
rect -17433 -20337 -17421 -20303
rect -17535 -20495 -17421 -20337
rect -17535 -20529 -17523 -20495
rect -17433 -20529 -17421 -20495
rect -17182 -20379 -16982 -20188
rect -16551 -20126 -15470 -20113
rect -16551 -20160 -15967 -20126
rect -15741 -20160 -15521 -20126
rect -15487 -20160 -15470 -20126
rect -16551 -20179 -15470 -20160
rect -16551 -20182 -16378 -20179
rect -16551 -20379 -16482 -20182
rect -15983 -20275 -12700 -20227
rect -15983 -20311 -15470 -20275
rect -17182 -20448 -16482 -20379
rect -16131 -20385 -16011 -20325
rect -16131 -20428 -16087 -20385
rect -17535 -20535 -17421 -20529
rect -17677 -20625 -17665 -20591
rect -17575 -20625 -17563 -20591
rect -24128 -20715 -21061 -20699
rect -24128 -20725 -21558 -20715
rect -24128 -20733 -23005 -20725
rect -24128 -20791 -24046 -20733
rect -22893 -20749 -21558 -20725
rect -21332 -20749 -21112 -20715
rect -21078 -20749 -21061 -20715
rect -22893 -20768 -21061 -20749
rect -17828 -20722 -17762 -20710
rect -24395 -20828 -24303 -20827
rect -24515 -20839 -24302 -20828
rect -24515 -20864 -24389 -20839
rect -24823 -21104 -24711 -21096
rect -24515 -21104 -24508 -20864
rect -24823 -21200 -24815 -21104
rect -24719 -21200 -24508 -21104
rect -24823 -21208 -24711 -21200
rect -24515 -21433 -24508 -21200
rect -24461 -20873 -24389 -20864
rect -24309 -20873 -24302 -20839
rect -24461 -21031 -24302 -20873
rect -24461 -21065 -24389 -21031
rect -24309 -21065 -24302 -21031
rect -24461 -21223 -24302 -21065
rect -24461 -21257 -24389 -21223
rect -24309 -21257 -24302 -21223
rect -24461 -21415 -24302 -21257
rect -24273 -20839 -23999 -20791
rect -18578 -20816 -18572 -20814
rect -24273 -20935 -24039 -20839
rect -24273 -20969 -24267 -20935
rect -24187 -20969 -24039 -20935
rect -24273 -21127 -24181 -20969
rect -24273 -21161 -24267 -21127
rect -24187 -21161 -24181 -21127
rect -24273 -21319 -24181 -21161
rect -24153 -21060 -24079 -21045
rect -24153 -21094 -24134 -21060
rect -24099 -21094 -24079 -21060
rect -24153 -21255 -24079 -21094
rect -24051 -21215 -24039 -20969
rect -24005 -21215 -23999 -20839
rect -24051 -21227 -23999 -21215
rect -23853 -20839 -23730 -20827
rect -23853 -21215 -23847 -20839
rect -23813 -20865 -23730 -20839
rect -23813 -21200 -23775 -20865
rect -23741 -20994 -23730 -20865
rect -21588 -20864 -18572 -20816
rect -21588 -20900 -21075 -20864
rect -18578 -20866 -18572 -20864
rect -18520 -20866 -18514 -20814
rect -18102 -20869 -18004 -20857
rect -17828 -20869 -17820 -20722
rect -21736 -20974 -21616 -20914
rect -23741 -21095 -23329 -20994
rect -23228 -21095 -23222 -20994
rect -21736 -21022 -21692 -20974
rect -21934 -21074 -21928 -21022
rect -21876 -21065 -21692 -21022
rect -21658 -21037 -21616 -20974
rect -21588 -20922 -21136 -20900
rect -21588 -20999 -21524 -20922
rect -21490 -20999 -21332 -20922
rect -21298 -20928 -21136 -20922
rect -21298 -20940 -21130 -20928
rect -21298 -20999 -21170 -20940
rect -21588 -21005 -21170 -20999
rect -21658 -21043 -21378 -21037
rect -21658 -21065 -21620 -21043
rect -21876 -21074 -21620 -21065
rect -23741 -21200 -23730 -21095
rect -21736 -21122 -21620 -21074
rect -21586 -21122 -21428 -21043
rect -21394 -21122 -21378 -21043
rect -21736 -21128 -21378 -21122
rect -21332 -21116 -21170 -21005
rect -21136 -21116 -21130 -20940
rect -21332 -21128 -21130 -21116
rect -21089 -20940 -20939 -20928
rect -21089 -21116 -21082 -20940
rect -21048 -20965 -20649 -20940
rect -21048 -21097 -20980 -20965
rect -20946 -21029 -20649 -20965
rect -20560 -21029 -20554 -20940
rect -18102 -20943 -18090 -20869
rect -18016 -20943 -17820 -20869
rect -18102 -20955 -18004 -20943
rect -20946 -21097 -20939 -21029
rect -17828 -21079 -17820 -20943
rect -17769 -21079 -17762 -20722
rect -17677 -20783 -17563 -20625
rect -17282 -20543 -17216 -20527
rect -17282 -20577 -17266 -20543
rect -17232 -20577 -17216 -20543
rect -17677 -20817 -17665 -20783
rect -17575 -20817 -17563 -20783
rect -17677 -20975 -17563 -20817
rect -17677 -21009 -17665 -20975
rect -17575 -21009 -17563 -20975
rect -17677 -21015 -17563 -21009
rect -17535 -20687 -17421 -20681
rect -17535 -20721 -17523 -20687
rect -17433 -20721 -17421 -20687
rect -17535 -20879 -17421 -20721
rect -17535 -20913 -17523 -20879
rect -17433 -20913 -17421 -20879
rect -17828 -21091 -17762 -21079
rect -17535 -21071 -17421 -20913
rect -21048 -21116 -20939 -21097
rect -17535 -21105 -17523 -21071
rect -17433 -21105 -17421 -21071
rect -17535 -21111 -17421 -21105
rect -17387 -20686 -17321 -20627
rect -17387 -20720 -17371 -20686
rect -17337 -20720 -17321 -20686
rect -21089 -21128 -20939 -21116
rect -23813 -21215 -23730 -21200
rect -23853 -21227 -23730 -21215
rect -22729 -21175 -21075 -21159
rect -22729 -21209 -21572 -21175
rect -21346 -21209 -21126 -21175
rect -21092 -21209 -21075 -21175
rect -22729 -21228 -21075 -21209
rect -18053 -21176 -17992 -21170
rect -24153 -21265 -23852 -21255
rect -24153 -21299 -24010 -21265
rect -23975 -21299 -23852 -21265
rect -24153 -21305 -23852 -21299
rect -24273 -21353 -24267 -21319
rect -24187 -21353 -24181 -21319
rect -24273 -21369 -24181 -21353
rect -24152 -21349 -24017 -21333
rect -24461 -21433 -24389 -21415
rect -24515 -21449 -24389 -21433
rect -24309 -21449 -24302 -21415
rect -24515 -21462 -24302 -21449
rect -24152 -21383 -24134 -21349
rect -24099 -21383 -24017 -21349
rect -24152 -21497 -24017 -21383
rect -24936 -21569 -24924 -21497
rect -24852 -21569 -24017 -21497
rect -23988 -21650 -23852 -21305
rect -24936 -21739 -24913 -21650
rect -24823 -21739 -23852 -21650
rect -24126 -21963 -23005 -21957
rect -22729 -21963 -22660 -21228
rect -17992 -21178 -17900 -21176
rect -17387 -21178 -17321 -20720
rect -17992 -21237 -17321 -21178
rect -18053 -21243 -17992 -21237
rect -17964 -21244 -17321 -21237
rect -17282 -21274 -17216 -20577
rect -17182 -20585 -16982 -20448
rect -16345 -20480 -16339 -20428
rect -16287 -20476 -16087 -20428
rect -16053 -20448 -16011 -20385
rect -15983 -20333 -15531 -20311
rect -15983 -20410 -15919 -20333
rect -15885 -20410 -15727 -20333
rect -15693 -20339 -15531 -20333
rect -15693 -20351 -15525 -20339
rect -15693 -20410 -15565 -20351
rect -15983 -20416 -15565 -20410
rect -16053 -20454 -15773 -20448
rect -16053 -20476 -16015 -20454
rect -16287 -20480 -16015 -20476
rect -16924 -20508 -16850 -20496
rect -17188 -20591 -16988 -20585
rect -17188 -20625 -17176 -20591
rect -17000 -20625 -16988 -20591
rect -17188 -20631 -16988 -20625
rect -16924 -20707 -16917 -20508
rect -16856 -20707 -16850 -20508
rect -16131 -20533 -16015 -20480
rect -15981 -20533 -15823 -20454
rect -15789 -20533 -15773 -20454
rect -16131 -20539 -15773 -20533
rect -15727 -20527 -15565 -20416
rect -15531 -20527 -15525 -20351
rect -15727 -20539 -15525 -20527
rect -15484 -20351 -15334 -20339
rect -15484 -20527 -15477 -20351
rect -15443 -20369 -15334 -20351
rect -15443 -20376 -15058 -20369
rect -15443 -20508 -15375 -20376
rect -15341 -20458 -15058 -20376
rect -14969 -20458 -14963 -20369
rect -15341 -20508 -15334 -20458
rect -15443 -20527 -15334 -20508
rect -15484 -20539 -15334 -20527
rect -16430 -20573 -15470 -20570
rect -16924 -20719 -16850 -20707
rect -16531 -20586 -15470 -20573
rect -16531 -20620 -15967 -20586
rect -15741 -20620 -15521 -20586
rect -15487 -20620 -15470 -20586
rect -16531 -20639 -15470 -20620
rect -16531 -20642 -16390 -20639
rect -16916 -20995 -16854 -20719
rect -16531 -20763 -16462 -20642
rect -16647 -20832 -16462 -20763
rect -15997 -20735 -12822 -20687
rect -15997 -20771 -15484 -20735
rect -16930 -21013 -16836 -20995
rect -16930 -21075 -16916 -21013
rect -16854 -21075 -16836 -21013
rect -16930 -21091 -16836 -21075
rect -18692 -21294 -18640 -21288
rect -21586 -21344 -18692 -21296
rect -21586 -21380 -21073 -21344
rect -17968 -21322 -17216 -21274
rect -18692 -21352 -18640 -21346
rect -17974 -21340 -17216 -21322
rect -21734 -21454 -21614 -21394
rect -21734 -21503 -21690 -21454
rect -21930 -21555 -21924 -21503
rect -21872 -21545 -21690 -21503
rect -21656 -21517 -21614 -21454
rect -21586 -21402 -21134 -21380
rect -21586 -21479 -21522 -21402
rect -21488 -21479 -21330 -21402
rect -21296 -21408 -21134 -21402
rect -17974 -21404 -17968 -21340
rect -17904 -21404 -17886 -21340
rect -21296 -21420 -21128 -21408
rect -21296 -21479 -21168 -21420
rect -21586 -21485 -21168 -21479
rect -21656 -21523 -21376 -21517
rect -21656 -21545 -21618 -21523
rect -21872 -21555 -21618 -21545
rect -21734 -21602 -21618 -21555
rect -21584 -21602 -21426 -21523
rect -21392 -21602 -21376 -21523
rect -21734 -21608 -21376 -21602
rect -21330 -21596 -21168 -21485
rect -21134 -21596 -21128 -21420
rect -21330 -21608 -21128 -21596
rect -21087 -21420 -20937 -21408
rect -17974 -21410 -17886 -21404
rect -21087 -21596 -21080 -21420
rect -21046 -21421 -20937 -21420
rect -21046 -21445 -20655 -21421
rect -21046 -21577 -20978 -21445
rect -20944 -21510 -20655 -21445
rect -20566 -21510 -20560 -21421
rect -17535 -21465 -16984 -21463
rect -20944 -21577 -20937 -21510
rect -21046 -21596 -20937 -21577
rect -21087 -21608 -20937 -21596
rect -17535 -21511 -16983 -21465
rect -17535 -21545 -17523 -21511
rect -17433 -21516 -16983 -21511
rect -17433 -21545 -16982 -21516
rect -17535 -21558 -16982 -21545
rect -16647 -21558 -16578 -20832
rect -16145 -20845 -16025 -20785
rect -16145 -20893 -16101 -20845
rect -16343 -20945 -16337 -20893
rect -16285 -20936 -16101 -20893
rect -16067 -20908 -16025 -20845
rect -15997 -20793 -15545 -20771
rect -15997 -20870 -15933 -20793
rect -15899 -20870 -15741 -20793
rect -15707 -20799 -15545 -20793
rect -15707 -20811 -15539 -20799
rect -15707 -20870 -15579 -20811
rect -15997 -20876 -15579 -20870
rect -16067 -20914 -15787 -20908
rect -16067 -20936 -16029 -20914
rect -16285 -20945 -16029 -20936
rect -16145 -20993 -16029 -20945
rect -15995 -20993 -15837 -20914
rect -15803 -20993 -15787 -20914
rect -16145 -20999 -15787 -20993
rect -15741 -20987 -15579 -20876
rect -15545 -20987 -15539 -20811
rect -15741 -20999 -15539 -20987
rect -15498 -20811 -15348 -20799
rect -15498 -20987 -15491 -20811
rect -15457 -20836 -15058 -20811
rect -15457 -20968 -15389 -20836
rect -15355 -20900 -15058 -20836
rect -14969 -20900 -14963 -20811
rect -15355 -20968 -15348 -20900
rect -15457 -20987 -15348 -20968
rect -15498 -20999 -15348 -20987
rect -16430 -21031 -15484 -21030
rect -17535 -21588 -16578 -21558
rect -17677 -21607 -17563 -21601
rect -24126 -22032 -22660 -21963
rect -22539 -21655 -21073 -21639
rect -22539 -21689 -21570 -21655
rect -21344 -21689 -21124 -21655
rect -21090 -21689 -21073 -21655
rect -22539 -21708 -21073 -21689
rect -17677 -21641 -17665 -21607
rect -17575 -21641 -17563 -21607
rect -24126 -22035 -23005 -22032
rect -24126 -22094 -24044 -22035
rect -24396 -22131 -24304 -22130
rect -24516 -22142 -24303 -22131
rect -24516 -22167 -24390 -22142
rect -24813 -22412 -24701 -22404
rect -24516 -22412 -24509 -22167
rect -24813 -22508 -24805 -22412
rect -24709 -22508 -24509 -22412
rect -24813 -22509 -24509 -22508
rect -24813 -22516 -24701 -22509
rect -24516 -22736 -24509 -22509
rect -24462 -22176 -24390 -22167
rect -24310 -22176 -24303 -22142
rect -24462 -22334 -24303 -22176
rect -24462 -22368 -24390 -22334
rect -24310 -22368 -24303 -22334
rect -24462 -22526 -24303 -22368
rect -24462 -22560 -24390 -22526
rect -24310 -22560 -24303 -22526
rect -24462 -22718 -24303 -22560
rect -24274 -22142 -24000 -22094
rect -24274 -22238 -24040 -22142
rect -24274 -22272 -24268 -22238
rect -24188 -22272 -24040 -22238
rect -24274 -22430 -24182 -22272
rect -24274 -22464 -24268 -22430
rect -24188 -22464 -24182 -22430
rect -24274 -22622 -24182 -22464
rect -24154 -22363 -24080 -22348
rect -24154 -22397 -24135 -22363
rect -24100 -22397 -24080 -22363
rect -24154 -22558 -24080 -22397
rect -24052 -22518 -24040 -22272
rect -24006 -22518 -24000 -22142
rect -24052 -22530 -24000 -22518
rect -23854 -22142 -23731 -22130
rect -23854 -22518 -23848 -22142
rect -23814 -22168 -23731 -22142
rect -23814 -22503 -23776 -22168
rect -23742 -22288 -23731 -22168
rect -23742 -22389 -23332 -22288
rect -23231 -22389 -23225 -22288
rect -23742 -22503 -23731 -22389
rect -23814 -22518 -23731 -22503
rect -23854 -22530 -23731 -22518
rect -24154 -22568 -23853 -22558
rect -24154 -22602 -24011 -22568
rect -23976 -22602 -23853 -22568
rect -24154 -22608 -23853 -22602
rect -24274 -22656 -24268 -22622
rect -24188 -22656 -24182 -22622
rect -24274 -22672 -24182 -22656
rect -24153 -22652 -24018 -22636
rect -24462 -22736 -24390 -22718
rect -24516 -22752 -24390 -22736
rect -24310 -22752 -24303 -22718
rect -24516 -22765 -24303 -22752
rect -24153 -22686 -24135 -22652
rect -24100 -22686 -24018 -22652
rect -24153 -22798 -24018 -22686
rect -24936 -22870 -24890 -22798
rect -24818 -22870 -24018 -22798
rect -23989 -22951 -23853 -22608
rect -24936 -23040 -24913 -22951
rect -24819 -23040 -23853 -22951
rect -24134 -23269 -23005 -23262
rect -22539 -23269 -22470 -21708
rect -17677 -21799 -17563 -21641
rect -17677 -21833 -17665 -21799
rect -17575 -21833 -17563 -21799
rect -17677 -21991 -17563 -21833
rect -17535 -21703 -17421 -21588
rect -17535 -21737 -17523 -21703
rect -17433 -21737 -17421 -21703
rect -17535 -21895 -17421 -21737
rect -17535 -21929 -17523 -21895
rect -17433 -21929 -17421 -21895
rect -17182 -21627 -16578 -21588
rect -16524 -21046 -15484 -21031
rect -16524 -21080 -15981 -21046
rect -15755 -21080 -15535 -21046
rect -15501 -21080 -15484 -21046
rect -16524 -21099 -15484 -21080
rect -17535 -21935 -17421 -21929
rect -17677 -22025 -17665 -21991
rect -17575 -22025 -17563 -21991
rect -17828 -22122 -17762 -22110
rect -18100 -22273 -18002 -22261
rect -17828 -22273 -17820 -22122
rect -18100 -22347 -18088 -22273
rect -18014 -22347 -17820 -22273
rect -18100 -22359 -18002 -22347
rect -17828 -22479 -17820 -22347
rect -17769 -22479 -17762 -22122
rect -17677 -22183 -17563 -22025
rect -17282 -21943 -17216 -21927
rect -17282 -21977 -17266 -21943
rect -17232 -21977 -17216 -21943
rect -17677 -22217 -17665 -22183
rect -17575 -22217 -17563 -22183
rect -17677 -22375 -17563 -22217
rect -17677 -22409 -17665 -22375
rect -17575 -22409 -17563 -22375
rect -17677 -22415 -17563 -22409
rect -17535 -22087 -17421 -22081
rect -17535 -22121 -17523 -22087
rect -17433 -22121 -17421 -22087
rect -17535 -22279 -17421 -22121
rect -17535 -22313 -17523 -22279
rect -17433 -22313 -17421 -22279
rect -17828 -22491 -17762 -22479
rect -17535 -22471 -17421 -22313
rect -17535 -22505 -17523 -22471
rect -17433 -22505 -17421 -22471
rect -17535 -22511 -17421 -22505
rect -17387 -22086 -17321 -22027
rect -17387 -22120 -17371 -22086
rect -17337 -22120 -17321 -22086
rect -17387 -22600 -17321 -22120
rect -18067 -22666 -18061 -22600
rect -17995 -22666 -17321 -22600
rect -17282 -22706 -17216 -21977
rect -17182 -21985 -16982 -21627
rect -16924 -21908 -16850 -21896
rect -17188 -21991 -16988 -21985
rect -17188 -22025 -17176 -21991
rect -17000 -22025 -16988 -21991
rect -17188 -22031 -16988 -22025
rect -16924 -22107 -16917 -21908
rect -16856 -21983 -16850 -21908
rect -16738 -21983 -16646 -21969
rect -16856 -22047 -16726 -21983
rect -16662 -22047 -16646 -21983
rect -16856 -22107 -16850 -22047
rect -16738 -22061 -16646 -22047
rect -16924 -22119 -16850 -22107
rect -17964 -22724 -17216 -22706
rect -18080 -22745 -17216 -22724
rect -18080 -22834 -18071 -22745
rect -17982 -22772 -17216 -22745
rect -17982 -22834 -17876 -22772
rect -18080 -22846 -17952 -22834
rect -17535 -22865 -16984 -22863
rect -17535 -22911 -16983 -22865
rect -17535 -22945 -17523 -22911
rect -17433 -22916 -16983 -22911
rect -17433 -22945 -16982 -22916
rect -17535 -22953 -16982 -22945
rect -16524 -22953 -16442 -21099
rect -15995 -21215 -12966 -21167
rect -15995 -21251 -15482 -21215
rect -16143 -21325 -16023 -21265
rect -16143 -21374 -16099 -21325
rect -16339 -21426 -16333 -21374
rect -16281 -21416 -16099 -21374
rect -16065 -21388 -16023 -21325
rect -15995 -21273 -15543 -21251
rect -15995 -21350 -15931 -21273
rect -15897 -21350 -15739 -21273
rect -15705 -21279 -15543 -21273
rect -15705 -21291 -15537 -21279
rect -15705 -21350 -15577 -21291
rect -15995 -21356 -15577 -21350
rect -16065 -21394 -15785 -21388
rect -16065 -21416 -16027 -21394
rect -16281 -21426 -16027 -21416
rect -16143 -21473 -16027 -21426
rect -15993 -21473 -15835 -21394
rect -15801 -21473 -15785 -21394
rect -16143 -21479 -15785 -21473
rect -15739 -21467 -15577 -21356
rect -15543 -21467 -15537 -21291
rect -15739 -21479 -15537 -21467
rect -15496 -21291 -15346 -21279
rect -15496 -21467 -15489 -21291
rect -15455 -21292 -15346 -21291
rect -15455 -21316 -15064 -21292
rect -15455 -21448 -15387 -21316
rect -15353 -21381 -15064 -21316
rect -14975 -21381 -14969 -21292
rect -15353 -21448 -15346 -21381
rect -15455 -21467 -15346 -21448
rect -15496 -21479 -15346 -21467
rect -16402 -21526 -15482 -21510
rect -16402 -21560 -15979 -21526
rect -15753 -21560 -15533 -21526
rect -15499 -21560 -15482 -21526
rect -16402 -21579 -15482 -21560
rect -17535 -22988 -16442 -22953
rect -24134 -23338 -22470 -23269
rect -17677 -23007 -17563 -23001
rect -17677 -23041 -17665 -23007
rect -17575 -23041 -17563 -23007
rect -17677 -23199 -17563 -23041
rect -17677 -23233 -17665 -23199
rect -17575 -23233 -17563 -23199
rect -24134 -23340 -23005 -23338
rect -24134 -23403 -24052 -23340
rect -17677 -23391 -17563 -23233
rect -17535 -23103 -17421 -22988
rect -17535 -23137 -17523 -23103
rect -17433 -23137 -17421 -23103
rect -17535 -23295 -17421 -23137
rect -17535 -23329 -17523 -23295
rect -17433 -23329 -17421 -23295
rect -17182 -23043 -16442 -22988
rect -17535 -23335 -17421 -23329
rect -24396 -23440 -24304 -23439
rect -24516 -23451 -24303 -23440
rect -24516 -23476 -24390 -23451
rect -24833 -23718 -24721 -23710
rect -24516 -23718 -24509 -23476
rect -24833 -23814 -24825 -23718
rect -24729 -23814 -24509 -23718
rect -24833 -23822 -24721 -23814
rect -24516 -24045 -24509 -23814
rect -24462 -23485 -24390 -23476
rect -24310 -23485 -24303 -23451
rect -24462 -23643 -24303 -23485
rect -24462 -23677 -24390 -23643
rect -24310 -23677 -24303 -23643
rect -24462 -23835 -24303 -23677
rect -24462 -23869 -24390 -23835
rect -24310 -23869 -24303 -23835
rect -24462 -24027 -24303 -23869
rect -24274 -23451 -24000 -23403
rect -17677 -23425 -17665 -23391
rect -17575 -23425 -17563 -23391
rect -24274 -23547 -24040 -23451
rect -24274 -23581 -24268 -23547
rect -24188 -23581 -24040 -23547
rect -24274 -23739 -24182 -23581
rect -24274 -23773 -24268 -23739
rect -24188 -23773 -24182 -23739
rect -24274 -23931 -24182 -23773
rect -24154 -23672 -24080 -23657
rect -24154 -23706 -24135 -23672
rect -24100 -23706 -24080 -23672
rect -24154 -23867 -24080 -23706
rect -24052 -23827 -24040 -23581
rect -24006 -23827 -24000 -23451
rect -24052 -23839 -24000 -23827
rect -23854 -23451 -23731 -23439
rect -23854 -23827 -23848 -23451
rect -23814 -23477 -23731 -23451
rect -23814 -23812 -23776 -23477
rect -23742 -23604 -23731 -23477
rect -17828 -23522 -17762 -23510
rect -23742 -23705 -23372 -23604
rect -23271 -23705 -23265 -23604
rect -18102 -23675 -18004 -23663
rect -17828 -23675 -17820 -23522
rect -23742 -23812 -23731 -23705
rect -18102 -23749 -18090 -23675
rect -18016 -23749 -17820 -23675
rect -18102 -23761 -18004 -23749
rect -23814 -23827 -23731 -23812
rect -23854 -23839 -23731 -23827
rect -24154 -23877 -23853 -23867
rect -24154 -23911 -24011 -23877
rect -23976 -23911 -23853 -23877
rect -17828 -23879 -17820 -23749
rect -17769 -23879 -17762 -23522
rect -17677 -23583 -17563 -23425
rect -17282 -23343 -17216 -23327
rect -17282 -23377 -17266 -23343
rect -17232 -23377 -17216 -23343
rect -17677 -23617 -17665 -23583
rect -17575 -23617 -17563 -23583
rect -17677 -23775 -17563 -23617
rect -17677 -23809 -17665 -23775
rect -17575 -23809 -17563 -23775
rect -17677 -23815 -17563 -23809
rect -17535 -23487 -17421 -23481
rect -17535 -23521 -17523 -23487
rect -17433 -23521 -17421 -23487
rect -17535 -23679 -17421 -23521
rect -17535 -23713 -17523 -23679
rect -17433 -23713 -17421 -23679
rect -17828 -23891 -17762 -23879
rect -17535 -23871 -17421 -23713
rect -17535 -23905 -17523 -23871
rect -17433 -23905 -17421 -23871
rect -17535 -23911 -17421 -23905
rect -17387 -23486 -17321 -23427
rect -17387 -23520 -17371 -23486
rect -17337 -23520 -17321 -23486
rect -24154 -23917 -23853 -23911
rect -24274 -23965 -24268 -23931
rect -24188 -23965 -24182 -23931
rect -24274 -23981 -24182 -23965
rect -24153 -23961 -24018 -23945
rect -24462 -24045 -24390 -24027
rect -24516 -24061 -24390 -24045
rect -24310 -24061 -24303 -24027
rect -24516 -24074 -24303 -24061
rect -24153 -23995 -24135 -23961
rect -24100 -23995 -24018 -23961
rect -24153 -24108 -24018 -23995
rect -24936 -24180 -24926 -24108
rect -24854 -24180 -24018 -24108
rect -24934 -24261 -24778 -24252
rect -23989 -24261 -23853 -23917
rect -17387 -23953 -17321 -23520
rect -18050 -23986 -17962 -23978
rect -18050 -24058 -18042 -23986
rect -17970 -24000 -17900 -23986
rect -17381 -24000 -17328 -23953
rect -17970 -24053 -17328 -24000
rect -17970 -24058 -17900 -24053
rect -18050 -24066 -17962 -24058
rect -17282 -24096 -17216 -23377
rect -17182 -23385 -16982 -23043
rect -16924 -23308 -16850 -23296
rect -17188 -23391 -16988 -23385
rect -17188 -23425 -17176 -23391
rect -17000 -23425 -16988 -23391
rect -17188 -23431 -16988 -23425
rect -16924 -23507 -16917 -23308
rect -16856 -23367 -16850 -23308
rect -16706 -23367 -16596 -23349
rect -16856 -23445 -16688 -23367
rect -16610 -23445 -16596 -23367
rect -16856 -23507 -16850 -23445
rect -16706 -23459 -16596 -23445
rect -16924 -23519 -16850 -23507
rect -17964 -24102 -17216 -24096
rect -18084 -24131 -17216 -24102
rect -18084 -24220 -18063 -24131
rect -17974 -24162 -17216 -24131
rect -17974 -24220 -17880 -24162
rect -18084 -24246 -17958 -24220
rect -24936 -24350 -24907 -24261
rect -24813 -24350 -23853 -24261
rect -17535 -24265 -16984 -24263
rect -17535 -24283 -16983 -24265
rect -16393 -24283 -16324 -21579
rect -17535 -24311 -16324 -24283
rect -17535 -24345 -17523 -24311
rect -17433 -24345 -16324 -24311
rect -24934 -24360 -24778 -24350
rect -17535 -24367 -16324 -24345
rect -17535 -24388 -16982 -24367
rect -17677 -24407 -17563 -24401
rect -17677 -24441 -17665 -24407
rect -17575 -24441 -17563 -24407
rect -17677 -24599 -17563 -24441
rect -17677 -24633 -17665 -24599
rect -17575 -24633 -17563 -24599
rect -17677 -24791 -17563 -24633
rect -17535 -24503 -17421 -24388
rect -17535 -24537 -17523 -24503
rect -17433 -24537 -17421 -24503
rect -17535 -24695 -17421 -24537
rect -17535 -24729 -17523 -24695
rect -17433 -24729 -17421 -24695
rect -17535 -24735 -17421 -24729
rect -17677 -24825 -17665 -24791
rect -17575 -24825 -17563 -24791
rect -17828 -24922 -17762 -24910
rect -18096 -25055 -17998 -25043
rect -17828 -25055 -17820 -24922
rect -18096 -25129 -18084 -25055
rect -18010 -25129 -17820 -25055
rect -18096 -25141 -17998 -25129
rect -17828 -25279 -17820 -25129
rect -17769 -25279 -17762 -24922
rect -17677 -24983 -17563 -24825
rect -17282 -24743 -17216 -24727
rect -17282 -24777 -17266 -24743
rect -17232 -24777 -17216 -24743
rect -17677 -25017 -17665 -24983
rect -17575 -25017 -17563 -24983
rect -17677 -25175 -17563 -25017
rect -17677 -25209 -17665 -25175
rect -17575 -25209 -17563 -25175
rect -17677 -25215 -17563 -25209
rect -17535 -24887 -17421 -24881
rect -17535 -24921 -17523 -24887
rect -17433 -24921 -17421 -24887
rect -17535 -25079 -17421 -24921
rect -17535 -25113 -17523 -25079
rect -17433 -25113 -17421 -25079
rect -17828 -25291 -17762 -25279
rect -17535 -25271 -17421 -25113
rect -17535 -25305 -17523 -25271
rect -17433 -25305 -17421 -25271
rect -17535 -25311 -17421 -25305
rect -17387 -24886 -17321 -24827
rect -17387 -24920 -17371 -24886
rect -17337 -24920 -17321 -24886
rect -17964 -25350 -17878 -25344
rect -17964 -25422 -17956 -25350
rect -17884 -25360 -17878 -25350
rect -17387 -25360 -17321 -24920
rect -17884 -25422 -17321 -25360
rect -17964 -25426 -17321 -25422
rect -17964 -25428 -17878 -25426
rect -17282 -25480 -17216 -24777
rect -17182 -24785 -16982 -24388
rect -16924 -24708 -16850 -24696
rect -17188 -24791 -16988 -24785
rect -17188 -24825 -17176 -24791
rect -17000 -24825 -16988 -24791
rect -17188 -24831 -16988 -24825
rect -16924 -24907 -16917 -24708
rect -16856 -24775 -16850 -24708
rect -16704 -24775 -16598 -24759
rect -16856 -24849 -16688 -24775
rect -16614 -24849 -16598 -24775
rect -16856 -24907 -16850 -24849
rect -16704 -24865 -16598 -24849
rect -16924 -24919 -16850 -24907
rect -13014 -25106 -12966 -21215
rect -12870 -22284 -12822 -20735
rect -12748 -22092 -12700 -20275
rect -12499 -21118 -12471 -19996
rect -12399 -20000 -12293 -19996
rect -12191 -20000 -12173 -19966
rect -12399 -20158 -12173 -20000
rect -11923 -19966 -11776 -19954
rect -11923 -20000 -11902 -19966
rect -11835 -20000 -11776 -19966
rect -12399 -20192 -12293 -20158
rect -12191 -20192 -12173 -20158
rect -12399 -20208 -12173 -20192
rect -12135 -20062 -11956 -20046
rect -12135 -20096 -12109 -20062
rect -11985 -20096 -11956 -20062
rect -12399 -20910 -12365 -20208
rect -12135 -20254 -11956 -20096
rect -11923 -20158 -11776 -20000
rect -11541 -19967 -11332 -19830
rect -11541 -20001 -11411 -19967
rect -11448 -20032 -11411 -20001
rect -11356 -20032 -11332 -19967
rect -11278 -19966 -10999 -19957
rect -11278 -20000 -11262 -19966
rect -11156 -19995 -10999 -19966
rect -11156 -20000 -11068 -19995
rect -11278 -20012 -11068 -20000
rect -11448 -20043 -11332 -20032
rect -11289 -20062 -11221 -20046
rect -11289 -20096 -11277 -20062
rect -11243 -20096 -11221 -20062
rect -11923 -20192 -11902 -20158
rect -11835 -20192 -11776 -20158
rect -11923 -20208 -11776 -20192
rect -11601 -20134 -11331 -20117
rect -11601 -20214 -11582 -20134
rect -11514 -20214 -11331 -20134
rect -11601 -20232 -11331 -20214
rect -12135 -20288 -12110 -20254
rect -11986 -20288 -11956 -20254
rect -12320 -20350 -12173 -20334
rect -12320 -20384 -12293 -20350
rect -12191 -20384 -12173 -20350
rect -12320 -20542 -12173 -20384
rect -12320 -20576 -12293 -20542
rect -12191 -20576 -12173 -20542
rect -12320 -20734 -12173 -20576
rect -12320 -20768 -12294 -20734
rect -12192 -20768 -12173 -20734
rect -12320 -20784 -12173 -20768
rect -12135 -20446 -11956 -20288
rect -11601 -20334 -11502 -20302
rect -12135 -20480 -12110 -20446
rect -11986 -20480 -11956 -20446
rect -12135 -20638 -11956 -20480
rect -12135 -20672 -12110 -20638
rect -11986 -20672 -11956 -20638
rect -12135 -20830 -11956 -20672
rect -11912 -20350 -11820 -20334
rect -11912 -20384 -11895 -20350
rect -11835 -20384 -11820 -20350
rect -11912 -20542 -11820 -20384
rect -11912 -20576 -11878 -20542
rect -11835 -20576 -11820 -20542
rect -11912 -20734 -11820 -20576
rect -11912 -20768 -11895 -20734
rect -11835 -20768 -11820 -20734
rect -11912 -20784 -11820 -20768
rect -11601 -20448 -11583 -20334
rect -11530 -20448 -11502 -20334
rect -12135 -20864 -12110 -20830
rect -11986 -20864 -11956 -20830
rect -12399 -20926 -12173 -20910
rect -12399 -20960 -12296 -20926
rect -12194 -20960 -12173 -20926
rect -12399 -21118 -12173 -20960
rect -12135 -21022 -11956 -20864
rect -12135 -21056 -12110 -21022
rect -11986 -21056 -11956 -21022
rect -12135 -21072 -11956 -21056
rect -11923 -20926 -11776 -20910
rect -11923 -20960 -11901 -20926
rect -11835 -20960 -11776 -20926
rect -12499 -21152 -12296 -21118
rect -12194 -21152 -12173 -21118
rect -12499 -21164 -12173 -21152
rect -11923 -21118 -11776 -20960
rect -11601 -20921 -11502 -20448
rect -11601 -21054 -11575 -20921
rect -11522 -21054 -11502 -20921
rect -11601 -21091 -11502 -21054
rect -11417 -21105 -11331 -20232
rect -11289 -20254 -11221 -20096
rect -11090 -20143 -11068 -20012
rect -11192 -20158 -11068 -20143
rect -11192 -20192 -11176 -20158
rect -11142 -20192 -11068 -20158
rect -11192 -20208 -11068 -20192
rect -11289 -20288 -11277 -20254
rect -11243 -20288 -11221 -20254
rect -11289 -20446 -11221 -20288
rect -11289 -20480 -11277 -20446
rect -11243 -20480 -11221 -20446
rect -11289 -20496 -11221 -20480
rect -11188 -20350 -11124 -20334
rect -11188 -20384 -11176 -20350
rect -11142 -20384 -11124 -20350
rect -11188 -20542 -11124 -20384
rect -11188 -20576 -11176 -20542
rect -11142 -20576 -11124 -20542
rect -11289 -20638 -11221 -20622
rect -11289 -20672 -11276 -20638
rect -11242 -20672 -11221 -20638
rect -11289 -20830 -11221 -20672
rect -11188 -20734 -11124 -20576
rect -11188 -20768 -11176 -20734
rect -11142 -20768 -11124 -20734
rect -11188 -20781 -11124 -20768
rect -11090 -20598 -11068 -20208
rect -11022 -20598 -10999 -19995
rect -11090 -20658 -11079 -20598
rect -11019 -20658 -10999 -20598
rect -11289 -20864 -11277 -20830
rect -11243 -20864 -11221 -20830
rect -11289 -21022 -11221 -20864
rect -11090 -20909 -11068 -20658
rect -11193 -20926 -11068 -20909
rect -11193 -20960 -11176 -20926
rect -11142 -20960 -11068 -20926
rect -11193 -20974 -11068 -20960
rect -11289 -21056 -11277 -21022
rect -11243 -21056 -11221 -21022
rect -11289 -21072 -11221 -21056
rect -11090 -21104 -11068 -20974
rect -11923 -21152 -11901 -21118
rect -11799 -21152 -11776 -21118
rect -11923 -21164 -11776 -21152
rect -11462 -21310 -11319 -21105
rect -11278 -21118 -11068 -21104
rect -11022 -21118 -10999 -20658
rect -11278 -21152 -11262 -21118
rect -11156 -21152 -10999 -21118
rect -11278 -21159 -10999 -21152
rect -12618 -21367 -12524 -21354
rect -12618 -21437 -12609 -21367
rect -12539 -21379 -11485 -21367
rect -12539 -21437 -11559 -21379
rect -12618 -21441 -11559 -21437
rect -11497 -21441 -11485 -21379
rect -12618 -21447 -11485 -21441
rect -12618 -21448 -12524 -21447
rect -11434 -21489 -11347 -21310
rect -12612 -21518 -11347 -21489
rect -12640 -21527 -11347 -21518
rect -12640 -21616 -12628 -21527
rect -12539 -21576 -11347 -21527
rect -12539 -21616 -12482 -21576
rect -12640 -21624 -12518 -21616
rect -12750 -22098 -12698 -22092
rect -12750 -22156 -12698 -22150
rect -12878 -22336 -12872 -22284
rect -12820 -22336 -12814 -22284
rect -11459 -22334 -10606 -22245
rect -11459 -22409 -11370 -22334
rect -12499 -22545 -12173 -22533
rect -12499 -22575 -12293 -22545
rect -12499 -23697 -12471 -22575
rect -12399 -22579 -12293 -22575
rect -12191 -22579 -12173 -22545
rect -12399 -22737 -12173 -22579
rect -11923 -22545 -11776 -22533
rect -11923 -22579 -11902 -22545
rect -11835 -22579 -11776 -22545
rect -12399 -22771 -12293 -22737
rect -12191 -22771 -12173 -22737
rect -12399 -22787 -12173 -22771
rect -12135 -22641 -11956 -22625
rect -12135 -22675 -12109 -22641
rect -11985 -22675 -11956 -22641
rect -12399 -23489 -12365 -22787
rect -12135 -22833 -11956 -22675
rect -11923 -22737 -11776 -22579
rect -11541 -22546 -11332 -22409
rect -11541 -22580 -11411 -22546
rect -11448 -22611 -11411 -22580
rect -11356 -22611 -11332 -22546
rect -11278 -22545 -10999 -22536
rect -11278 -22579 -11262 -22545
rect -11156 -22574 -10999 -22545
rect -11156 -22579 -11068 -22574
rect -11278 -22591 -11068 -22579
rect -11448 -22622 -11332 -22611
rect -11289 -22641 -11221 -22625
rect -11289 -22675 -11277 -22641
rect -11243 -22675 -11221 -22641
rect -11923 -22771 -11902 -22737
rect -11835 -22771 -11776 -22737
rect -11923 -22787 -11776 -22771
rect -11601 -22713 -11331 -22696
rect -11601 -22793 -11582 -22713
rect -11514 -22793 -11331 -22713
rect -11601 -22811 -11331 -22793
rect -12135 -22867 -12110 -22833
rect -11986 -22867 -11956 -22833
rect -12320 -22929 -12173 -22913
rect -12320 -22963 -12293 -22929
rect -12191 -22963 -12173 -22929
rect -12320 -23121 -12173 -22963
rect -12320 -23155 -12293 -23121
rect -12191 -23155 -12173 -23121
rect -12320 -23313 -12173 -23155
rect -12320 -23347 -12294 -23313
rect -12192 -23347 -12173 -23313
rect -12320 -23363 -12173 -23347
rect -12135 -23025 -11956 -22867
rect -11601 -22913 -11502 -22881
rect -12135 -23059 -12110 -23025
rect -11986 -23059 -11956 -23025
rect -12135 -23217 -11956 -23059
rect -12135 -23251 -12110 -23217
rect -11986 -23251 -11956 -23217
rect -12135 -23409 -11956 -23251
rect -11912 -22929 -11820 -22913
rect -11912 -22963 -11895 -22929
rect -11835 -22963 -11820 -22929
rect -11912 -23121 -11820 -22963
rect -11912 -23155 -11878 -23121
rect -11835 -23155 -11820 -23121
rect -11912 -23313 -11820 -23155
rect -11912 -23347 -11895 -23313
rect -11835 -23347 -11820 -23313
rect -11912 -23363 -11820 -23347
rect -11601 -23027 -11583 -22913
rect -11530 -23027 -11502 -22913
rect -12135 -23443 -12110 -23409
rect -11986 -23443 -11956 -23409
rect -12399 -23505 -12173 -23489
rect -12399 -23539 -12296 -23505
rect -12194 -23539 -12173 -23505
rect -12399 -23697 -12173 -23539
rect -12135 -23601 -11956 -23443
rect -12135 -23635 -12110 -23601
rect -11986 -23635 -11956 -23601
rect -12135 -23651 -11956 -23635
rect -11923 -23505 -11776 -23489
rect -11923 -23539 -11901 -23505
rect -11835 -23539 -11776 -23505
rect -12499 -23731 -12296 -23697
rect -12194 -23731 -12173 -23697
rect -12499 -23743 -12173 -23731
rect -11923 -23697 -11776 -23539
rect -11601 -23500 -11502 -23027
rect -11601 -23633 -11575 -23500
rect -11522 -23633 -11502 -23500
rect -11601 -23670 -11502 -23633
rect -11417 -23684 -11331 -22811
rect -11289 -22833 -11221 -22675
rect -11090 -22722 -11068 -22591
rect -11192 -22737 -11068 -22722
rect -11192 -22771 -11176 -22737
rect -11142 -22771 -11068 -22737
rect -11192 -22787 -11068 -22771
rect -11289 -22867 -11277 -22833
rect -11243 -22867 -11221 -22833
rect -11289 -23025 -11221 -22867
rect -11289 -23059 -11277 -23025
rect -11243 -23059 -11221 -23025
rect -11289 -23075 -11221 -23059
rect -11188 -22929 -11124 -22913
rect -11188 -22963 -11176 -22929
rect -11142 -22963 -11124 -22929
rect -11188 -23121 -11124 -22963
rect -11188 -23155 -11176 -23121
rect -11142 -23155 -11124 -23121
rect -11289 -23217 -11221 -23201
rect -11289 -23251 -11276 -23217
rect -11242 -23251 -11221 -23217
rect -11289 -23409 -11221 -23251
rect -11188 -23313 -11124 -23155
rect -11188 -23347 -11176 -23313
rect -11142 -23347 -11124 -23313
rect -11188 -23360 -11124 -23347
rect -11090 -23177 -11068 -22787
rect -11022 -23177 -10999 -22574
rect -11090 -23237 -11079 -23177
rect -11019 -23237 -10999 -23177
rect -11289 -23443 -11277 -23409
rect -11243 -23443 -11221 -23409
rect -11289 -23601 -11221 -23443
rect -11090 -23488 -11068 -23237
rect -11193 -23505 -11068 -23488
rect -11193 -23539 -11176 -23505
rect -11142 -23539 -11068 -23505
rect -11193 -23553 -11068 -23539
rect -11289 -23635 -11277 -23601
rect -11243 -23635 -11221 -23601
rect -11289 -23651 -11221 -23635
rect -11090 -23683 -11068 -23553
rect -11923 -23731 -11901 -23697
rect -11799 -23731 -11776 -23697
rect -11923 -23743 -11776 -23731
rect -11462 -23889 -11319 -23684
rect -11278 -23697 -11068 -23683
rect -11022 -23697 -10999 -23237
rect -11278 -23731 -11262 -23697
rect -11156 -23731 -10999 -23697
rect -11278 -23738 -10999 -23731
rect -12688 -23949 -12602 -23946
rect -12688 -23951 -11482 -23949
rect -12688 -23952 -12676 -23951
rect -12736 -24014 -12676 -23952
rect -12613 -23960 -11482 -23951
rect -12613 -24014 -11563 -23960
rect -12736 -24016 -11563 -24014
rect -12612 -24029 -11563 -24016
rect -11494 -24029 -11482 -23960
rect -12612 -24035 -11482 -24029
rect -11435 -24076 -11346 -23889
rect -12738 -24092 -11346 -24076
rect -12738 -24163 -12685 -24092
rect -12614 -24163 -11346 -24092
rect -12738 -24164 -11346 -24163
rect -12612 -24165 -11346 -24164
rect -10695 -24593 -10606 -22334
rect -6030 -24356 -5982 -18656
rect -6032 -24362 -5980 -24356
rect -5852 -24358 -5804 -18176
rect -5700 -22398 -5652 -17716
rect -5584 -20422 -5536 -17256
rect -5592 -20474 -5586 -20422
rect -5534 -20474 -5528 -20422
rect -5702 -22404 -5650 -22398
rect -5702 -22462 -5650 -22456
rect -5860 -24410 -5854 -24358
rect -5802 -24410 -5796 -24358
rect -6032 -24420 -5980 -24414
rect -5396 -24593 -5307 -17252
rect -5234 -17314 -5186 -16776
rect -4932 -16814 -4888 -16723
rect -4854 -16745 -4816 -16723
rect -4782 -16745 -4624 -16666
rect -4590 -16745 -4574 -16666
rect -4854 -16751 -4574 -16745
rect -4528 -16672 -4326 -16660
rect -4854 -16814 -4812 -16751
rect -4528 -16783 -4366 -16672
rect -4932 -16874 -4812 -16814
rect -4784 -16789 -4366 -16783
rect -4784 -16866 -4720 -16789
rect -4686 -16866 -4528 -16789
rect -4494 -16848 -4366 -16789
rect -4332 -16848 -4326 -16672
rect -4494 -16860 -4326 -16848
rect -4285 -16672 -4135 -16660
rect -4285 -16848 -4278 -16672
rect -4244 -16691 -4135 -16672
rect -4244 -16823 -4176 -16691
rect -4142 -16823 -4135 -16691
rect -4244 -16848 -4135 -16823
rect -4285 -16860 -4135 -16848
rect -2216 -16714 -2096 -16658
rect -2216 -16805 -2172 -16714
rect -2138 -16777 -2096 -16714
rect -2068 -16536 -1555 -16520
rect -2068 -16570 -2052 -16536
rect -1826 -16570 -1606 -16536
rect -1572 -16570 -1555 -16536
rect -2068 -16640 -1555 -16570
rect -1516 -16531 -1419 -16489
rect -1516 -16628 -1288 -16531
rect -1191 -16628 -1185 -16531
rect -2068 -16662 -1616 -16640
rect -2068 -16739 -2004 -16662
rect -1970 -16739 -1812 -16662
rect -1778 -16668 -1616 -16662
rect -1516 -16668 -1419 -16628
rect -1778 -16680 -1610 -16668
rect -1778 -16739 -1650 -16680
rect -2068 -16745 -1650 -16739
rect -2138 -16783 -1858 -16777
rect -2138 -16805 -2100 -16783
rect -4494 -16866 -4332 -16860
rect -4784 -16888 -4332 -16866
rect -2216 -16862 -2100 -16805
rect -2066 -16862 -1908 -16783
rect -1874 -16862 -1858 -16783
rect -2216 -16868 -1858 -16862
rect -1812 -16856 -1650 -16745
rect -1616 -16856 -1610 -16680
rect -1812 -16868 -1610 -16856
rect -1569 -16680 -1419 -16668
rect -1569 -16856 -1562 -16680
rect -1528 -16705 -1419 -16680
rect -1528 -16837 -1460 -16705
rect -1426 -16837 -1419 -16705
rect -116 -16706 -57 -12682
rect 59 -16557 125 -12549
rect 229 -16409 295 -12387
rect 407 -15427 473 -11789
rect 407 -15499 473 -15493
rect 229 -16475 1433 -16409
rect 59 -16623 1287 -16557
rect -116 -16765 1137 -16706
rect -1528 -16856 -1419 -16837
rect -1569 -16868 -1419 -16856
rect -5048 -16958 -4864 -16903
rect -5048 -17021 -5000 -16958
rect -4937 -17000 -4864 -16958
rect -4784 -16972 -3774 -16888
rect -4056 -16980 -3774 -16972
rect -2332 -16915 -1555 -16899
rect -2332 -16949 -2052 -16915
rect -1826 -16949 -1606 -16915
rect -1572 -16949 -1555 -16915
rect -2332 -16958 -1555 -16949
rect -4937 -17019 -4271 -17000
rect -4937 -17021 -4768 -17019
rect -5048 -17053 -4768 -17021
rect -4542 -17053 -4322 -17019
rect -4288 -17053 -4271 -17019
rect -5048 -17069 -4271 -17053
rect -4056 -17064 -2524 -16980
rect -3958 -17069 -3774 -17064
rect -4932 -17106 -4574 -17100
rect -4932 -17163 -4816 -17106
rect -4932 -17254 -4888 -17163
rect -4854 -17185 -4816 -17163
rect -4782 -17185 -4624 -17106
rect -4590 -17185 -4574 -17106
rect -4854 -17191 -4574 -17185
rect -4528 -17112 -4326 -17100
rect -4854 -17254 -4812 -17191
rect -4528 -17223 -4366 -17112
rect -4932 -17310 -4812 -17254
rect -5236 -17320 -5184 -17314
rect -5236 -17378 -5184 -17372
rect -5048 -17344 -4812 -17310
rect -5048 -17448 -5020 -17344
rect -4916 -17448 -4812 -17344
rect -4784 -17229 -4366 -17223
rect -4784 -17306 -4720 -17229
rect -4686 -17306 -4528 -17229
rect -4494 -17288 -4366 -17229
rect -4332 -17288 -4326 -17112
rect -4494 -17300 -4326 -17288
rect -4285 -17112 -4135 -17100
rect -4285 -17288 -4278 -17112
rect -4244 -17131 -4135 -17112
rect -4244 -17263 -4176 -17131
rect -4142 -17263 -4135 -17131
rect -4244 -17288 -4135 -17263
rect -4285 -17300 -4135 -17288
rect -4494 -17306 -4332 -17300
rect -4784 -17328 -4332 -17306
rect -4784 -17398 -4271 -17328
rect -4784 -17432 -4768 -17398
rect -4542 -17432 -4322 -17398
rect -4288 -17432 -4271 -17398
rect -4784 -17448 -4271 -17432
rect -4232 -17340 -4135 -17300
rect -4232 -17437 -4004 -17340
rect -3907 -17437 -3901 -17340
rect -5048 -17479 -4812 -17448
rect -4232 -17479 -4135 -17437
rect -5048 -17480 -4574 -17479
rect -4932 -17485 -4574 -17480
rect -4932 -17542 -4816 -17485
rect -4932 -17633 -4888 -17542
rect -4854 -17564 -4816 -17542
rect -4782 -17564 -4624 -17485
rect -4590 -17564 -4574 -17485
rect -4854 -17570 -4574 -17564
rect -4528 -17491 -4326 -17479
rect -4854 -17633 -4812 -17570
rect -4528 -17602 -4366 -17491
rect -4932 -17693 -4812 -17633
rect -4784 -17608 -4366 -17602
rect -4784 -17685 -4720 -17608
rect -4686 -17685 -4528 -17608
rect -4494 -17667 -4366 -17608
rect -4332 -17667 -4326 -17491
rect -4494 -17679 -4326 -17667
rect -4285 -17491 -4135 -17479
rect -4285 -17667 -4278 -17491
rect -4244 -17510 -4135 -17491
rect -4244 -17642 -4176 -17510
rect -4142 -17642 -4135 -17510
rect -4244 -17667 -4135 -17642
rect -4285 -17679 -4135 -17667
rect -4494 -17685 -4332 -17679
rect -4784 -17707 -4332 -17685
rect -5048 -17780 -4864 -17722
rect -5048 -17841 -4979 -17780
rect -4918 -17819 -4864 -17780
rect -4784 -17791 -2674 -17707
rect -4918 -17838 -4271 -17819
rect -4918 -17841 -4768 -17838
rect -5048 -17872 -4768 -17841
rect -4542 -17872 -4322 -17838
rect -4288 -17872 -4271 -17838
rect -5048 -17888 -4271 -17872
rect -3958 -17888 -3774 -17791
rect -4932 -17925 -4574 -17919
rect -4932 -17982 -4816 -17925
rect -4932 -18073 -4888 -17982
rect -4854 -18004 -4816 -17982
rect -4782 -18004 -4624 -17925
rect -4590 -18004 -4574 -17925
rect -4854 -18010 -4574 -18004
rect -4528 -17931 -4326 -17919
rect -4854 -18073 -4812 -18010
rect -4528 -18042 -4366 -17931
rect -4932 -18129 -4812 -18073
rect -5048 -18163 -4812 -18129
rect -5048 -18267 -5020 -18163
rect -4916 -18267 -4812 -18163
rect -4784 -18048 -4366 -18042
rect -4784 -18125 -4720 -18048
rect -4686 -18125 -4528 -18048
rect -4494 -18107 -4366 -18048
rect -4332 -18107 -4326 -17931
rect -4494 -18119 -4326 -18107
rect -4285 -17931 -4135 -17919
rect -4285 -18107 -4278 -17931
rect -4244 -17950 -4135 -17931
rect -4244 -18082 -4176 -17950
rect -4142 -18082 -4135 -17950
rect -4244 -18107 -4135 -18082
rect -4285 -18119 -4135 -18107
rect -4494 -18125 -4332 -18119
rect -4784 -18147 -4332 -18125
rect -4784 -18217 -4271 -18147
rect -4784 -18251 -4768 -18217
rect -4542 -18251 -4322 -18217
rect -4288 -18251 -4271 -18217
rect -4784 -18267 -4271 -18251
rect -4232 -18159 -4135 -18119
rect -4232 -18256 -4004 -18159
rect -3907 -18256 -3901 -18159
rect -5048 -18298 -4812 -18267
rect -4232 -18298 -4135 -18256
rect -5048 -18299 -4574 -18298
rect -4932 -18304 -4574 -18299
rect -4932 -18361 -4816 -18304
rect -4932 -18452 -4888 -18361
rect -4854 -18383 -4816 -18361
rect -4782 -18383 -4624 -18304
rect -4590 -18383 -4574 -18304
rect -4854 -18389 -4574 -18383
rect -4528 -18310 -4326 -18298
rect -4854 -18452 -4812 -18389
rect -4528 -18421 -4366 -18310
rect -4932 -18512 -4812 -18452
rect -4784 -18427 -4366 -18421
rect -4784 -18504 -4720 -18427
rect -4686 -18504 -4528 -18427
rect -4494 -18486 -4366 -18427
rect -4332 -18486 -4326 -18310
rect -4494 -18498 -4326 -18486
rect -4285 -18310 -4135 -18298
rect -4285 -18486 -4278 -18310
rect -4244 -18329 -4135 -18310
rect -4244 -18461 -4176 -18329
rect -4142 -18461 -4135 -18329
rect -4244 -18486 -4135 -18461
rect -4285 -18498 -4135 -18486
rect -4494 -18504 -4332 -18498
rect -4784 -18526 -4332 -18504
rect -5048 -18582 -4864 -18541
rect -5048 -18654 -5006 -18582
rect -4934 -18638 -4864 -18582
rect -4784 -18610 -2830 -18526
rect -4934 -18654 -4271 -18638
rect -5048 -18657 -4271 -18654
rect -5048 -18691 -4768 -18657
rect -4542 -18691 -4322 -18657
rect -4288 -18691 -4271 -18657
rect -5048 -18707 -4271 -18691
rect -3958 -18707 -3774 -18610
rect -4932 -18744 -4574 -18738
rect -4932 -18801 -4816 -18744
rect -4932 -18892 -4888 -18801
rect -4854 -18823 -4816 -18801
rect -4782 -18823 -4624 -18744
rect -4590 -18823 -4574 -18744
rect -4854 -18829 -4574 -18823
rect -4528 -18750 -4326 -18738
rect -4854 -18892 -4812 -18829
rect -4528 -18861 -4366 -18750
rect -4932 -18948 -4812 -18892
rect -5048 -18982 -4812 -18948
rect -5048 -19086 -5020 -18982
rect -4916 -19086 -4812 -18982
rect -4784 -18867 -4366 -18861
rect -4784 -18944 -4720 -18867
rect -4686 -18944 -4528 -18867
rect -4494 -18926 -4366 -18867
rect -4332 -18926 -4326 -18750
rect -4494 -18938 -4326 -18926
rect -4285 -18750 -4135 -18738
rect -4285 -18926 -4278 -18750
rect -4244 -18769 -4135 -18750
rect -4244 -18901 -4176 -18769
rect -4142 -18901 -4135 -18769
rect -4244 -18926 -4135 -18901
rect -4285 -18938 -4135 -18926
rect -4494 -18944 -4332 -18938
rect -4784 -18966 -4332 -18944
rect -4784 -19036 -4271 -18966
rect -4784 -19070 -4768 -19036
rect -4542 -19070 -4322 -19036
rect -4288 -19070 -4271 -19036
rect -4784 -19086 -4271 -19070
rect -4232 -18978 -4135 -18938
rect -4232 -19075 -4004 -18978
rect -3907 -19075 -3901 -18978
rect -5048 -19117 -4812 -19086
rect -4232 -19117 -4135 -19075
rect -5048 -19118 -4574 -19117
rect -4932 -19123 -4574 -19118
rect -4932 -19180 -4816 -19123
rect -4932 -19271 -4888 -19180
rect -4854 -19202 -4816 -19180
rect -4782 -19202 -4624 -19123
rect -4590 -19202 -4574 -19123
rect -4854 -19208 -4574 -19202
rect -4528 -19129 -4326 -19117
rect -4854 -19271 -4812 -19208
rect -4528 -19240 -4366 -19129
rect -4932 -19331 -4812 -19271
rect -4784 -19246 -4366 -19240
rect -4784 -19323 -4720 -19246
rect -4686 -19323 -4528 -19246
rect -4494 -19305 -4366 -19246
rect -4332 -19305 -4326 -19129
rect -4494 -19317 -4326 -19305
rect -4285 -19129 -4135 -19117
rect -4285 -19305 -4278 -19129
rect -4244 -19148 -4135 -19129
rect -4244 -19280 -4176 -19148
rect -4142 -19280 -4135 -19148
rect -4244 -19305 -4135 -19280
rect -4285 -19317 -4135 -19305
rect -4494 -19323 -4332 -19317
rect -4784 -19345 -4332 -19323
rect -5048 -19430 -4864 -19360
rect -4784 -19429 -2998 -19345
rect -5048 -19502 -5014 -19430
rect -4942 -19457 -4864 -19430
rect -4942 -19476 -4271 -19457
rect -4942 -19502 -4768 -19476
rect -5048 -19510 -4768 -19502
rect -4542 -19510 -4322 -19476
rect -4288 -19510 -4271 -19476
rect -5048 -19526 -4271 -19510
rect -3958 -19526 -3774 -19429
rect -4932 -19563 -4574 -19557
rect -4932 -19620 -4816 -19563
rect -4932 -19711 -4888 -19620
rect -4854 -19642 -4816 -19620
rect -4782 -19642 -4624 -19563
rect -4590 -19642 -4574 -19563
rect -4854 -19648 -4574 -19642
rect -4528 -19569 -4326 -19557
rect -4854 -19711 -4812 -19648
rect -4528 -19680 -4366 -19569
rect -4932 -19767 -4812 -19711
rect -5048 -19801 -4812 -19767
rect -5048 -19905 -5020 -19801
rect -4916 -19905 -4812 -19801
rect -4784 -19686 -4366 -19680
rect -4784 -19763 -4720 -19686
rect -4686 -19763 -4528 -19686
rect -4494 -19745 -4366 -19686
rect -4332 -19745 -4326 -19569
rect -4494 -19757 -4326 -19745
rect -4285 -19569 -4135 -19557
rect -4285 -19745 -4278 -19569
rect -4244 -19588 -4135 -19569
rect -4244 -19720 -4176 -19588
rect -4142 -19720 -4135 -19588
rect -4244 -19745 -4135 -19720
rect -4285 -19757 -4135 -19745
rect -4494 -19763 -4332 -19757
rect -4784 -19785 -4332 -19763
rect -4784 -19855 -4271 -19785
rect -4784 -19889 -4768 -19855
rect -4542 -19889 -4322 -19855
rect -4288 -19889 -4271 -19855
rect -4784 -19905 -4271 -19889
rect -4232 -19797 -4135 -19757
rect -4232 -19894 -4004 -19797
rect -3907 -19894 -3901 -19797
rect -5048 -19936 -4812 -19905
rect -4232 -19936 -4135 -19894
rect -5048 -19937 -4574 -19936
rect -4932 -19942 -4574 -19937
rect -4932 -19999 -4816 -19942
rect -5174 -20056 -5074 -20044
rect -5174 -20128 -5166 -20056
rect -5094 -20128 -5074 -20056
rect -5174 -20134 -5074 -20128
rect -4932 -20090 -4888 -19999
rect -4854 -20021 -4816 -19999
rect -4782 -20021 -4624 -19942
rect -4590 -20021 -4574 -19942
rect -4854 -20027 -4574 -20021
rect -4528 -19948 -4326 -19936
rect -4854 -20090 -4812 -20027
rect -4528 -20059 -4366 -19948
rect -5166 -20202 -5094 -20134
rect -4932 -20150 -4812 -20090
rect -4784 -20065 -4366 -20059
rect -4784 -20142 -4720 -20065
rect -4686 -20142 -4528 -20065
rect -4494 -20124 -4366 -20065
rect -4332 -20124 -4326 -19948
rect -4494 -20136 -4326 -20124
rect -4285 -19948 -4135 -19936
rect -4285 -20124 -4278 -19948
rect -4244 -19967 -4135 -19948
rect -4244 -20099 -4176 -19967
rect -4142 -20099 -4135 -19967
rect -4244 -20124 -4135 -20099
rect -4285 -20136 -4135 -20124
rect -4494 -20142 -4332 -20136
rect -4784 -20164 -4332 -20142
rect -5048 -20202 -4864 -20179
rect -5166 -20274 -4864 -20202
rect -4784 -20248 -3176 -20164
rect -5048 -20276 -4864 -20274
rect -5048 -20295 -4271 -20276
rect -5048 -20329 -4768 -20295
rect -4542 -20329 -4322 -20295
rect -4288 -20329 -4271 -20295
rect -5048 -20345 -4271 -20329
rect -3958 -20345 -3774 -20248
rect -4932 -20382 -4574 -20376
rect -4932 -20439 -4816 -20382
rect -4932 -20530 -4888 -20439
rect -4854 -20461 -4816 -20439
rect -4782 -20461 -4624 -20382
rect -4590 -20461 -4574 -20382
rect -4854 -20467 -4574 -20461
rect -4528 -20388 -4326 -20376
rect -4854 -20530 -4812 -20467
rect -4528 -20499 -4366 -20388
rect -4932 -20586 -4812 -20530
rect -5048 -20620 -4812 -20586
rect -5048 -20724 -5020 -20620
rect -4916 -20724 -4812 -20620
rect -4784 -20505 -4366 -20499
rect -4784 -20582 -4720 -20505
rect -4686 -20582 -4528 -20505
rect -4494 -20564 -4366 -20505
rect -4332 -20564 -4326 -20388
rect -4494 -20576 -4326 -20564
rect -4285 -20388 -4135 -20376
rect -4285 -20564 -4278 -20388
rect -4244 -20407 -4135 -20388
rect -4244 -20539 -4176 -20407
rect -4142 -20539 -4135 -20407
rect -4244 -20564 -4135 -20539
rect -4285 -20576 -4135 -20564
rect -4494 -20582 -4332 -20576
rect -4784 -20604 -4332 -20582
rect -4784 -20674 -4271 -20604
rect -4784 -20708 -4768 -20674
rect -4542 -20708 -4322 -20674
rect -4288 -20708 -4271 -20674
rect -4784 -20724 -4271 -20708
rect -4232 -20616 -4135 -20576
rect -4232 -20713 -4004 -20616
rect -3907 -20713 -3901 -20616
rect -5048 -20755 -4812 -20724
rect -4232 -20755 -4135 -20713
rect -5048 -20756 -4574 -20755
rect -4932 -20761 -4574 -20756
rect -4932 -20818 -4816 -20761
rect -4932 -20909 -4888 -20818
rect -4854 -20840 -4816 -20818
rect -4782 -20840 -4624 -20761
rect -4590 -20840 -4574 -20761
rect -4854 -20846 -4574 -20840
rect -4528 -20767 -4326 -20755
rect -4854 -20909 -4812 -20846
rect -4528 -20878 -4366 -20767
rect -4932 -20969 -4812 -20909
rect -4784 -20884 -4366 -20878
rect -4784 -20961 -4720 -20884
rect -4686 -20961 -4528 -20884
rect -4494 -20943 -4366 -20884
rect -4332 -20943 -4326 -20767
rect -4494 -20955 -4326 -20943
rect -4285 -20767 -4135 -20755
rect -4285 -20943 -4278 -20767
rect -4244 -20786 -4135 -20767
rect -4244 -20918 -4176 -20786
rect -4142 -20918 -4135 -20786
rect -4244 -20943 -4135 -20918
rect -4285 -20955 -4135 -20943
rect -4494 -20961 -4332 -20955
rect -4784 -20983 -4332 -20961
rect -4784 -21046 -3774 -20983
rect -4784 -21067 -3906 -21046
rect -3958 -21130 -3906 -21067
rect -3822 -21130 -3774 -21046
rect -3958 -21164 -3774 -21130
rect -5130 -21525 -5047 -21519
rect -5130 -22437 -5047 -21608
rect -5140 -22520 -5047 -22437
rect -10695 -24682 -5298 -24593
rect -5396 -24688 -5307 -24682
rect -5130 -24796 -5047 -22520
rect -10647 -24879 -5047 -24796
rect -10647 -24987 -10563 -24879
rect -11457 -25070 -10563 -24987
rect -6038 -25036 -6032 -24984
rect -5980 -25036 -5974 -24984
rect -13016 -25112 -12964 -25106
rect -13016 -25170 -12964 -25164
rect -11457 -25177 -11374 -25070
rect -10479 -25107 -10393 -25096
rect -17982 -25546 -17216 -25480
rect -12499 -25313 -12173 -25301
rect -12499 -25343 -12293 -25313
rect -17982 -25553 -17878 -25546
rect -17982 -25642 -17976 -25553
rect -17887 -25642 -17878 -25553
rect -17982 -25650 -17878 -25642
rect -12499 -26465 -12471 -25343
rect -12399 -25347 -12293 -25343
rect -12191 -25347 -12173 -25313
rect -12399 -25505 -12173 -25347
rect -11923 -25313 -11776 -25301
rect -11923 -25347 -11902 -25313
rect -11835 -25347 -11776 -25313
rect -12399 -25539 -12293 -25505
rect -12191 -25539 -12173 -25505
rect -12399 -25555 -12173 -25539
rect -12135 -25409 -11956 -25393
rect -12135 -25443 -12109 -25409
rect -11985 -25443 -11956 -25409
rect -12399 -26257 -12365 -25555
rect -12135 -25601 -11956 -25443
rect -11923 -25505 -11776 -25347
rect -11541 -25314 -11332 -25177
rect -11541 -25348 -11411 -25314
rect -11448 -25379 -11411 -25348
rect -11356 -25379 -11332 -25314
rect -11278 -25313 -10999 -25304
rect -11278 -25347 -11262 -25313
rect -11156 -25342 -10999 -25313
rect -11156 -25347 -11068 -25342
rect -11278 -25359 -11068 -25347
rect -11448 -25390 -11332 -25379
rect -11289 -25409 -11221 -25393
rect -11289 -25443 -11277 -25409
rect -11243 -25443 -11221 -25409
rect -11923 -25539 -11902 -25505
rect -11835 -25539 -11776 -25505
rect -11923 -25555 -11776 -25539
rect -11601 -25481 -11331 -25464
rect -11601 -25561 -11582 -25481
rect -11514 -25561 -11331 -25481
rect -11601 -25579 -11331 -25561
rect -12135 -25635 -12110 -25601
rect -11986 -25635 -11956 -25601
rect -12320 -25697 -12173 -25681
rect -12320 -25731 -12293 -25697
rect -12191 -25731 -12173 -25697
rect -12320 -25889 -12173 -25731
rect -12320 -25923 -12293 -25889
rect -12191 -25923 -12173 -25889
rect -12320 -26081 -12173 -25923
rect -12320 -26115 -12294 -26081
rect -12192 -26115 -12173 -26081
rect -12320 -26131 -12173 -26115
rect -12135 -25793 -11956 -25635
rect -11601 -25681 -11502 -25649
rect -12135 -25827 -12110 -25793
rect -11986 -25827 -11956 -25793
rect -12135 -25985 -11956 -25827
rect -12135 -26019 -12110 -25985
rect -11986 -26019 -11956 -25985
rect -12135 -26177 -11956 -26019
rect -11912 -25697 -11820 -25681
rect -11912 -25731 -11895 -25697
rect -11835 -25731 -11820 -25697
rect -11912 -25889 -11820 -25731
rect -11912 -25923 -11878 -25889
rect -11835 -25923 -11820 -25889
rect -11912 -26081 -11820 -25923
rect -11912 -26115 -11895 -26081
rect -11835 -26115 -11820 -26081
rect -11912 -26131 -11820 -26115
rect -11601 -25795 -11583 -25681
rect -11530 -25795 -11502 -25681
rect -12135 -26211 -12110 -26177
rect -11986 -26211 -11956 -26177
rect -12399 -26273 -12173 -26257
rect -12399 -26307 -12296 -26273
rect -12194 -26307 -12173 -26273
rect -12399 -26465 -12173 -26307
rect -12135 -26369 -11956 -26211
rect -12135 -26403 -12110 -26369
rect -11986 -26403 -11956 -26369
rect -12135 -26419 -11956 -26403
rect -11923 -26273 -11776 -26257
rect -11923 -26307 -11901 -26273
rect -11835 -26307 -11776 -26273
rect -12499 -26499 -12296 -26465
rect -12194 -26499 -12173 -26465
rect -12499 -26511 -12173 -26499
rect -11923 -26465 -11776 -26307
rect -11601 -26268 -11502 -25795
rect -11601 -26401 -11575 -26268
rect -11522 -26401 -11502 -26268
rect -11601 -26438 -11502 -26401
rect -11417 -26452 -11331 -25579
rect -11289 -25601 -11221 -25443
rect -11090 -25490 -11068 -25359
rect -11192 -25505 -11068 -25490
rect -11192 -25539 -11176 -25505
rect -11142 -25539 -11068 -25505
rect -11192 -25555 -11068 -25539
rect -11289 -25635 -11277 -25601
rect -11243 -25635 -11221 -25601
rect -11289 -25793 -11221 -25635
rect -11289 -25827 -11277 -25793
rect -11243 -25827 -11221 -25793
rect -11289 -25843 -11221 -25827
rect -11188 -25697 -11124 -25681
rect -11188 -25731 -11176 -25697
rect -11142 -25731 -11124 -25697
rect -11188 -25889 -11124 -25731
rect -11188 -25923 -11176 -25889
rect -11142 -25923 -11124 -25889
rect -11289 -25985 -11221 -25969
rect -11289 -26019 -11276 -25985
rect -11242 -26019 -11221 -25985
rect -11289 -26177 -11221 -26019
rect -11188 -26081 -11124 -25923
rect -11188 -26115 -11176 -26081
rect -11142 -26115 -11124 -26081
rect -11188 -26128 -11124 -26115
rect -11090 -25945 -11068 -25555
rect -11022 -25945 -10999 -25342
rect -11090 -26005 -11079 -25945
rect -11019 -26005 -10999 -25945
rect -11289 -26211 -11277 -26177
rect -11243 -26211 -11221 -26177
rect -11289 -26369 -11221 -26211
rect -11090 -26256 -11068 -26005
rect -11193 -26273 -11068 -26256
rect -11193 -26307 -11176 -26273
rect -11142 -26307 -11068 -26273
rect -11193 -26321 -11068 -26307
rect -11289 -26403 -11277 -26369
rect -11243 -26403 -11221 -26369
rect -11289 -26419 -11221 -26403
rect -11090 -26451 -11068 -26321
rect -11923 -26499 -11901 -26465
rect -11799 -26499 -11776 -26465
rect -11923 -26511 -11776 -26499
rect -11462 -26657 -11319 -26452
rect -11278 -26465 -11068 -26451
rect -11022 -26465 -10999 -26005
rect -11278 -26499 -11262 -26465
rect -11156 -26499 -10999 -26465
rect -11278 -26506 -10999 -26499
rect -12612 -26742 -11480 -26736
rect -12770 -26744 -11480 -26742
rect -12770 -26805 -12743 -26744
rect -12682 -26748 -11480 -26744
rect -12682 -26805 -11564 -26748
rect -12770 -26806 -11564 -26805
rect -12612 -26820 -11564 -26806
rect -11492 -26820 -11480 -26748
rect -12612 -26832 -11480 -26820
rect -11436 -26917 -11344 -26657
rect -12612 -26934 -11344 -26917
rect -12794 -26998 -12748 -26934
rect -12684 -26998 -11344 -26934
rect -12612 -27009 -11344 -26998
rect -10479 -27674 -10393 -25193
rect -11454 -27760 -10393 -27674
rect -10152 -25530 -10048 -25524
rect -11454 -27810 -11368 -27760
rect -12499 -27946 -12173 -27934
rect -12499 -27976 -12293 -27946
rect -12499 -29098 -12471 -27976
rect -12399 -27980 -12293 -27976
rect -12191 -27980 -12173 -27946
rect -12399 -28138 -12173 -27980
rect -11923 -27946 -11776 -27934
rect -11923 -27980 -11902 -27946
rect -11835 -27980 -11776 -27946
rect -12399 -28172 -12293 -28138
rect -12191 -28172 -12173 -28138
rect -12399 -28188 -12173 -28172
rect -12135 -28042 -11956 -28026
rect -12135 -28076 -12109 -28042
rect -11985 -28076 -11956 -28042
rect -12399 -28890 -12365 -28188
rect -12135 -28234 -11956 -28076
rect -11923 -28138 -11776 -27980
rect -11541 -27947 -11332 -27810
rect -11541 -27981 -11411 -27947
rect -11448 -28012 -11411 -27981
rect -11356 -28012 -11332 -27947
rect -11278 -27946 -10999 -27937
rect -11278 -27980 -11262 -27946
rect -11156 -27975 -10999 -27946
rect -10152 -27954 -10048 -25634
rect -11156 -27980 -11068 -27975
rect -11278 -27992 -11068 -27980
rect -11448 -28023 -11332 -28012
rect -11289 -28042 -11221 -28026
rect -11289 -28076 -11277 -28042
rect -11243 -28076 -11221 -28042
rect -11923 -28172 -11902 -28138
rect -11835 -28172 -11776 -28138
rect -11923 -28188 -11776 -28172
rect -11601 -28114 -11331 -28097
rect -11601 -28194 -11582 -28114
rect -11514 -28194 -11331 -28114
rect -11601 -28212 -11331 -28194
rect -12135 -28268 -12110 -28234
rect -11986 -28268 -11956 -28234
rect -12320 -28330 -12173 -28314
rect -12320 -28364 -12293 -28330
rect -12191 -28364 -12173 -28330
rect -12320 -28522 -12173 -28364
rect -12320 -28556 -12293 -28522
rect -12191 -28556 -12173 -28522
rect -12320 -28714 -12173 -28556
rect -12320 -28748 -12294 -28714
rect -12192 -28748 -12173 -28714
rect -12320 -28764 -12173 -28748
rect -12135 -28426 -11956 -28268
rect -11601 -28314 -11502 -28282
rect -12135 -28460 -12110 -28426
rect -11986 -28460 -11956 -28426
rect -12135 -28618 -11956 -28460
rect -12135 -28652 -12110 -28618
rect -11986 -28652 -11956 -28618
rect -12135 -28810 -11956 -28652
rect -11912 -28330 -11820 -28314
rect -11912 -28364 -11895 -28330
rect -11835 -28364 -11820 -28330
rect -11912 -28522 -11820 -28364
rect -11912 -28556 -11878 -28522
rect -11835 -28556 -11820 -28522
rect -11912 -28714 -11820 -28556
rect -11912 -28748 -11895 -28714
rect -11835 -28748 -11820 -28714
rect -11912 -28764 -11820 -28748
rect -11601 -28428 -11583 -28314
rect -11530 -28428 -11502 -28314
rect -12135 -28844 -12110 -28810
rect -11986 -28844 -11956 -28810
rect -12399 -28906 -12173 -28890
rect -12399 -28940 -12296 -28906
rect -12194 -28940 -12173 -28906
rect -12399 -29098 -12173 -28940
rect -12135 -29002 -11956 -28844
rect -12135 -29036 -12110 -29002
rect -11986 -29036 -11956 -29002
rect -12135 -29052 -11956 -29036
rect -11923 -28906 -11776 -28890
rect -11923 -28940 -11901 -28906
rect -11835 -28940 -11776 -28906
rect -12499 -29132 -12296 -29098
rect -12194 -29132 -12173 -29098
rect -12499 -29144 -12173 -29132
rect -11923 -29098 -11776 -28940
rect -11601 -28901 -11502 -28428
rect -11601 -29034 -11575 -28901
rect -11522 -29034 -11502 -28901
rect -11601 -29071 -11502 -29034
rect -11417 -29085 -11331 -28212
rect -11289 -28234 -11221 -28076
rect -11090 -28123 -11068 -27992
rect -11192 -28138 -11068 -28123
rect -11192 -28172 -11176 -28138
rect -11142 -28172 -11068 -28138
rect -11192 -28188 -11068 -28172
rect -11289 -28268 -11277 -28234
rect -11243 -28268 -11221 -28234
rect -11289 -28426 -11221 -28268
rect -11289 -28460 -11277 -28426
rect -11243 -28460 -11221 -28426
rect -11289 -28476 -11221 -28460
rect -11188 -28330 -11124 -28314
rect -11188 -28364 -11176 -28330
rect -11142 -28364 -11124 -28330
rect -11188 -28522 -11124 -28364
rect -11188 -28556 -11176 -28522
rect -11142 -28556 -11124 -28522
rect -11289 -28618 -11221 -28602
rect -11289 -28652 -11276 -28618
rect -11242 -28652 -11221 -28618
rect -11289 -28810 -11221 -28652
rect -11188 -28714 -11124 -28556
rect -11188 -28748 -11176 -28714
rect -11142 -28748 -11124 -28714
rect -11188 -28761 -11124 -28748
rect -11090 -28578 -11068 -28188
rect -11022 -28578 -10999 -27975
rect -11090 -28638 -11079 -28578
rect -11019 -28638 -10999 -28578
rect -11289 -28844 -11277 -28810
rect -11243 -28844 -11221 -28810
rect -11289 -29002 -11221 -28844
rect -11090 -28889 -11068 -28638
rect -11193 -28906 -11068 -28889
rect -11193 -28940 -11176 -28906
rect -11142 -28940 -11068 -28906
rect -11193 -28954 -11068 -28940
rect -11289 -29036 -11277 -29002
rect -11243 -29036 -11221 -29002
rect -11289 -29052 -11221 -29036
rect -11090 -29084 -11068 -28954
rect -11923 -29132 -11901 -29098
rect -11799 -29132 -11776 -29098
rect -11923 -29144 -11776 -29132
rect -11462 -29290 -11319 -29085
rect -11278 -29098 -11068 -29084
rect -11022 -29098 -10999 -28638
rect -11278 -29132 -11262 -29098
rect -11156 -29132 -10999 -29098
rect -11278 -29139 -10999 -29132
rect -10366 -28058 -10048 -27954
rect -12612 -29374 -11488 -29373
rect -12758 -29446 -12724 -29374
rect -12652 -29385 -11488 -29374
rect -12652 -29446 -11562 -29385
rect -12612 -29453 -11562 -29446
rect -11494 -29453 -11488 -29385
rect -12612 -29465 -11488 -29453
rect -11437 -29520 -11343 -29290
rect -12772 -29537 -11343 -29520
rect -12772 -29626 -12727 -29537
rect -12638 -29614 -11343 -29537
rect -12638 -29626 -12432 -29614
rect -10366 -30233 -10262 -28058
rect -11452 -30337 -10262 -30233
rect -11452 -30419 -11348 -30337
rect -12499 -30555 -12173 -30543
rect -12499 -30585 -12293 -30555
rect -12499 -31707 -12471 -30585
rect -12399 -30589 -12293 -30585
rect -12191 -30589 -12173 -30555
rect -12399 -30747 -12173 -30589
rect -11923 -30555 -11776 -30543
rect -11923 -30589 -11902 -30555
rect -11835 -30589 -11776 -30555
rect -12399 -30781 -12293 -30747
rect -12191 -30781 -12173 -30747
rect -12399 -30797 -12173 -30781
rect -12135 -30651 -11956 -30635
rect -12135 -30685 -12109 -30651
rect -11985 -30685 -11956 -30651
rect -12399 -31499 -12365 -30797
rect -12135 -30843 -11956 -30685
rect -11923 -30747 -11776 -30589
rect -11541 -30556 -11332 -30419
rect -11541 -30590 -11411 -30556
rect -11448 -30621 -11411 -30590
rect -11356 -30621 -11332 -30556
rect -11278 -30555 -10999 -30546
rect -11278 -30589 -11262 -30555
rect -11156 -30584 -10999 -30555
rect -11156 -30589 -11068 -30584
rect -11278 -30601 -11068 -30589
rect -11448 -30632 -11332 -30621
rect -11289 -30651 -11221 -30635
rect -11289 -30685 -11277 -30651
rect -11243 -30685 -11221 -30651
rect -11923 -30781 -11902 -30747
rect -11835 -30781 -11776 -30747
rect -11923 -30797 -11776 -30781
rect -11601 -30723 -11331 -30706
rect -11601 -30803 -11582 -30723
rect -11514 -30803 -11331 -30723
rect -11601 -30821 -11331 -30803
rect -12135 -30877 -12110 -30843
rect -11986 -30877 -11956 -30843
rect -12320 -30939 -12173 -30923
rect -12320 -30973 -12293 -30939
rect -12191 -30973 -12173 -30939
rect -12320 -31131 -12173 -30973
rect -12320 -31165 -12293 -31131
rect -12191 -31165 -12173 -31131
rect -12320 -31323 -12173 -31165
rect -12320 -31357 -12294 -31323
rect -12192 -31357 -12173 -31323
rect -12320 -31373 -12173 -31357
rect -12135 -31035 -11956 -30877
rect -11601 -30923 -11502 -30891
rect -12135 -31069 -12110 -31035
rect -11986 -31069 -11956 -31035
rect -12135 -31227 -11956 -31069
rect -12135 -31261 -12110 -31227
rect -11986 -31261 -11956 -31227
rect -12135 -31419 -11956 -31261
rect -11912 -30939 -11820 -30923
rect -11912 -30973 -11895 -30939
rect -11835 -30973 -11820 -30939
rect -11912 -31131 -11820 -30973
rect -11912 -31165 -11878 -31131
rect -11835 -31165 -11820 -31131
rect -11912 -31323 -11820 -31165
rect -11912 -31357 -11895 -31323
rect -11835 -31357 -11820 -31323
rect -11912 -31373 -11820 -31357
rect -11601 -31037 -11583 -30923
rect -11530 -31037 -11502 -30923
rect -12135 -31453 -12110 -31419
rect -11986 -31453 -11956 -31419
rect -12399 -31515 -12173 -31499
rect -12399 -31549 -12296 -31515
rect -12194 -31549 -12173 -31515
rect -12399 -31707 -12173 -31549
rect -12135 -31611 -11956 -31453
rect -12135 -31645 -12110 -31611
rect -11986 -31645 -11956 -31611
rect -12135 -31661 -11956 -31645
rect -11923 -31515 -11776 -31499
rect -11923 -31549 -11901 -31515
rect -11835 -31549 -11776 -31515
rect -12499 -31741 -12296 -31707
rect -12194 -31741 -12173 -31707
rect -12499 -31753 -12173 -31741
rect -11923 -31707 -11776 -31549
rect -11601 -31510 -11502 -31037
rect -11601 -31643 -11575 -31510
rect -11522 -31643 -11502 -31510
rect -11601 -31680 -11502 -31643
rect -11417 -31694 -11331 -30821
rect -11289 -30843 -11221 -30685
rect -11090 -30732 -11068 -30601
rect -11192 -30747 -11068 -30732
rect -11192 -30781 -11176 -30747
rect -11142 -30781 -11068 -30747
rect -11192 -30797 -11068 -30781
rect -11289 -30877 -11277 -30843
rect -11243 -30877 -11221 -30843
rect -11289 -31035 -11221 -30877
rect -11289 -31069 -11277 -31035
rect -11243 -31069 -11221 -31035
rect -11289 -31085 -11221 -31069
rect -11188 -30939 -11124 -30923
rect -11188 -30973 -11176 -30939
rect -11142 -30973 -11124 -30939
rect -11188 -31131 -11124 -30973
rect -11188 -31165 -11176 -31131
rect -11142 -31165 -11124 -31131
rect -11289 -31227 -11221 -31211
rect -11289 -31261 -11276 -31227
rect -11242 -31261 -11221 -31227
rect -11289 -31419 -11221 -31261
rect -11188 -31323 -11124 -31165
rect -11188 -31357 -11176 -31323
rect -11142 -31357 -11124 -31323
rect -11188 -31370 -11124 -31357
rect -11090 -31187 -11068 -30797
rect -11022 -31187 -10999 -30584
rect -11090 -31247 -11079 -31187
rect -11019 -31247 -10999 -31187
rect -11289 -31453 -11277 -31419
rect -11243 -31453 -11221 -31419
rect -11289 -31611 -11221 -31453
rect -11090 -31498 -11068 -31247
rect -11193 -31515 -11068 -31498
rect -11193 -31549 -11176 -31515
rect -11142 -31549 -11068 -31515
rect -11193 -31563 -11068 -31549
rect -11289 -31645 -11277 -31611
rect -11243 -31645 -11221 -31611
rect -11289 -31661 -11221 -31645
rect -11090 -31693 -11068 -31563
rect -11923 -31741 -11901 -31707
rect -11799 -31741 -11776 -31707
rect -11923 -31753 -11776 -31741
rect -11462 -31899 -11319 -31694
rect -11278 -31707 -11068 -31693
rect -11022 -31707 -10999 -31247
rect -11278 -31741 -11262 -31707
rect -11156 -31741 -10999 -31707
rect -11278 -31748 -10999 -31741
rect -12834 -31918 -12670 -31900
rect -12834 -31990 -12758 -31918
rect -12686 -31927 -12478 -31918
rect -11576 -31927 -11487 -31915
rect -12686 -31990 -11564 -31927
rect -12612 -31998 -11564 -31990
rect -11493 -31998 -11487 -31927
rect -11576 -32010 -11487 -31998
rect -12612 -32048 -11576 -32047
rect -11432 -32048 -11348 -31899
rect -12838 -32087 -12674 -32086
rect -12612 -32087 -11348 -32048
rect -12838 -32176 -12791 -32087
rect -12702 -32132 -11348 -32087
rect -12702 -32133 -11576 -32132
rect -12702 -32176 -12464 -32133
rect -11497 -33009 -9857 -32916
rect -9764 -33009 -9758 -32916
rect -11497 -33039 -11360 -33009
rect -12501 -33175 -12175 -33163
rect -12501 -33205 -12295 -33175
rect -12501 -34327 -12473 -33205
rect -12401 -33209 -12295 -33205
rect -12193 -33209 -12175 -33175
rect -12401 -33367 -12175 -33209
rect -11925 -33175 -11778 -33163
rect -11925 -33209 -11904 -33175
rect -11837 -33209 -11778 -33175
rect -12401 -33401 -12295 -33367
rect -12193 -33401 -12175 -33367
rect -12401 -33417 -12175 -33401
rect -12137 -33271 -11958 -33255
rect -12137 -33305 -12111 -33271
rect -11987 -33305 -11958 -33271
rect -12401 -34119 -12367 -33417
rect -12137 -33463 -11958 -33305
rect -11925 -33367 -11778 -33209
rect -11543 -33176 -11334 -33039
rect -6030 -33110 -5982 -25036
rect -5860 -25086 -5854 -25034
rect -5802 -25086 -5796 -25034
rect -5852 -25742 -5804 -25086
rect -5860 -25794 -5854 -25742
rect -5802 -25794 -5796 -25742
rect -6032 -33116 -5980 -33110
rect -11543 -33210 -11413 -33176
rect -11450 -33241 -11413 -33210
rect -11358 -33241 -11334 -33176
rect -11280 -33175 -11001 -33166
rect -6032 -33174 -5980 -33168
rect -11280 -33209 -11264 -33175
rect -11158 -33204 -11001 -33175
rect -11158 -33209 -11070 -33204
rect -11280 -33221 -11070 -33209
rect -11450 -33252 -11334 -33241
rect -11291 -33271 -11223 -33255
rect -11291 -33305 -11279 -33271
rect -11245 -33305 -11223 -33271
rect -11925 -33401 -11904 -33367
rect -11837 -33401 -11778 -33367
rect -11925 -33417 -11778 -33401
rect -11603 -33343 -11333 -33326
rect -11603 -33423 -11584 -33343
rect -11516 -33423 -11333 -33343
rect -11603 -33441 -11333 -33423
rect -12137 -33497 -12112 -33463
rect -11988 -33497 -11958 -33463
rect -12322 -33559 -12175 -33543
rect -12322 -33593 -12295 -33559
rect -12193 -33593 -12175 -33559
rect -12322 -33751 -12175 -33593
rect -12322 -33785 -12295 -33751
rect -12193 -33785 -12175 -33751
rect -12322 -33943 -12175 -33785
rect -12322 -33977 -12296 -33943
rect -12194 -33977 -12175 -33943
rect -12322 -33993 -12175 -33977
rect -12137 -33655 -11958 -33497
rect -11603 -33543 -11504 -33511
rect -12137 -33689 -12112 -33655
rect -11988 -33689 -11958 -33655
rect -12137 -33847 -11958 -33689
rect -12137 -33881 -12112 -33847
rect -11988 -33881 -11958 -33847
rect -12137 -34039 -11958 -33881
rect -11914 -33559 -11822 -33543
rect -11914 -33593 -11897 -33559
rect -11837 -33593 -11822 -33559
rect -11914 -33751 -11822 -33593
rect -11914 -33785 -11880 -33751
rect -11837 -33785 -11822 -33751
rect -11914 -33943 -11822 -33785
rect -11914 -33977 -11897 -33943
rect -11837 -33977 -11822 -33943
rect -11914 -33993 -11822 -33977
rect -11603 -33657 -11585 -33543
rect -11532 -33657 -11504 -33543
rect -12137 -34073 -12112 -34039
rect -11988 -34073 -11958 -34039
rect -12401 -34135 -12175 -34119
rect -12401 -34169 -12298 -34135
rect -12196 -34169 -12175 -34135
rect -12401 -34327 -12175 -34169
rect -12137 -34231 -11958 -34073
rect -12137 -34265 -12112 -34231
rect -11988 -34265 -11958 -34231
rect -12137 -34281 -11958 -34265
rect -11925 -34135 -11778 -34119
rect -11925 -34169 -11903 -34135
rect -11837 -34169 -11778 -34135
rect -12501 -34361 -12298 -34327
rect -12196 -34361 -12175 -34327
rect -12501 -34373 -12175 -34361
rect -11925 -34327 -11778 -34169
rect -11603 -34130 -11504 -33657
rect -11603 -34263 -11577 -34130
rect -11524 -34263 -11504 -34130
rect -11603 -34300 -11504 -34263
rect -11419 -34314 -11333 -33441
rect -11291 -33463 -11223 -33305
rect -11092 -33352 -11070 -33221
rect -11194 -33367 -11070 -33352
rect -11194 -33401 -11178 -33367
rect -11144 -33401 -11070 -33367
rect -11194 -33417 -11070 -33401
rect -11291 -33497 -11279 -33463
rect -11245 -33497 -11223 -33463
rect -11291 -33655 -11223 -33497
rect -11291 -33689 -11279 -33655
rect -11245 -33689 -11223 -33655
rect -11291 -33705 -11223 -33689
rect -11190 -33559 -11126 -33543
rect -11190 -33593 -11178 -33559
rect -11144 -33593 -11126 -33559
rect -11190 -33751 -11126 -33593
rect -11190 -33785 -11178 -33751
rect -11144 -33785 -11126 -33751
rect -11291 -33847 -11223 -33831
rect -11291 -33881 -11278 -33847
rect -11244 -33881 -11223 -33847
rect -11291 -34039 -11223 -33881
rect -11190 -33943 -11126 -33785
rect -11190 -33977 -11178 -33943
rect -11144 -33977 -11126 -33943
rect -11190 -33990 -11126 -33977
rect -11092 -33807 -11070 -33417
rect -11024 -33807 -11001 -33204
rect -3260 -33272 -3176 -20248
rect -3082 -25874 -2998 -19429
rect -2914 -22526 -2830 -18610
rect -2751 -21748 -2680 -17791
rect -2608 -17980 -2524 -17064
rect -2332 -17021 -2291 -16958
rect -2228 -16968 -1555 -16958
rect -2228 -17021 -2148 -16968
rect -1242 -16996 -1058 -16899
rect 816 -16996 900 -16992
rect -2332 -17065 -2148 -17021
rect -2068 -17080 914 -16996
rect -2216 -17154 -2096 -17094
rect -2216 -17245 -2172 -17154
rect -2138 -17217 -2096 -17154
rect -2068 -17102 -1616 -17080
rect 674 -17086 758 -17080
rect -2068 -17179 -2004 -17102
rect -1970 -17179 -1812 -17102
rect -1778 -17108 -1616 -17102
rect -1778 -17120 -1610 -17108
rect -1778 -17179 -1650 -17120
rect -2068 -17185 -1650 -17179
rect -2138 -17223 -1858 -17217
rect -2138 -17245 -2100 -17223
rect -2216 -17302 -2100 -17245
rect -2066 -17302 -1908 -17223
rect -1874 -17302 -1858 -17223
rect -2216 -17307 -1858 -17302
rect -2332 -17308 -1858 -17307
rect -1812 -17296 -1650 -17185
rect -1616 -17296 -1610 -17120
rect -1812 -17308 -1610 -17296
rect -1569 -17120 -1419 -17108
rect -1569 -17296 -1562 -17120
rect -1528 -17145 -1419 -17120
rect -1528 -17277 -1460 -17145
rect -1426 -17277 -1419 -17145
rect -1528 -17296 -1419 -17277
rect -1569 -17308 -1419 -17296
rect -2332 -17339 -2096 -17308
rect -2332 -17443 -2304 -17339
rect -2200 -17443 -2096 -17339
rect -2332 -17477 -2096 -17443
rect -2216 -17533 -2096 -17477
rect -2216 -17624 -2172 -17533
rect -2138 -17596 -2096 -17533
rect -2068 -17355 -1555 -17339
rect -2068 -17389 -2052 -17355
rect -1826 -17389 -1606 -17355
rect -1572 -17389 -1555 -17355
rect -2068 -17459 -1555 -17389
rect -1516 -17350 -1419 -17308
rect -1516 -17447 -1288 -17350
rect -1191 -17447 -1185 -17350
rect -2068 -17481 -1616 -17459
rect -2068 -17558 -2004 -17481
rect -1970 -17558 -1812 -17481
rect -1778 -17487 -1616 -17481
rect -1516 -17487 -1419 -17447
rect -1778 -17499 -1610 -17487
rect -1778 -17558 -1650 -17499
rect -2068 -17564 -1650 -17558
rect -2138 -17602 -1858 -17596
rect -2138 -17624 -2100 -17602
rect -2216 -17681 -2100 -17624
rect -2066 -17681 -1908 -17602
rect -1874 -17681 -1858 -17602
rect -2216 -17687 -1858 -17681
rect -1812 -17675 -1650 -17564
rect -1616 -17675 -1610 -17499
rect -1812 -17687 -1610 -17675
rect -1569 -17499 -1419 -17487
rect -1569 -17675 -1562 -17499
rect -1528 -17524 -1419 -17499
rect -1528 -17656 -1460 -17524
rect -1426 -17656 -1419 -17524
rect -1528 -17675 -1419 -17656
rect -1569 -17687 -1419 -17675
rect -2332 -17734 -1555 -17718
rect -2332 -17768 -2052 -17734
rect -1826 -17768 -1606 -17734
rect -1572 -17768 -1555 -17734
rect -2332 -17780 -1555 -17768
rect -2332 -17841 -2269 -17780
rect -2208 -17787 -1555 -17780
rect -2208 -17841 -2148 -17787
rect -1242 -17815 -1058 -17718
rect 816 -17812 900 -17080
rect 674 -17815 758 -17812
rect -2332 -17884 -2148 -17841
rect -2068 -17899 758 -17815
rect -2608 -18070 -2524 -18064
rect -2216 -17973 -2096 -17913
rect -2216 -18064 -2172 -17973
rect -2138 -18036 -2096 -17973
rect -2068 -17921 -1616 -17899
rect -2068 -17998 -2004 -17921
rect -1970 -17998 -1812 -17921
rect -1778 -17927 -1616 -17921
rect -1778 -17939 -1610 -17927
rect -1778 -17998 -1650 -17939
rect -2068 -18004 -1650 -17998
rect -2138 -18042 -1858 -18036
rect -2138 -18064 -2100 -18042
rect -2216 -18121 -2100 -18064
rect -2066 -18121 -1908 -18042
rect -1874 -18121 -1858 -18042
rect -2216 -18126 -1858 -18121
rect -2332 -18127 -1858 -18126
rect -1812 -18115 -1650 -18004
rect -1616 -18115 -1610 -17939
rect -1812 -18127 -1610 -18115
rect -1569 -17939 -1419 -17927
rect -1569 -18115 -1562 -17939
rect -1528 -17964 -1419 -17939
rect -1528 -18096 -1460 -17964
rect -1426 -18096 -1419 -17964
rect -1528 -18115 -1419 -18096
rect -1569 -18127 -1419 -18115
rect -2332 -18158 -2096 -18127
rect -2332 -18262 -2304 -18158
rect -2200 -18262 -2096 -18158
rect -2332 -18296 -2096 -18262
rect -2216 -18352 -2096 -18296
rect -2216 -18443 -2172 -18352
rect -2138 -18415 -2096 -18352
rect -2068 -18174 -1555 -18158
rect -2068 -18208 -2052 -18174
rect -1826 -18208 -1606 -18174
rect -1572 -18208 -1555 -18174
rect -2068 -18278 -1555 -18208
rect -1516 -18169 -1419 -18127
rect -1516 -18266 -1288 -18169
rect -1191 -18266 -1185 -18169
rect -2068 -18300 -1616 -18278
rect -2068 -18377 -2004 -18300
rect -1970 -18377 -1812 -18300
rect -1778 -18306 -1616 -18300
rect -1516 -18306 -1419 -18266
rect -1778 -18318 -1610 -18306
rect -1778 -18377 -1650 -18318
rect -2068 -18383 -1650 -18377
rect -2138 -18421 -1858 -18415
rect -2138 -18443 -2100 -18421
rect -2216 -18500 -2100 -18443
rect -2066 -18500 -1908 -18421
rect -1874 -18500 -1858 -18421
rect -2216 -18506 -1858 -18500
rect -1812 -18494 -1650 -18383
rect -1616 -18494 -1610 -18318
rect -1812 -18506 -1610 -18494
rect -1569 -18318 -1419 -18306
rect -1569 -18494 -1562 -18318
rect -1528 -18343 -1419 -18318
rect -1528 -18475 -1460 -18343
rect -1426 -18475 -1419 -18343
rect -1528 -18494 -1419 -18475
rect -1569 -18506 -1419 -18494
rect -2332 -18553 -1555 -18537
rect -2332 -18582 -2052 -18553
rect -2332 -18654 -2294 -18582
rect -2222 -18587 -2052 -18582
rect -1826 -18587 -1606 -18553
rect -1572 -18587 -1555 -18553
rect -2222 -18606 -1555 -18587
rect -2222 -18654 -2148 -18606
rect -1242 -18634 -1058 -18537
rect -2332 -18703 -2148 -18654
rect -2068 -18718 574 -18634
rect -2216 -18792 -2096 -18732
rect -2216 -18883 -2172 -18792
rect -2138 -18855 -2096 -18792
rect -2068 -18740 -1616 -18718
rect -2068 -18817 -2004 -18740
rect -1970 -18817 -1812 -18740
rect -1778 -18746 -1616 -18740
rect -1778 -18758 -1610 -18746
rect -1778 -18817 -1650 -18758
rect -2068 -18823 -1650 -18817
rect -2138 -18861 -1858 -18855
rect -2138 -18883 -2100 -18861
rect -2216 -18940 -2100 -18883
rect -2066 -18940 -1908 -18861
rect -1874 -18940 -1858 -18861
rect -2216 -18945 -1858 -18940
rect -2332 -18946 -1858 -18945
rect -1812 -18934 -1650 -18823
rect -1616 -18934 -1610 -18758
rect -1812 -18946 -1610 -18934
rect -1569 -18758 -1419 -18746
rect -1569 -18934 -1562 -18758
rect -1528 -18783 -1419 -18758
rect -1528 -18915 -1460 -18783
rect -1426 -18915 -1419 -18783
rect -1528 -18934 -1419 -18915
rect -1569 -18946 -1419 -18934
rect -2332 -18977 -2096 -18946
rect -2332 -19081 -2304 -18977
rect -2200 -19081 -2096 -18977
rect -2332 -19115 -2096 -19081
rect -2216 -19171 -2096 -19115
rect -2216 -19262 -2172 -19171
rect -2138 -19234 -2096 -19171
rect -2068 -18993 -1555 -18977
rect -2068 -19027 -2052 -18993
rect -1826 -19027 -1606 -18993
rect -1572 -19027 -1555 -18993
rect -2068 -19097 -1555 -19027
rect -1516 -18988 -1419 -18946
rect -1516 -19085 -1288 -18988
rect -1191 -19085 -1185 -18988
rect -2068 -19119 -1616 -19097
rect -2068 -19196 -2004 -19119
rect -1970 -19196 -1812 -19119
rect -1778 -19125 -1616 -19119
rect -1516 -19125 -1419 -19085
rect -1778 -19137 -1610 -19125
rect -1778 -19196 -1650 -19137
rect -2068 -19202 -1650 -19196
rect -2138 -19240 -1858 -19234
rect -2138 -19262 -2100 -19240
rect -2216 -19319 -2100 -19262
rect -2066 -19319 -1908 -19240
rect -1874 -19319 -1858 -19240
rect -2216 -19325 -1858 -19319
rect -1812 -19313 -1650 -19202
rect -1616 -19313 -1610 -19137
rect -1812 -19325 -1610 -19313
rect -1569 -19137 -1419 -19125
rect -1569 -19313 -1562 -19137
rect -1528 -19162 -1419 -19137
rect -1528 -19294 -1460 -19162
rect -1426 -19294 -1419 -19162
rect -1528 -19313 -1419 -19294
rect -1569 -19325 -1419 -19313
rect -2332 -19372 -1555 -19356
rect -2332 -19406 -2052 -19372
rect -1826 -19406 -1606 -19372
rect -1572 -19406 -1555 -19372
rect -2332 -19425 -1555 -19406
rect -2332 -19430 -2148 -19425
rect -2332 -19502 -2300 -19430
rect -2228 -19502 -2148 -19430
rect -1242 -19453 -1058 -19356
rect -2332 -19522 -2148 -19502
rect -2068 -19537 404 -19453
rect -2216 -19611 -2096 -19551
rect -2216 -19702 -2172 -19611
rect -2138 -19674 -2096 -19611
rect -2068 -19559 -1616 -19537
rect -2068 -19636 -2004 -19559
rect -1970 -19636 -1812 -19559
rect -1778 -19565 -1616 -19559
rect -1778 -19577 -1610 -19565
rect -1778 -19636 -1650 -19577
rect -2068 -19642 -1650 -19636
rect -2138 -19680 -1858 -19674
rect -2138 -19702 -2100 -19680
rect -2216 -19759 -2100 -19702
rect -2066 -19759 -1908 -19680
rect -1874 -19759 -1858 -19680
rect -2216 -19764 -1858 -19759
rect -2332 -19765 -1858 -19764
rect -1812 -19753 -1650 -19642
rect -1616 -19753 -1610 -19577
rect -1812 -19765 -1610 -19753
rect -1569 -19577 -1419 -19565
rect -1569 -19753 -1562 -19577
rect -1528 -19602 -1419 -19577
rect -1528 -19734 -1460 -19602
rect -1426 -19734 -1419 -19602
rect -1528 -19753 -1419 -19734
rect -1569 -19765 -1419 -19753
rect -2332 -19796 -2096 -19765
rect -2332 -19900 -2304 -19796
rect -2200 -19900 -2096 -19796
rect -2332 -19934 -2096 -19900
rect -2216 -19990 -2096 -19934
rect -2426 -20128 -2420 -20056
rect -2348 -20128 -2342 -20056
rect -2216 -20081 -2172 -19990
rect -2138 -20053 -2096 -19990
rect -2068 -19812 -1555 -19796
rect -2068 -19846 -2052 -19812
rect -1826 -19846 -1606 -19812
rect -1572 -19846 -1555 -19812
rect -2068 -19916 -1555 -19846
rect -1516 -19807 -1419 -19765
rect -413 -19617 -347 -19611
rect -1516 -19904 -1288 -19807
rect -1191 -19904 -1185 -19807
rect -2068 -19938 -1616 -19916
rect -2068 -20015 -2004 -19938
rect -1970 -20015 -1812 -19938
rect -1778 -19944 -1616 -19938
rect -1516 -19944 -1419 -19904
rect -1778 -19956 -1610 -19944
rect -1778 -20015 -1650 -19956
rect -2068 -20021 -1650 -20015
rect -2138 -20059 -1858 -20053
rect -2138 -20081 -2100 -20059
rect -2420 -20170 -2348 -20128
rect -2216 -20138 -2100 -20081
rect -2066 -20138 -1908 -20059
rect -1874 -20138 -1858 -20059
rect -2216 -20144 -1858 -20138
rect -1812 -20132 -1650 -20021
rect -1616 -20132 -1610 -19956
rect -1812 -20144 -1610 -20132
rect -1569 -19956 -1419 -19944
rect -1569 -20132 -1562 -19956
rect -1528 -19981 -1419 -19956
rect -1528 -20113 -1460 -19981
rect -1426 -20113 -1419 -19981
rect -1528 -20132 -1419 -20113
rect -1569 -20144 -1419 -20132
rect -2420 -20175 -2320 -20170
rect -2420 -20191 -1555 -20175
rect -2420 -20225 -2052 -20191
rect -1826 -20225 -1606 -20191
rect -1572 -20225 -1555 -20191
rect -2420 -20244 -1555 -20225
rect -2420 -20304 -2148 -20244
rect -1242 -20259 -1058 -20175
rect -1243 -20272 -1058 -20259
rect -2332 -20341 -2148 -20304
rect -2068 -20356 -614 -20272
rect -2216 -20411 -2096 -20370
rect -2310 -20417 -2096 -20411
rect -2194 -20430 -2096 -20417
rect -2194 -20521 -2172 -20430
rect -2138 -20493 -2096 -20430
rect -2068 -20378 -1616 -20356
rect -2068 -20455 -2004 -20378
rect -1970 -20455 -1812 -20378
rect -1778 -20384 -1616 -20378
rect -1778 -20396 -1610 -20384
rect -1778 -20455 -1650 -20396
rect -2068 -20461 -1650 -20455
rect -2138 -20499 -1858 -20493
rect -2138 -20521 -2100 -20499
rect -2194 -20533 -2100 -20521
rect -2310 -20539 -2100 -20533
rect -2216 -20578 -2100 -20539
rect -2066 -20578 -1908 -20499
rect -1874 -20578 -1858 -20499
rect -2216 -20584 -1858 -20578
rect -1812 -20572 -1650 -20461
rect -1616 -20572 -1610 -20396
rect -1812 -20584 -1610 -20572
rect -1569 -20396 -1419 -20384
rect -1569 -20572 -1562 -20396
rect -1528 -20421 -1419 -20396
rect -1528 -20553 -1460 -20421
rect -1426 -20440 -1419 -20421
rect -1426 -20537 -1288 -20440
rect -1191 -20537 -1185 -20440
rect -1426 -20553 -1419 -20537
rect -1528 -20572 -1419 -20553
rect -1569 -20584 -1419 -20572
rect -2216 -20615 -2153 -20584
rect -2216 -20631 -1555 -20615
rect -2216 -20665 -2052 -20631
rect -1826 -20665 -1606 -20631
rect -1572 -20665 -1555 -20631
rect -2216 -20684 -1555 -20665
rect -2751 -21825 -2680 -21819
rect -2914 -22616 -2830 -22610
rect -3082 -25964 -2998 -25958
rect -3260 -33362 -3176 -33356
rect -698 -33494 -614 -20356
rect -698 -33584 -614 -33578
rect -11092 -33867 -11081 -33807
rect -11021 -33867 -11001 -33807
rect -413 -33801 -347 -19683
rect 320 -26064 404 -19537
rect 490 -22696 574 -18718
rect 674 -21872 758 -17899
rect 816 -17902 900 -17896
rect 674 -21962 758 -21956
rect 484 -22780 490 -22696
rect 574 -22780 580 -22696
rect 320 -26154 404 -26148
rect 1078 -29278 1137 -16765
rect 1221 -21389 1287 -16623
rect 1367 -20217 1433 -16475
rect 1367 -20289 1433 -20283
rect 3886 -21046 3970 -1635
rect 4164 -1602 4248 -1596
rect 4164 -13666 4248 -1686
rect 4158 -13750 4164 -13666
rect 4248 -13750 4254 -13666
rect 3880 -21130 3886 -21046
rect 3970 -21130 3976 -21046
rect 1215 -21455 1221 -21389
rect 1287 -21455 1293 -21389
rect 4427 -28308 4493 -1375
rect 4573 -28064 4639 -1204
rect 4838 -17961 4904 -1014
rect 4948 -15747 5014 -851
rect 5096 -13052 5162 -684
rect 5261 -6685 5327 -487
rect 5419 -6437 5485 -298
rect 5658 -545 7357 -501
rect 5658 -579 5721 -545
rect 5812 -579 6161 -545
rect 6252 -579 6601 -545
rect 6692 -579 7357 -545
rect 5658 -591 7357 -579
rect 5658 -617 5872 -591
rect 5558 -649 5627 -643
rect 5558 -891 5577 -718
rect 5611 -891 5627 -718
rect 5658 -651 5664 -617
rect 5743 -621 5872 -617
rect 6098 -617 6312 -591
rect 5743 -651 5749 -621
rect 5998 -649 6067 -643
rect 5658 -809 5749 -651
rect 5658 -843 5664 -809
rect 5743 -843 5749 -809
rect 5658 -859 5749 -843
rect 5781 -713 5970 -649
rect 5781 -747 5787 -713
rect 5864 -747 5970 -713
rect 5558 -993 5627 -891
rect 5781 -905 5970 -747
rect 5658 -939 5787 -905
rect 5864 -939 5970 -905
rect 5558 -1111 5628 -993
rect 5658 -1067 5970 -939
rect 5658 -1101 5670 -1067
rect 5846 -1101 5970 -1067
rect 5658 -1107 5858 -1101
rect 5558 -1145 5577 -1111
rect 5611 -1145 5628 -1111
rect 5558 -1162 5628 -1145
rect 5559 -1239 5628 -1162
rect 5558 -1298 5628 -1239
rect 5658 -1155 5858 -1148
rect 5658 -1189 5670 -1155
rect 5846 -1189 5858 -1155
rect 5886 -1162 5970 -1101
rect 5658 -1257 5858 -1189
rect 5658 -1291 5689 -1257
rect 5821 -1291 5858 -1257
rect 5658 -1298 5858 -1291
rect 5901 -1214 5970 -1162
rect 5559 -1414 5628 -1298
rect 5703 -1300 5823 -1298
rect 5703 -1352 5734 -1300
rect 5786 -1352 5823 -1300
rect 5901 -1304 5970 -1283
rect 5998 -891 6017 -718
rect 6051 -891 6067 -718
rect 6098 -651 6104 -617
rect 6183 -621 6312 -617
rect 6538 -604 7357 -591
rect 6538 -617 6752 -604
rect 6183 -651 6189 -621
rect 6438 -649 6507 -643
rect 6098 -809 6189 -651
rect 6098 -843 6104 -809
rect 6183 -843 6189 -809
rect 6098 -859 6189 -843
rect 6221 -713 6410 -649
rect 6221 -747 6227 -713
rect 6304 -747 6410 -713
rect 5998 -1111 6067 -891
rect 6221 -905 6410 -747
rect 6098 -939 6227 -905
rect 6304 -939 6410 -905
rect 6098 -1067 6410 -939
rect 6098 -1101 6110 -1067
rect 6286 -1101 6410 -1067
rect 6098 -1107 6298 -1101
rect 5998 -1145 6017 -1111
rect 6051 -1145 6067 -1111
rect 5703 -1383 5823 -1352
rect 5559 -1483 5901 -1414
rect 5559 -1495 5628 -1483
rect 5832 -4076 5901 -1483
rect 5998 -1747 6067 -1145
rect 6098 -1155 6298 -1148
rect 6098 -1189 6110 -1155
rect 6286 -1189 6298 -1155
rect 6326 -1162 6410 -1101
rect 6098 -1257 6298 -1189
rect 6098 -1291 6129 -1257
rect 6261 -1291 6298 -1257
rect 6098 -1298 6172 -1291
rect 6143 -1333 6172 -1298
rect 6224 -1298 6298 -1291
rect 6341 -1216 6410 -1162
rect 6341 -1298 6410 -1285
rect 6438 -891 6457 -718
rect 6491 -891 6507 -718
rect 6538 -651 6544 -617
rect 6623 -621 6752 -617
rect 6623 -651 6629 -621
rect 6538 -809 6629 -651
rect 6538 -843 6544 -809
rect 6623 -843 6629 -809
rect 6538 -859 6629 -843
rect 6661 -713 6850 -649
rect 6661 -747 6667 -713
rect 6744 -747 6850 -713
rect 6438 -1111 6507 -891
rect 6661 -905 6850 -747
rect 6538 -939 6667 -905
rect 6744 -939 6850 -905
rect 6538 -1067 6850 -939
rect 6538 -1101 6550 -1067
rect 6726 -1101 6850 -1067
rect 6538 -1107 6738 -1101
rect 6438 -1145 6457 -1111
rect 6491 -1145 6507 -1111
rect 6224 -1333 6263 -1298
rect 6143 -1358 6263 -1333
rect 5992 -1753 6073 -1747
rect 5992 -1822 5998 -1753
rect 6067 -1756 6073 -1753
rect 6067 -1822 6085 -1756
rect 5992 -1828 6073 -1822
rect 5998 -3982 6067 -1828
rect 6438 -1888 6507 -1145
rect 6538 -1155 6738 -1148
rect 6538 -1189 6550 -1155
rect 6726 -1189 6738 -1155
rect 6766 -1162 6850 -1101
rect 6538 -1257 6738 -1189
rect 6781 -1207 6850 -1162
rect 7254 -1201 7357 -604
rect 11860 -1201 12409 -1200
rect 12750 -1201 13092 -1200
rect 6538 -1291 6569 -1257
rect 6701 -1291 6738 -1257
rect 6538 -1298 6612 -1291
rect 6580 -1324 6612 -1298
rect 6664 -1298 6738 -1291
rect 6780 -1238 6850 -1207
rect 7137 -1202 7964 -1201
rect 8085 -1202 8912 -1201
rect 9021 -1202 9848 -1201
rect 9952 -1202 10779 -1201
rect 7137 -1217 10780 -1202
rect 6664 -1324 6700 -1298
rect 6580 -1367 6700 -1324
rect 6438 -1963 6507 -1957
rect 6780 -1850 6849 -1238
rect 7137 -1252 7389 -1217
rect 7677 -1252 8337 -1217
rect 8625 -1252 9273 -1217
rect 9561 -1252 10204 -1217
rect 10492 -1252 10780 -1217
rect 7137 -1313 10780 -1252
rect 10879 -1217 13092 -1201
rect 10879 -1252 11131 -1217
rect 11419 -1252 13092 -1217
rect 10879 -1313 13092 -1252
rect 7138 -1324 10780 -1313
rect 7138 -1434 7150 -1324
rect 7184 -1434 7342 -1324
rect 7376 -1434 7534 -1324
rect 7568 -1434 7726 -1324
rect 7760 -1434 7918 -1324
rect 7952 -1434 8098 -1324
rect 8132 -1434 8290 -1324
rect 8324 -1434 8482 -1324
rect 8516 -1434 8674 -1324
rect 8708 -1434 8866 -1324
rect 8900 -1434 9034 -1324
rect 9068 -1434 9226 -1324
rect 9260 -1434 9418 -1324
rect 9452 -1434 9610 -1324
rect 9644 -1434 9802 -1324
rect 9836 -1434 9965 -1324
rect 9999 -1434 10157 -1324
rect 10191 -1434 10349 -1324
rect 10383 -1434 10541 -1324
rect 10575 -1434 10733 -1324
rect 10767 -1434 10780 -1324
rect 7138 -1443 10780 -1434
rect 10880 -1324 13092 -1313
rect 10880 -1434 10892 -1324
rect 10926 -1434 11084 -1324
rect 11118 -1434 11276 -1324
rect 11310 -1434 11468 -1324
rect 11502 -1434 11660 -1324
rect 11694 -1434 13092 -1324
rect 10880 -1443 13092 -1434
rect 7138 -1512 8001 -1497
rect 7138 -1624 7245 -1512
rect 7280 -1624 7438 -1512
rect 7473 -1624 7630 -1512
rect 7665 -1624 7822 -1512
rect 7857 -1624 8001 -1512
rect 7138 -1631 8001 -1624
rect 8086 -1512 8949 -1497
rect 8086 -1624 8193 -1512
rect 8228 -1624 8386 -1512
rect 8421 -1624 8578 -1512
rect 8613 -1624 8770 -1512
rect 8805 -1624 8949 -1512
rect 8086 -1631 8949 -1624
rect 9022 -1512 9885 -1497
rect 9022 -1624 9129 -1512
rect 9164 -1624 9322 -1512
rect 9357 -1624 9514 -1512
rect 9549 -1624 9706 -1512
rect 9741 -1624 9885 -1512
rect 9022 -1631 9885 -1624
rect 9953 -1512 10816 -1497
rect 9953 -1624 10060 -1512
rect 10095 -1624 10253 -1512
rect 10288 -1624 10445 -1512
rect 10480 -1624 10637 -1512
rect 10672 -1624 10816 -1512
rect 9953 -1631 10816 -1624
rect 10880 -1512 11743 -1497
rect 10880 -1624 10987 -1512
rect 11022 -1624 11180 -1512
rect 11215 -1624 11372 -1512
rect 11407 -1624 11564 -1512
rect 11599 -1624 11743 -1512
rect 10880 -1631 11743 -1624
rect 7106 -1662 7158 -1661
rect 7102 -1667 7248 -1662
rect 7102 -1719 7106 -1667
rect 7158 -1678 7248 -1667
rect 7158 -1712 7198 -1678
rect 7232 -1712 7248 -1678
rect 7158 -1719 7248 -1712
rect 7102 -1728 7248 -1719
rect 7304 -1678 7441 -1662
rect 7304 -1712 7390 -1678
rect 7424 -1712 7441 -1678
rect 7304 -1728 7441 -1712
rect 7491 -1678 7632 -1663
rect 7491 -1712 7582 -1678
rect 7616 -1712 7632 -1678
rect 7304 -1756 7370 -1728
rect 7097 -1761 7370 -1756
rect 7097 -1813 7113 -1761
rect 7165 -1813 7370 -1761
rect 7491 -1729 7632 -1712
rect 7661 -1678 7825 -1662
rect 7661 -1712 7774 -1678
rect 7808 -1712 7825 -1678
rect 7661 -1728 7825 -1712
rect 7491 -1765 7557 -1729
rect 7594 -1730 7628 -1729
rect 7097 -1822 7370 -1813
rect 7409 -1850 7557 -1765
rect 6780 -1916 7327 -1850
rect 7393 -1916 7557 -1850
rect 6780 -3879 6849 -1916
rect 7661 -1944 7727 -1728
rect 7102 -2010 7727 -1944
rect 7106 -2211 7172 -2010
rect 7891 -2038 8001 -1631
rect 8050 -1668 8196 -1662
rect 8050 -1720 8069 -1668
rect 8122 -1678 8196 -1668
rect 8122 -1712 8146 -1678
rect 8180 -1712 8196 -1678
rect 8122 -1720 8196 -1712
rect 8050 -1728 8196 -1720
rect 8252 -1678 8389 -1662
rect 8252 -1712 8338 -1678
rect 8372 -1712 8389 -1678
rect 8252 -1728 8389 -1712
rect 8439 -1678 8580 -1663
rect 8439 -1712 8530 -1678
rect 8564 -1712 8580 -1678
rect 8252 -1756 8318 -1728
rect 8050 -1760 8318 -1756
rect 8050 -1812 8057 -1760
rect 8109 -1812 8318 -1760
rect 8439 -1729 8580 -1712
rect 8609 -1678 8773 -1662
rect 8609 -1712 8722 -1678
rect 8756 -1712 8773 -1678
rect 8609 -1728 8773 -1712
rect 8439 -1765 8505 -1729
rect 8542 -1730 8576 -1729
rect 8050 -1822 8318 -1812
rect 8357 -1843 8505 -1765
rect 8357 -1850 8424 -1843
rect 8050 -1895 8424 -1850
rect 8493 -1895 8505 -1843
rect 8050 -1916 8505 -1895
rect 8609 -1944 8675 -1728
rect 7106 -2283 7172 -2277
rect 7214 -2050 7413 -2038
rect 7214 -2062 7372 -2050
rect 7214 -2813 7298 -2062
rect 7333 -2813 7372 -2062
rect 7214 -2991 7227 -2813
rect 7406 -2826 7413 -2050
rect 7405 -2978 7413 -2826
rect 7750 -2050 8001 -2038
rect 7750 -2826 7756 -2050
rect 7790 -2053 8001 -2050
rect 8050 -2010 8675 -1944
rect 7790 -2468 8000 -2053
rect 8050 -2315 8116 -2010
rect 8839 -2038 8949 -1631
rect 8986 -1667 9132 -1662
rect 8986 -1719 9002 -1667
rect 9055 -1678 9132 -1667
rect 9055 -1712 9082 -1678
rect 9116 -1712 9132 -1678
rect 9055 -1719 9132 -1712
rect 8986 -1728 9132 -1719
rect 9188 -1678 9325 -1662
rect 9188 -1712 9274 -1678
rect 9308 -1712 9325 -1678
rect 9188 -1728 9325 -1712
rect 9375 -1678 9516 -1663
rect 9375 -1712 9466 -1678
rect 9500 -1712 9516 -1678
rect 9188 -1756 9254 -1728
rect 8986 -1765 9254 -1756
rect 9375 -1729 9516 -1712
rect 9545 -1678 9709 -1662
rect 9545 -1712 9658 -1678
rect 9692 -1712 9709 -1678
rect 9545 -1728 9709 -1712
rect 9375 -1765 9441 -1729
rect 9478 -1730 9512 -1729
rect 8986 -1817 9000 -1765
rect 9052 -1817 9254 -1765
rect 8986 -1822 9254 -1817
rect 9293 -1850 9441 -1765
rect 8986 -1856 9441 -1850
rect 8986 -1909 8989 -1856
rect 9042 -1909 9441 -1856
rect 8986 -1916 9441 -1909
rect 9545 -1944 9611 -1728
rect 8050 -2387 8116 -2381
rect 8162 -2050 8361 -2038
rect 8162 -2062 8320 -2050
rect 7790 -2534 7872 -2468
rect 7938 -2534 8000 -2468
rect 7790 -2826 8000 -2534
rect 7750 -2838 8000 -2826
rect 8162 -2813 8246 -2062
rect 8281 -2813 8320 -2062
rect 8354 -2826 8361 -2050
rect 7102 -3637 7168 -3631
rect 7102 -3794 7168 -3703
rect 7214 -3742 7298 -2991
rect 7333 -3742 7372 -2991
rect 7214 -3754 7372 -3742
rect 7406 -3754 7413 -2978
rect 7214 -3766 7413 -3754
rect 7750 -2978 8000 -2966
rect 7750 -3754 7756 -2978
rect 7790 -3261 8000 -2978
rect 7790 -3327 7853 -3261
rect 7919 -3327 8000 -3261
rect 7790 -3751 8000 -3327
rect 8340 -2978 8361 -2826
rect 8698 -2050 8949 -2038
rect 8698 -2826 8704 -2050
rect 8738 -2053 8949 -2050
rect 8986 -2009 9611 -1944
rect 8738 -2214 8948 -2053
rect 9052 -2010 9611 -2009
rect 9775 -1966 9885 -1631
rect 10706 -1662 10816 -1631
rect 9917 -1667 10063 -1662
rect 9917 -1719 9933 -1667
rect 9986 -1678 10063 -1667
rect 9986 -1712 10013 -1678
rect 10047 -1712 10063 -1678
rect 9986 -1719 10063 -1712
rect 9917 -1728 10063 -1719
rect 10119 -1678 10256 -1662
rect 10119 -1712 10205 -1678
rect 10239 -1712 10256 -1678
rect 10119 -1728 10256 -1712
rect 10306 -1678 10447 -1663
rect 10306 -1712 10397 -1678
rect 10431 -1712 10447 -1678
rect 10119 -1756 10185 -1728
rect 9917 -1765 10185 -1756
rect 10306 -1729 10447 -1712
rect 10476 -1678 10640 -1662
rect 10476 -1712 10589 -1678
rect 10623 -1712 10640 -1678
rect 10476 -1728 10640 -1712
rect 10706 -1678 10990 -1662
rect 10706 -1712 10940 -1678
rect 10974 -1712 10990 -1678
rect 10706 -1728 10990 -1712
rect 11046 -1678 11183 -1662
rect 11046 -1712 11132 -1678
rect 11166 -1712 11183 -1678
rect 11046 -1728 11183 -1712
rect 11233 -1678 11374 -1663
rect 11233 -1712 11324 -1678
rect 11358 -1712 11374 -1678
rect 10306 -1765 10372 -1729
rect 10409 -1730 10443 -1729
rect 9917 -1817 9935 -1765
rect 9987 -1817 10185 -1765
rect 9917 -1822 10185 -1817
rect 10224 -1812 10372 -1765
rect 10224 -1850 10262 -1812
rect 9917 -1881 10262 -1850
rect 10331 -1881 10372 -1812
rect 9917 -1916 10372 -1881
rect 10476 -1944 10542 -1728
rect 9775 -2032 9798 -1966
rect 9864 -2032 9885 -1966
rect 9775 -2038 9885 -2032
rect 8986 -2093 9052 -2075
rect 9098 -2050 9297 -2038
rect 9098 -2062 9256 -2050
rect 8738 -2280 8818 -2214
rect 8884 -2280 8948 -2214
rect 8738 -2826 8948 -2280
rect 8698 -2838 8948 -2826
rect 9098 -2813 9182 -2062
rect 9217 -2813 9256 -2062
rect 9290 -2826 9297 -2050
rect 8162 -3742 8246 -2991
rect 8281 -3742 8320 -2991
rect 7790 -3754 8001 -3751
rect 7750 -3766 8001 -3754
rect 7102 -3860 7727 -3794
rect 6774 -3948 6780 -3879
rect 6849 -3888 6855 -3879
rect 6849 -3948 7557 -3888
rect 6780 -3954 7557 -3948
rect 5998 -4046 6066 -3982
rect 5999 -4048 6066 -4046
rect 6132 -4048 7370 -3982
rect 7409 -4039 7557 -3954
rect 7304 -4076 7370 -4048
rect 7491 -4075 7557 -4039
rect 7594 -4075 7628 -4074
rect 5832 -4142 6941 -4076
rect 7007 -4092 7248 -4076
rect 7007 -4126 7198 -4092
rect 7232 -4126 7248 -4092
rect 7007 -4142 7248 -4126
rect 7304 -4092 7441 -4076
rect 7304 -4126 7390 -4092
rect 7424 -4126 7441 -4092
rect 7304 -4142 7441 -4126
rect 7491 -4092 7632 -4075
rect 7491 -4126 7582 -4092
rect 7616 -4126 7632 -4092
rect 7491 -4141 7632 -4126
rect 7661 -4076 7727 -3860
rect 7661 -4092 7825 -4076
rect 7661 -4126 7774 -4092
rect 7808 -4126 7825 -4092
rect 7661 -4142 7825 -4126
rect 5832 -4152 5901 -4142
rect 7891 -4173 8001 -3766
rect 8050 -3758 8116 -3752
rect 8162 -3754 8320 -3742
rect 8354 -3754 8361 -2978
rect 8162 -3766 8361 -3754
rect 8698 -2978 8948 -2966
rect 8698 -3754 8704 -2978
rect 8738 -3671 8948 -2978
rect 9276 -2978 9297 -2826
rect 9634 -2050 9885 -2038
rect 9634 -2826 9640 -2050
rect 9674 -2053 9885 -2050
rect 9917 -2010 10542 -1944
rect 9674 -2826 9884 -2053
rect 9917 -2105 9983 -2010
rect 10706 -2038 10816 -1728
rect 11046 -1756 11112 -1728
rect 10844 -1822 10860 -1756
rect 10926 -1822 11112 -1756
rect 11233 -1729 11374 -1712
rect 11403 -1678 11567 -1662
rect 11403 -1712 11516 -1678
rect 11550 -1712 11567 -1678
rect 11403 -1728 11567 -1712
rect 11233 -1765 11299 -1729
rect 11336 -1730 11370 -1729
rect 11151 -1850 11299 -1765
rect 10844 -1916 10858 -1850
rect 10924 -1916 11299 -1850
rect 11403 -1944 11469 -1728
rect 10844 -2010 10850 -1944
rect 10915 -2010 11469 -1944
rect 11633 -2038 11743 -1631
rect 9917 -2177 9983 -2171
rect 10029 -2050 10228 -2038
rect 10029 -2062 10187 -2050
rect 9634 -2838 9884 -2826
rect 10029 -2813 10113 -2062
rect 10148 -2813 10187 -2062
rect 10221 -2826 10228 -2050
rect 8738 -3737 8837 -3671
rect 8903 -3737 8948 -3671
rect 8738 -3751 8948 -3737
rect 8989 -3417 9055 -3411
rect 8738 -3754 8949 -3751
rect 8698 -3766 8949 -3754
rect 8116 -3824 8675 -3794
rect 8050 -3860 8675 -3824
rect 8050 -3895 8505 -3888
rect 8050 -3954 8401 -3895
rect 8357 -3959 8401 -3954
rect 8465 -3959 8505 -3895
rect 8050 -3991 8318 -3982
rect 8050 -4043 8079 -3991
rect 8131 -4043 8318 -3991
rect 8357 -4039 8505 -3959
rect 8050 -4048 8318 -4043
rect 8252 -4076 8318 -4048
rect 8439 -4075 8505 -4039
rect 8542 -4075 8576 -4074
rect 8050 -4085 8196 -4076
rect 8050 -4137 8063 -4085
rect 8128 -4092 8196 -4085
rect 8128 -4126 8146 -4092
rect 8180 -4126 8196 -4092
rect 8128 -4137 8196 -4126
rect 8050 -4142 8196 -4137
rect 8252 -4092 8389 -4076
rect 8252 -4126 8338 -4092
rect 8372 -4126 8389 -4092
rect 8252 -4142 8389 -4126
rect 8439 -4092 8580 -4075
rect 8439 -4126 8530 -4092
rect 8564 -4126 8580 -4092
rect 8439 -4141 8580 -4126
rect 8609 -4076 8675 -3860
rect 8609 -4092 8773 -4076
rect 8609 -4126 8722 -4092
rect 8756 -4126 8773 -4092
rect 8609 -4142 8773 -4126
rect 8839 -4173 8949 -3766
rect 8989 -3794 9055 -3483
rect 9098 -3742 9182 -2991
rect 9217 -3742 9256 -2991
rect 9098 -3754 9256 -3742
rect 9290 -3754 9297 -2978
rect 9098 -3766 9297 -3754
rect 9634 -2978 9884 -2966
rect 9634 -3754 9640 -2978
rect 9674 -3751 9884 -2978
rect 10206 -2977 10228 -2826
rect 10565 -2050 10816 -2038
rect 10565 -2826 10571 -2050
rect 10605 -2053 10816 -2050
rect 10956 -2050 11155 -2038
rect 10605 -2826 10815 -2053
rect 10565 -2838 10815 -2826
rect 10956 -2062 11114 -2050
rect 10956 -2813 11040 -2062
rect 11075 -2813 11114 -2062
rect 11148 -2826 11155 -2050
rect 9917 -3539 9983 -3533
rect 9674 -3754 9885 -3751
rect 9634 -3765 9885 -3754
rect 9634 -3766 9807 -3765
rect 8986 -3860 9611 -3794
rect 8986 -3954 8993 -3888
rect 9059 -3954 9441 -3888
rect 8986 -4048 9001 -3982
rect 9067 -4048 9254 -3982
rect 9293 -4039 9441 -3954
rect 9188 -4076 9254 -4048
rect 9375 -4075 9441 -4039
rect 9478 -4075 9512 -4074
rect 8986 -4085 9132 -4076
rect 8986 -4137 8992 -4085
rect 9057 -4092 9132 -4085
rect 9057 -4126 9082 -4092
rect 9116 -4126 9132 -4092
rect 9057 -4137 9132 -4126
rect 8986 -4142 9132 -4137
rect 9188 -4092 9325 -4076
rect 9188 -4126 9274 -4092
rect 9308 -4126 9325 -4092
rect 9188 -4142 9325 -4126
rect 9375 -4092 9516 -4075
rect 9375 -4126 9466 -4092
rect 9500 -4126 9516 -4092
rect 9375 -4141 9516 -4126
rect 9545 -4076 9611 -3860
rect 9775 -3829 9807 -3766
rect 9873 -3829 9885 -3765
rect 9545 -4092 9709 -4076
rect 9545 -4126 9658 -4092
rect 9692 -4126 9709 -4092
rect 9545 -4142 9709 -4126
rect 9775 -4173 9885 -3829
rect 9917 -3793 9983 -3605
rect 10029 -3741 10113 -2990
rect 10148 -3741 10187 -2990
rect 10029 -3753 10187 -3741
rect 10221 -3753 10228 -2977
rect 10029 -3765 10228 -3753
rect 10565 -2977 10815 -2965
rect 10565 -3753 10571 -2977
rect 10605 -3750 10815 -2977
rect 11134 -2978 11155 -2826
rect 11492 -2050 11743 -2038
rect 11492 -2826 11498 -2050
rect 11532 -2053 11743 -2050
rect 11860 -1667 13092 -1443
rect 11860 -1870 12189 -1667
rect 12410 -1870 13092 -1667
rect 11532 -2809 11742 -2053
rect 11860 -2368 13092 -1870
rect 11799 -2376 13092 -2368
rect 11799 -2427 11811 -2376
rect 12168 -2385 13092 -2376
rect 12168 -2427 12180 -2385
rect 11799 -2434 12180 -2427
rect 11860 -2472 11903 -2434
rect 12726 -2519 13092 -2385
rect 11875 -2531 12689 -2519
rect 12726 -2526 13137 -2519
rect 11875 -2621 11881 -2531
rect 11915 -2621 12073 -2531
rect 12107 -2621 12265 -2531
rect 12299 -2621 12457 -2531
rect 12491 -2621 12649 -2531
rect 12683 -2621 12689 -2531
rect 11875 -2633 12689 -2621
rect 12923 -2563 13137 -2526
rect 12923 -2597 12986 -2563
rect 13077 -2597 13137 -2563
rect 12923 -2635 13137 -2597
rect 11779 -2673 12209 -2661
rect 11779 -2763 11785 -2673
rect 11819 -2763 11977 -2673
rect 12011 -2763 12169 -2673
rect 12203 -2763 12209 -2673
rect 11779 -2775 12209 -2763
rect 12355 -2667 12827 -2661
rect 12355 -2673 12892 -2667
rect 12355 -2763 12361 -2673
rect 12395 -2763 12553 -2673
rect 12587 -2763 12745 -2673
rect 12779 -2683 12892 -2673
rect 12779 -2763 12842 -2683
rect 12355 -2775 12842 -2763
rect 11532 -2825 12263 -2809
rect 11532 -2826 12170 -2825
rect 11492 -2838 12170 -2826
rect 11737 -2859 12170 -2838
rect 12204 -2859 12263 -2825
rect 11737 -2875 12263 -2859
rect 12702 -2909 12842 -2775
rect 12876 -2909 12892 -2683
rect 12923 -2669 12929 -2635
rect 13008 -2639 13137 -2635
rect 13008 -2669 13014 -2639
rect 12923 -2827 13014 -2669
rect 12923 -2861 12929 -2827
rect 13008 -2861 13014 -2827
rect 12923 -2877 13014 -2861
rect 13046 -2731 13235 -2667
rect 13046 -2765 13052 -2731
rect 13129 -2765 13235 -2731
rect 11703 -2930 12363 -2914
rect 11703 -2964 12313 -2930
rect 12347 -2964 12363 -2930
rect 11703 -2966 12363 -2964
rect 10956 -3742 11040 -2991
rect 11075 -3742 11114 -2991
rect 10605 -3753 10816 -3750
rect 10565 -3765 10816 -3753
rect 9917 -3859 10542 -3793
rect 9917 -3895 10372 -3887
rect 9917 -3953 10264 -3895
rect 10224 -3955 10264 -3953
rect 10324 -3955 10372 -3895
rect 9917 -4047 9937 -3981
rect 10003 -4047 10185 -3981
rect 10224 -4038 10372 -3955
rect 10119 -4075 10185 -4047
rect 10306 -4074 10372 -4038
rect 10409 -4074 10443 -4073
rect 9917 -4085 10063 -4075
rect 9917 -4137 9951 -4085
rect 10016 -4091 10063 -4085
rect 10047 -4125 10063 -4091
rect 10016 -4137 10063 -4125
rect 9917 -4141 10063 -4137
rect 10119 -4091 10256 -4075
rect 10119 -4125 10205 -4091
rect 10239 -4125 10256 -4091
rect 10119 -4141 10256 -4125
rect 10306 -4091 10447 -4074
rect 10306 -4125 10397 -4091
rect 10431 -4125 10447 -4091
rect 10306 -4140 10447 -4125
rect 10476 -4075 10542 -3859
rect 10476 -4091 10640 -4075
rect 10476 -4125 10589 -4091
rect 10623 -4125 10640 -4091
rect 10476 -4141 10640 -4125
rect 10706 -4076 10816 -3765
rect 10956 -3754 11114 -3742
rect 11148 -3754 11155 -2978
rect 10956 -3766 11155 -3754
rect 11492 -2978 12363 -2966
rect 11492 -3754 11498 -2978
rect 11532 -2980 12363 -2978
rect 11532 -3011 11815 -2980
rect 11532 -3751 11742 -3011
rect 12259 -3014 12305 -3008
rect 12702 -3014 12892 -2909
rect 13046 -2923 13235 -2765
rect 12259 -3020 12892 -3014
rect 12259 -3196 12265 -3020
rect 12299 -3129 12892 -3020
rect 12923 -2957 13052 -2923
rect 13129 -2934 13235 -2923
rect 13129 -2957 15683 -2934
rect 12923 -3000 15683 -2957
rect 12923 -3085 13235 -3000
rect 12923 -3119 12935 -3085
rect 13111 -3119 13235 -3085
rect 12923 -3125 13123 -3119
rect 12299 -3163 12842 -3129
rect 12876 -3163 12892 -3129
rect 12299 -3180 12892 -3163
rect 12923 -3173 13123 -3166
rect 12299 -3196 12827 -3180
rect 12259 -3208 12827 -3196
rect 12305 -3212 12827 -3208
rect 12923 -3207 12935 -3173
rect 13111 -3207 13123 -3173
rect 13151 -3180 13235 -3119
rect 12305 -3213 12825 -3212
rect 12305 -3214 12774 -3213
rect 12171 -3279 12394 -3272
rect 12171 -3327 12183 -3279
rect 12074 -3340 12183 -3327
rect 12382 -3327 12394 -3279
rect 12923 -3275 13123 -3207
rect 12923 -3309 12954 -3275
rect 13086 -3309 13123 -3275
rect 12921 -3316 13123 -3309
rect 12382 -3340 12473 -3327
rect 12074 -3443 12233 -3340
rect 12352 -3443 12473 -3340
rect 12921 -3365 13121 -3316
rect 12921 -3387 12960 -3365
rect 12074 -3517 12473 -3443
rect 12923 -3484 12960 -3387
rect 13079 -3387 13121 -3365
rect 13079 -3484 13113 -3387
rect 12923 -3542 13113 -3484
rect 11532 -3754 11743 -3751
rect 11492 -3766 11743 -3754
rect 10844 -3860 10850 -3794
rect 10916 -3860 11469 -3794
rect 10844 -3954 10888 -3888
rect 10954 -3954 11299 -3888
rect 10844 -4048 10859 -3982
rect 10925 -4048 11112 -3982
rect 11151 -4039 11299 -3954
rect 11046 -4076 11112 -4048
rect 11233 -4075 11299 -4039
rect 11336 -4075 11370 -4074
rect 10706 -4092 10990 -4076
rect 10706 -4126 10940 -4092
rect 10974 -4126 10990 -4092
rect 10706 -4142 10990 -4126
rect 11046 -4092 11183 -4076
rect 11046 -4126 11132 -4092
rect 11166 -4126 11183 -4092
rect 11046 -4142 11183 -4126
rect 11233 -4092 11374 -4075
rect 11233 -4126 11324 -4092
rect 11358 -4126 11374 -4092
rect 11233 -4141 11374 -4126
rect 11403 -4076 11469 -3860
rect 11403 -4092 11567 -4076
rect 11403 -4126 11516 -4092
rect 11550 -4126 11567 -4092
rect 11403 -4142 11567 -4126
rect 10706 -4172 10816 -4142
rect 7138 -4180 8001 -4173
rect 7138 -4292 7245 -4180
rect 7280 -4292 7438 -4180
rect 7473 -4292 7630 -4180
rect 7665 -4292 7822 -4180
rect 7857 -4292 8001 -4180
rect 7138 -4307 8001 -4292
rect 8086 -4180 8949 -4173
rect 8086 -4292 8193 -4180
rect 8228 -4292 8386 -4180
rect 8421 -4292 8578 -4180
rect 8613 -4292 8770 -4180
rect 8805 -4292 8949 -4180
rect 8086 -4307 8949 -4292
rect 9022 -4180 9885 -4173
rect 9022 -4292 9129 -4180
rect 9164 -4292 9322 -4180
rect 9357 -4292 9514 -4180
rect 9549 -4292 9706 -4180
rect 9741 -4292 9885 -4180
rect 9022 -4307 9885 -4292
rect 9953 -4179 10816 -4172
rect 11633 -4173 11743 -3766
rect 9953 -4291 10060 -4179
rect 10095 -4291 10253 -4179
rect 10288 -4291 10445 -4179
rect 10480 -4291 10637 -4179
rect 10672 -4291 10816 -4179
rect 9953 -4306 10816 -4291
rect 10880 -4180 11743 -4173
rect 10880 -4292 10987 -4180
rect 11022 -4292 11180 -4180
rect 11215 -4292 11372 -4180
rect 11407 -4292 11564 -4180
rect 11599 -4292 11743 -4180
rect 10880 -4307 11743 -4292
rect 7137 -4369 10779 -4360
rect 11883 -4361 12147 -4350
rect 7137 -4370 9965 -4369
rect 7137 -4480 7150 -4370
rect 7184 -4480 7342 -4370
rect 7376 -4480 7534 -4370
rect 7568 -4480 7726 -4370
rect 7760 -4480 7918 -4370
rect 7952 -4480 8098 -4370
rect 8132 -4480 8290 -4370
rect 8324 -4480 8482 -4370
rect 8516 -4480 8674 -4370
rect 8708 -4480 8866 -4370
rect 8900 -4480 9034 -4370
rect 9068 -4480 9226 -4370
rect 9260 -4480 9418 -4370
rect 9452 -4480 9610 -4370
rect 9644 -4480 9802 -4370
rect 9836 -4479 9965 -4370
rect 9999 -4479 10157 -4369
rect 10191 -4479 10349 -4369
rect 10383 -4479 10541 -4369
rect 10575 -4479 10733 -4369
rect 10767 -4479 10779 -4369
rect 9836 -4480 10779 -4479
rect 7137 -4551 10779 -4480
rect 10880 -4370 11894 -4361
rect 10880 -4480 10892 -4370
rect 10926 -4480 11084 -4370
rect 11118 -4480 11276 -4370
rect 11310 -4480 11468 -4370
rect 11502 -4480 11660 -4370
rect 11694 -4480 11894 -4370
rect 10880 -4491 11894 -4480
rect 7137 -4552 10204 -4551
rect 7137 -4587 7389 -4552
rect 7677 -4587 8337 -4552
rect 8625 -4587 9273 -4552
rect 9561 -4586 10204 -4552
rect 10492 -4586 10779 -4551
rect 9561 -4587 10779 -4586
rect 7137 -4601 10779 -4587
rect 7137 -4603 7964 -4601
rect 8085 -4603 8912 -4601
rect 9021 -4603 9848 -4601
rect 9952 -4602 10779 -4601
rect 10879 -4552 11894 -4491
rect 10879 -4587 11131 -4552
rect 11419 -4587 11894 -4552
rect 10879 -4603 11894 -4587
rect 12136 -4603 12147 -4361
rect 11883 -4614 12147 -4603
rect 5658 -4973 7357 -4929
rect 5658 -5007 5721 -4973
rect 5812 -5007 6161 -4973
rect 6252 -5007 6601 -4973
rect 6692 -5007 7357 -4973
rect 5658 -5019 7357 -5007
rect 5658 -5045 5872 -5019
rect 5558 -5077 5627 -5071
rect 5558 -5319 5577 -5146
rect 5611 -5319 5627 -5146
rect 5658 -5079 5664 -5045
rect 5743 -5049 5872 -5045
rect 6098 -5045 6312 -5019
rect 5743 -5079 5749 -5049
rect 5998 -5077 6067 -5071
rect 5658 -5237 5749 -5079
rect 5658 -5271 5664 -5237
rect 5743 -5271 5749 -5237
rect 5658 -5287 5749 -5271
rect 5781 -5141 5970 -5077
rect 5781 -5175 5787 -5141
rect 5864 -5175 5970 -5141
rect 5558 -5421 5627 -5319
rect 5781 -5333 5970 -5175
rect 5658 -5367 5787 -5333
rect 5864 -5367 5970 -5333
rect 5558 -5539 5628 -5421
rect 5658 -5495 5970 -5367
rect 5658 -5529 5670 -5495
rect 5846 -5529 5970 -5495
rect 5658 -5535 5858 -5529
rect 5558 -5573 5577 -5539
rect 5611 -5573 5628 -5539
rect 5558 -5590 5628 -5573
rect 5559 -5667 5628 -5590
rect 5558 -5726 5628 -5667
rect 5658 -5583 5858 -5576
rect 5658 -5617 5670 -5583
rect 5846 -5617 5858 -5583
rect 5886 -5590 5970 -5529
rect 5658 -5685 5858 -5617
rect 5658 -5719 5689 -5685
rect 5821 -5719 5858 -5685
rect 5658 -5726 5858 -5719
rect 5901 -5642 5970 -5590
rect 5559 -5842 5628 -5726
rect 5703 -5728 5823 -5726
rect 5703 -5780 5734 -5728
rect 5786 -5780 5823 -5728
rect 5901 -5732 5970 -5711
rect 5998 -5319 6017 -5146
rect 6051 -5319 6067 -5146
rect 6098 -5079 6104 -5045
rect 6183 -5049 6312 -5045
rect 6538 -5032 7357 -5019
rect 6538 -5045 6752 -5032
rect 6183 -5079 6189 -5049
rect 6438 -5077 6507 -5071
rect 6098 -5237 6189 -5079
rect 6098 -5271 6104 -5237
rect 6183 -5271 6189 -5237
rect 6098 -5287 6189 -5271
rect 6221 -5141 6410 -5077
rect 6221 -5175 6227 -5141
rect 6304 -5175 6410 -5141
rect 5998 -5539 6067 -5319
rect 6221 -5333 6410 -5175
rect 6098 -5367 6227 -5333
rect 6304 -5367 6410 -5333
rect 6098 -5495 6410 -5367
rect 6098 -5529 6110 -5495
rect 6286 -5529 6410 -5495
rect 6098 -5535 6298 -5529
rect 5998 -5573 6017 -5539
rect 6051 -5573 6067 -5539
rect 5703 -5811 5823 -5780
rect 5559 -5911 5901 -5842
rect 5559 -5923 5628 -5911
rect 5413 -6503 5419 -6437
rect 5485 -6503 5491 -6437
rect 5261 -6751 5492 -6685
rect 5426 -11065 5492 -6751
rect 5832 -8504 5901 -5911
rect 5998 -6175 6067 -5573
rect 6098 -5583 6298 -5576
rect 6098 -5617 6110 -5583
rect 6286 -5617 6298 -5583
rect 6326 -5590 6410 -5529
rect 6098 -5685 6298 -5617
rect 6098 -5719 6129 -5685
rect 6261 -5719 6298 -5685
rect 6098 -5726 6172 -5719
rect 6143 -5761 6172 -5726
rect 6224 -5726 6298 -5719
rect 6341 -5644 6410 -5590
rect 6341 -5726 6410 -5713
rect 6438 -5319 6457 -5146
rect 6491 -5319 6507 -5146
rect 6538 -5079 6544 -5045
rect 6623 -5049 6752 -5045
rect 6623 -5079 6629 -5049
rect 6538 -5237 6629 -5079
rect 6538 -5271 6544 -5237
rect 6623 -5271 6629 -5237
rect 6538 -5287 6629 -5271
rect 6661 -5141 6850 -5077
rect 6661 -5175 6667 -5141
rect 6744 -5175 6850 -5141
rect 6438 -5539 6507 -5319
rect 6661 -5333 6850 -5175
rect 6538 -5367 6667 -5333
rect 6744 -5367 6850 -5333
rect 6538 -5495 6850 -5367
rect 6538 -5529 6550 -5495
rect 6726 -5529 6850 -5495
rect 6538 -5535 6738 -5529
rect 6438 -5573 6457 -5539
rect 6491 -5573 6507 -5539
rect 6224 -5761 6263 -5726
rect 6143 -5786 6263 -5761
rect 5992 -6181 6073 -6175
rect 5992 -6250 5998 -6181
rect 6067 -6184 6073 -6181
rect 6067 -6250 6085 -6184
rect 5992 -6256 6073 -6250
rect 5998 -8410 6067 -6256
rect 6438 -6316 6507 -5573
rect 6538 -5583 6738 -5576
rect 6538 -5617 6550 -5583
rect 6726 -5617 6738 -5583
rect 6766 -5590 6850 -5529
rect 6538 -5685 6738 -5617
rect 6781 -5635 6850 -5590
rect 7254 -5629 7357 -5032
rect 11860 -5629 12409 -5628
rect 12750 -5629 13092 -5628
rect 6538 -5719 6569 -5685
rect 6701 -5719 6738 -5685
rect 6538 -5726 6612 -5719
rect 6580 -5752 6612 -5726
rect 6664 -5726 6738 -5719
rect 6780 -5666 6850 -5635
rect 7137 -5630 7964 -5629
rect 8085 -5630 8912 -5629
rect 9021 -5630 9848 -5629
rect 9952 -5630 10779 -5629
rect 7137 -5645 10780 -5630
rect 6664 -5752 6700 -5726
rect 6580 -5795 6700 -5752
rect 6438 -6391 6507 -6385
rect 6780 -6278 6849 -5666
rect 7137 -5680 7389 -5645
rect 7677 -5680 8337 -5645
rect 8625 -5680 9273 -5645
rect 9561 -5680 10204 -5645
rect 10492 -5680 10780 -5645
rect 7137 -5741 10780 -5680
rect 10879 -5645 13092 -5629
rect 10879 -5680 11131 -5645
rect 11419 -5680 13092 -5645
rect 10879 -5741 13092 -5680
rect 7138 -5752 10780 -5741
rect 7138 -5862 7150 -5752
rect 7184 -5862 7342 -5752
rect 7376 -5862 7534 -5752
rect 7568 -5862 7726 -5752
rect 7760 -5862 7918 -5752
rect 7952 -5862 8098 -5752
rect 8132 -5862 8290 -5752
rect 8324 -5862 8482 -5752
rect 8516 -5862 8674 -5752
rect 8708 -5862 8866 -5752
rect 8900 -5862 9034 -5752
rect 9068 -5862 9226 -5752
rect 9260 -5862 9418 -5752
rect 9452 -5862 9610 -5752
rect 9644 -5862 9802 -5752
rect 9836 -5862 9965 -5752
rect 9999 -5862 10157 -5752
rect 10191 -5862 10349 -5752
rect 10383 -5862 10541 -5752
rect 10575 -5862 10733 -5752
rect 10767 -5862 10780 -5752
rect 7138 -5871 10780 -5862
rect 10880 -5752 13092 -5741
rect 10880 -5862 10892 -5752
rect 10926 -5862 11084 -5752
rect 11118 -5862 11276 -5752
rect 11310 -5862 11468 -5752
rect 11502 -5862 11660 -5752
rect 11694 -5862 13092 -5752
rect 10880 -5871 13092 -5862
rect 7138 -5940 8001 -5925
rect 7138 -6052 7245 -5940
rect 7280 -6052 7438 -5940
rect 7473 -6052 7630 -5940
rect 7665 -6052 7822 -5940
rect 7857 -6052 8001 -5940
rect 7138 -6059 8001 -6052
rect 8086 -5940 8949 -5925
rect 8086 -6052 8193 -5940
rect 8228 -6052 8386 -5940
rect 8421 -6052 8578 -5940
rect 8613 -6052 8770 -5940
rect 8805 -6052 8949 -5940
rect 8086 -6059 8949 -6052
rect 9022 -5940 9885 -5925
rect 9022 -6052 9129 -5940
rect 9164 -6052 9322 -5940
rect 9357 -6052 9514 -5940
rect 9549 -6052 9706 -5940
rect 9741 -6052 9885 -5940
rect 9022 -6059 9885 -6052
rect 9953 -5940 10816 -5925
rect 9953 -6052 10060 -5940
rect 10095 -6052 10253 -5940
rect 10288 -6052 10445 -5940
rect 10480 -6052 10637 -5940
rect 10672 -6052 10816 -5940
rect 9953 -6059 10816 -6052
rect 10880 -5940 11743 -5925
rect 10880 -6052 10987 -5940
rect 11022 -6052 11180 -5940
rect 11215 -6052 11372 -5940
rect 11407 -6052 11564 -5940
rect 11599 -6052 11743 -5940
rect 10880 -6059 11743 -6052
rect 7106 -6090 7158 -6089
rect 7102 -6095 7248 -6090
rect 7102 -6147 7106 -6095
rect 7158 -6106 7248 -6095
rect 7158 -6140 7198 -6106
rect 7232 -6140 7248 -6106
rect 7158 -6147 7248 -6140
rect 7102 -6156 7248 -6147
rect 7304 -6106 7441 -6090
rect 7304 -6140 7390 -6106
rect 7424 -6140 7441 -6106
rect 7304 -6156 7441 -6140
rect 7491 -6106 7632 -6091
rect 7491 -6140 7582 -6106
rect 7616 -6140 7632 -6106
rect 7304 -6184 7370 -6156
rect 7097 -6189 7370 -6184
rect 7097 -6241 7113 -6189
rect 7165 -6241 7370 -6189
rect 7491 -6157 7632 -6140
rect 7661 -6106 7825 -6090
rect 7661 -6140 7774 -6106
rect 7808 -6140 7825 -6106
rect 7661 -6156 7825 -6140
rect 7491 -6193 7557 -6157
rect 7594 -6158 7628 -6157
rect 7097 -6250 7370 -6241
rect 7409 -6278 7557 -6193
rect 6780 -6344 7327 -6278
rect 7393 -6344 7557 -6278
rect 6780 -8307 6849 -6344
rect 7661 -6372 7727 -6156
rect 7102 -6438 7727 -6372
rect 7106 -6639 7172 -6438
rect 7891 -6466 8001 -6059
rect 8050 -6096 8196 -6090
rect 8050 -6148 8069 -6096
rect 8122 -6106 8196 -6096
rect 8122 -6140 8146 -6106
rect 8180 -6140 8196 -6106
rect 8122 -6148 8196 -6140
rect 8050 -6156 8196 -6148
rect 8252 -6106 8389 -6090
rect 8252 -6140 8338 -6106
rect 8372 -6140 8389 -6106
rect 8252 -6156 8389 -6140
rect 8439 -6106 8580 -6091
rect 8439 -6140 8530 -6106
rect 8564 -6140 8580 -6106
rect 8252 -6184 8318 -6156
rect 8050 -6188 8318 -6184
rect 8050 -6240 8057 -6188
rect 8109 -6240 8318 -6188
rect 8439 -6157 8580 -6140
rect 8609 -6106 8773 -6090
rect 8609 -6140 8722 -6106
rect 8756 -6140 8773 -6106
rect 8609 -6156 8773 -6140
rect 8439 -6193 8505 -6157
rect 8542 -6158 8576 -6157
rect 8050 -6250 8318 -6240
rect 8357 -6271 8505 -6193
rect 8357 -6278 8424 -6271
rect 8050 -6323 8424 -6278
rect 8493 -6323 8505 -6271
rect 8050 -6344 8505 -6323
rect 8609 -6372 8675 -6156
rect 7106 -6711 7172 -6705
rect 7214 -6478 7413 -6466
rect 7214 -6490 7372 -6478
rect 7214 -7241 7298 -6490
rect 7333 -7241 7372 -6490
rect 7214 -7419 7227 -7241
rect 7406 -7254 7413 -6478
rect 7405 -7406 7413 -7254
rect 7750 -6478 8001 -6466
rect 7750 -7254 7756 -6478
rect 7790 -6481 8001 -6478
rect 8050 -6438 8675 -6372
rect 7790 -6896 8000 -6481
rect 8050 -6743 8116 -6438
rect 8839 -6466 8949 -6059
rect 8986 -6095 9132 -6090
rect 8986 -6147 9002 -6095
rect 9055 -6106 9132 -6095
rect 9055 -6140 9082 -6106
rect 9116 -6140 9132 -6106
rect 9055 -6147 9132 -6140
rect 8986 -6156 9132 -6147
rect 9188 -6106 9325 -6090
rect 9188 -6140 9274 -6106
rect 9308 -6140 9325 -6106
rect 9188 -6156 9325 -6140
rect 9375 -6106 9516 -6091
rect 9375 -6140 9466 -6106
rect 9500 -6140 9516 -6106
rect 9188 -6184 9254 -6156
rect 8986 -6193 9254 -6184
rect 9375 -6157 9516 -6140
rect 9545 -6106 9709 -6090
rect 9545 -6140 9658 -6106
rect 9692 -6140 9709 -6106
rect 9545 -6156 9709 -6140
rect 9375 -6193 9441 -6157
rect 9478 -6158 9512 -6157
rect 8986 -6245 9000 -6193
rect 9052 -6245 9254 -6193
rect 8986 -6250 9254 -6245
rect 9293 -6278 9441 -6193
rect 8986 -6284 9441 -6278
rect 8986 -6337 8989 -6284
rect 9042 -6337 9441 -6284
rect 8986 -6344 9441 -6337
rect 9545 -6372 9611 -6156
rect 8050 -6815 8116 -6809
rect 8162 -6478 8361 -6466
rect 8162 -6490 8320 -6478
rect 7790 -6962 7872 -6896
rect 7938 -6962 8000 -6896
rect 7790 -7254 8000 -6962
rect 7750 -7266 8000 -7254
rect 8162 -7241 8246 -6490
rect 8281 -7241 8320 -6490
rect 8354 -7254 8361 -6478
rect 7102 -8065 7168 -8059
rect 7102 -8222 7168 -8131
rect 7214 -8170 7298 -7419
rect 7333 -8170 7372 -7419
rect 7214 -8182 7372 -8170
rect 7406 -8182 7413 -7406
rect 7214 -8194 7413 -8182
rect 7750 -7406 8000 -7394
rect 7750 -8182 7756 -7406
rect 7790 -7689 8000 -7406
rect 7790 -7755 7853 -7689
rect 7919 -7755 8000 -7689
rect 7790 -8179 8000 -7755
rect 8340 -7406 8361 -7254
rect 8698 -6478 8949 -6466
rect 8698 -7254 8704 -6478
rect 8738 -6481 8949 -6478
rect 8986 -6437 9611 -6372
rect 8738 -6642 8948 -6481
rect 9052 -6438 9611 -6437
rect 9775 -6394 9885 -6059
rect 10706 -6090 10816 -6059
rect 9917 -6095 10063 -6090
rect 9917 -6147 9933 -6095
rect 9986 -6106 10063 -6095
rect 9986 -6140 10013 -6106
rect 10047 -6140 10063 -6106
rect 9986 -6147 10063 -6140
rect 9917 -6156 10063 -6147
rect 10119 -6106 10256 -6090
rect 10119 -6140 10205 -6106
rect 10239 -6140 10256 -6106
rect 10119 -6156 10256 -6140
rect 10306 -6106 10447 -6091
rect 10306 -6140 10397 -6106
rect 10431 -6140 10447 -6106
rect 10119 -6184 10185 -6156
rect 9917 -6193 10185 -6184
rect 10306 -6157 10447 -6140
rect 10476 -6106 10640 -6090
rect 10476 -6140 10589 -6106
rect 10623 -6140 10640 -6106
rect 10476 -6156 10640 -6140
rect 10706 -6106 10990 -6090
rect 10706 -6140 10940 -6106
rect 10974 -6140 10990 -6106
rect 10706 -6156 10990 -6140
rect 11046 -6106 11183 -6090
rect 11046 -6140 11132 -6106
rect 11166 -6140 11183 -6106
rect 11046 -6156 11183 -6140
rect 11233 -6106 11374 -6091
rect 11233 -6140 11324 -6106
rect 11358 -6140 11374 -6106
rect 10306 -6193 10372 -6157
rect 10409 -6158 10443 -6157
rect 9917 -6245 9935 -6193
rect 9987 -6245 10185 -6193
rect 9917 -6250 10185 -6245
rect 10224 -6240 10372 -6193
rect 10224 -6278 10262 -6240
rect 9917 -6309 10262 -6278
rect 10331 -6309 10372 -6240
rect 9917 -6344 10372 -6309
rect 10476 -6372 10542 -6156
rect 9775 -6460 9798 -6394
rect 9864 -6460 9885 -6394
rect 9775 -6466 9885 -6460
rect 8986 -6521 9052 -6503
rect 9098 -6478 9297 -6466
rect 9098 -6490 9256 -6478
rect 8738 -6708 8818 -6642
rect 8884 -6708 8948 -6642
rect 8738 -7254 8948 -6708
rect 8698 -7266 8948 -7254
rect 9098 -7241 9182 -6490
rect 9217 -7241 9256 -6490
rect 9290 -7254 9297 -6478
rect 8162 -8170 8246 -7419
rect 8281 -8170 8320 -7419
rect 7790 -8182 8001 -8179
rect 7750 -8194 8001 -8182
rect 7102 -8288 7727 -8222
rect 6774 -8376 6780 -8307
rect 6849 -8316 6855 -8307
rect 6849 -8376 7557 -8316
rect 6780 -8382 7557 -8376
rect 5998 -8474 6066 -8410
rect 5999 -8476 6066 -8474
rect 6132 -8476 7370 -8410
rect 7409 -8467 7557 -8382
rect 7304 -8504 7370 -8476
rect 7491 -8503 7557 -8467
rect 7594 -8503 7628 -8502
rect 5832 -8570 6941 -8504
rect 7007 -8520 7248 -8504
rect 7007 -8554 7198 -8520
rect 7232 -8554 7248 -8520
rect 7007 -8570 7248 -8554
rect 7304 -8520 7441 -8504
rect 7304 -8554 7390 -8520
rect 7424 -8554 7441 -8520
rect 7304 -8570 7441 -8554
rect 7491 -8520 7632 -8503
rect 7491 -8554 7582 -8520
rect 7616 -8554 7632 -8520
rect 7491 -8569 7632 -8554
rect 7661 -8504 7727 -8288
rect 7661 -8520 7825 -8504
rect 7661 -8554 7774 -8520
rect 7808 -8554 7825 -8520
rect 7661 -8570 7825 -8554
rect 5832 -8580 5901 -8570
rect 7891 -8601 8001 -8194
rect 8050 -8186 8116 -8180
rect 8162 -8182 8320 -8170
rect 8354 -8182 8361 -7406
rect 8162 -8194 8361 -8182
rect 8698 -7406 8948 -7394
rect 8698 -8182 8704 -7406
rect 8738 -8099 8948 -7406
rect 9276 -7406 9297 -7254
rect 9634 -6478 9885 -6466
rect 9634 -7254 9640 -6478
rect 9674 -6481 9885 -6478
rect 9917 -6438 10542 -6372
rect 9674 -7254 9884 -6481
rect 9917 -6533 9983 -6438
rect 10706 -6466 10816 -6156
rect 11046 -6184 11112 -6156
rect 10844 -6250 10860 -6184
rect 10926 -6250 11112 -6184
rect 11233 -6157 11374 -6140
rect 11403 -6106 11567 -6090
rect 11403 -6140 11516 -6106
rect 11550 -6140 11567 -6106
rect 11403 -6156 11567 -6140
rect 11233 -6193 11299 -6157
rect 11336 -6158 11370 -6157
rect 11151 -6278 11299 -6193
rect 10844 -6344 10858 -6278
rect 10924 -6344 11299 -6278
rect 11403 -6372 11469 -6156
rect 10844 -6438 10850 -6372
rect 10915 -6438 11469 -6372
rect 11633 -6466 11743 -6059
rect 9917 -6605 9983 -6599
rect 10029 -6478 10228 -6466
rect 10029 -6490 10187 -6478
rect 9634 -7266 9884 -7254
rect 10029 -7241 10113 -6490
rect 10148 -7241 10187 -6490
rect 10221 -7254 10228 -6478
rect 8738 -8165 8837 -8099
rect 8903 -8165 8948 -8099
rect 8738 -8179 8948 -8165
rect 8989 -7845 9055 -7839
rect 8738 -8182 8949 -8179
rect 8698 -8194 8949 -8182
rect 8116 -8252 8675 -8222
rect 8050 -8288 8675 -8252
rect 8050 -8323 8505 -8316
rect 8050 -8382 8401 -8323
rect 8357 -8387 8401 -8382
rect 8465 -8387 8505 -8323
rect 8050 -8419 8318 -8410
rect 8050 -8471 8079 -8419
rect 8131 -8471 8318 -8419
rect 8357 -8467 8505 -8387
rect 8050 -8476 8318 -8471
rect 8252 -8504 8318 -8476
rect 8439 -8503 8505 -8467
rect 8542 -8503 8576 -8502
rect 8050 -8513 8196 -8504
rect 8050 -8565 8063 -8513
rect 8128 -8520 8196 -8513
rect 8128 -8554 8146 -8520
rect 8180 -8554 8196 -8520
rect 8128 -8565 8196 -8554
rect 8050 -8570 8196 -8565
rect 8252 -8520 8389 -8504
rect 8252 -8554 8338 -8520
rect 8372 -8554 8389 -8520
rect 8252 -8570 8389 -8554
rect 8439 -8520 8580 -8503
rect 8439 -8554 8530 -8520
rect 8564 -8554 8580 -8520
rect 8439 -8569 8580 -8554
rect 8609 -8504 8675 -8288
rect 8609 -8520 8773 -8504
rect 8609 -8554 8722 -8520
rect 8756 -8554 8773 -8520
rect 8609 -8570 8773 -8554
rect 8839 -8601 8949 -8194
rect 8989 -8222 9055 -7911
rect 9098 -8170 9182 -7419
rect 9217 -8170 9256 -7419
rect 9098 -8182 9256 -8170
rect 9290 -8182 9297 -7406
rect 9098 -8194 9297 -8182
rect 9634 -7406 9884 -7394
rect 9634 -8182 9640 -7406
rect 9674 -8179 9884 -7406
rect 10206 -7405 10228 -7254
rect 10565 -6478 10816 -6466
rect 10565 -7254 10571 -6478
rect 10605 -6481 10816 -6478
rect 10956 -6478 11155 -6466
rect 10605 -7254 10815 -6481
rect 10565 -7266 10815 -7254
rect 10956 -6490 11114 -6478
rect 10956 -7241 11040 -6490
rect 11075 -7241 11114 -6490
rect 11148 -7254 11155 -6478
rect 9917 -7967 9983 -7961
rect 9674 -8182 9885 -8179
rect 9634 -8193 9885 -8182
rect 9634 -8194 9807 -8193
rect 8986 -8288 9611 -8222
rect 8986 -8382 8993 -8316
rect 9059 -8382 9441 -8316
rect 8986 -8476 9001 -8410
rect 9067 -8476 9254 -8410
rect 9293 -8467 9441 -8382
rect 9188 -8504 9254 -8476
rect 9375 -8503 9441 -8467
rect 9478 -8503 9512 -8502
rect 8986 -8513 9132 -8504
rect 8986 -8565 8992 -8513
rect 9057 -8520 9132 -8513
rect 9057 -8554 9082 -8520
rect 9116 -8554 9132 -8520
rect 9057 -8565 9132 -8554
rect 8986 -8570 9132 -8565
rect 9188 -8520 9325 -8504
rect 9188 -8554 9274 -8520
rect 9308 -8554 9325 -8520
rect 9188 -8570 9325 -8554
rect 9375 -8520 9516 -8503
rect 9375 -8554 9466 -8520
rect 9500 -8554 9516 -8520
rect 9375 -8569 9516 -8554
rect 9545 -8504 9611 -8288
rect 9775 -8257 9807 -8194
rect 9873 -8257 9885 -8193
rect 9545 -8520 9709 -8504
rect 9545 -8554 9658 -8520
rect 9692 -8554 9709 -8520
rect 9545 -8570 9709 -8554
rect 9775 -8601 9885 -8257
rect 9917 -8221 9983 -8033
rect 10029 -8169 10113 -7418
rect 10148 -8169 10187 -7418
rect 10029 -8181 10187 -8169
rect 10221 -8181 10228 -7405
rect 10029 -8193 10228 -8181
rect 10565 -7405 10815 -7393
rect 10565 -8181 10571 -7405
rect 10605 -8178 10815 -7405
rect 11134 -7406 11155 -7254
rect 11492 -6478 11743 -6466
rect 11492 -7254 11498 -6478
rect 11532 -6481 11743 -6478
rect 11860 -6095 13092 -5871
rect 11860 -6298 12189 -6095
rect 12410 -6298 13092 -6095
rect 11532 -7237 11742 -6481
rect 11860 -6796 13092 -6298
rect 11799 -6804 13092 -6796
rect 11799 -6855 11811 -6804
rect 12168 -6813 13092 -6804
rect 12168 -6855 12180 -6813
rect 11799 -6862 12180 -6855
rect 11860 -6900 11903 -6862
rect 12726 -6947 13092 -6813
rect 11875 -6959 12689 -6947
rect 12726 -6954 13137 -6947
rect 11875 -7049 11881 -6959
rect 11915 -7049 12073 -6959
rect 12107 -7049 12265 -6959
rect 12299 -7049 12457 -6959
rect 12491 -7049 12649 -6959
rect 12683 -7049 12689 -6959
rect 11875 -7061 12689 -7049
rect 12923 -6991 13137 -6954
rect 12923 -7025 12986 -6991
rect 13077 -7025 13137 -6991
rect 12923 -7063 13137 -7025
rect 11779 -7101 12209 -7089
rect 11779 -7191 11785 -7101
rect 11819 -7191 11977 -7101
rect 12011 -7191 12169 -7101
rect 12203 -7191 12209 -7101
rect 11779 -7203 12209 -7191
rect 12355 -7095 12827 -7089
rect 12355 -7101 12892 -7095
rect 12355 -7191 12361 -7101
rect 12395 -7191 12553 -7101
rect 12587 -7191 12745 -7101
rect 12779 -7111 12892 -7101
rect 12779 -7191 12842 -7111
rect 12355 -7203 12842 -7191
rect 11532 -7253 12263 -7237
rect 11532 -7254 12170 -7253
rect 11492 -7266 12170 -7254
rect 11737 -7287 12170 -7266
rect 12204 -7287 12263 -7253
rect 11737 -7303 12263 -7287
rect 12702 -7337 12842 -7203
rect 12876 -7337 12892 -7111
rect 12923 -7097 12929 -7063
rect 13008 -7067 13137 -7063
rect 13008 -7097 13014 -7067
rect 12923 -7255 13014 -7097
rect 12923 -7289 12929 -7255
rect 13008 -7289 13014 -7255
rect 12923 -7305 13014 -7289
rect 13046 -7159 13235 -7095
rect 13046 -7193 13052 -7159
rect 13129 -7193 13235 -7159
rect 11703 -7358 12363 -7342
rect 11703 -7392 12313 -7358
rect 12347 -7392 12363 -7358
rect 11703 -7394 12363 -7392
rect 10956 -8170 11040 -7419
rect 11075 -8170 11114 -7419
rect 10605 -8181 10816 -8178
rect 10565 -8193 10816 -8181
rect 9917 -8287 10542 -8221
rect 9917 -8323 10372 -8315
rect 9917 -8381 10264 -8323
rect 10224 -8383 10264 -8381
rect 10324 -8383 10372 -8323
rect 9917 -8475 9937 -8409
rect 10003 -8475 10185 -8409
rect 10224 -8466 10372 -8383
rect 10119 -8503 10185 -8475
rect 10306 -8502 10372 -8466
rect 10409 -8502 10443 -8501
rect 9917 -8513 10063 -8503
rect 9917 -8565 9951 -8513
rect 10016 -8519 10063 -8513
rect 10047 -8553 10063 -8519
rect 10016 -8565 10063 -8553
rect 9917 -8569 10063 -8565
rect 10119 -8519 10256 -8503
rect 10119 -8553 10205 -8519
rect 10239 -8553 10256 -8519
rect 10119 -8569 10256 -8553
rect 10306 -8519 10447 -8502
rect 10306 -8553 10397 -8519
rect 10431 -8553 10447 -8519
rect 10306 -8568 10447 -8553
rect 10476 -8503 10542 -8287
rect 10476 -8519 10640 -8503
rect 10476 -8553 10589 -8519
rect 10623 -8553 10640 -8519
rect 10476 -8569 10640 -8553
rect 10706 -8504 10816 -8193
rect 10956 -8182 11114 -8170
rect 11148 -8182 11155 -7406
rect 10956 -8194 11155 -8182
rect 11492 -7406 12363 -7394
rect 11492 -8182 11498 -7406
rect 11532 -7408 12363 -7406
rect 11532 -7439 11815 -7408
rect 11532 -8179 11742 -7439
rect 12259 -7442 12305 -7436
rect 12702 -7442 12892 -7337
rect 13046 -7351 13235 -7193
rect 12259 -7448 12892 -7442
rect 12259 -7624 12265 -7448
rect 12299 -7557 12892 -7448
rect 12923 -7385 13052 -7351
rect 13129 -7385 13235 -7351
rect 12923 -7415 13235 -7385
rect 12923 -7481 15547 -7415
rect 12923 -7513 13235 -7481
rect 12923 -7547 12935 -7513
rect 13111 -7547 13235 -7513
rect 12923 -7553 13123 -7547
rect 12299 -7591 12842 -7557
rect 12876 -7591 12892 -7557
rect 12299 -7608 12892 -7591
rect 12923 -7601 13123 -7594
rect 12299 -7624 12827 -7608
rect 12259 -7636 12827 -7624
rect 12305 -7640 12827 -7636
rect 12923 -7635 12935 -7601
rect 13111 -7635 13123 -7601
rect 13151 -7608 13235 -7547
rect 12305 -7641 12825 -7640
rect 12305 -7642 12774 -7641
rect 12171 -7707 12394 -7700
rect 12171 -7755 12183 -7707
rect 12074 -7768 12183 -7755
rect 12382 -7755 12394 -7707
rect 12923 -7703 13123 -7635
rect 12923 -7737 12954 -7703
rect 13086 -7737 13123 -7703
rect 12921 -7744 13123 -7737
rect 12382 -7768 12473 -7755
rect 12074 -7871 12233 -7768
rect 12352 -7871 12473 -7768
rect 12921 -7793 13121 -7744
rect 12921 -7815 12960 -7793
rect 12074 -7945 12473 -7871
rect 12923 -7912 12960 -7815
rect 13079 -7815 13121 -7793
rect 13079 -7912 13113 -7815
rect 12923 -7970 13113 -7912
rect 11532 -8182 11743 -8179
rect 11492 -8194 11743 -8182
rect 10844 -8288 10850 -8222
rect 10916 -8288 11469 -8222
rect 10844 -8382 10888 -8316
rect 10954 -8382 11299 -8316
rect 10844 -8476 10859 -8410
rect 10925 -8476 11112 -8410
rect 11151 -8467 11299 -8382
rect 11046 -8504 11112 -8476
rect 11233 -8503 11299 -8467
rect 11336 -8503 11370 -8502
rect 10706 -8520 10990 -8504
rect 10706 -8554 10940 -8520
rect 10974 -8554 10990 -8520
rect 10706 -8570 10990 -8554
rect 11046 -8520 11183 -8504
rect 11046 -8554 11132 -8520
rect 11166 -8554 11183 -8520
rect 11046 -8570 11183 -8554
rect 11233 -8520 11374 -8503
rect 11233 -8554 11324 -8520
rect 11358 -8554 11374 -8520
rect 11233 -8569 11374 -8554
rect 11403 -8504 11469 -8288
rect 11403 -8520 11567 -8504
rect 11403 -8554 11516 -8520
rect 11550 -8554 11567 -8520
rect 11403 -8570 11567 -8554
rect 10706 -8600 10816 -8570
rect 7138 -8608 8001 -8601
rect 7138 -8720 7245 -8608
rect 7280 -8720 7438 -8608
rect 7473 -8720 7630 -8608
rect 7665 -8720 7822 -8608
rect 7857 -8720 8001 -8608
rect 7138 -8735 8001 -8720
rect 8086 -8608 8949 -8601
rect 8086 -8720 8193 -8608
rect 8228 -8720 8386 -8608
rect 8421 -8720 8578 -8608
rect 8613 -8720 8770 -8608
rect 8805 -8720 8949 -8608
rect 8086 -8735 8949 -8720
rect 9022 -8608 9885 -8601
rect 9022 -8720 9129 -8608
rect 9164 -8720 9322 -8608
rect 9357 -8720 9514 -8608
rect 9549 -8720 9706 -8608
rect 9741 -8720 9885 -8608
rect 9022 -8735 9885 -8720
rect 9953 -8607 10816 -8600
rect 11633 -8601 11743 -8194
rect 9953 -8719 10060 -8607
rect 10095 -8719 10253 -8607
rect 10288 -8719 10445 -8607
rect 10480 -8719 10637 -8607
rect 10672 -8719 10816 -8607
rect 9953 -8734 10816 -8719
rect 10880 -8608 11743 -8601
rect 10880 -8720 10987 -8608
rect 11022 -8720 11180 -8608
rect 11215 -8720 11372 -8608
rect 11407 -8720 11564 -8608
rect 11599 -8720 11743 -8608
rect 10880 -8735 11743 -8720
rect 7137 -8797 10779 -8788
rect 11883 -8789 12147 -8778
rect 7137 -8798 9965 -8797
rect 7137 -8908 7150 -8798
rect 7184 -8908 7342 -8798
rect 7376 -8908 7534 -8798
rect 7568 -8908 7726 -8798
rect 7760 -8908 7918 -8798
rect 7952 -8908 8098 -8798
rect 8132 -8908 8290 -8798
rect 8324 -8908 8482 -8798
rect 8516 -8908 8674 -8798
rect 8708 -8908 8866 -8798
rect 8900 -8908 9034 -8798
rect 9068 -8908 9226 -8798
rect 9260 -8908 9418 -8798
rect 9452 -8908 9610 -8798
rect 9644 -8908 9802 -8798
rect 9836 -8907 9965 -8798
rect 9999 -8907 10157 -8797
rect 10191 -8907 10349 -8797
rect 10383 -8907 10541 -8797
rect 10575 -8907 10733 -8797
rect 10767 -8907 10779 -8797
rect 9836 -8908 10779 -8907
rect 7137 -8979 10779 -8908
rect 10880 -8798 11894 -8789
rect 10880 -8908 10892 -8798
rect 10926 -8908 11084 -8798
rect 11118 -8908 11276 -8798
rect 11310 -8908 11468 -8798
rect 11502 -8908 11660 -8798
rect 11694 -8908 11894 -8798
rect 10880 -8919 11894 -8908
rect 7137 -8980 10204 -8979
rect 7137 -9015 7389 -8980
rect 7677 -9015 8337 -8980
rect 8625 -9015 9273 -8980
rect 9561 -9014 10204 -8980
rect 10492 -9014 10779 -8979
rect 9561 -9015 10779 -9014
rect 7137 -9029 10779 -9015
rect 7137 -9031 7964 -9029
rect 8085 -9031 8912 -9029
rect 9021 -9031 9848 -9029
rect 9952 -9030 10779 -9029
rect 10879 -8980 11894 -8919
rect 10879 -9015 11131 -8980
rect 11419 -9015 11894 -8980
rect 10879 -9031 11894 -9015
rect 12136 -9031 12147 -8789
rect 11883 -9042 12147 -9031
rect 5658 -9601 7357 -9557
rect 5658 -9635 5721 -9601
rect 5812 -9635 6161 -9601
rect 6252 -9635 6601 -9601
rect 6692 -9635 7357 -9601
rect 5658 -9647 7357 -9635
rect 5658 -9673 5872 -9647
rect 5558 -9705 5627 -9699
rect 5558 -9947 5577 -9774
rect 5611 -9947 5627 -9774
rect 5658 -9707 5664 -9673
rect 5743 -9677 5872 -9673
rect 6098 -9673 6312 -9647
rect 5743 -9707 5749 -9677
rect 5998 -9705 6067 -9699
rect 5658 -9865 5749 -9707
rect 5658 -9899 5664 -9865
rect 5743 -9899 5749 -9865
rect 5658 -9915 5749 -9899
rect 5781 -9769 5970 -9705
rect 5781 -9803 5787 -9769
rect 5864 -9803 5970 -9769
rect 5558 -10049 5627 -9947
rect 5781 -9961 5970 -9803
rect 5658 -9995 5787 -9961
rect 5864 -9995 5970 -9961
rect 5558 -10167 5628 -10049
rect 5658 -10123 5970 -9995
rect 5658 -10157 5670 -10123
rect 5846 -10157 5970 -10123
rect 5658 -10163 5858 -10157
rect 5558 -10201 5577 -10167
rect 5611 -10201 5628 -10167
rect 5558 -10218 5628 -10201
rect 5559 -10295 5628 -10218
rect 5558 -10354 5628 -10295
rect 5658 -10211 5858 -10204
rect 5658 -10245 5670 -10211
rect 5846 -10245 5858 -10211
rect 5886 -10218 5970 -10157
rect 5658 -10313 5858 -10245
rect 5658 -10347 5689 -10313
rect 5821 -10347 5858 -10313
rect 5658 -10354 5858 -10347
rect 5901 -10270 5970 -10218
rect 5559 -10470 5628 -10354
rect 5703 -10356 5823 -10354
rect 5703 -10408 5734 -10356
rect 5786 -10408 5823 -10356
rect 5901 -10360 5970 -10339
rect 5998 -9947 6017 -9774
rect 6051 -9947 6067 -9774
rect 6098 -9707 6104 -9673
rect 6183 -9677 6312 -9673
rect 6538 -9660 7357 -9647
rect 6538 -9673 6752 -9660
rect 6183 -9707 6189 -9677
rect 6438 -9705 6507 -9699
rect 6098 -9865 6189 -9707
rect 6098 -9899 6104 -9865
rect 6183 -9899 6189 -9865
rect 6098 -9915 6189 -9899
rect 6221 -9769 6410 -9705
rect 6221 -9803 6227 -9769
rect 6304 -9803 6410 -9769
rect 5998 -10167 6067 -9947
rect 6221 -9961 6410 -9803
rect 6098 -9995 6227 -9961
rect 6304 -9995 6410 -9961
rect 6098 -10123 6410 -9995
rect 6098 -10157 6110 -10123
rect 6286 -10157 6410 -10123
rect 6098 -10163 6298 -10157
rect 5998 -10201 6017 -10167
rect 6051 -10201 6067 -10167
rect 5703 -10439 5823 -10408
rect 5559 -10539 5901 -10470
rect 5559 -10551 5628 -10539
rect 5426 -11137 5492 -11131
rect 5096 -13118 5354 -13052
rect 5420 -13118 5426 -13052
rect 5832 -13132 5901 -10539
rect 5998 -10803 6067 -10201
rect 6098 -10211 6298 -10204
rect 6098 -10245 6110 -10211
rect 6286 -10245 6298 -10211
rect 6326 -10218 6410 -10157
rect 6098 -10313 6298 -10245
rect 6098 -10347 6129 -10313
rect 6261 -10347 6298 -10313
rect 6098 -10354 6172 -10347
rect 6143 -10389 6172 -10354
rect 6224 -10354 6298 -10347
rect 6341 -10272 6410 -10218
rect 6341 -10354 6410 -10341
rect 6438 -9947 6457 -9774
rect 6491 -9947 6507 -9774
rect 6538 -9707 6544 -9673
rect 6623 -9677 6752 -9673
rect 6623 -9707 6629 -9677
rect 6538 -9865 6629 -9707
rect 6538 -9899 6544 -9865
rect 6623 -9899 6629 -9865
rect 6538 -9915 6629 -9899
rect 6661 -9769 6850 -9705
rect 6661 -9803 6667 -9769
rect 6744 -9803 6850 -9769
rect 6438 -10167 6507 -9947
rect 6661 -9961 6850 -9803
rect 6538 -9995 6667 -9961
rect 6744 -9995 6850 -9961
rect 6538 -10123 6850 -9995
rect 6538 -10157 6550 -10123
rect 6726 -10157 6850 -10123
rect 6538 -10163 6738 -10157
rect 6438 -10201 6457 -10167
rect 6491 -10201 6507 -10167
rect 6224 -10389 6263 -10354
rect 6143 -10414 6263 -10389
rect 5992 -10809 6073 -10803
rect 5992 -10878 5998 -10809
rect 6067 -10812 6073 -10809
rect 6067 -10878 6085 -10812
rect 5992 -10884 6073 -10878
rect 5998 -13038 6067 -10884
rect 6438 -10944 6507 -10201
rect 6538 -10211 6738 -10204
rect 6538 -10245 6550 -10211
rect 6726 -10245 6738 -10211
rect 6766 -10218 6850 -10157
rect 6538 -10313 6738 -10245
rect 6781 -10263 6850 -10218
rect 7254 -10257 7357 -9660
rect 11860 -10257 12409 -10256
rect 12750 -10257 13092 -10256
rect 6538 -10347 6569 -10313
rect 6701 -10347 6738 -10313
rect 6538 -10354 6612 -10347
rect 6580 -10380 6612 -10354
rect 6664 -10354 6738 -10347
rect 6780 -10294 6850 -10263
rect 7137 -10258 7964 -10257
rect 8085 -10258 8912 -10257
rect 9021 -10258 9848 -10257
rect 9952 -10258 10779 -10257
rect 7137 -10273 10780 -10258
rect 6664 -10380 6700 -10354
rect 6580 -10423 6700 -10380
rect 6438 -11019 6507 -11013
rect 6780 -10906 6849 -10294
rect 7137 -10308 7389 -10273
rect 7677 -10308 8337 -10273
rect 8625 -10308 9273 -10273
rect 9561 -10308 10204 -10273
rect 10492 -10308 10780 -10273
rect 7137 -10369 10780 -10308
rect 10879 -10273 13092 -10257
rect 10879 -10308 11131 -10273
rect 11419 -10308 13092 -10273
rect 10879 -10369 13092 -10308
rect 7138 -10380 10780 -10369
rect 7138 -10490 7150 -10380
rect 7184 -10490 7342 -10380
rect 7376 -10490 7534 -10380
rect 7568 -10490 7726 -10380
rect 7760 -10490 7918 -10380
rect 7952 -10490 8098 -10380
rect 8132 -10490 8290 -10380
rect 8324 -10490 8482 -10380
rect 8516 -10490 8674 -10380
rect 8708 -10490 8866 -10380
rect 8900 -10490 9034 -10380
rect 9068 -10490 9226 -10380
rect 9260 -10490 9418 -10380
rect 9452 -10490 9610 -10380
rect 9644 -10490 9802 -10380
rect 9836 -10490 9965 -10380
rect 9999 -10490 10157 -10380
rect 10191 -10490 10349 -10380
rect 10383 -10490 10541 -10380
rect 10575 -10490 10733 -10380
rect 10767 -10490 10780 -10380
rect 7138 -10499 10780 -10490
rect 10880 -10380 13092 -10369
rect 10880 -10490 10892 -10380
rect 10926 -10490 11084 -10380
rect 11118 -10490 11276 -10380
rect 11310 -10490 11468 -10380
rect 11502 -10490 11660 -10380
rect 11694 -10490 13092 -10380
rect 10880 -10499 13092 -10490
rect 7138 -10568 8001 -10553
rect 7138 -10680 7245 -10568
rect 7280 -10680 7438 -10568
rect 7473 -10680 7630 -10568
rect 7665 -10680 7822 -10568
rect 7857 -10680 8001 -10568
rect 7138 -10687 8001 -10680
rect 8086 -10568 8949 -10553
rect 8086 -10680 8193 -10568
rect 8228 -10680 8386 -10568
rect 8421 -10680 8578 -10568
rect 8613 -10680 8770 -10568
rect 8805 -10680 8949 -10568
rect 8086 -10687 8949 -10680
rect 9022 -10568 9885 -10553
rect 9022 -10680 9129 -10568
rect 9164 -10680 9322 -10568
rect 9357 -10680 9514 -10568
rect 9549 -10680 9706 -10568
rect 9741 -10680 9885 -10568
rect 9022 -10687 9885 -10680
rect 9953 -10568 10816 -10553
rect 9953 -10680 10060 -10568
rect 10095 -10680 10253 -10568
rect 10288 -10680 10445 -10568
rect 10480 -10680 10637 -10568
rect 10672 -10680 10816 -10568
rect 9953 -10687 10816 -10680
rect 10880 -10568 11743 -10553
rect 10880 -10680 10987 -10568
rect 11022 -10680 11180 -10568
rect 11215 -10680 11372 -10568
rect 11407 -10680 11564 -10568
rect 11599 -10680 11743 -10568
rect 10880 -10687 11743 -10680
rect 7106 -10718 7158 -10717
rect 7102 -10723 7248 -10718
rect 7102 -10775 7106 -10723
rect 7158 -10734 7248 -10723
rect 7158 -10768 7198 -10734
rect 7232 -10768 7248 -10734
rect 7158 -10775 7248 -10768
rect 7102 -10784 7248 -10775
rect 7304 -10734 7441 -10718
rect 7304 -10768 7390 -10734
rect 7424 -10768 7441 -10734
rect 7304 -10784 7441 -10768
rect 7491 -10734 7632 -10719
rect 7491 -10768 7582 -10734
rect 7616 -10768 7632 -10734
rect 7304 -10812 7370 -10784
rect 7097 -10817 7370 -10812
rect 7097 -10869 7113 -10817
rect 7165 -10869 7370 -10817
rect 7491 -10785 7632 -10768
rect 7661 -10734 7825 -10718
rect 7661 -10768 7774 -10734
rect 7808 -10768 7825 -10734
rect 7661 -10784 7825 -10768
rect 7491 -10821 7557 -10785
rect 7594 -10786 7628 -10785
rect 7097 -10878 7370 -10869
rect 7409 -10906 7557 -10821
rect 6780 -10972 7327 -10906
rect 7393 -10972 7557 -10906
rect 6780 -12935 6849 -10972
rect 7661 -11000 7727 -10784
rect 7102 -11066 7727 -11000
rect 7106 -11267 7172 -11066
rect 7891 -11094 8001 -10687
rect 8050 -10724 8196 -10718
rect 8050 -10776 8069 -10724
rect 8122 -10734 8196 -10724
rect 8122 -10768 8146 -10734
rect 8180 -10768 8196 -10734
rect 8122 -10776 8196 -10768
rect 8050 -10784 8196 -10776
rect 8252 -10734 8389 -10718
rect 8252 -10768 8338 -10734
rect 8372 -10768 8389 -10734
rect 8252 -10784 8389 -10768
rect 8439 -10734 8580 -10719
rect 8439 -10768 8530 -10734
rect 8564 -10768 8580 -10734
rect 8252 -10812 8318 -10784
rect 8050 -10816 8318 -10812
rect 8050 -10868 8057 -10816
rect 8109 -10868 8318 -10816
rect 8439 -10785 8580 -10768
rect 8609 -10734 8773 -10718
rect 8609 -10768 8722 -10734
rect 8756 -10768 8773 -10734
rect 8609 -10784 8773 -10768
rect 8439 -10821 8505 -10785
rect 8542 -10786 8576 -10785
rect 8050 -10878 8318 -10868
rect 8357 -10899 8505 -10821
rect 8357 -10906 8424 -10899
rect 8050 -10951 8424 -10906
rect 8493 -10951 8505 -10899
rect 8050 -10972 8505 -10951
rect 8609 -11000 8675 -10784
rect 7106 -11339 7172 -11333
rect 7214 -11106 7413 -11094
rect 7214 -11118 7372 -11106
rect 7214 -11869 7298 -11118
rect 7333 -11869 7372 -11118
rect 7214 -12047 7227 -11869
rect 7406 -11882 7413 -11106
rect 7405 -12034 7413 -11882
rect 7750 -11106 8001 -11094
rect 7750 -11882 7756 -11106
rect 7790 -11109 8001 -11106
rect 8050 -11066 8675 -11000
rect 7790 -11524 8000 -11109
rect 8050 -11371 8116 -11066
rect 8839 -11094 8949 -10687
rect 8986 -10723 9132 -10718
rect 8986 -10775 9002 -10723
rect 9055 -10734 9132 -10723
rect 9055 -10768 9082 -10734
rect 9116 -10768 9132 -10734
rect 9055 -10775 9132 -10768
rect 8986 -10784 9132 -10775
rect 9188 -10734 9325 -10718
rect 9188 -10768 9274 -10734
rect 9308 -10768 9325 -10734
rect 9188 -10784 9325 -10768
rect 9375 -10734 9516 -10719
rect 9375 -10768 9466 -10734
rect 9500 -10768 9516 -10734
rect 9188 -10812 9254 -10784
rect 8986 -10821 9254 -10812
rect 9375 -10785 9516 -10768
rect 9545 -10734 9709 -10718
rect 9545 -10768 9658 -10734
rect 9692 -10768 9709 -10734
rect 9545 -10784 9709 -10768
rect 9375 -10821 9441 -10785
rect 9478 -10786 9512 -10785
rect 8986 -10873 9000 -10821
rect 9052 -10873 9254 -10821
rect 8986 -10878 9254 -10873
rect 9293 -10906 9441 -10821
rect 8986 -10912 9441 -10906
rect 8986 -10965 8989 -10912
rect 9042 -10965 9441 -10912
rect 8986 -10972 9441 -10965
rect 9545 -11000 9611 -10784
rect 8050 -11443 8116 -11437
rect 8162 -11106 8361 -11094
rect 8162 -11118 8320 -11106
rect 7790 -11590 7872 -11524
rect 7938 -11590 8000 -11524
rect 7790 -11882 8000 -11590
rect 7750 -11894 8000 -11882
rect 8162 -11869 8246 -11118
rect 8281 -11869 8320 -11118
rect 8354 -11882 8361 -11106
rect 7102 -12693 7168 -12687
rect 7102 -12850 7168 -12759
rect 7214 -12798 7298 -12047
rect 7333 -12798 7372 -12047
rect 7214 -12810 7372 -12798
rect 7406 -12810 7413 -12034
rect 7214 -12822 7413 -12810
rect 7750 -12034 8000 -12022
rect 7750 -12810 7756 -12034
rect 7790 -12317 8000 -12034
rect 7790 -12383 7853 -12317
rect 7919 -12383 8000 -12317
rect 7790 -12807 8000 -12383
rect 8340 -12034 8361 -11882
rect 8698 -11106 8949 -11094
rect 8698 -11882 8704 -11106
rect 8738 -11109 8949 -11106
rect 8986 -11065 9611 -11000
rect 8738 -11270 8948 -11109
rect 9052 -11066 9611 -11065
rect 9775 -11022 9885 -10687
rect 10706 -10718 10816 -10687
rect 9917 -10723 10063 -10718
rect 9917 -10775 9933 -10723
rect 9986 -10734 10063 -10723
rect 9986 -10768 10013 -10734
rect 10047 -10768 10063 -10734
rect 9986 -10775 10063 -10768
rect 9917 -10784 10063 -10775
rect 10119 -10734 10256 -10718
rect 10119 -10768 10205 -10734
rect 10239 -10768 10256 -10734
rect 10119 -10784 10256 -10768
rect 10306 -10734 10447 -10719
rect 10306 -10768 10397 -10734
rect 10431 -10768 10447 -10734
rect 10119 -10812 10185 -10784
rect 9917 -10821 10185 -10812
rect 10306 -10785 10447 -10768
rect 10476 -10734 10640 -10718
rect 10476 -10768 10589 -10734
rect 10623 -10768 10640 -10734
rect 10476 -10784 10640 -10768
rect 10706 -10734 10990 -10718
rect 10706 -10768 10940 -10734
rect 10974 -10768 10990 -10734
rect 10706 -10784 10990 -10768
rect 11046 -10734 11183 -10718
rect 11046 -10768 11132 -10734
rect 11166 -10768 11183 -10734
rect 11046 -10784 11183 -10768
rect 11233 -10734 11374 -10719
rect 11233 -10768 11324 -10734
rect 11358 -10768 11374 -10734
rect 10306 -10821 10372 -10785
rect 10409 -10786 10443 -10785
rect 9917 -10873 9935 -10821
rect 9987 -10873 10185 -10821
rect 9917 -10878 10185 -10873
rect 10224 -10868 10372 -10821
rect 10224 -10906 10262 -10868
rect 9917 -10937 10262 -10906
rect 10331 -10937 10372 -10868
rect 9917 -10972 10372 -10937
rect 10476 -11000 10542 -10784
rect 9775 -11088 9798 -11022
rect 9864 -11088 9885 -11022
rect 9775 -11094 9885 -11088
rect 8986 -11149 9052 -11131
rect 9098 -11106 9297 -11094
rect 9098 -11118 9256 -11106
rect 8738 -11336 8818 -11270
rect 8884 -11336 8948 -11270
rect 8738 -11882 8948 -11336
rect 8698 -11894 8948 -11882
rect 9098 -11869 9182 -11118
rect 9217 -11869 9256 -11118
rect 9290 -11882 9297 -11106
rect 8162 -12798 8246 -12047
rect 8281 -12798 8320 -12047
rect 7790 -12810 8001 -12807
rect 7750 -12822 8001 -12810
rect 7102 -12916 7727 -12850
rect 6774 -13004 6780 -12935
rect 6849 -12944 6855 -12935
rect 6849 -13004 7557 -12944
rect 6780 -13010 7557 -13004
rect 5998 -13102 6066 -13038
rect 5999 -13104 6066 -13102
rect 6132 -13104 7370 -13038
rect 7409 -13095 7557 -13010
rect 7304 -13132 7370 -13104
rect 7491 -13131 7557 -13095
rect 7594 -13131 7628 -13130
rect 5832 -13198 6941 -13132
rect 7007 -13148 7248 -13132
rect 7007 -13182 7198 -13148
rect 7232 -13182 7248 -13148
rect 7007 -13198 7248 -13182
rect 7304 -13148 7441 -13132
rect 7304 -13182 7390 -13148
rect 7424 -13182 7441 -13148
rect 7304 -13198 7441 -13182
rect 7491 -13148 7632 -13131
rect 7491 -13182 7582 -13148
rect 7616 -13182 7632 -13148
rect 7491 -13197 7632 -13182
rect 7661 -13132 7727 -12916
rect 7661 -13148 7825 -13132
rect 7661 -13182 7774 -13148
rect 7808 -13182 7825 -13148
rect 7661 -13198 7825 -13182
rect 5832 -13208 5901 -13198
rect 7891 -13229 8001 -12822
rect 8050 -12814 8116 -12808
rect 8162 -12810 8320 -12798
rect 8354 -12810 8361 -12034
rect 8162 -12822 8361 -12810
rect 8698 -12034 8948 -12022
rect 8698 -12810 8704 -12034
rect 8738 -12727 8948 -12034
rect 9276 -12034 9297 -11882
rect 9634 -11106 9885 -11094
rect 9634 -11882 9640 -11106
rect 9674 -11109 9885 -11106
rect 9917 -11066 10542 -11000
rect 9674 -11882 9884 -11109
rect 9917 -11161 9983 -11066
rect 10706 -11094 10816 -10784
rect 11046 -10812 11112 -10784
rect 10844 -10878 10860 -10812
rect 10926 -10878 11112 -10812
rect 11233 -10785 11374 -10768
rect 11403 -10734 11567 -10718
rect 11403 -10768 11516 -10734
rect 11550 -10768 11567 -10734
rect 11403 -10784 11567 -10768
rect 11233 -10821 11299 -10785
rect 11336 -10786 11370 -10785
rect 11151 -10906 11299 -10821
rect 10844 -10972 10858 -10906
rect 10924 -10972 11299 -10906
rect 11403 -11000 11469 -10784
rect 10844 -11066 10850 -11000
rect 10915 -11066 11469 -11000
rect 11633 -11094 11743 -10687
rect 9917 -11233 9983 -11227
rect 10029 -11106 10228 -11094
rect 10029 -11118 10187 -11106
rect 9634 -11894 9884 -11882
rect 10029 -11869 10113 -11118
rect 10148 -11869 10187 -11118
rect 10221 -11882 10228 -11106
rect 8738 -12793 8837 -12727
rect 8903 -12793 8948 -12727
rect 8738 -12807 8948 -12793
rect 8989 -12473 9055 -12467
rect 8738 -12810 8949 -12807
rect 8698 -12822 8949 -12810
rect 8116 -12880 8675 -12850
rect 8050 -12916 8675 -12880
rect 8050 -12951 8505 -12944
rect 8050 -13010 8401 -12951
rect 8357 -13015 8401 -13010
rect 8465 -13015 8505 -12951
rect 8050 -13047 8318 -13038
rect 8050 -13099 8079 -13047
rect 8131 -13099 8318 -13047
rect 8357 -13095 8505 -13015
rect 8050 -13104 8318 -13099
rect 8252 -13132 8318 -13104
rect 8439 -13131 8505 -13095
rect 8542 -13131 8576 -13130
rect 8050 -13141 8196 -13132
rect 8050 -13193 8063 -13141
rect 8128 -13148 8196 -13141
rect 8128 -13182 8146 -13148
rect 8180 -13182 8196 -13148
rect 8128 -13193 8196 -13182
rect 8050 -13198 8196 -13193
rect 8252 -13148 8389 -13132
rect 8252 -13182 8338 -13148
rect 8372 -13182 8389 -13148
rect 8252 -13198 8389 -13182
rect 8439 -13148 8580 -13131
rect 8439 -13182 8530 -13148
rect 8564 -13182 8580 -13148
rect 8439 -13197 8580 -13182
rect 8609 -13132 8675 -12916
rect 8609 -13148 8773 -13132
rect 8609 -13182 8722 -13148
rect 8756 -13182 8773 -13148
rect 8609 -13198 8773 -13182
rect 8839 -13229 8949 -12822
rect 8989 -12850 9055 -12539
rect 9098 -12798 9182 -12047
rect 9217 -12798 9256 -12047
rect 9098 -12810 9256 -12798
rect 9290 -12810 9297 -12034
rect 9098 -12822 9297 -12810
rect 9634 -12034 9884 -12022
rect 9634 -12810 9640 -12034
rect 9674 -12807 9884 -12034
rect 10206 -12033 10228 -11882
rect 10565 -11106 10816 -11094
rect 10565 -11882 10571 -11106
rect 10605 -11109 10816 -11106
rect 10956 -11106 11155 -11094
rect 10605 -11882 10815 -11109
rect 10565 -11894 10815 -11882
rect 10956 -11118 11114 -11106
rect 10956 -11869 11040 -11118
rect 11075 -11869 11114 -11118
rect 11148 -11882 11155 -11106
rect 9917 -12595 9983 -12589
rect 9674 -12810 9885 -12807
rect 9634 -12821 9885 -12810
rect 9634 -12822 9807 -12821
rect 8986 -12916 9611 -12850
rect 8986 -13010 8993 -12944
rect 9059 -13010 9441 -12944
rect 8986 -13104 9001 -13038
rect 9067 -13104 9254 -13038
rect 9293 -13095 9441 -13010
rect 9188 -13132 9254 -13104
rect 9375 -13131 9441 -13095
rect 9478 -13131 9512 -13130
rect 8986 -13141 9132 -13132
rect 8986 -13193 8992 -13141
rect 9057 -13148 9132 -13141
rect 9057 -13182 9082 -13148
rect 9116 -13182 9132 -13148
rect 9057 -13193 9132 -13182
rect 8986 -13198 9132 -13193
rect 9188 -13148 9325 -13132
rect 9188 -13182 9274 -13148
rect 9308 -13182 9325 -13148
rect 9188 -13198 9325 -13182
rect 9375 -13148 9516 -13131
rect 9375 -13182 9466 -13148
rect 9500 -13182 9516 -13148
rect 9375 -13197 9516 -13182
rect 9545 -13132 9611 -12916
rect 9775 -12885 9807 -12822
rect 9873 -12885 9885 -12821
rect 9545 -13148 9709 -13132
rect 9545 -13182 9658 -13148
rect 9692 -13182 9709 -13148
rect 9545 -13198 9709 -13182
rect 9775 -13229 9885 -12885
rect 9917 -12849 9983 -12661
rect 10029 -12797 10113 -12046
rect 10148 -12797 10187 -12046
rect 10029 -12809 10187 -12797
rect 10221 -12809 10228 -12033
rect 10029 -12821 10228 -12809
rect 10565 -12033 10815 -12021
rect 10565 -12809 10571 -12033
rect 10605 -12806 10815 -12033
rect 11134 -12034 11155 -11882
rect 11492 -11106 11743 -11094
rect 11492 -11882 11498 -11106
rect 11532 -11109 11743 -11106
rect 11860 -10723 13092 -10499
rect 11860 -10926 12189 -10723
rect 12410 -10926 13092 -10723
rect 11532 -11865 11742 -11109
rect 11860 -11424 13092 -10926
rect 11799 -11432 13092 -11424
rect 11799 -11483 11811 -11432
rect 12168 -11441 13092 -11432
rect 12168 -11483 12180 -11441
rect 11799 -11490 12180 -11483
rect 11860 -11528 11903 -11490
rect 12726 -11575 13092 -11441
rect 11875 -11587 12689 -11575
rect 12726 -11582 13137 -11575
rect 11875 -11677 11881 -11587
rect 11915 -11677 12073 -11587
rect 12107 -11677 12265 -11587
rect 12299 -11677 12457 -11587
rect 12491 -11677 12649 -11587
rect 12683 -11677 12689 -11587
rect 11875 -11689 12689 -11677
rect 12923 -11619 13137 -11582
rect 12923 -11653 12986 -11619
rect 13077 -11653 13137 -11619
rect 12923 -11691 13137 -11653
rect 11779 -11729 12209 -11717
rect 11779 -11819 11785 -11729
rect 11819 -11819 11977 -11729
rect 12011 -11819 12169 -11729
rect 12203 -11819 12209 -11729
rect 11779 -11831 12209 -11819
rect 12355 -11723 12827 -11717
rect 12355 -11729 12892 -11723
rect 12355 -11819 12361 -11729
rect 12395 -11819 12553 -11729
rect 12587 -11819 12745 -11729
rect 12779 -11739 12892 -11729
rect 12779 -11819 12842 -11739
rect 12355 -11831 12842 -11819
rect 11532 -11881 12263 -11865
rect 11532 -11882 12170 -11881
rect 11492 -11894 12170 -11882
rect 11737 -11915 12170 -11894
rect 12204 -11915 12263 -11881
rect 11737 -11931 12263 -11915
rect 12702 -11965 12842 -11831
rect 12876 -11965 12892 -11739
rect 12923 -11725 12929 -11691
rect 13008 -11695 13137 -11691
rect 13008 -11725 13014 -11695
rect 12923 -11883 13014 -11725
rect 12923 -11917 12929 -11883
rect 13008 -11917 13014 -11883
rect 12923 -11933 13014 -11917
rect 13046 -11787 13235 -11723
rect 13046 -11821 13052 -11787
rect 13129 -11821 13235 -11787
rect 11703 -11986 12363 -11970
rect 11703 -12020 12313 -11986
rect 12347 -12020 12363 -11986
rect 11703 -12022 12363 -12020
rect 10956 -12798 11040 -12047
rect 11075 -12798 11114 -12047
rect 10605 -12809 10816 -12806
rect 10565 -12821 10816 -12809
rect 9917 -12915 10542 -12849
rect 9917 -12951 10372 -12943
rect 9917 -13009 10264 -12951
rect 10224 -13011 10264 -13009
rect 10324 -13011 10372 -12951
rect 9917 -13103 9937 -13037
rect 10003 -13103 10185 -13037
rect 10224 -13094 10372 -13011
rect 10119 -13131 10185 -13103
rect 10306 -13130 10372 -13094
rect 10409 -13130 10443 -13129
rect 9917 -13141 10063 -13131
rect 9917 -13193 9951 -13141
rect 10016 -13147 10063 -13141
rect 10047 -13181 10063 -13147
rect 10016 -13193 10063 -13181
rect 9917 -13197 10063 -13193
rect 10119 -13147 10256 -13131
rect 10119 -13181 10205 -13147
rect 10239 -13181 10256 -13147
rect 10119 -13197 10256 -13181
rect 10306 -13147 10447 -13130
rect 10306 -13181 10397 -13147
rect 10431 -13181 10447 -13147
rect 10306 -13196 10447 -13181
rect 10476 -13131 10542 -12915
rect 10476 -13147 10640 -13131
rect 10476 -13181 10589 -13147
rect 10623 -13181 10640 -13147
rect 10476 -13197 10640 -13181
rect 10706 -13132 10816 -12821
rect 10956 -12810 11114 -12798
rect 11148 -12810 11155 -12034
rect 10956 -12822 11155 -12810
rect 11492 -12034 12363 -12022
rect 11492 -12810 11498 -12034
rect 11532 -12036 12363 -12034
rect 11532 -12067 11815 -12036
rect 11532 -12807 11742 -12067
rect 12259 -12070 12305 -12064
rect 12702 -12070 12892 -11965
rect 13046 -11946 13235 -11821
rect 13046 -11979 15435 -11946
rect 12259 -12076 12892 -12070
rect 12259 -12252 12265 -12076
rect 12299 -12185 12892 -12076
rect 12923 -12013 13052 -11979
rect 13129 -12012 15435 -11979
rect 13129 -12013 13235 -12012
rect 12923 -12141 13235 -12013
rect 12923 -12175 12935 -12141
rect 13111 -12175 13235 -12141
rect 12923 -12181 13123 -12175
rect 12299 -12219 12842 -12185
rect 12876 -12219 12892 -12185
rect 12299 -12236 12892 -12219
rect 12923 -12229 13123 -12222
rect 12299 -12252 12827 -12236
rect 12259 -12264 12827 -12252
rect 12305 -12268 12827 -12264
rect 12923 -12263 12935 -12229
rect 13111 -12263 13123 -12229
rect 13151 -12236 13235 -12175
rect 12305 -12269 12825 -12268
rect 12305 -12270 12774 -12269
rect 12171 -12335 12394 -12328
rect 12171 -12383 12183 -12335
rect 12074 -12396 12183 -12383
rect 12382 -12383 12394 -12335
rect 12923 -12331 13123 -12263
rect 12923 -12365 12954 -12331
rect 13086 -12365 13123 -12331
rect 12921 -12372 13123 -12365
rect 12382 -12396 12473 -12383
rect 12074 -12499 12233 -12396
rect 12352 -12499 12473 -12396
rect 12921 -12421 13121 -12372
rect 12921 -12443 12960 -12421
rect 12074 -12573 12473 -12499
rect 12923 -12540 12960 -12443
rect 13079 -12443 13121 -12421
rect 13079 -12540 13113 -12443
rect 12923 -12598 13113 -12540
rect 11532 -12810 11743 -12807
rect 11492 -12822 11743 -12810
rect 10844 -12916 10850 -12850
rect 10916 -12916 11469 -12850
rect 10844 -13010 10888 -12944
rect 10954 -13010 11299 -12944
rect 10844 -13104 10859 -13038
rect 10925 -13104 11112 -13038
rect 11151 -13095 11299 -13010
rect 11046 -13132 11112 -13104
rect 11233 -13131 11299 -13095
rect 11336 -13131 11370 -13130
rect 10706 -13148 10990 -13132
rect 10706 -13182 10940 -13148
rect 10974 -13182 10990 -13148
rect 10706 -13198 10990 -13182
rect 11046 -13148 11183 -13132
rect 11046 -13182 11132 -13148
rect 11166 -13182 11183 -13148
rect 11046 -13198 11183 -13182
rect 11233 -13148 11374 -13131
rect 11233 -13182 11324 -13148
rect 11358 -13182 11374 -13148
rect 11233 -13197 11374 -13182
rect 11403 -13132 11469 -12916
rect 11403 -13148 11567 -13132
rect 11403 -13182 11516 -13148
rect 11550 -13182 11567 -13148
rect 11403 -13198 11567 -13182
rect 10706 -13228 10816 -13198
rect 7138 -13236 8001 -13229
rect 7138 -13348 7245 -13236
rect 7280 -13348 7438 -13236
rect 7473 -13348 7630 -13236
rect 7665 -13348 7822 -13236
rect 7857 -13348 8001 -13236
rect 7138 -13363 8001 -13348
rect 8086 -13236 8949 -13229
rect 8086 -13348 8193 -13236
rect 8228 -13348 8386 -13236
rect 8421 -13348 8578 -13236
rect 8613 -13348 8770 -13236
rect 8805 -13348 8949 -13236
rect 8086 -13363 8949 -13348
rect 9022 -13236 9885 -13229
rect 9022 -13348 9129 -13236
rect 9164 -13348 9322 -13236
rect 9357 -13348 9514 -13236
rect 9549 -13348 9706 -13236
rect 9741 -13348 9885 -13236
rect 9022 -13363 9885 -13348
rect 9953 -13235 10816 -13228
rect 11633 -13229 11743 -12822
rect 9953 -13347 10060 -13235
rect 10095 -13347 10253 -13235
rect 10288 -13347 10445 -13235
rect 10480 -13347 10637 -13235
rect 10672 -13347 10816 -13235
rect 9953 -13362 10816 -13347
rect 10880 -13236 11743 -13229
rect 10880 -13348 10987 -13236
rect 11022 -13348 11180 -13236
rect 11215 -13348 11372 -13236
rect 11407 -13348 11564 -13236
rect 11599 -13348 11743 -13236
rect 10880 -13363 11743 -13348
rect 7137 -13425 10779 -13416
rect 11883 -13417 12147 -13406
rect 7137 -13426 9965 -13425
rect 7137 -13536 7150 -13426
rect 7184 -13536 7342 -13426
rect 7376 -13536 7534 -13426
rect 7568 -13536 7726 -13426
rect 7760 -13536 7918 -13426
rect 7952 -13536 8098 -13426
rect 8132 -13536 8290 -13426
rect 8324 -13536 8482 -13426
rect 8516 -13536 8674 -13426
rect 8708 -13536 8866 -13426
rect 8900 -13536 9034 -13426
rect 9068 -13536 9226 -13426
rect 9260 -13536 9418 -13426
rect 9452 -13536 9610 -13426
rect 9644 -13536 9802 -13426
rect 9836 -13535 9965 -13426
rect 9999 -13535 10157 -13425
rect 10191 -13535 10349 -13425
rect 10383 -13535 10541 -13425
rect 10575 -13535 10733 -13425
rect 10767 -13535 10779 -13425
rect 9836 -13536 10779 -13535
rect 7137 -13607 10779 -13536
rect 10880 -13426 11894 -13417
rect 10880 -13536 10892 -13426
rect 10926 -13536 11084 -13426
rect 11118 -13536 11276 -13426
rect 11310 -13536 11468 -13426
rect 11502 -13536 11660 -13426
rect 11694 -13536 11894 -13426
rect 10880 -13547 11894 -13536
rect 7137 -13608 10204 -13607
rect 7137 -13643 7389 -13608
rect 7677 -13643 8337 -13608
rect 8625 -13643 9273 -13608
rect 9561 -13642 10204 -13608
rect 10492 -13642 10779 -13607
rect 9561 -13643 10779 -13642
rect 7137 -13657 10779 -13643
rect 7137 -13659 7964 -13657
rect 8085 -13659 8912 -13657
rect 9021 -13659 9848 -13657
rect 9952 -13658 10779 -13657
rect 10879 -13608 11894 -13547
rect 10879 -13643 11131 -13608
rect 11419 -13643 11894 -13608
rect 10879 -13659 11894 -13643
rect 12136 -13659 12147 -13417
rect 11883 -13670 12147 -13659
rect 5658 -14129 7357 -14085
rect 5658 -14163 5721 -14129
rect 5812 -14163 6161 -14129
rect 6252 -14163 6601 -14129
rect 6692 -14163 7357 -14129
rect 5658 -14175 7357 -14163
rect 5658 -14201 5872 -14175
rect 5558 -14233 5627 -14227
rect 5558 -14475 5577 -14302
rect 5611 -14475 5627 -14302
rect 5658 -14235 5664 -14201
rect 5743 -14205 5872 -14201
rect 6098 -14201 6312 -14175
rect 5743 -14235 5749 -14205
rect 5998 -14233 6067 -14227
rect 5658 -14393 5749 -14235
rect 5658 -14427 5664 -14393
rect 5743 -14427 5749 -14393
rect 5658 -14443 5749 -14427
rect 5781 -14297 5970 -14233
rect 5781 -14331 5787 -14297
rect 5864 -14331 5970 -14297
rect 5558 -14577 5627 -14475
rect 5781 -14489 5970 -14331
rect 5658 -14523 5787 -14489
rect 5864 -14523 5970 -14489
rect 5558 -14695 5628 -14577
rect 5658 -14651 5970 -14523
rect 5658 -14685 5670 -14651
rect 5846 -14685 5970 -14651
rect 5658 -14691 5858 -14685
rect 5558 -14729 5577 -14695
rect 5611 -14729 5628 -14695
rect 5558 -14746 5628 -14729
rect 5559 -14823 5628 -14746
rect 5558 -14882 5628 -14823
rect 5658 -14739 5858 -14732
rect 5658 -14773 5670 -14739
rect 5846 -14773 5858 -14739
rect 5886 -14746 5970 -14685
rect 5658 -14841 5858 -14773
rect 5658 -14875 5689 -14841
rect 5821 -14875 5858 -14841
rect 5658 -14882 5858 -14875
rect 5901 -14798 5970 -14746
rect 5559 -14998 5628 -14882
rect 5703 -14884 5823 -14882
rect 5703 -14936 5734 -14884
rect 5786 -14936 5823 -14884
rect 5901 -14888 5970 -14867
rect 5998 -14475 6017 -14302
rect 6051 -14475 6067 -14302
rect 6098 -14235 6104 -14201
rect 6183 -14205 6312 -14201
rect 6538 -14188 7357 -14175
rect 6538 -14201 6752 -14188
rect 6183 -14235 6189 -14205
rect 6438 -14233 6507 -14227
rect 6098 -14393 6189 -14235
rect 6098 -14427 6104 -14393
rect 6183 -14427 6189 -14393
rect 6098 -14443 6189 -14427
rect 6221 -14297 6410 -14233
rect 6221 -14331 6227 -14297
rect 6304 -14331 6410 -14297
rect 5998 -14695 6067 -14475
rect 6221 -14489 6410 -14331
rect 6098 -14523 6227 -14489
rect 6304 -14523 6410 -14489
rect 6098 -14651 6410 -14523
rect 6098 -14685 6110 -14651
rect 6286 -14685 6410 -14651
rect 6098 -14691 6298 -14685
rect 5998 -14729 6017 -14695
rect 6051 -14729 6067 -14695
rect 5703 -14967 5823 -14936
rect 5559 -15067 5901 -14998
rect 5559 -15079 5628 -15067
rect 4948 -15813 5473 -15747
rect 5407 -17552 5473 -15813
rect 5401 -17619 5407 -17552
rect 5473 -17619 5479 -17552
rect 5832 -17660 5901 -15067
rect 5998 -15331 6067 -14729
rect 6098 -14739 6298 -14732
rect 6098 -14773 6110 -14739
rect 6286 -14773 6298 -14739
rect 6326 -14746 6410 -14685
rect 6098 -14841 6298 -14773
rect 6098 -14875 6129 -14841
rect 6261 -14875 6298 -14841
rect 6098 -14882 6172 -14875
rect 6143 -14917 6172 -14882
rect 6224 -14882 6298 -14875
rect 6341 -14800 6410 -14746
rect 6341 -14882 6410 -14869
rect 6438 -14475 6457 -14302
rect 6491 -14475 6507 -14302
rect 6538 -14235 6544 -14201
rect 6623 -14205 6752 -14201
rect 6623 -14235 6629 -14205
rect 6538 -14393 6629 -14235
rect 6538 -14427 6544 -14393
rect 6623 -14427 6629 -14393
rect 6538 -14443 6629 -14427
rect 6661 -14297 6850 -14233
rect 6661 -14331 6667 -14297
rect 6744 -14331 6850 -14297
rect 6438 -14695 6507 -14475
rect 6661 -14489 6850 -14331
rect 6538 -14523 6667 -14489
rect 6744 -14523 6850 -14489
rect 6538 -14651 6850 -14523
rect 6538 -14685 6550 -14651
rect 6726 -14685 6850 -14651
rect 6538 -14691 6738 -14685
rect 6438 -14729 6457 -14695
rect 6491 -14729 6507 -14695
rect 6224 -14917 6263 -14882
rect 6143 -14942 6263 -14917
rect 5992 -15337 6073 -15331
rect 5992 -15406 5998 -15337
rect 6067 -15340 6073 -15337
rect 6067 -15406 6085 -15340
rect 5992 -15412 6073 -15406
rect 5998 -17566 6067 -15412
rect 6438 -15472 6507 -14729
rect 6538 -14739 6738 -14732
rect 6538 -14773 6550 -14739
rect 6726 -14773 6738 -14739
rect 6766 -14746 6850 -14685
rect 6538 -14841 6738 -14773
rect 6781 -14791 6850 -14746
rect 7254 -14785 7357 -14188
rect 11860 -14785 12409 -14784
rect 12750 -14785 13092 -14784
rect 6538 -14875 6569 -14841
rect 6701 -14875 6738 -14841
rect 6538 -14882 6612 -14875
rect 6580 -14908 6612 -14882
rect 6664 -14882 6738 -14875
rect 6780 -14822 6850 -14791
rect 7137 -14786 7964 -14785
rect 8085 -14786 8912 -14785
rect 9021 -14786 9848 -14785
rect 9952 -14786 10779 -14785
rect 7137 -14801 10780 -14786
rect 6664 -14908 6700 -14882
rect 6580 -14951 6700 -14908
rect 6438 -15547 6507 -15541
rect 6780 -15434 6849 -14822
rect 7137 -14836 7389 -14801
rect 7677 -14836 8337 -14801
rect 8625 -14836 9273 -14801
rect 9561 -14836 10204 -14801
rect 10492 -14836 10780 -14801
rect 7137 -14897 10780 -14836
rect 10879 -14801 13092 -14785
rect 10879 -14836 11131 -14801
rect 11419 -14836 13092 -14801
rect 10879 -14897 13092 -14836
rect 7138 -14908 10780 -14897
rect 7138 -15018 7150 -14908
rect 7184 -15018 7342 -14908
rect 7376 -15018 7534 -14908
rect 7568 -15018 7726 -14908
rect 7760 -15018 7918 -14908
rect 7952 -15018 8098 -14908
rect 8132 -15018 8290 -14908
rect 8324 -15018 8482 -14908
rect 8516 -15018 8674 -14908
rect 8708 -15018 8866 -14908
rect 8900 -15018 9034 -14908
rect 9068 -15018 9226 -14908
rect 9260 -15018 9418 -14908
rect 9452 -15018 9610 -14908
rect 9644 -15018 9802 -14908
rect 9836 -15018 9965 -14908
rect 9999 -15018 10157 -14908
rect 10191 -15018 10349 -14908
rect 10383 -15018 10541 -14908
rect 10575 -15018 10733 -14908
rect 10767 -15018 10780 -14908
rect 7138 -15027 10780 -15018
rect 10880 -14908 13092 -14897
rect 10880 -15018 10892 -14908
rect 10926 -15018 11084 -14908
rect 11118 -15018 11276 -14908
rect 11310 -15018 11468 -14908
rect 11502 -15018 11660 -14908
rect 11694 -15018 13092 -14908
rect 10880 -15027 13092 -15018
rect 7138 -15096 8001 -15081
rect 7138 -15208 7245 -15096
rect 7280 -15208 7438 -15096
rect 7473 -15208 7630 -15096
rect 7665 -15208 7822 -15096
rect 7857 -15208 8001 -15096
rect 7138 -15215 8001 -15208
rect 8086 -15096 8949 -15081
rect 8086 -15208 8193 -15096
rect 8228 -15208 8386 -15096
rect 8421 -15208 8578 -15096
rect 8613 -15208 8770 -15096
rect 8805 -15208 8949 -15096
rect 8086 -15215 8949 -15208
rect 9022 -15096 9885 -15081
rect 9022 -15208 9129 -15096
rect 9164 -15208 9322 -15096
rect 9357 -15208 9514 -15096
rect 9549 -15208 9706 -15096
rect 9741 -15208 9885 -15096
rect 9022 -15215 9885 -15208
rect 9953 -15096 10816 -15081
rect 9953 -15208 10060 -15096
rect 10095 -15208 10253 -15096
rect 10288 -15208 10445 -15096
rect 10480 -15208 10637 -15096
rect 10672 -15208 10816 -15096
rect 9953 -15215 10816 -15208
rect 10880 -15096 11743 -15081
rect 10880 -15208 10987 -15096
rect 11022 -15208 11180 -15096
rect 11215 -15208 11372 -15096
rect 11407 -15208 11564 -15096
rect 11599 -15208 11743 -15096
rect 10880 -15215 11743 -15208
rect 7106 -15246 7158 -15245
rect 7102 -15251 7248 -15246
rect 7102 -15303 7106 -15251
rect 7158 -15262 7248 -15251
rect 7158 -15296 7198 -15262
rect 7232 -15296 7248 -15262
rect 7158 -15303 7248 -15296
rect 7102 -15312 7248 -15303
rect 7304 -15262 7441 -15246
rect 7304 -15296 7390 -15262
rect 7424 -15296 7441 -15262
rect 7304 -15312 7441 -15296
rect 7491 -15262 7632 -15247
rect 7491 -15296 7582 -15262
rect 7616 -15296 7632 -15262
rect 7304 -15340 7370 -15312
rect 7097 -15345 7370 -15340
rect 7097 -15397 7113 -15345
rect 7165 -15397 7370 -15345
rect 7491 -15313 7632 -15296
rect 7661 -15262 7825 -15246
rect 7661 -15296 7774 -15262
rect 7808 -15296 7825 -15262
rect 7661 -15312 7825 -15296
rect 7491 -15349 7557 -15313
rect 7594 -15314 7628 -15313
rect 7097 -15406 7370 -15397
rect 7409 -15434 7557 -15349
rect 6780 -15500 7327 -15434
rect 7393 -15500 7557 -15434
rect 6780 -17463 6849 -15500
rect 7661 -15528 7727 -15312
rect 7102 -15594 7727 -15528
rect 7106 -15795 7172 -15594
rect 7891 -15622 8001 -15215
rect 8050 -15252 8196 -15246
rect 8050 -15304 8069 -15252
rect 8122 -15262 8196 -15252
rect 8122 -15296 8146 -15262
rect 8180 -15296 8196 -15262
rect 8122 -15304 8196 -15296
rect 8050 -15312 8196 -15304
rect 8252 -15262 8389 -15246
rect 8252 -15296 8338 -15262
rect 8372 -15296 8389 -15262
rect 8252 -15312 8389 -15296
rect 8439 -15262 8580 -15247
rect 8439 -15296 8530 -15262
rect 8564 -15296 8580 -15262
rect 8252 -15340 8318 -15312
rect 8050 -15344 8318 -15340
rect 8050 -15396 8057 -15344
rect 8109 -15396 8318 -15344
rect 8439 -15313 8580 -15296
rect 8609 -15262 8773 -15246
rect 8609 -15296 8722 -15262
rect 8756 -15296 8773 -15262
rect 8609 -15312 8773 -15296
rect 8439 -15349 8505 -15313
rect 8542 -15314 8576 -15313
rect 8050 -15406 8318 -15396
rect 8357 -15427 8505 -15349
rect 8357 -15434 8424 -15427
rect 8050 -15479 8424 -15434
rect 8493 -15479 8505 -15427
rect 8050 -15500 8505 -15479
rect 8609 -15528 8675 -15312
rect 7106 -15867 7172 -15861
rect 7214 -15634 7413 -15622
rect 7214 -15646 7372 -15634
rect 7214 -16397 7298 -15646
rect 7333 -16397 7372 -15646
rect 7214 -16575 7227 -16397
rect 7406 -16410 7413 -15634
rect 7405 -16562 7413 -16410
rect 7750 -15634 8001 -15622
rect 7750 -16410 7756 -15634
rect 7790 -15637 8001 -15634
rect 8050 -15594 8675 -15528
rect 7790 -16052 8000 -15637
rect 8050 -15899 8116 -15594
rect 8839 -15622 8949 -15215
rect 8986 -15251 9132 -15246
rect 8986 -15303 9002 -15251
rect 9055 -15262 9132 -15251
rect 9055 -15296 9082 -15262
rect 9116 -15296 9132 -15262
rect 9055 -15303 9132 -15296
rect 8986 -15312 9132 -15303
rect 9188 -15262 9325 -15246
rect 9188 -15296 9274 -15262
rect 9308 -15296 9325 -15262
rect 9188 -15312 9325 -15296
rect 9375 -15262 9516 -15247
rect 9375 -15296 9466 -15262
rect 9500 -15296 9516 -15262
rect 9188 -15340 9254 -15312
rect 8986 -15349 9254 -15340
rect 9375 -15313 9516 -15296
rect 9545 -15262 9709 -15246
rect 9545 -15296 9658 -15262
rect 9692 -15296 9709 -15262
rect 9545 -15312 9709 -15296
rect 9375 -15349 9441 -15313
rect 9478 -15314 9512 -15313
rect 8986 -15401 9000 -15349
rect 9052 -15401 9254 -15349
rect 8986 -15406 9254 -15401
rect 9293 -15434 9441 -15349
rect 8986 -15440 9441 -15434
rect 8986 -15493 8989 -15440
rect 9042 -15493 9441 -15440
rect 8986 -15500 9441 -15493
rect 9545 -15528 9611 -15312
rect 8050 -15971 8116 -15965
rect 8162 -15634 8361 -15622
rect 8162 -15646 8320 -15634
rect 7790 -16118 7872 -16052
rect 7938 -16118 8000 -16052
rect 7790 -16410 8000 -16118
rect 7750 -16422 8000 -16410
rect 8162 -16397 8246 -15646
rect 8281 -16397 8320 -15646
rect 8354 -16410 8361 -15634
rect 7102 -17221 7168 -17215
rect 7102 -17378 7168 -17287
rect 7214 -17326 7298 -16575
rect 7333 -17326 7372 -16575
rect 7214 -17338 7372 -17326
rect 7406 -17338 7413 -16562
rect 7214 -17350 7413 -17338
rect 7750 -16562 8000 -16550
rect 7750 -17338 7756 -16562
rect 7790 -16845 8000 -16562
rect 7790 -16911 7853 -16845
rect 7919 -16911 8000 -16845
rect 7790 -17335 8000 -16911
rect 8340 -16562 8361 -16410
rect 8698 -15634 8949 -15622
rect 8698 -16410 8704 -15634
rect 8738 -15637 8949 -15634
rect 8986 -15593 9611 -15528
rect 8738 -15798 8948 -15637
rect 9052 -15594 9611 -15593
rect 9775 -15550 9885 -15215
rect 10706 -15246 10816 -15215
rect 9917 -15251 10063 -15246
rect 9917 -15303 9933 -15251
rect 9986 -15262 10063 -15251
rect 9986 -15296 10013 -15262
rect 10047 -15296 10063 -15262
rect 9986 -15303 10063 -15296
rect 9917 -15312 10063 -15303
rect 10119 -15262 10256 -15246
rect 10119 -15296 10205 -15262
rect 10239 -15296 10256 -15262
rect 10119 -15312 10256 -15296
rect 10306 -15262 10447 -15247
rect 10306 -15296 10397 -15262
rect 10431 -15296 10447 -15262
rect 10119 -15340 10185 -15312
rect 9917 -15349 10185 -15340
rect 10306 -15313 10447 -15296
rect 10476 -15262 10640 -15246
rect 10476 -15296 10589 -15262
rect 10623 -15296 10640 -15262
rect 10476 -15312 10640 -15296
rect 10706 -15262 10990 -15246
rect 10706 -15296 10940 -15262
rect 10974 -15296 10990 -15262
rect 10706 -15312 10990 -15296
rect 11046 -15262 11183 -15246
rect 11046 -15296 11132 -15262
rect 11166 -15296 11183 -15262
rect 11046 -15312 11183 -15296
rect 11233 -15262 11374 -15247
rect 11233 -15296 11324 -15262
rect 11358 -15296 11374 -15262
rect 10306 -15349 10372 -15313
rect 10409 -15314 10443 -15313
rect 9917 -15401 9935 -15349
rect 9987 -15401 10185 -15349
rect 9917 -15406 10185 -15401
rect 10224 -15396 10372 -15349
rect 10224 -15434 10262 -15396
rect 9917 -15465 10262 -15434
rect 10331 -15465 10372 -15396
rect 9917 -15500 10372 -15465
rect 10476 -15528 10542 -15312
rect 9775 -15616 9798 -15550
rect 9864 -15616 9885 -15550
rect 9775 -15622 9885 -15616
rect 8986 -15677 9052 -15659
rect 9098 -15634 9297 -15622
rect 9098 -15646 9256 -15634
rect 8738 -15864 8818 -15798
rect 8884 -15864 8948 -15798
rect 8738 -16410 8948 -15864
rect 8698 -16422 8948 -16410
rect 9098 -16397 9182 -15646
rect 9217 -16397 9256 -15646
rect 9290 -16410 9297 -15634
rect 8162 -17326 8246 -16575
rect 8281 -17326 8320 -16575
rect 7790 -17338 8001 -17335
rect 7750 -17350 8001 -17338
rect 7102 -17444 7727 -17378
rect 6774 -17532 6780 -17463
rect 6849 -17472 6855 -17463
rect 6849 -17532 7557 -17472
rect 6780 -17538 7557 -17532
rect 5998 -17630 6066 -17566
rect 5999 -17632 6066 -17630
rect 6132 -17632 7370 -17566
rect 7409 -17623 7557 -17538
rect 7304 -17660 7370 -17632
rect 7491 -17659 7557 -17623
rect 7594 -17659 7628 -17658
rect 5832 -17726 6941 -17660
rect 7007 -17676 7248 -17660
rect 7007 -17710 7198 -17676
rect 7232 -17710 7248 -17676
rect 7007 -17726 7248 -17710
rect 7304 -17676 7441 -17660
rect 7304 -17710 7390 -17676
rect 7424 -17710 7441 -17676
rect 7304 -17726 7441 -17710
rect 7491 -17676 7632 -17659
rect 7491 -17710 7582 -17676
rect 7616 -17710 7632 -17676
rect 7491 -17725 7632 -17710
rect 7661 -17660 7727 -17444
rect 7661 -17676 7825 -17660
rect 7661 -17710 7774 -17676
rect 7808 -17710 7825 -17676
rect 7661 -17726 7825 -17710
rect 5832 -17736 5901 -17726
rect 7891 -17757 8001 -17350
rect 8050 -17342 8116 -17336
rect 8162 -17338 8320 -17326
rect 8354 -17338 8361 -16562
rect 8162 -17350 8361 -17338
rect 8698 -16562 8948 -16550
rect 8698 -17338 8704 -16562
rect 8738 -17255 8948 -16562
rect 9276 -16562 9297 -16410
rect 9634 -15634 9885 -15622
rect 9634 -16410 9640 -15634
rect 9674 -15637 9885 -15634
rect 9917 -15594 10542 -15528
rect 9674 -16410 9884 -15637
rect 9917 -15689 9983 -15594
rect 10706 -15622 10816 -15312
rect 11046 -15340 11112 -15312
rect 10844 -15406 10860 -15340
rect 10926 -15406 11112 -15340
rect 11233 -15313 11374 -15296
rect 11403 -15262 11567 -15246
rect 11403 -15296 11516 -15262
rect 11550 -15296 11567 -15262
rect 11403 -15312 11567 -15296
rect 11233 -15349 11299 -15313
rect 11336 -15314 11370 -15313
rect 11151 -15434 11299 -15349
rect 10844 -15500 10858 -15434
rect 10924 -15500 11299 -15434
rect 11403 -15528 11469 -15312
rect 10844 -15594 10850 -15528
rect 10915 -15594 11469 -15528
rect 11633 -15622 11743 -15215
rect 9917 -15761 9983 -15755
rect 10029 -15634 10228 -15622
rect 10029 -15646 10187 -15634
rect 9634 -16422 9884 -16410
rect 10029 -16397 10113 -15646
rect 10148 -16397 10187 -15646
rect 10221 -16410 10228 -15634
rect 8738 -17321 8837 -17255
rect 8903 -17321 8948 -17255
rect 8738 -17335 8948 -17321
rect 8989 -17001 9055 -16995
rect 8738 -17338 8949 -17335
rect 8698 -17350 8949 -17338
rect 8116 -17408 8675 -17378
rect 8050 -17444 8675 -17408
rect 8050 -17479 8505 -17472
rect 8050 -17538 8401 -17479
rect 8357 -17543 8401 -17538
rect 8465 -17543 8505 -17479
rect 8050 -17575 8318 -17566
rect 8050 -17627 8079 -17575
rect 8131 -17627 8318 -17575
rect 8357 -17623 8505 -17543
rect 8050 -17632 8318 -17627
rect 8252 -17660 8318 -17632
rect 8439 -17659 8505 -17623
rect 8542 -17659 8576 -17658
rect 8050 -17669 8196 -17660
rect 8050 -17721 8063 -17669
rect 8128 -17676 8196 -17669
rect 8128 -17710 8146 -17676
rect 8180 -17710 8196 -17676
rect 8128 -17721 8196 -17710
rect 8050 -17726 8196 -17721
rect 8252 -17676 8389 -17660
rect 8252 -17710 8338 -17676
rect 8372 -17710 8389 -17676
rect 8252 -17726 8389 -17710
rect 8439 -17676 8580 -17659
rect 8439 -17710 8530 -17676
rect 8564 -17710 8580 -17676
rect 8439 -17725 8580 -17710
rect 8609 -17660 8675 -17444
rect 8609 -17676 8773 -17660
rect 8609 -17710 8722 -17676
rect 8756 -17710 8773 -17676
rect 8609 -17726 8773 -17710
rect 8839 -17757 8949 -17350
rect 8989 -17378 9055 -17067
rect 9098 -17326 9182 -16575
rect 9217 -17326 9256 -16575
rect 9098 -17338 9256 -17326
rect 9290 -17338 9297 -16562
rect 9098 -17350 9297 -17338
rect 9634 -16562 9884 -16550
rect 9634 -17338 9640 -16562
rect 9674 -17335 9884 -16562
rect 10206 -16561 10228 -16410
rect 10565 -15634 10816 -15622
rect 10565 -16410 10571 -15634
rect 10605 -15637 10816 -15634
rect 10956 -15634 11155 -15622
rect 10605 -16410 10815 -15637
rect 10565 -16422 10815 -16410
rect 10956 -15646 11114 -15634
rect 10956 -16397 11040 -15646
rect 11075 -16397 11114 -15646
rect 11148 -16410 11155 -15634
rect 9917 -17123 9983 -17117
rect 9674 -17338 9885 -17335
rect 9634 -17349 9885 -17338
rect 9634 -17350 9807 -17349
rect 8986 -17444 9611 -17378
rect 8986 -17538 8993 -17472
rect 9059 -17538 9441 -17472
rect 8986 -17632 9001 -17566
rect 9067 -17632 9254 -17566
rect 9293 -17623 9441 -17538
rect 9188 -17660 9254 -17632
rect 9375 -17659 9441 -17623
rect 9478 -17659 9512 -17658
rect 8986 -17669 9132 -17660
rect 8986 -17721 8992 -17669
rect 9057 -17676 9132 -17669
rect 9057 -17710 9082 -17676
rect 9116 -17710 9132 -17676
rect 9057 -17721 9132 -17710
rect 8986 -17726 9132 -17721
rect 9188 -17676 9325 -17660
rect 9188 -17710 9274 -17676
rect 9308 -17710 9325 -17676
rect 9188 -17726 9325 -17710
rect 9375 -17676 9516 -17659
rect 9375 -17710 9466 -17676
rect 9500 -17710 9516 -17676
rect 9375 -17725 9516 -17710
rect 9545 -17660 9611 -17444
rect 9775 -17413 9807 -17350
rect 9873 -17413 9885 -17349
rect 9545 -17676 9709 -17660
rect 9545 -17710 9658 -17676
rect 9692 -17710 9709 -17676
rect 9545 -17726 9709 -17710
rect 9775 -17757 9885 -17413
rect 9917 -17377 9983 -17189
rect 10029 -17325 10113 -16574
rect 10148 -17325 10187 -16574
rect 10029 -17337 10187 -17325
rect 10221 -17337 10228 -16561
rect 10029 -17349 10228 -17337
rect 10565 -16561 10815 -16549
rect 10565 -17337 10571 -16561
rect 10605 -17334 10815 -16561
rect 11134 -16562 11155 -16410
rect 11492 -15634 11743 -15622
rect 11492 -16410 11498 -15634
rect 11532 -15637 11743 -15634
rect 11860 -15251 13092 -15027
rect 11860 -15454 12189 -15251
rect 12410 -15454 13092 -15251
rect 11532 -16393 11742 -15637
rect 11860 -15952 13092 -15454
rect 11799 -15960 13092 -15952
rect 11799 -16011 11811 -15960
rect 12168 -15969 13092 -15960
rect 12168 -16011 12180 -15969
rect 11799 -16018 12180 -16011
rect 11860 -16056 11903 -16018
rect 12726 -16103 13092 -15969
rect 11875 -16115 12689 -16103
rect 12726 -16110 13137 -16103
rect 11875 -16205 11881 -16115
rect 11915 -16205 12073 -16115
rect 12107 -16205 12265 -16115
rect 12299 -16205 12457 -16115
rect 12491 -16205 12649 -16115
rect 12683 -16205 12689 -16115
rect 11875 -16217 12689 -16205
rect 12923 -16147 13137 -16110
rect 12923 -16181 12986 -16147
rect 13077 -16181 13137 -16147
rect 12923 -16219 13137 -16181
rect 11779 -16257 12209 -16245
rect 11779 -16347 11785 -16257
rect 11819 -16347 11977 -16257
rect 12011 -16347 12169 -16257
rect 12203 -16347 12209 -16257
rect 11779 -16359 12209 -16347
rect 12355 -16251 12827 -16245
rect 12355 -16257 12892 -16251
rect 12355 -16347 12361 -16257
rect 12395 -16347 12553 -16257
rect 12587 -16347 12745 -16257
rect 12779 -16267 12892 -16257
rect 12779 -16347 12842 -16267
rect 12355 -16359 12842 -16347
rect 11532 -16409 12263 -16393
rect 11532 -16410 12170 -16409
rect 11492 -16422 12170 -16410
rect 11737 -16443 12170 -16422
rect 12204 -16443 12263 -16409
rect 11737 -16459 12263 -16443
rect 12702 -16493 12842 -16359
rect 12876 -16493 12892 -16267
rect 12923 -16253 12929 -16219
rect 13008 -16223 13137 -16219
rect 13008 -16253 13014 -16223
rect 12923 -16411 13014 -16253
rect 12923 -16445 12929 -16411
rect 13008 -16445 13014 -16411
rect 12923 -16461 13014 -16445
rect 13046 -16315 13235 -16251
rect 13046 -16349 13052 -16315
rect 13129 -16349 13235 -16315
rect 11703 -16514 12363 -16498
rect 11703 -16548 12313 -16514
rect 12347 -16548 12363 -16514
rect 11703 -16550 12363 -16548
rect 10956 -17326 11040 -16575
rect 11075 -17326 11114 -16575
rect 10605 -17337 10816 -17334
rect 10565 -17349 10816 -17337
rect 9917 -17443 10542 -17377
rect 9917 -17479 10372 -17471
rect 9917 -17537 10264 -17479
rect 10224 -17539 10264 -17537
rect 10324 -17539 10372 -17479
rect 9917 -17631 9937 -17565
rect 10003 -17631 10185 -17565
rect 10224 -17622 10372 -17539
rect 10119 -17659 10185 -17631
rect 10306 -17658 10372 -17622
rect 10409 -17658 10443 -17657
rect 9917 -17669 10063 -17659
rect 9917 -17721 9951 -17669
rect 10016 -17675 10063 -17669
rect 10047 -17709 10063 -17675
rect 10016 -17721 10063 -17709
rect 9917 -17725 10063 -17721
rect 10119 -17675 10256 -17659
rect 10119 -17709 10205 -17675
rect 10239 -17709 10256 -17675
rect 10119 -17725 10256 -17709
rect 10306 -17675 10447 -17658
rect 10306 -17709 10397 -17675
rect 10431 -17709 10447 -17675
rect 10306 -17724 10447 -17709
rect 10476 -17659 10542 -17443
rect 10476 -17675 10640 -17659
rect 10476 -17709 10589 -17675
rect 10623 -17709 10640 -17675
rect 10476 -17725 10640 -17709
rect 10706 -17660 10816 -17349
rect 10956 -17338 11114 -17326
rect 11148 -17338 11155 -16562
rect 10956 -17350 11155 -17338
rect 11492 -16562 12363 -16550
rect 11492 -17338 11498 -16562
rect 11532 -16564 12363 -16562
rect 11532 -16595 11815 -16564
rect 11532 -17335 11742 -16595
rect 12259 -16598 12305 -16592
rect 12702 -16598 12892 -16493
rect 13046 -16507 13235 -16349
rect 12259 -16604 12892 -16598
rect 12259 -16780 12265 -16604
rect 12299 -16713 12892 -16604
rect 12923 -16541 13052 -16507
rect 13129 -16518 13235 -16507
rect 13129 -16541 15223 -16518
rect 12923 -16584 15223 -16541
rect 12923 -16669 13235 -16584
rect 12923 -16703 12935 -16669
rect 13111 -16703 13235 -16669
rect 12923 -16709 13123 -16703
rect 12299 -16747 12842 -16713
rect 12876 -16747 12892 -16713
rect 12299 -16764 12892 -16747
rect 12923 -16757 13123 -16750
rect 12299 -16780 12827 -16764
rect 12259 -16792 12827 -16780
rect 12305 -16796 12827 -16792
rect 12923 -16791 12935 -16757
rect 13111 -16791 13123 -16757
rect 13151 -16764 13235 -16703
rect 12305 -16797 12825 -16796
rect 12305 -16798 12774 -16797
rect 12171 -16863 12394 -16856
rect 12171 -16911 12183 -16863
rect 12074 -16924 12183 -16911
rect 12382 -16911 12394 -16863
rect 12923 -16859 13123 -16791
rect 12923 -16893 12954 -16859
rect 13086 -16893 13123 -16859
rect 12921 -16900 13123 -16893
rect 12382 -16924 12473 -16911
rect 12074 -17027 12233 -16924
rect 12352 -17027 12473 -16924
rect 12921 -16949 13121 -16900
rect 12921 -16971 12960 -16949
rect 12074 -17101 12473 -17027
rect 12923 -17068 12960 -16971
rect 13079 -16971 13121 -16949
rect 13079 -17068 13113 -16971
rect 12923 -17126 13113 -17068
rect 11532 -17338 11743 -17335
rect 11492 -17350 11743 -17338
rect 10844 -17444 10850 -17378
rect 10916 -17444 11469 -17378
rect 10844 -17538 10888 -17472
rect 10954 -17538 11299 -17472
rect 10844 -17632 10859 -17566
rect 10925 -17632 11112 -17566
rect 11151 -17623 11299 -17538
rect 11046 -17660 11112 -17632
rect 11233 -17659 11299 -17623
rect 11336 -17659 11370 -17658
rect 10706 -17676 10990 -17660
rect 10706 -17710 10940 -17676
rect 10974 -17710 10990 -17676
rect 10706 -17726 10990 -17710
rect 11046 -17676 11183 -17660
rect 11046 -17710 11132 -17676
rect 11166 -17710 11183 -17676
rect 11046 -17726 11183 -17710
rect 11233 -17676 11374 -17659
rect 11233 -17710 11324 -17676
rect 11358 -17710 11374 -17676
rect 11233 -17725 11374 -17710
rect 11403 -17660 11469 -17444
rect 11403 -17676 11567 -17660
rect 11403 -17710 11516 -17676
rect 11550 -17710 11567 -17676
rect 11403 -17726 11567 -17710
rect 10706 -17756 10816 -17726
rect 7138 -17764 8001 -17757
rect 7138 -17876 7245 -17764
rect 7280 -17876 7438 -17764
rect 7473 -17876 7630 -17764
rect 7665 -17876 7822 -17764
rect 7857 -17876 8001 -17764
rect 7138 -17891 8001 -17876
rect 8086 -17764 8949 -17757
rect 8086 -17876 8193 -17764
rect 8228 -17876 8386 -17764
rect 8421 -17876 8578 -17764
rect 8613 -17876 8770 -17764
rect 8805 -17876 8949 -17764
rect 8086 -17891 8949 -17876
rect 9022 -17764 9885 -17757
rect 9022 -17876 9129 -17764
rect 9164 -17876 9322 -17764
rect 9357 -17876 9514 -17764
rect 9549 -17876 9706 -17764
rect 9741 -17876 9885 -17764
rect 9022 -17891 9885 -17876
rect 9953 -17763 10816 -17756
rect 11633 -17757 11743 -17350
rect 15157 -17570 15223 -16584
rect 15369 -17476 15435 -12012
rect 15481 -17382 15547 -7481
rect 15617 -17288 15683 -3000
rect 16145 -16814 16285 -16737
rect 16145 -16927 16211 -16814
rect 16145 -16995 16285 -16927
rect 16543 -16995 16590 -16737
rect 16249 -17061 16990 -17049
rect 16249 -17237 16255 -17061
rect 16289 -17237 16447 -17061
rect 16481 -17237 16990 -17061
rect 16249 -17249 16990 -17237
rect 15617 -17304 16719 -17288
rect 15617 -17338 16669 -17304
rect 16703 -17338 16719 -17304
rect 15617 -17354 16719 -17338
rect 15481 -17448 16244 -17382
rect 16177 -17476 16244 -17448
rect 15369 -17542 16144 -17476
rect 16177 -17542 16467 -17476
rect 16078 -17570 16144 -17542
rect 15157 -17586 16047 -17570
rect 15157 -17620 15997 -17586
rect 16031 -17620 16047 -17586
rect 15157 -17636 16047 -17620
rect 16078 -17586 16335 -17570
rect 16078 -17620 16285 -17586
rect 16319 -17620 16335 -17586
rect 16078 -17636 16335 -17620
rect 16401 -17586 16467 -17542
rect 16401 -17620 16417 -17586
rect 16451 -17620 16467 -17586
rect 16401 -17636 16467 -17620
rect 16830 -17569 16990 -17249
rect 16830 -17667 17258 -17569
rect 9953 -17875 10060 -17763
rect 10095 -17875 10253 -17763
rect 10288 -17875 10445 -17763
rect 10480 -17875 10637 -17763
rect 10672 -17875 10816 -17763
rect 9953 -17890 10816 -17875
rect 10880 -17764 11743 -17757
rect 10880 -17876 10987 -17764
rect 11022 -17876 11180 -17764
rect 11215 -17876 11372 -17764
rect 11407 -17876 11564 -17764
rect 11599 -17876 11743 -17764
rect 10880 -17891 11743 -17876
rect 15617 -17679 16007 -17667
rect 7137 -17953 10779 -17944
rect 11883 -17945 12147 -17934
rect 7137 -17954 9965 -17953
rect 4838 -18027 5471 -17961
rect 4745 -21389 4811 -21383
rect 4811 -21455 5319 -21389
rect 4745 -21461 4811 -21455
rect 5253 -24739 5319 -21455
rect 5405 -24649 5471 -18027
rect 7137 -18064 7150 -17954
rect 7184 -18064 7342 -17954
rect 7376 -18064 7534 -17954
rect 7568 -18064 7726 -17954
rect 7760 -18064 7918 -17954
rect 7952 -18064 8098 -17954
rect 8132 -18064 8290 -17954
rect 8324 -18064 8482 -17954
rect 8516 -18064 8674 -17954
rect 8708 -18064 8866 -17954
rect 8900 -18064 9034 -17954
rect 9068 -18064 9226 -17954
rect 9260 -18064 9418 -17954
rect 9452 -18064 9610 -17954
rect 9644 -18064 9802 -17954
rect 9836 -18063 9965 -17954
rect 9999 -18063 10157 -17953
rect 10191 -18063 10349 -17953
rect 10383 -18063 10541 -17953
rect 10575 -18063 10733 -17953
rect 10767 -18063 10779 -17953
rect 9836 -18064 10779 -18063
rect 7137 -18135 10779 -18064
rect 10880 -17954 11894 -17945
rect 10880 -18064 10892 -17954
rect 10926 -18064 11084 -17954
rect 11118 -18064 11276 -17954
rect 11310 -18064 11468 -17954
rect 11502 -18064 11660 -17954
rect 11694 -18064 11894 -17954
rect 10880 -18075 11894 -18064
rect 7137 -18136 10204 -18135
rect 7137 -18171 7389 -18136
rect 7677 -18171 8337 -18136
rect 8625 -18171 9273 -18136
rect 9561 -18170 10204 -18136
rect 10492 -18170 10779 -18135
rect 9561 -18171 10779 -18170
rect 7137 -18185 10779 -18171
rect 7137 -18187 7964 -18185
rect 8085 -18187 8912 -18185
rect 9021 -18187 9848 -18185
rect 9952 -18186 10779 -18185
rect 10879 -18136 11894 -18075
rect 10879 -18171 11131 -18136
rect 11419 -18171 11894 -18136
rect 10879 -18187 11894 -18171
rect 12136 -18187 12147 -17945
rect 11883 -18198 12147 -18187
rect 15617 -18033 15703 -17679
rect 15737 -18033 15775 -17679
rect 15809 -18033 15967 -17679
rect 16001 -18033 16007 -17679
rect 15617 -18045 16007 -18033
rect 16153 -17679 16583 -17667
rect 16153 -18033 16159 -17679
rect 16193 -18033 16351 -17679
rect 16385 -18033 16543 -17679
rect 16577 -18033 16583 -17679
rect 16153 -18045 16583 -18033
rect 16729 -17679 17258 -17667
rect 16729 -18033 16735 -17679
rect 16769 -18033 16927 -17679
rect 16961 -18033 17258 -17679
rect 16729 -18045 17258 -18033
rect 15617 -18501 15763 -18045
rect 16941 -18046 17258 -18045
rect 15538 -18514 15763 -18501
rect 5658 -18657 7357 -18613
rect 5658 -18691 5721 -18657
rect 5812 -18691 6161 -18657
rect 6252 -18691 6601 -18657
rect 6692 -18691 7357 -18657
rect 15538 -18658 15551 -18514
rect 15695 -18658 15763 -18514
rect 15865 -18155 16295 -18143
rect 15865 -18511 15871 -18155
rect 15905 -18511 16063 -18155
rect 16097 -18511 16255 -18155
rect 16289 -18511 16295 -18155
rect 15865 -18523 16295 -18511
rect 16441 -18155 16871 -18143
rect 16441 -18511 16447 -18155
rect 16481 -18511 16639 -18155
rect 16673 -18511 16831 -18155
rect 16865 -18511 16871 -18155
rect 16441 -18523 16871 -18511
rect 17192 -18518 17258 -18046
rect 17515 -18021 17672 -18008
rect 17515 -18154 17526 -18021
rect 17659 -18148 17672 -18021
rect 18096 -18148 18310 -18143
rect 17659 -18154 18377 -18148
rect 17515 -18155 18377 -18154
rect 17293 -18162 18377 -18155
rect 17293 -18209 17322 -18162
rect 17891 -18187 18377 -18162
rect 17891 -18209 18159 -18187
rect 17293 -18221 18159 -18209
rect 18250 -18221 18377 -18187
rect 17293 -18247 18377 -18221
rect 17293 -18275 17927 -18247
rect 18096 -18259 18310 -18247
rect 17293 -18281 17928 -18275
rect 17293 -18361 17306 -18281
rect 17340 -18361 17498 -18281
rect 17532 -18361 17690 -18281
rect 17724 -18361 17882 -18281
rect 17916 -18361 17928 -18281
rect 17293 -18367 17928 -18361
rect 17996 -18307 18065 -18291
rect 17293 -18368 17927 -18367
rect 17996 -18397 18015 -18307
rect 17386 -18403 18015 -18397
rect 17386 -18483 17402 -18403
rect 17436 -18483 17594 -18403
rect 17628 -18483 17786 -18403
rect 17820 -18483 18015 -18403
rect 17386 -18489 18015 -18483
rect 17192 -18536 17422 -18518
rect 17192 -18571 17372 -18536
rect 17406 -18571 17422 -18536
rect 15538 -18671 15763 -18658
rect 5658 -18703 7357 -18691
rect 5658 -18729 5872 -18703
rect 5558 -18761 5627 -18755
rect 5558 -19003 5577 -18830
rect 5611 -19003 5627 -18830
rect 5658 -18763 5664 -18729
rect 5743 -18733 5872 -18729
rect 6098 -18729 6312 -18703
rect 5743 -18763 5749 -18733
rect 5998 -18761 6067 -18755
rect 5658 -18921 5749 -18763
rect 5658 -18955 5664 -18921
rect 5743 -18955 5749 -18921
rect 5658 -18971 5749 -18955
rect 5781 -18825 5970 -18761
rect 5781 -18859 5787 -18825
rect 5864 -18859 5970 -18825
rect 5558 -19105 5627 -19003
rect 5781 -19017 5970 -18859
rect 5658 -19051 5787 -19017
rect 5864 -19051 5970 -19017
rect 5558 -19223 5628 -19105
rect 5658 -19179 5970 -19051
rect 5658 -19213 5670 -19179
rect 5846 -19213 5970 -19179
rect 5658 -19219 5858 -19213
rect 5558 -19257 5577 -19223
rect 5611 -19257 5628 -19223
rect 5558 -19274 5628 -19257
rect 5559 -19351 5628 -19274
rect 5558 -19410 5628 -19351
rect 5658 -19267 5858 -19260
rect 5658 -19301 5670 -19267
rect 5846 -19301 5858 -19267
rect 5886 -19274 5970 -19213
rect 5658 -19369 5858 -19301
rect 5658 -19403 5689 -19369
rect 5821 -19403 5858 -19369
rect 5658 -19410 5858 -19403
rect 5901 -19326 5970 -19274
rect 5559 -19526 5628 -19410
rect 5703 -19412 5823 -19410
rect 5703 -19464 5734 -19412
rect 5786 -19464 5823 -19412
rect 5901 -19416 5970 -19395
rect 5998 -19003 6017 -18830
rect 6051 -19003 6067 -18830
rect 6098 -18763 6104 -18729
rect 6183 -18733 6312 -18729
rect 6538 -18716 7357 -18703
rect 6538 -18729 6752 -18716
rect 6183 -18763 6189 -18733
rect 6438 -18761 6507 -18755
rect 6098 -18921 6189 -18763
rect 6098 -18955 6104 -18921
rect 6183 -18955 6189 -18921
rect 6098 -18971 6189 -18955
rect 6221 -18825 6410 -18761
rect 6221 -18859 6227 -18825
rect 6304 -18859 6410 -18825
rect 5998 -19223 6067 -19003
rect 6221 -19017 6410 -18859
rect 6098 -19051 6227 -19017
rect 6304 -19051 6410 -19017
rect 6098 -19179 6410 -19051
rect 6098 -19213 6110 -19179
rect 6286 -19213 6410 -19179
rect 6098 -19219 6298 -19213
rect 5998 -19257 6017 -19223
rect 6051 -19257 6067 -19223
rect 5703 -19495 5823 -19464
rect 5559 -19595 5901 -19526
rect 5559 -19607 5628 -19595
rect 5832 -22188 5901 -19595
rect 5998 -19859 6067 -19257
rect 6098 -19267 6298 -19260
rect 6098 -19301 6110 -19267
rect 6286 -19301 6298 -19267
rect 6326 -19274 6410 -19213
rect 6098 -19369 6298 -19301
rect 6098 -19403 6129 -19369
rect 6261 -19403 6298 -19369
rect 6098 -19410 6172 -19403
rect 6143 -19445 6172 -19410
rect 6224 -19410 6298 -19403
rect 6341 -19328 6410 -19274
rect 6341 -19410 6410 -19397
rect 6438 -19003 6457 -18830
rect 6491 -19003 6507 -18830
rect 6538 -18763 6544 -18729
rect 6623 -18733 6752 -18729
rect 6623 -18763 6629 -18733
rect 6538 -18921 6629 -18763
rect 6538 -18955 6544 -18921
rect 6623 -18955 6629 -18921
rect 6538 -18971 6629 -18955
rect 6661 -18825 6850 -18761
rect 6661 -18859 6667 -18825
rect 6744 -18859 6850 -18825
rect 6438 -19223 6507 -19003
rect 6661 -19017 6850 -18859
rect 6538 -19051 6667 -19017
rect 6744 -19051 6850 -19017
rect 6538 -19179 6850 -19051
rect 6538 -19213 6550 -19179
rect 6726 -19213 6850 -19179
rect 6538 -19219 6738 -19213
rect 6438 -19257 6457 -19223
rect 6491 -19257 6507 -19223
rect 6224 -19445 6263 -19410
rect 6143 -19470 6263 -19445
rect 5992 -19865 6073 -19859
rect 5992 -19934 5998 -19865
rect 6067 -19868 6073 -19865
rect 6067 -19934 6085 -19868
rect 5992 -19940 6073 -19934
rect 5998 -22094 6067 -19940
rect 6438 -20000 6507 -19257
rect 6538 -19267 6738 -19260
rect 6538 -19301 6550 -19267
rect 6726 -19301 6738 -19267
rect 6766 -19274 6850 -19213
rect 6538 -19369 6738 -19301
rect 6781 -19319 6850 -19274
rect 7254 -19313 7357 -18716
rect 15617 -19127 15763 -18671
rect 15865 -18661 16295 -18649
rect 15865 -19017 15871 -18661
rect 15905 -19017 16063 -18661
rect 16097 -19017 16255 -18661
rect 16289 -19017 16295 -18661
rect 15865 -19029 16295 -19017
rect 16441 -18661 16871 -18649
rect 17192 -18653 17422 -18571
rect 17450 -18536 17710 -18517
rect 17450 -18571 17661 -18536
rect 17695 -18571 17710 -18536
rect 17450 -18591 17710 -18571
rect 17786 -18533 18015 -18489
rect 18049 -18533 18065 -18307
rect 18096 -18293 18102 -18259
rect 18181 -18263 18310 -18259
rect 18181 -18293 18187 -18263
rect 18096 -18451 18187 -18293
rect 18096 -18485 18102 -18451
rect 18181 -18485 18187 -18451
rect 18096 -18501 18187 -18485
rect 18219 -18355 18408 -18291
rect 18219 -18389 18225 -18355
rect 18302 -18389 18408 -18355
rect 16441 -19017 16447 -18661
rect 16481 -19017 16639 -18661
rect 16673 -19017 16831 -18661
rect 16865 -19017 16871 -18661
rect 17450 -18660 17500 -18591
rect 17786 -18619 18065 -18533
rect 18219 -18547 18408 -18389
rect 17450 -18682 17456 -18660
rect 16441 -19029 16871 -19017
rect 17192 -18695 17456 -18682
rect 17490 -18695 17500 -18660
rect 17528 -18631 18065 -18619
rect 17528 -18665 17540 -18631
rect 17916 -18665 18065 -18631
rect 17528 -18671 18065 -18665
rect 17192 -18818 17500 -18695
rect 17996 -18753 18065 -18671
rect 18096 -18581 18225 -18547
rect 18302 -18581 18408 -18547
rect 18096 -18709 18408 -18581
rect 18096 -18743 18108 -18709
rect 18284 -18743 18408 -18709
rect 18096 -18749 18296 -18743
rect 17996 -18787 18015 -18753
rect 18049 -18787 18065 -18753
rect 17996 -18804 18065 -18787
rect 18096 -18797 18296 -18790
rect 15617 -19139 16007 -19127
rect 11860 -19313 12409 -19312
rect 12750 -19313 13092 -19312
rect 6538 -19403 6569 -19369
rect 6701 -19403 6738 -19369
rect 6538 -19410 6612 -19403
rect 6580 -19436 6612 -19410
rect 6664 -19410 6738 -19403
rect 6780 -19350 6850 -19319
rect 7137 -19314 7964 -19313
rect 8085 -19314 8912 -19313
rect 9021 -19314 9848 -19313
rect 9952 -19314 10779 -19313
rect 7137 -19329 10780 -19314
rect 6664 -19436 6700 -19410
rect 6580 -19479 6700 -19436
rect 6438 -20075 6507 -20069
rect 6780 -19962 6849 -19350
rect 7137 -19364 7389 -19329
rect 7677 -19364 8337 -19329
rect 8625 -19364 9273 -19329
rect 9561 -19364 10204 -19329
rect 10492 -19364 10780 -19329
rect 7137 -19425 10780 -19364
rect 10879 -19329 13092 -19313
rect 10879 -19364 11131 -19329
rect 11419 -19364 13092 -19329
rect 10879 -19425 13092 -19364
rect 7138 -19436 10780 -19425
rect 7138 -19546 7150 -19436
rect 7184 -19546 7342 -19436
rect 7376 -19546 7534 -19436
rect 7568 -19546 7726 -19436
rect 7760 -19546 7918 -19436
rect 7952 -19546 8098 -19436
rect 8132 -19546 8290 -19436
rect 8324 -19546 8482 -19436
rect 8516 -19546 8674 -19436
rect 8708 -19546 8866 -19436
rect 8900 -19546 9034 -19436
rect 9068 -19546 9226 -19436
rect 9260 -19546 9418 -19436
rect 9452 -19546 9610 -19436
rect 9644 -19546 9802 -19436
rect 9836 -19546 9965 -19436
rect 9999 -19546 10157 -19436
rect 10191 -19546 10349 -19436
rect 10383 -19546 10541 -19436
rect 10575 -19546 10733 -19436
rect 10767 -19546 10780 -19436
rect 7138 -19555 10780 -19546
rect 10880 -19436 13092 -19425
rect 10880 -19546 10892 -19436
rect 10926 -19546 11084 -19436
rect 11118 -19546 11276 -19436
rect 11310 -19546 11468 -19436
rect 11502 -19546 11660 -19436
rect 11694 -19546 13092 -19436
rect 15617 -19493 15703 -19139
rect 15737 -19493 15775 -19139
rect 15809 -19493 15967 -19139
rect 16001 -19493 16007 -19139
rect 15617 -19505 16007 -19493
rect 16153 -19139 16583 -19127
rect 16153 -19493 16159 -19139
rect 16193 -19493 16351 -19139
rect 16385 -19493 16543 -19139
rect 16577 -19493 16583 -19139
rect 16153 -19505 16583 -19493
rect 16729 -19128 16967 -19127
rect 17192 -19128 17258 -18818
rect 17528 -18823 17928 -18817
rect 17528 -18857 17540 -18823
rect 17916 -18857 17928 -18823
rect 17528 -18869 17928 -18857
rect 18096 -18831 18108 -18797
rect 18284 -18831 18296 -18797
rect 18324 -18804 18408 -18743
rect 18096 -18869 18296 -18831
rect 17528 -18895 17977 -18869
rect 17528 -18929 17555 -18895
rect 17890 -18929 17977 -18895
rect 17528 -18940 17977 -18929
rect 18048 -18899 18296 -18869
rect 18048 -18933 18127 -18899
rect 18259 -18933 18296 -18899
rect 18048 -18940 18296 -18933
rect 16729 -19139 17258 -19128
rect 16729 -19493 16735 -19139
rect 16769 -19493 16927 -19139
rect 16961 -19493 17258 -19139
rect 16729 -19505 17258 -19493
rect 15617 -19506 15763 -19505
rect 10880 -19555 13092 -19546
rect 7138 -19624 8001 -19609
rect 7138 -19736 7245 -19624
rect 7280 -19736 7438 -19624
rect 7473 -19736 7630 -19624
rect 7665 -19736 7822 -19624
rect 7857 -19736 8001 -19624
rect 7138 -19743 8001 -19736
rect 8086 -19624 8949 -19609
rect 8086 -19736 8193 -19624
rect 8228 -19736 8386 -19624
rect 8421 -19736 8578 -19624
rect 8613 -19736 8770 -19624
rect 8805 -19736 8949 -19624
rect 8086 -19743 8949 -19736
rect 9022 -19624 9885 -19609
rect 9022 -19736 9129 -19624
rect 9164 -19736 9322 -19624
rect 9357 -19736 9514 -19624
rect 9549 -19736 9706 -19624
rect 9741 -19736 9885 -19624
rect 9022 -19743 9885 -19736
rect 9953 -19624 10816 -19609
rect 9953 -19736 10060 -19624
rect 10095 -19736 10253 -19624
rect 10288 -19736 10445 -19624
rect 10480 -19736 10637 -19624
rect 10672 -19736 10816 -19624
rect 9953 -19743 10816 -19736
rect 10880 -19624 11743 -19609
rect 10880 -19736 10987 -19624
rect 11022 -19736 11180 -19624
rect 11215 -19736 11372 -19624
rect 11407 -19736 11564 -19624
rect 11599 -19736 11743 -19624
rect 10880 -19743 11743 -19736
rect 7106 -19774 7158 -19773
rect 7102 -19779 7248 -19774
rect 7102 -19831 7106 -19779
rect 7158 -19790 7248 -19779
rect 7158 -19824 7198 -19790
rect 7232 -19824 7248 -19790
rect 7158 -19831 7248 -19824
rect 7102 -19840 7248 -19831
rect 7304 -19790 7441 -19774
rect 7304 -19824 7390 -19790
rect 7424 -19824 7441 -19790
rect 7304 -19840 7441 -19824
rect 7491 -19790 7632 -19775
rect 7491 -19824 7582 -19790
rect 7616 -19824 7632 -19790
rect 7304 -19868 7370 -19840
rect 7097 -19873 7370 -19868
rect 7097 -19925 7113 -19873
rect 7165 -19925 7370 -19873
rect 7491 -19841 7632 -19824
rect 7661 -19790 7825 -19774
rect 7661 -19824 7774 -19790
rect 7808 -19824 7825 -19790
rect 7661 -19840 7825 -19824
rect 7491 -19877 7557 -19841
rect 7594 -19842 7628 -19841
rect 7097 -19934 7370 -19925
rect 7409 -19962 7557 -19877
rect 6780 -20028 7327 -19962
rect 7393 -20028 7557 -19962
rect 6780 -21991 6849 -20028
rect 7661 -20056 7727 -19840
rect 7102 -20122 7727 -20056
rect 7106 -20323 7172 -20122
rect 7891 -20150 8001 -19743
rect 8050 -19780 8196 -19774
rect 8050 -19832 8069 -19780
rect 8122 -19790 8196 -19780
rect 8122 -19824 8146 -19790
rect 8180 -19824 8196 -19790
rect 8122 -19832 8196 -19824
rect 8050 -19840 8196 -19832
rect 8252 -19790 8389 -19774
rect 8252 -19824 8338 -19790
rect 8372 -19824 8389 -19790
rect 8252 -19840 8389 -19824
rect 8439 -19790 8580 -19775
rect 8439 -19824 8530 -19790
rect 8564 -19824 8580 -19790
rect 8252 -19868 8318 -19840
rect 8050 -19872 8318 -19868
rect 8050 -19924 8057 -19872
rect 8109 -19924 8318 -19872
rect 8439 -19841 8580 -19824
rect 8609 -19790 8773 -19774
rect 8609 -19824 8722 -19790
rect 8756 -19824 8773 -19790
rect 8609 -19840 8773 -19824
rect 8439 -19877 8505 -19841
rect 8542 -19842 8576 -19841
rect 8050 -19934 8318 -19924
rect 8357 -19955 8505 -19877
rect 8357 -19962 8424 -19955
rect 8050 -20007 8424 -19962
rect 8493 -20007 8505 -19955
rect 8050 -20028 8505 -20007
rect 8609 -20056 8675 -19840
rect 7106 -20395 7172 -20389
rect 7214 -20162 7413 -20150
rect 7214 -20174 7372 -20162
rect 7214 -20925 7298 -20174
rect 7333 -20925 7372 -20174
rect 7214 -21103 7227 -20925
rect 7406 -20938 7413 -20162
rect 7405 -21090 7413 -20938
rect 7750 -20162 8001 -20150
rect 7750 -20938 7756 -20162
rect 7790 -20165 8001 -20162
rect 8050 -20122 8675 -20056
rect 7790 -20580 8000 -20165
rect 8050 -20427 8116 -20122
rect 8839 -20150 8949 -19743
rect 8986 -19779 9132 -19774
rect 8986 -19831 9002 -19779
rect 9055 -19790 9132 -19779
rect 9055 -19824 9082 -19790
rect 9116 -19824 9132 -19790
rect 9055 -19831 9132 -19824
rect 8986 -19840 9132 -19831
rect 9188 -19790 9325 -19774
rect 9188 -19824 9274 -19790
rect 9308 -19824 9325 -19790
rect 9188 -19840 9325 -19824
rect 9375 -19790 9516 -19775
rect 9375 -19824 9466 -19790
rect 9500 -19824 9516 -19790
rect 9188 -19868 9254 -19840
rect 8986 -19877 9254 -19868
rect 9375 -19841 9516 -19824
rect 9545 -19790 9709 -19774
rect 9545 -19824 9658 -19790
rect 9692 -19824 9709 -19790
rect 9545 -19840 9709 -19824
rect 9375 -19877 9441 -19841
rect 9478 -19842 9512 -19841
rect 8986 -19929 9000 -19877
rect 9052 -19929 9254 -19877
rect 8986 -19934 9254 -19929
rect 9293 -19962 9441 -19877
rect 8986 -19968 9441 -19962
rect 8986 -20021 8989 -19968
rect 9042 -20021 9441 -19968
rect 8986 -20028 9441 -20021
rect 9545 -20056 9611 -19840
rect 8050 -20499 8116 -20493
rect 8162 -20162 8361 -20150
rect 8162 -20174 8320 -20162
rect 7790 -20646 7872 -20580
rect 7938 -20646 8000 -20580
rect 7790 -20938 8000 -20646
rect 7750 -20950 8000 -20938
rect 8162 -20925 8246 -20174
rect 8281 -20925 8320 -20174
rect 8354 -20938 8361 -20162
rect 7102 -21749 7168 -21743
rect 7102 -21906 7168 -21815
rect 7214 -21854 7298 -21103
rect 7333 -21854 7372 -21103
rect 7214 -21866 7372 -21854
rect 7406 -21866 7413 -21090
rect 7214 -21878 7413 -21866
rect 7750 -21090 8000 -21078
rect 7750 -21866 7756 -21090
rect 7790 -21373 8000 -21090
rect 7790 -21439 7853 -21373
rect 7919 -21439 8000 -21373
rect 7790 -21863 8000 -21439
rect 8340 -21090 8361 -20938
rect 8698 -20162 8949 -20150
rect 8698 -20938 8704 -20162
rect 8738 -20165 8949 -20162
rect 8986 -20121 9611 -20056
rect 8738 -20326 8948 -20165
rect 9052 -20122 9611 -20121
rect 9775 -20078 9885 -19743
rect 10706 -19774 10816 -19743
rect 9917 -19779 10063 -19774
rect 9917 -19831 9933 -19779
rect 9986 -19790 10063 -19779
rect 9986 -19824 10013 -19790
rect 10047 -19824 10063 -19790
rect 9986 -19831 10063 -19824
rect 9917 -19840 10063 -19831
rect 10119 -19790 10256 -19774
rect 10119 -19824 10205 -19790
rect 10239 -19824 10256 -19790
rect 10119 -19840 10256 -19824
rect 10306 -19790 10447 -19775
rect 10306 -19824 10397 -19790
rect 10431 -19824 10447 -19790
rect 10119 -19868 10185 -19840
rect 9917 -19877 10185 -19868
rect 10306 -19841 10447 -19824
rect 10476 -19790 10640 -19774
rect 10476 -19824 10589 -19790
rect 10623 -19824 10640 -19790
rect 10476 -19840 10640 -19824
rect 10706 -19790 10990 -19774
rect 10706 -19824 10940 -19790
rect 10974 -19824 10990 -19790
rect 10706 -19840 10990 -19824
rect 11046 -19790 11183 -19774
rect 11046 -19824 11132 -19790
rect 11166 -19824 11183 -19790
rect 11046 -19840 11183 -19824
rect 11233 -19790 11374 -19775
rect 11233 -19824 11324 -19790
rect 11358 -19824 11374 -19790
rect 10306 -19877 10372 -19841
rect 10409 -19842 10443 -19841
rect 9917 -19929 9935 -19877
rect 9987 -19929 10185 -19877
rect 9917 -19934 10185 -19929
rect 10224 -19924 10372 -19877
rect 10224 -19962 10262 -19924
rect 9917 -19993 10262 -19962
rect 10331 -19993 10372 -19924
rect 9917 -20028 10372 -19993
rect 10476 -20056 10542 -19840
rect 9775 -20144 9798 -20078
rect 9864 -20144 9885 -20078
rect 9775 -20150 9885 -20144
rect 8986 -20205 9052 -20187
rect 9098 -20162 9297 -20150
rect 9098 -20174 9256 -20162
rect 8738 -20392 8818 -20326
rect 8884 -20392 8948 -20326
rect 8738 -20938 8948 -20392
rect 8698 -20950 8948 -20938
rect 9098 -20925 9182 -20174
rect 9217 -20925 9256 -20174
rect 9290 -20938 9297 -20162
rect 8162 -21854 8246 -21103
rect 8281 -21854 8320 -21103
rect 7790 -21866 8001 -21863
rect 7750 -21878 8001 -21866
rect 7102 -21972 7727 -21906
rect 6774 -22060 6780 -21991
rect 6849 -22000 6855 -21991
rect 6849 -22060 7557 -22000
rect 6780 -22066 7557 -22060
rect 5998 -22158 6066 -22094
rect 5999 -22160 6066 -22158
rect 6132 -22160 7370 -22094
rect 7409 -22151 7557 -22066
rect 7304 -22188 7370 -22160
rect 7491 -22187 7557 -22151
rect 7594 -22187 7628 -22186
rect 5832 -22254 6941 -22188
rect 7007 -22204 7248 -22188
rect 7007 -22238 7198 -22204
rect 7232 -22238 7248 -22204
rect 7007 -22254 7248 -22238
rect 7304 -22204 7441 -22188
rect 7304 -22238 7390 -22204
rect 7424 -22238 7441 -22204
rect 7304 -22254 7441 -22238
rect 7491 -22204 7632 -22187
rect 7491 -22238 7582 -22204
rect 7616 -22238 7632 -22204
rect 7491 -22253 7632 -22238
rect 7661 -22188 7727 -21972
rect 7661 -22204 7825 -22188
rect 7661 -22238 7774 -22204
rect 7808 -22238 7825 -22204
rect 7661 -22254 7825 -22238
rect 5832 -22264 5901 -22254
rect 7891 -22285 8001 -21878
rect 8050 -21870 8116 -21864
rect 8162 -21866 8320 -21854
rect 8354 -21866 8361 -21090
rect 8162 -21878 8361 -21866
rect 8698 -21090 8948 -21078
rect 8698 -21866 8704 -21090
rect 8738 -21783 8948 -21090
rect 9276 -21090 9297 -20938
rect 9634 -20162 9885 -20150
rect 9634 -20938 9640 -20162
rect 9674 -20165 9885 -20162
rect 9917 -20122 10542 -20056
rect 9674 -20938 9884 -20165
rect 9917 -20217 9983 -20122
rect 10706 -20150 10816 -19840
rect 11046 -19868 11112 -19840
rect 10844 -19934 10860 -19868
rect 10926 -19934 11112 -19868
rect 11233 -19841 11374 -19824
rect 11403 -19790 11567 -19774
rect 11403 -19824 11516 -19790
rect 11550 -19824 11567 -19790
rect 11403 -19840 11567 -19824
rect 11233 -19877 11299 -19841
rect 11336 -19842 11370 -19841
rect 11151 -19962 11299 -19877
rect 10844 -20028 10858 -19962
rect 10924 -20028 11299 -19962
rect 11403 -20056 11469 -19840
rect 10844 -20122 10850 -20056
rect 10915 -20122 11469 -20056
rect 11633 -20150 11743 -19743
rect 9917 -20289 9983 -20283
rect 10029 -20162 10228 -20150
rect 10029 -20174 10187 -20162
rect 9634 -20950 9884 -20938
rect 10029 -20925 10113 -20174
rect 10148 -20925 10187 -20174
rect 10221 -20938 10228 -20162
rect 8738 -21849 8837 -21783
rect 8903 -21849 8948 -21783
rect 8738 -21863 8948 -21849
rect 8989 -21529 9055 -21523
rect 8738 -21866 8949 -21863
rect 8698 -21878 8949 -21866
rect 8116 -21936 8675 -21906
rect 8050 -21972 8675 -21936
rect 8050 -22007 8505 -22000
rect 8050 -22066 8401 -22007
rect 8357 -22071 8401 -22066
rect 8465 -22071 8505 -22007
rect 8050 -22103 8318 -22094
rect 8050 -22155 8079 -22103
rect 8131 -22155 8318 -22103
rect 8357 -22151 8505 -22071
rect 8050 -22160 8318 -22155
rect 8252 -22188 8318 -22160
rect 8439 -22187 8505 -22151
rect 8542 -22187 8576 -22186
rect 8050 -22197 8196 -22188
rect 8050 -22249 8063 -22197
rect 8128 -22204 8196 -22197
rect 8128 -22238 8146 -22204
rect 8180 -22238 8196 -22204
rect 8128 -22249 8196 -22238
rect 8050 -22254 8196 -22249
rect 8252 -22204 8389 -22188
rect 8252 -22238 8338 -22204
rect 8372 -22238 8389 -22204
rect 8252 -22254 8389 -22238
rect 8439 -22204 8580 -22187
rect 8439 -22238 8530 -22204
rect 8564 -22238 8580 -22204
rect 8439 -22253 8580 -22238
rect 8609 -22188 8675 -21972
rect 8609 -22204 8773 -22188
rect 8609 -22238 8722 -22204
rect 8756 -22238 8773 -22204
rect 8609 -22254 8773 -22238
rect 8839 -22285 8949 -21878
rect 8989 -21906 9055 -21595
rect 9098 -21854 9182 -21103
rect 9217 -21854 9256 -21103
rect 9098 -21866 9256 -21854
rect 9290 -21866 9297 -21090
rect 9098 -21878 9297 -21866
rect 9634 -21090 9884 -21078
rect 9634 -21866 9640 -21090
rect 9674 -21863 9884 -21090
rect 10206 -21089 10228 -20938
rect 10565 -20162 10816 -20150
rect 10565 -20938 10571 -20162
rect 10605 -20165 10816 -20162
rect 10956 -20162 11155 -20150
rect 10605 -20938 10815 -20165
rect 10565 -20950 10815 -20938
rect 10956 -20174 11114 -20162
rect 10956 -20925 11040 -20174
rect 11075 -20925 11114 -20174
rect 11148 -20938 11155 -20162
rect 9917 -21651 9983 -21645
rect 9674 -21866 9885 -21863
rect 9634 -21877 9885 -21866
rect 9634 -21878 9807 -21877
rect 8986 -21972 9611 -21906
rect 8986 -22066 8993 -22000
rect 9059 -22066 9441 -22000
rect 8986 -22160 9001 -22094
rect 9067 -22160 9254 -22094
rect 9293 -22151 9441 -22066
rect 9188 -22188 9254 -22160
rect 9375 -22187 9441 -22151
rect 9478 -22187 9512 -22186
rect 8986 -22197 9132 -22188
rect 8986 -22249 8992 -22197
rect 9057 -22204 9132 -22197
rect 9057 -22238 9082 -22204
rect 9116 -22238 9132 -22204
rect 9057 -22249 9132 -22238
rect 8986 -22254 9132 -22249
rect 9188 -22204 9325 -22188
rect 9188 -22238 9274 -22204
rect 9308 -22238 9325 -22204
rect 9188 -22254 9325 -22238
rect 9375 -22204 9516 -22187
rect 9375 -22238 9466 -22204
rect 9500 -22238 9516 -22204
rect 9375 -22253 9516 -22238
rect 9545 -22188 9611 -21972
rect 9775 -21941 9807 -21878
rect 9873 -21941 9885 -21877
rect 9545 -22204 9709 -22188
rect 9545 -22238 9658 -22204
rect 9692 -22238 9709 -22204
rect 9545 -22254 9709 -22238
rect 9775 -22285 9885 -21941
rect 9917 -21905 9983 -21717
rect 10029 -21853 10113 -21102
rect 10148 -21853 10187 -21102
rect 10029 -21865 10187 -21853
rect 10221 -21865 10228 -21089
rect 10029 -21877 10228 -21865
rect 10565 -21089 10815 -21077
rect 10565 -21865 10571 -21089
rect 10605 -21862 10815 -21089
rect 11134 -21090 11155 -20938
rect 11492 -20162 11743 -20150
rect 11492 -20938 11498 -20162
rect 11532 -20165 11743 -20162
rect 11860 -19779 13092 -19555
rect 11860 -19982 12189 -19779
rect 12410 -19982 13092 -19779
rect 11532 -20921 11742 -20165
rect 11860 -20480 13092 -19982
rect 11799 -20488 13092 -20480
rect 11799 -20539 11811 -20488
rect 12168 -20497 13092 -20488
rect 12168 -20539 12180 -20497
rect 11799 -20546 12180 -20539
rect 11860 -20584 11903 -20546
rect 12726 -20631 13092 -20497
rect 15066 -19552 16047 -19536
rect 15066 -19586 15997 -19552
rect 16031 -19586 16047 -19552
rect 15066 -19602 16047 -19586
rect 16078 -19552 16335 -19536
rect 16078 -19586 16285 -19552
rect 16319 -19586 16335 -19552
rect 16078 -19602 16335 -19586
rect 16401 -19552 16467 -19536
rect 16401 -19586 16417 -19552
rect 16451 -19586 16467 -19552
rect 11875 -20643 12689 -20631
rect 12726 -20638 13137 -20631
rect 11875 -20733 11881 -20643
rect 11915 -20733 12073 -20643
rect 12107 -20733 12265 -20643
rect 12299 -20733 12457 -20643
rect 12491 -20733 12649 -20643
rect 12683 -20733 12689 -20643
rect 11875 -20745 12689 -20733
rect 12923 -20675 13137 -20638
rect 12923 -20709 12986 -20675
rect 13077 -20709 13137 -20675
rect 12923 -20747 13137 -20709
rect 11779 -20785 12209 -20773
rect 11779 -20875 11785 -20785
rect 11819 -20875 11977 -20785
rect 12011 -20875 12169 -20785
rect 12203 -20875 12209 -20785
rect 11779 -20887 12209 -20875
rect 12355 -20779 12827 -20773
rect 12355 -20785 12892 -20779
rect 12355 -20875 12361 -20785
rect 12395 -20875 12553 -20785
rect 12587 -20875 12745 -20785
rect 12779 -20795 12892 -20785
rect 12779 -20875 12842 -20795
rect 12355 -20887 12842 -20875
rect 11532 -20937 12263 -20921
rect 11532 -20938 12170 -20937
rect 11492 -20950 12170 -20938
rect 11737 -20971 12170 -20950
rect 12204 -20971 12263 -20937
rect 11737 -20987 12263 -20971
rect 12702 -21021 12842 -20887
rect 12876 -21021 12892 -20795
rect 12923 -20781 12929 -20747
rect 13008 -20751 13137 -20747
rect 13008 -20781 13014 -20751
rect 12923 -20939 13014 -20781
rect 12923 -20973 12929 -20939
rect 13008 -20973 13014 -20939
rect 12923 -20989 13014 -20973
rect 13046 -20843 13235 -20779
rect 13046 -20877 13052 -20843
rect 13129 -20877 13235 -20843
rect 11703 -21042 12363 -21026
rect 11703 -21076 12313 -21042
rect 12347 -21076 12363 -21042
rect 11703 -21078 12363 -21076
rect 10956 -21854 11040 -21103
rect 11075 -21854 11114 -21103
rect 10605 -21865 10816 -21862
rect 10565 -21877 10816 -21865
rect 9917 -21971 10542 -21905
rect 9917 -22007 10372 -21999
rect 9917 -22065 10264 -22007
rect 10224 -22067 10264 -22065
rect 10324 -22067 10372 -22007
rect 9917 -22159 9937 -22093
rect 10003 -22159 10185 -22093
rect 10224 -22150 10372 -22067
rect 10119 -22187 10185 -22159
rect 10306 -22186 10372 -22150
rect 10409 -22186 10443 -22185
rect 9917 -22197 10063 -22187
rect 9917 -22249 9951 -22197
rect 10016 -22203 10063 -22197
rect 10047 -22237 10063 -22203
rect 10016 -22249 10063 -22237
rect 9917 -22253 10063 -22249
rect 10119 -22203 10256 -22187
rect 10119 -22237 10205 -22203
rect 10239 -22237 10256 -22203
rect 10119 -22253 10256 -22237
rect 10306 -22203 10447 -22186
rect 10306 -22237 10397 -22203
rect 10431 -22237 10447 -22203
rect 10306 -22252 10447 -22237
rect 10476 -22187 10542 -21971
rect 10476 -22203 10640 -22187
rect 10476 -22237 10589 -22203
rect 10623 -22237 10640 -22203
rect 10476 -22253 10640 -22237
rect 10706 -22188 10816 -21877
rect 10956 -21866 11114 -21854
rect 11148 -21866 11155 -21090
rect 10956 -21878 11155 -21866
rect 11492 -21090 12363 -21078
rect 11492 -21866 11498 -21090
rect 11532 -21092 12363 -21090
rect 11532 -21123 11815 -21092
rect 11532 -21863 11742 -21123
rect 12259 -21126 12305 -21120
rect 12702 -21126 12892 -21021
rect 13046 -21035 13235 -20877
rect 12259 -21132 12892 -21126
rect 12259 -21308 12265 -21132
rect 12299 -21241 12892 -21132
rect 12923 -21069 13052 -21035
rect 13129 -21039 13235 -21035
rect 15066 -21039 15132 -19602
rect 16078 -19630 16144 -19602
rect 16401 -19630 16467 -19586
rect 13129 -21069 15132 -21039
rect 12923 -21105 15132 -21069
rect 15261 -19696 16144 -19630
rect 16177 -19696 16467 -19630
rect 16830 -19607 17258 -19505
rect 12923 -21197 13235 -21105
rect 12923 -21231 12935 -21197
rect 13111 -21231 13235 -21197
rect 12923 -21237 13123 -21231
rect 12299 -21275 12842 -21241
rect 12876 -21275 12892 -21241
rect 12299 -21292 12892 -21275
rect 12923 -21285 13123 -21278
rect 12299 -21308 12827 -21292
rect 12259 -21320 12827 -21308
rect 12305 -21324 12827 -21320
rect 12923 -21319 12935 -21285
rect 13111 -21319 13123 -21285
rect 13151 -21292 13235 -21231
rect 12305 -21325 12825 -21324
rect 12305 -21326 12774 -21325
rect 12171 -21391 12394 -21384
rect 12171 -21439 12183 -21391
rect 12074 -21452 12183 -21439
rect 12382 -21439 12394 -21391
rect 12923 -21387 13123 -21319
rect 12923 -21421 12954 -21387
rect 13086 -21421 13123 -21387
rect 12921 -21428 13123 -21421
rect 12382 -21452 12473 -21439
rect 12074 -21555 12233 -21452
rect 12352 -21555 12473 -21452
rect 12921 -21477 13121 -21428
rect 12921 -21499 12960 -21477
rect 12074 -21629 12473 -21555
rect 12923 -21596 12960 -21499
rect 13079 -21499 13121 -21477
rect 13079 -21596 13113 -21499
rect 12923 -21654 13113 -21596
rect 11532 -21866 11743 -21863
rect 11492 -21878 11743 -21866
rect 10844 -21972 10850 -21906
rect 10916 -21972 11469 -21906
rect 10844 -22066 10888 -22000
rect 10954 -22066 11299 -22000
rect 10844 -22160 10859 -22094
rect 10925 -22160 11112 -22094
rect 11151 -22151 11299 -22066
rect 11046 -22188 11112 -22160
rect 11233 -22187 11299 -22151
rect 11336 -22187 11370 -22186
rect 10706 -22204 10990 -22188
rect 10706 -22238 10940 -22204
rect 10974 -22238 10990 -22204
rect 10706 -22254 10990 -22238
rect 11046 -22204 11183 -22188
rect 11046 -22238 11132 -22204
rect 11166 -22238 11183 -22204
rect 11046 -22254 11183 -22238
rect 11233 -22204 11374 -22187
rect 11233 -22238 11324 -22204
rect 11358 -22238 11374 -22204
rect 11233 -22253 11374 -22238
rect 11403 -22188 11469 -21972
rect 11403 -22204 11567 -22188
rect 11403 -22238 11516 -22204
rect 11550 -22238 11567 -22204
rect 11403 -22254 11567 -22238
rect 10706 -22284 10816 -22254
rect 7138 -22292 8001 -22285
rect 7138 -22404 7245 -22292
rect 7280 -22404 7438 -22292
rect 7473 -22404 7630 -22292
rect 7665 -22404 7822 -22292
rect 7857 -22404 8001 -22292
rect 7138 -22419 8001 -22404
rect 8086 -22292 8949 -22285
rect 8086 -22404 8193 -22292
rect 8228 -22404 8386 -22292
rect 8421 -22404 8578 -22292
rect 8613 -22404 8770 -22292
rect 8805 -22404 8949 -22292
rect 8086 -22419 8949 -22404
rect 9022 -22292 9885 -22285
rect 9022 -22404 9129 -22292
rect 9164 -22404 9322 -22292
rect 9357 -22404 9514 -22292
rect 9549 -22404 9706 -22292
rect 9741 -22404 9885 -22292
rect 9022 -22419 9885 -22404
rect 9953 -22291 10816 -22284
rect 11633 -22285 11743 -21878
rect 9953 -22403 10060 -22291
rect 10095 -22403 10253 -22291
rect 10288 -22403 10445 -22291
rect 10480 -22403 10637 -22291
rect 10672 -22403 10816 -22291
rect 9953 -22418 10816 -22403
rect 10880 -22292 11743 -22285
rect 10880 -22404 10987 -22292
rect 11022 -22404 11180 -22292
rect 11215 -22404 11372 -22292
rect 11407 -22404 11564 -22292
rect 11599 -22404 11743 -22292
rect 10880 -22419 11743 -22404
rect 7137 -22481 10779 -22472
rect 11883 -22473 12147 -22462
rect 7137 -22482 9965 -22481
rect 7137 -22592 7150 -22482
rect 7184 -22592 7342 -22482
rect 7376 -22592 7534 -22482
rect 7568 -22592 7726 -22482
rect 7760 -22592 7918 -22482
rect 7952 -22592 8098 -22482
rect 8132 -22592 8290 -22482
rect 8324 -22592 8482 -22482
rect 8516 -22592 8674 -22482
rect 8708 -22592 8866 -22482
rect 8900 -22592 9034 -22482
rect 9068 -22592 9226 -22482
rect 9260 -22592 9418 -22482
rect 9452 -22592 9610 -22482
rect 9644 -22592 9802 -22482
rect 9836 -22591 9965 -22482
rect 9999 -22591 10157 -22481
rect 10191 -22591 10349 -22481
rect 10383 -22591 10541 -22481
rect 10575 -22591 10733 -22481
rect 10767 -22591 10779 -22481
rect 9836 -22592 10779 -22591
rect 7137 -22663 10779 -22592
rect 10880 -22482 11894 -22473
rect 10880 -22592 10892 -22482
rect 10926 -22592 11084 -22482
rect 11118 -22592 11276 -22482
rect 11310 -22592 11468 -22482
rect 11502 -22592 11660 -22482
rect 11694 -22592 11894 -22482
rect 10880 -22603 11894 -22592
rect 7137 -22664 10204 -22663
rect 7137 -22699 7389 -22664
rect 7677 -22699 8337 -22664
rect 8625 -22699 9273 -22664
rect 9561 -22698 10204 -22664
rect 10492 -22698 10779 -22663
rect 9561 -22699 10779 -22698
rect 7137 -22713 10779 -22699
rect 7137 -22715 7964 -22713
rect 8085 -22715 8912 -22713
rect 9021 -22715 9848 -22713
rect 9952 -22714 10779 -22713
rect 10879 -22664 11894 -22603
rect 10879 -22699 11131 -22664
rect 11419 -22699 11894 -22664
rect 10879 -22715 11894 -22699
rect 12136 -22715 12147 -22473
rect 11883 -22726 12147 -22715
rect 5658 -23185 7357 -23141
rect 5658 -23219 5721 -23185
rect 5812 -23219 6161 -23185
rect 6252 -23219 6601 -23185
rect 6692 -23219 7357 -23185
rect 5658 -23231 7357 -23219
rect 5658 -23257 5872 -23231
rect 5558 -23289 5627 -23283
rect 5558 -23531 5577 -23358
rect 5611 -23531 5627 -23358
rect 5658 -23291 5664 -23257
rect 5743 -23261 5872 -23257
rect 6098 -23257 6312 -23231
rect 5743 -23291 5749 -23261
rect 5998 -23289 6067 -23283
rect 5658 -23449 5749 -23291
rect 5658 -23483 5664 -23449
rect 5743 -23483 5749 -23449
rect 5658 -23499 5749 -23483
rect 5781 -23353 5970 -23289
rect 5781 -23387 5787 -23353
rect 5864 -23387 5970 -23353
rect 5558 -23633 5627 -23531
rect 5781 -23545 5970 -23387
rect 5658 -23579 5787 -23545
rect 5864 -23579 5970 -23545
rect 5558 -23751 5628 -23633
rect 5658 -23707 5970 -23579
rect 5658 -23741 5670 -23707
rect 5846 -23741 5970 -23707
rect 5658 -23747 5858 -23741
rect 5558 -23785 5577 -23751
rect 5611 -23785 5628 -23751
rect 5558 -23802 5628 -23785
rect 5559 -23879 5628 -23802
rect 5558 -23938 5628 -23879
rect 5658 -23795 5858 -23788
rect 5658 -23829 5670 -23795
rect 5846 -23829 5858 -23795
rect 5886 -23802 5970 -23741
rect 5658 -23897 5858 -23829
rect 5658 -23931 5689 -23897
rect 5821 -23931 5858 -23897
rect 5658 -23938 5858 -23931
rect 5901 -23854 5970 -23802
rect 5559 -24054 5628 -23938
rect 5703 -23940 5823 -23938
rect 5703 -23992 5734 -23940
rect 5786 -23992 5823 -23940
rect 5901 -23944 5970 -23923
rect 5998 -23531 6017 -23358
rect 6051 -23531 6067 -23358
rect 6098 -23291 6104 -23257
rect 6183 -23261 6312 -23257
rect 6538 -23244 7357 -23231
rect 6538 -23257 6752 -23244
rect 6183 -23291 6189 -23261
rect 6438 -23289 6507 -23283
rect 6098 -23449 6189 -23291
rect 6098 -23483 6104 -23449
rect 6183 -23483 6189 -23449
rect 6098 -23499 6189 -23483
rect 6221 -23353 6410 -23289
rect 6221 -23387 6227 -23353
rect 6304 -23387 6410 -23353
rect 5998 -23751 6067 -23531
rect 6221 -23545 6410 -23387
rect 6098 -23579 6227 -23545
rect 6304 -23579 6410 -23545
rect 6098 -23707 6410 -23579
rect 6098 -23741 6110 -23707
rect 6286 -23741 6410 -23707
rect 6098 -23747 6298 -23741
rect 5998 -23785 6017 -23751
rect 6051 -23785 6067 -23751
rect 5703 -24023 5823 -23992
rect 5559 -24123 5901 -24054
rect 5559 -24135 5628 -24123
rect 5732 -24649 5798 -24643
rect 5405 -24715 5732 -24649
rect 5732 -24721 5798 -24715
rect 5253 -24745 5383 -24739
rect 5253 -24811 5317 -24745
rect 5317 -24817 5383 -24811
rect 5832 -26716 5901 -24123
rect 5998 -24387 6067 -23785
rect 6098 -23795 6298 -23788
rect 6098 -23829 6110 -23795
rect 6286 -23829 6298 -23795
rect 6326 -23802 6410 -23741
rect 6098 -23897 6298 -23829
rect 6098 -23931 6129 -23897
rect 6261 -23931 6298 -23897
rect 6098 -23938 6172 -23931
rect 6143 -23973 6172 -23938
rect 6224 -23938 6298 -23931
rect 6341 -23856 6410 -23802
rect 6341 -23938 6410 -23925
rect 6438 -23531 6457 -23358
rect 6491 -23531 6507 -23358
rect 6538 -23291 6544 -23257
rect 6623 -23261 6752 -23257
rect 6623 -23291 6629 -23261
rect 6538 -23449 6629 -23291
rect 6538 -23483 6544 -23449
rect 6623 -23483 6629 -23449
rect 6538 -23499 6629 -23483
rect 6661 -23353 6850 -23289
rect 6661 -23387 6667 -23353
rect 6744 -23387 6850 -23353
rect 6438 -23751 6507 -23531
rect 6661 -23545 6850 -23387
rect 6538 -23579 6667 -23545
rect 6744 -23579 6850 -23545
rect 6538 -23707 6850 -23579
rect 6538 -23741 6550 -23707
rect 6726 -23741 6850 -23707
rect 6538 -23747 6738 -23741
rect 6438 -23785 6457 -23751
rect 6491 -23785 6507 -23751
rect 6224 -23973 6263 -23938
rect 6143 -23998 6263 -23973
rect 5992 -24393 6073 -24387
rect 5992 -24462 5998 -24393
rect 6067 -24396 6073 -24393
rect 6067 -24462 6085 -24396
rect 5992 -24468 6073 -24462
rect 5998 -26622 6067 -24468
rect 6438 -24528 6507 -23785
rect 6538 -23795 6738 -23788
rect 6538 -23829 6550 -23795
rect 6726 -23829 6738 -23795
rect 6766 -23802 6850 -23741
rect 6538 -23897 6738 -23829
rect 6781 -23847 6850 -23802
rect 7254 -23841 7357 -23244
rect 11860 -23841 12409 -23840
rect 12750 -23841 13092 -23840
rect 6538 -23931 6569 -23897
rect 6701 -23931 6738 -23897
rect 6538 -23938 6612 -23931
rect 6580 -23964 6612 -23938
rect 6664 -23938 6738 -23931
rect 6780 -23878 6850 -23847
rect 7137 -23842 7964 -23841
rect 8085 -23842 8912 -23841
rect 9021 -23842 9848 -23841
rect 9952 -23842 10779 -23841
rect 7137 -23857 10780 -23842
rect 6664 -23964 6700 -23938
rect 6580 -24007 6700 -23964
rect 6438 -24603 6507 -24597
rect 6780 -24490 6849 -23878
rect 7137 -23892 7389 -23857
rect 7677 -23892 8337 -23857
rect 8625 -23892 9273 -23857
rect 9561 -23892 10204 -23857
rect 10492 -23892 10780 -23857
rect 7137 -23953 10780 -23892
rect 10879 -23857 13092 -23841
rect 10879 -23892 11131 -23857
rect 11419 -23892 13092 -23857
rect 10879 -23953 13092 -23892
rect 7138 -23964 10780 -23953
rect 7138 -24074 7150 -23964
rect 7184 -24074 7342 -23964
rect 7376 -24074 7534 -23964
rect 7568 -24074 7726 -23964
rect 7760 -24074 7918 -23964
rect 7952 -24074 8098 -23964
rect 8132 -24074 8290 -23964
rect 8324 -24074 8482 -23964
rect 8516 -24074 8674 -23964
rect 8708 -24074 8866 -23964
rect 8900 -24074 9034 -23964
rect 9068 -24074 9226 -23964
rect 9260 -24074 9418 -23964
rect 9452 -24074 9610 -23964
rect 9644 -24074 9802 -23964
rect 9836 -24074 9965 -23964
rect 9999 -24074 10157 -23964
rect 10191 -24074 10349 -23964
rect 10383 -24074 10541 -23964
rect 10575 -24074 10733 -23964
rect 10767 -24074 10780 -23964
rect 7138 -24083 10780 -24074
rect 10880 -23964 13092 -23953
rect 10880 -24074 10892 -23964
rect 10926 -24074 11084 -23964
rect 11118 -24074 11276 -23964
rect 11310 -24074 11468 -23964
rect 11502 -24074 11660 -23964
rect 11694 -24074 13092 -23964
rect 10880 -24083 13092 -24074
rect 7138 -24152 8001 -24137
rect 7138 -24264 7245 -24152
rect 7280 -24264 7438 -24152
rect 7473 -24264 7630 -24152
rect 7665 -24264 7822 -24152
rect 7857 -24264 8001 -24152
rect 7138 -24271 8001 -24264
rect 8086 -24152 8949 -24137
rect 8086 -24264 8193 -24152
rect 8228 -24264 8386 -24152
rect 8421 -24264 8578 -24152
rect 8613 -24264 8770 -24152
rect 8805 -24264 8949 -24152
rect 8086 -24271 8949 -24264
rect 9022 -24152 9885 -24137
rect 9022 -24264 9129 -24152
rect 9164 -24264 9322 -24152
rect 9357 -24264 9514 -24152
rect 9549 -24264 9706 -24152
rect 9741 -24264 9885 -24152
rect 9022 -24271 9885 -24264
rect 9953 -24152 10816 -24137
rect 9953 -24264 10060 -24152
rect 10095 -24264 10253 -24152
rect 10288 -24264 10445 -24152
rect 10480 -24264 10637 -24152
rect 10672 -24264 10816 -24152
rect 9953 -24271 10816 -24264
rect 10880 -24152 11743 -24137
rect 10880 -24264 10987 -24152
rect 11022 -24264 11180 -24152
rect 11215 -24264 11372 -24152
rect 11407 -24264 11564 -24152
rect 11599 -24264 11743 -24152
rect 10880 -24271 11743 -24264
rect 7106 -24302 7158 -24301
rect 7102 -24307 7248 -24302
rect 7102 -24359 7106 -24307
rect 7158 -24318 7248 -24307
rect 7158 -24352 7198 -24318
rect 7232 -24352 7248 -24318
rect 7158 -24359 7248 -24352
rect 7102 -24368 7248 -24359
rect 7304 -24318 7441 -24302
rect 7304 -24352 7390 -24318
rect 7424 -24352 7441 -24318
rect 7304 -24368 7441 -24352
rect 7491 -24318 7632 -24303
rect 7491 -24352 7582 -24318
rect 7616 -24352 7632 -24318
rect 7304 -24396 7370 -24368
rect 7097 -24401 7370 -24396
rect 7097 -24453 7113 -24401
rect 7165 -24453 7370 -24401
rect 7491 -24369 7632 -24352
rect 7661 -24318 7825 -24302
rect 7661 -24352 7774 -24318
rect 7808 -24352 7825 -24318
rect 7661 -24368 7825 -24352
rect 7491 -24405 7557 -24369
rect 7594 -24370 7628 -24369
rect 7097 -24462 7370 -24453
rect 7409 -24490 7557 -24405
rect 6780 -24556 7327 -24490
rect 7393 -24556 7557 -24490
rect 6780 -26519 6849 -24556
rect 7661 -24584 7727 -24368
rect 7102 -24650 7727 -24584
rect 7106 -24851 7172 -24650
rect 7891 -24678 8001 -24271
rect 8050 -24308 8196 -24302
rect 8050 -24360 8069 -24308
rect 8122 -24318 8196 -24308
rect 8122 -24352 8146 -24318
rect 8180 -24352 8196 -24318
rect 8122 -24360 8196 -24352
rect 8050 -24368 8196 -24360
rect 8252 -24318 8389 -24302
rect 8252 -24352 8338 -24318
rect 8372 -24352 8389 -24318
rect 8252 -24368 8389 -24352
rect 8439 -24318 8580 -24303
rect 8439 -24352 8530 -24318
rect 8564 -24352 8580 -24318
rect 8252 -24396 8318 -24368
rect 8050 -24400 8318 -24396
rect 8050 -24452 8057 -24400
rect 8109 -24452 8318 -24400
rect 8439 -24369 8580 -24352
rect 8609 -24318 8773 -24302
rect 8609 -24352 8722 -24318
rect 8756 -24352 8773 -24318
rect 8609 -24368 8773 -24352
rect 8439 -24405 8505 -24369
rect 8542 -24370 8576 -24369
rect 8050 -24462 8318 -24452
rect 8357 -24483 8505 -24405
rect 8357 -24490 8424 -24483
rect 8050 -24535 8424 -24490
rect 8493 -24535 8505 -24483
rect 8050 -24556 8505 -24535
rect 8609 -24584 8675 -24368
rect 7106 -24923 7172 -24917
rect 7214 -24690 7413 -24678
rect 7214 -24702 7372 -24690
rect 7214 -25453 7298 -24702
rect 7333 -25453 7372 -24702
rect 7214 -25631 7227 -25453
rect 7406 -25466 7413 -24690
rect 7405 -25618 7413 -25466
rect 7750 -24690 8001 -24678
rect 7750 -25466 7756 -24690
rect 7790 -24693 8001 -24690
rect 8050 -24650 8675 -24584
rect 7790 -25108 8000 -24693
rect 8050 -24955 8116 -24650
rect 8839 -24678 8949 -24271
rect 8986 -24307 9132 -24302
rect 8986 -24359 9002 -24307
rect 9055 -24318 9132 -24307
rect 9055 -24352 9082 -24318
rect 9116 -24352 9132 -24318
rect 9055 -24359 9132 -24352
rect 8986 -24368 9132 -24359
rect 9188 -24318 9325 -24302
rect 9188 -24352 9274 -24318
rect 9308 -24352 9325 -24318
rect 9188 -24368 9325 -24352
rect 9375 -24318 9516 -24303
rect 9375 -24352 9466 -24318
rect 9500 -24352 9516 -24318
rect 9188 -24396 9254 -24368
rect 8986 -24405 9254 -24396
rect 9375 -24369 9516 -24352
rect 9545 -24318 9709 -24302
rect 9545 -24352 9658 -24318
rect 9692 -24352 9709 -24318
rect 9545 -24368 9709 -24352
rect 9375 -24405 9441 -24369
rect 9478 -24370 9512 -24369
rect 8986 -24457 9000 -24405
rect 9052 -24457 9254 -24405
rect 8986 -24462 9254 -24457
rect 9293 -24490 9441 -24405
rect 8986 -24496 9441 -24490
rect 8986 -24549 8989 -24496
rect 9042 -24549 9441 -24496
rect 8986 -24556 9441 -24549
rect 9545 -24584 9611 -24368
rect 8050 -25027 8116 -25021
rect 8162 -24690 8361 -24678
rect 8162 -24702 8320 -24690
rect 7790 -25174 7872 -25108
rect 7938 -25174 8000 -25108
rect 7790 -25466 8000 -25174
rect 7750 -25478 8000 -25466
rect 8162 -25453 8246 -24702
rect 8281 -25453 8320 -24702
rect 8354 -25466 8361 -24690
rect 7102 -26277 7168 -26271
rect 7102 -26434 7168 -26343
rect 7214 -26382 7298 -25631
rect 7333 -26382 7372 -25631
rect 7214 -26394 7372 -26382
rect 7406 -26394 7413 -25618
rect 7214 -26406 7413 -26394
rect 7750 -25618 8000 -25606
rect 7750 -26394 7756 -25618
rect 7790 -25901 8000 -25618
rect 7790 -25967 7853 -25901
rect 7919 -25967 8000 -25901
rect 7790 -26391 8000 -25967
rect 8340 -25618 8361 -25466
rect 8698 -24690 8949 -24678
rect 8698 -25466 8704 -24690
rect 8738 -24693 8949 -24690
rect 8986 -24649 9611 -24584
rect 8738 -24854 8948 -24693
rect 9052 -24650 9611 -24649
rect 9775 -24606 9885 -24271
rect 10706 -24302 10816 -24271
rect 9917 -24307 10063 -24302
rect 9917 -24359 9933 -24307
rect 9986 -24318 10063 -24307
rect 9986 -24352 10013 -24318
rect 10047 -24352 10063 -24318
rect 9986 -24359 10063 -24352
rect 9917 -24368 10063 -24359
rect 10119 -24318 10256 -24302
rect 10119 -24352 10205 -24318
rect 10239 -24352 10256 -24318
rect 10119 -24368 10256 -24352
rect 10306 -24318 10447 -24303
rect 10306 -24352 10397 -24318
rect 10431 -24352 10447 -24318
rect 10119 -24396 10185 -24368
rect 9917 -24405 10185 -24396
rect 10306 -24369 10447 -24352
rect 10476 -24318 10640 -24302
rect 10476 -24352 10589 -24318
rect 10623 -24352 10640 -24318
rect 10476 -24368 10640 -24352
rect 10706 -24318 10990 -24302
rect 10706 -24352 10940 -24318
rect 10974 -24352 10990 -24318
rect 10706 -24368 10990 -24352
rect 11046 -24318 11183 -24302
rect 11046 -24352 11132 -24318
rect 11166 -24352 11183 -24318
rect 11046 -24368 11183 -24352
rect 11233 -24318 11374 -24303
rect 11233 -24352 11324 -24318
rect 11358 -24352 11374 -24318
rect 10306 -24405 10372 -24369
rect 10409 -24370 10443 -24369
rect 9917 -24457 9935 -24405
rect 9987 -24457 10185 -24405
rect 9917 -24462 10185 -24457
rect 10224 -24452 10372 -24405
rect 10224 -24490 10262 -24452
rect 9917 -24521 10262 -24490
rect 10331 -24521 10372 -24452
rect 9917 -24556 10372 -24521
rect 10476 -24584 10542 -24368
rect 9775 -24672 9798 -24606
rect 9864 -24672 9885 -24606
rect 9775 -24678 9885 -24672
rect 8986 -24733 9052 -24715
rect 9098 -24690 9297 -24678
rect 9098 -24702 9256 -24690
rect 8738 -24920 8818 -24854
rect 8884 -24920 8948 -24854
rect 8738 -25466 8948 -24920
rect 8698 -25478 8948 -25466
rect 9098 -25453 9182 -24702
rect 9217 -25453 9256 -24702
rect 9290 -25466 9297 -24690
rect 8162 -26382 8246 -25631
rect 8281 -26382 8320 -25631
rect 7790 -26394 8001 -26391
rect 7750 -26406 8001 -26394
rect 7102 -26500 7727 -26434
rect 6774 -26588 6780 -26519
rect 6849 -26528 6855 -26519
rect 6849 -26588 7557 -26528
rect 6780 -26594 7557 -26588
rect 5998 -26686 6066 -26622
rect 5999 -26688 6066 -26686
rect 6132 -26688 7370 -26622
rect 7409 -26679 7557 -26594
rect 7304 -26716 7370 -26688
rect 7491 -26715 7557 -26679
rect 7594 -26715 7628 -26714
rect 5832 -26782 6941 -26716
rect 7007 -26732 7248 -26716
rect 7007 -26766 7198 -26732
rect 7232 -26766 7248 -26732
rect 7007 -26782 7248 -26766
rect 7304 -26732 7441 -26716
rect 7304 -26766 7390 -26732
rect 7424 -26766 7441 -26732
rect 7304 -26782 7441 -26766
rect 7491 -26732 7632 -26715
rect 7491 -26766 7582 -26732
rect 7616 -26766 7632 -26732
rect 7491 -26781 7632 -26766
rect 7661 -26716 7727 -26500
rect 7661 -26732 7825 -26716
rect 7661 -26766 7774 -26732
rect 7808 -26766 7825 -26732
rect 7661 -26782 7825 -26766
rect 5832 -26792 5901 -26782
rect 7891 -26813 8001 -26406
rect 8050 -26398 8116 -26392
rect 8162 -26394 8320 -26382
rect 8354 -26394 8361 -25618
rect 8162 -26406 8361 -26394
rect 8698 -25618 8948 -25606
rect 8698 -26394 8704 -25618
rect 8738 -26311 8948 -25618
rect 9276 -25618 9297 -25466
rect 9634 -24690 9885 -24678
rect 9634 -25466 9640 -24690
rect 9674 -24693 9885 -24690
rect 9917 -24650 10542 -24584
rect 9674 -25466 9884 -24693
rect 9917 -24745 9983 -24650
rect 10706 -24678 10816 -24368
rect 11046 -24396 11112 -24368
rect 10844 -24462 10860 -24396
rect 10926 -24462 11112 -24396
rect 11233 -24369 11374 -24352
rect 11403 -24318 11567 -24302
rect 11403 -24352 11516 -24318
rect 11550 -24352 11567 -24318
rect 11403 -24368 11567 -24352
rect 11233 -24405 11299 -24369
rect 11336 -24370 11370 -24369
rect 11151 -24490 11299 -24405
rect 10844 -24556 10858 -24490
rect 10924 -24556 11299 -24490
rect 11403 -24584 11469 -24368
rect 10844 -24650 10850 -24584
rect 10915 -24650 11469 -24584
rect 11633 -24678 11743 -24271
rect 9917 -24817 9983 -24811
rect 10029 -24690 10228 -24678
rect 10029 -24702 10187 -24690
rect 9634 -25478 9884 -25466
rect 10029 -25453 10113 -24702
rect 10148 -25453 10187 -24702
rect 10221 -25466 10228 -24690
rect 8738 -26377 8837 -26311
rect 8903 -26377 8948 -26311
rect 8738 -26391 8948 -26377
rect 8989 -26057 9055 -26051
rect 8738 -26394 8949 -26391
rect 8698 -26406 8949 -26394
rect 8116 -26464 8675 -26434
rect 8050 -26500 8675 -26464
rect 8050 -26535 8505 -26528
rect 8050 -26594 8401 -26535
rect 8357 -26599 8401 -26594
rect 8465 -26599 8505 -26535
rect 8050 -26631 8318 -26622
rect 8050 -26683 8079 -26631
rect 8131 -26683 8318 -26631
rect 8357 -26679 8505 -26599
rect 8050 -26688 8318 -26683
rect 8252 -26716 8318 -26688
rect 8439 -26715 8505 -26679
rect 8542 -26715 8576 -26714
rect 8050 -26725 8196 -26716
rect 8050 -26777 8063 -26725
rect 8128 -26732 8196 -26725
rect 8128 -26766 8146 -26732
rect 8180 -26766 8196 -26732
rect 8128 -26777 8196 -26766
rect 8050 -26782 8196 -26777
rect 8252 -26732 8389 -26716
rect 8252 -26766 8338 -26732
rect 8372 -26766 8389 -26732
rect 8252 -26782 8389 -26766
rect 8439 -26732 8580 -26715
rect 8439 -26766 8530 -26732
rect 8564 -26766 8580 -26732
rect 8439 -26781 8580 -26766
rect 8609 -26716 8675 -26500
rect 8609 -26732 8773 -26716
rect 8609 -26766 8722 -26732
rect 8756 -26766 8773 -26732
rect 8609 -26782 8773 -26766
rect 8839 -26813 8949 -26406
rect 8989 -26434 9055 -26123
rect 9098 -26382 9182 -25631
rect 9217 -26382 9256 -25631
rect 9098 -26394 9256 -26382
rect 9290 -26394 9297 -25618
rect 9098 -26406 9297 -26394
rect 9634 -25618 9884 -25606
rect 9634 -26394 9640 -25618
rect 9674 -26391 9884 -25618
rect 10206 -25617 10228 -25466
rect 10565 -24690 10816 -24678
rect 10565 -25466 10571 -24690
rect 10605 -24693 10816 -24690
rect 10956 -24690 11155 -24678
rect 10605 -25466 10815 -24693
rect 10565 -25478 10815 -25466
rect 10956 -24702 11114 -24690
rect 10956 -25453 11040 -24702
rect 11075 -25453 11114 -24702
rect 11148 -25466 11155 -24690
rect 9917 -26179 9983 -26173
rect 9674 -26394 9885 -26391
rect 9634 -26405 9885 -26394
rect 9634 -26406 9807 -26405
rect 8986 -26500 9611 -26434
rect 8986 -26594 8993 -26528
rect 9059 -26594 9441 -26528
rect 8986 -26688 9001 -26622
rect 9067 -26688 9254 -26622
rect 9293 -26679 9441 -26594
rect 9188 -26716 9254 -26688
rect 9375 -26715 9441 -26679
rect 9478 -26715 9512 -26714
rect 8986 -26725 9132 -26716
rect 8986 -26777 8992 -26725
rect 9057 -26732 9132 -26725
rect 9057 -26766 9082 -26732
rect 9116 -26766 9132 -26732
rect 9057 -26777 9132 -26766
rect 8986 -26782 9132 -26777
rect 9188 -26732 9325 -26716
rect 9188 -26766 9274 -26732
rect 9308 -26766 9325 -26732
rect 9188 -26782 9325 -26766
rect 9375 -26732 9516 -26715
rect 9375 -26766 9466 -26732
rect 9500 -26766 9516 -26732
rect 9375 -26781 9516 -26766
rect 9545 -26716 9611 -26500
rect 9775 -26469 9807 -26406
rect 9873 -26469 9885 -26405
rect 9545 -26732 9709 -26716
rect 9545 -26766 9658 -26732
rect 9692 -26766 9709 -26732
rect 9545 -26782 9709 -26766
rect 9775 -26813 9885 -26469
rect 9917 -26433 9983 -26245
rect 10029 -26381 10113 -25630
rect 10148 -26381 10187 -25630
rect 10029 -26393 10187 -26381
rect 10221 -26393 10228 -25617
rect 10029 -26405 10228 -26393
rect 10565 -25617 10815 -25605
rect 10565 -26393 10571 -25617
rect 10605 -26390 10815 -25617
rect 11134 -25618 11155 -25466
rect 11492 -24690 11743 -24678
rect 11492 -25466 11498 -24690
rect 11532 -24693 11743 -24690
rect 11860 -24307 13092 -24083
rect 11860 -24510 12189 -24307
rect 12410 -24510 13092 -24307
rect 11532 -25449 11742 -24693
rect 11860 -25008 13092 -24510
rect 11799 -25016 13092 -25008
rect 11799 -25067 11811 -25016
rect 12168 -25025 13092 -25016
rect 12168 -25067 12180 -25025
rect 11799 -25074 12180 -25067
rect 11860 -25112 11903 -25074
rect 12726 -25159 13092 -25025
rect 11875 -25171 12689 -25159
rect 12726 -25166 13137 -25159
rect 11875 -25261 11881 -25171
rect 11915 -25261 12073 -25171
rect 12107 -25261 12265 -25171
rect 12299 -25261 12457 -25171
rect 12491 -25261 12649 -25171
rect 12683 -25261 12689 -25171
rect 11875 -25273 12689 -25261
rect 12923 -25203 13137 -25166
rect 12923 -25237 12986 -25203
rect 13077 -25237 13137 -25203
rect 12923 -25275 13137 -25237
rect 11779 -25313 12209 -25301
rect 11779 -25403 11785 -25313
rect 11819 -25403 11977 -25313
rect 12011 -25403 12169 -25313
rect 12203 -25403 12209 -25313
rect 11779 -25415 12209 -25403
rect 12355 -25307 12827 -25301
rect 12355 -25313 12892 -25307
rect 12355 -25403 12361 -25313
rect 12395 -25403 12553 -25313
rect 12587 -25403 12745 -25313
rect 12779 -25323 12892 -25313
rect 12779 -25403 12842 -25323
rect 12355 -25415 12842 -25403
rect 11532 -25465 12263 -25449
rect 11532 -25466 12170 -25465
rect 11492 -25478 12170 -25466
rect 11737 -25499 12170 -25478
rect 12204 -25499 12263 -25465
rect 11737 -25515 12263 -25499
rect 12702 -25549 12842 -25415
rect 12876 -25549 12892 -25323
rect 12923 -25309 12929 -25275
rect 13008 -25279 13137 -25275
rect 13008 -25309 13014 -25279
rect 12923 -25467 13014 -25309
rect 12923 -25501 12929 -25467
rect 13008 -25501 13014 -25467
rect 12923 -25517 13014 -25501
rect 13046 -25371 13235 -25307
rect 13046 -25405 13052 -25371
rect 13129 -25405 13235 -25371
rect 13046 -25506 13235 -25405
rect 15261 -25506 15327 -19696
rect 16177 -19724 16244 -19696
rect 11703 -25570 12363 -25554
rect 11703 -25604 12313 -25570
rect 12347 -25604 12363 -25570
rect 11703 -25606 12363 -25604
rect 10956 -26382 11040 -25631
rect 11075 -26382 11114 -25631
rect 10605 -26393 10816 -26390
rect 10565 -26405 10816 -26393
rect 9917 -26499 10542 -26433
rect 9917 -26535 10372 -26527
rect 9917 -26593 10264 -26535
rect 10224 -26595 10264 -26593
rect 10324 -26595 10372 -26535
rect 9917 -26687 9937 -26621
rect 10003 -26687 10185 -26621
rect 10224 -26678 10372 -26595
rect 10119 -26715 10185 -26687
rect 10306 -26714 10372 -26678
rect 10409 -26714 10443 -26713
rect 9917 -26725 10063 -26715
rect 9917 -26777 9951 -26725
rect 10016 -26731 10063 -26725
rect 10047 -26765 10063 -26731
rect 10016 -26777 10063 -26765
rect 9917 -26781 10063 -26777
rect 10119 -26731 10256 -26715
rect 10119 -26765 10205 -26731
rect 10239 -26765 10256 -26731
rect 10119 -26781 10256 -26765
rect 10306 -26731 10447 -26714
rect 10306 -26765 10397 -26731
rect 10431 -26765 10447 -26731
rect 10306 -26780 10447 -26765
rect 10476 -26715 10542 -26499
rect 10476 -26731 10640 -26715
rect 10476 -26765 10589 -26731
rect 10623 -26765 10640 -26731
rect 10476 -26781 10640 -26765
rect 10706 -26716 10816 -26405
rect 10956 -26394 11114 -26382
rect 11148 -26394 11155 -25618
rect 10956 -26406 11155 -26394
rect 11492 -25618 12363 -25606
rect 11492 -26394 11498 -25618
rect 11532 -25620 12363 -25618
rect 11532 -25651 11815 -25620
rect 11532 -26391 11742 -25651
rect 12259 -25654 12305 -25648
rect 12702 -25654 12892 -25549
rect 13046 -25563 15327 -25506
rect 12259 -25660 12892 -25654
rect 12259 -25836 12265 -25660
rect 12299 -25769 12892 -25660
rect 12923 -25597 13052 -25563
rect 13129 -25572 15327 -25563
rect 15447 -19790 16244 -19724
rect 13129 -25597 13235 -25572
rect 12923 -25725 13235 -25597
rect 12923 -25759 12935 -25725
rect 13111 -25759 13235 -25725
rect 12923 -25765 13123 -25759
rect 12299 -25803 12842 -25769
rect 12876 -25803 12892 -25769
rect 12299 -25820 12892 -25803
rect 12923 -25813 13123 -25806
rect 12299 -25836 12827 -25820
rect 12259 -25848 12827 -25836
rect 12305 -25852 12827 -25848
rect 12923 -25847 12935 -25813
rect 13111 -25847 13123 -25813
rect 13151 -25820 13235 -25759
rect 12305 -25853 12825 -25852
rect 12305 -25854 12774 -25853
rect 12171 -25919 12394 -25912
rect 12171 -25967 12183 -25919
rect 12074 -25980 12183 -25967
rect 12382 -25967 12394 -25919
rect 12923 -25915 13123 -25847
rect 12923 -25949 12954 -25915
rect 13086 -25949 13123 -25915
rect 12921 -25956 13123 -25949
rect 12382 -25980 12473 -25967
rect 12074 -26083 12233 -25980
rect 12352 -26083 12473 -25980
rect 12921 -26005 13121 -25956
rect 12921 -26027 12960 -26005
rect 12074 -26157 12473 -26083
rect 12923 -26124 12960 -26027
rect 13079 -26027 13121 -26005
rect 13079 -26124 13113 -26027
rect 12923 -26182 13113 -26124
rect 11532 -26394 11743 -26391
rect 11492 -26406 11743 -26394
rect 10844 -26500 10850 -26434
rect 10916 -26500 11469 -26434
rect 10844 -26594 10888 -26528
rect 10954 -26594 11299 -26528
rect 10844 -26688 10859 -26622
rect 10925 -26688 11112 -26622
rect 11151 -26679 11299 -26594
rect 11046 -26716 11112 -26688
rect 11233 -26715 11299 -26679
rect 11336 -26715 11370 -26714
rect 10706 -26732 10990 -26716
rect 10706 -26766 10940 -26732
rect 10974 -26766 10990 -26732
rect 10706 -26782 10990 -26766
rect 11046 -26732 11183 -26716
rect 11046 -26766 11132 -26732
rect 11166 -26766 11183 -26732
rect 11046 -26782 11183 -26766
rect 11233 -26732 11374 -26715
rect 11233 -26766 11324 -26732
rect 11358 -26766 11374 -26732
rect 11233 -26781 11374 -26766
rect 11403 -26716 11469 -26500
rect 11403 -26732 11567 -26716
rect 11403 -26766 11516 -26732
rect 11550 -26766 11567 -26732
rect 11403 -26782 11567 -26766
rect 10706 -26812 10816 -26782
rect 7138 -26820 8001 -26813
rect 7138 -26932 7245 -26820
rect 7280 -26932 7438 -26820
rect 7473 -26932 7630 -26820
rect 7665 -26932 7822 -26820
rect 7857 -26932 8001 -26820
rect 7138 -26947 8001 -26932
rect 8086 -26820 8949 -26813
rect 8086 -26932 8193 -26820
rect 8228 -26932 8386 -26820
rect 8421 -26932 8578 -26820
rect 8613 -26932 8770 -26820
rect 8805 -26932 8949 -26820
rect 8086 -26947 8949 -26932
rect 9022 -26820 9885 -26813
rect 9022 -26932 9129 -26820
rect 9164 -26932 9322 -26820
rect 9357 -26932 9514 -26820
rect 9549 -26932 9706 -26820
rect 9741 -26932 9885 -26820
rect 9022 -26947 9885 -26932
rect 9953 -26819 10816 -26812
rect 11633 -26813 11743 -26406
rect 9953 -26931 10060 -26819
rect 10095 -26931 10253 -26819
rect 10288 -26931 10445 -26819
rect 10480 -26931 10637 -26819
rect 10672 -26931 10816 -26819
rect 9953 -26946 10816 -26931
rect 10880 -26820 11743 -26813
rect 10880 -26932 10987 -26820
rect 11022 -26932 11180 -26820
rect 11215 -26932 11372 -26820
rect 11407 -26932 11564 -26820
rect 11599 -26932 11743 -26820
rect 10880 -26947 11743 -26932
rect 7137 -27009 10779 -27000
rect 11883 -27001 12147 -26990
rect 7137 -27010 9965 -27009
rect 7137 -27120 7150 -27010
rect 7184 -27120 7342 -27010
rect 7376 -27120 7534 -27010
rect 7568 -27120 7726 -27010
rect 7760 -27120 7918 -27010
rect 7952 -27120 8098 -27010
rect 8132 -27120 8290 -27010
rect 8324 -27120 8482 -27010
rect 8516 -27120 8674 -27010
rect 8708 -27120 8866 -27010
rect 8900 -27120 9034 -27010
rect 9068 -27120 9226 -27010
rect 9260 -27120 9418 -27010
rect 9452 -27120 9610 -27010
rect 9644 -27120 9802 -27010
rect 9836 -27119 9965 -27010
rect 9999 -27119 10157 -27009
rect 10191 -27119 10349 -27009
rect 10383 -27119 10541 -27009
rect 10575 -27119 10733 -27009
rect 10767 -27119 10779 -27009
rect 9836 -27120 10779 -27119
rect 7137 -27191 10779 -27120
rect 10880 -27010 11894 -27001
rect 10880 -27120 10892 -27010
rect 10926 -27120 11084 -27010
rect 11118 -27120 11276 -27010
rect 11310 -27120 11468 -27010
rect 11502 -27120 11660 -27010
rect 11694 -27120 11894 -27010
rect 10880 -27131 11894 -27120
rect 7137 -27192 10204 -27191
rect 7137 -27227 7389 -27192
rect 7677 -27227 8337 -27192
rect 8625 -27227 9273 -27192
rect 9561 -27226 10204 -27192
rect 10492 -27226 10779 -27191
rect 9561 -27227 10779 -27226
rect 7137 -27241 10779 -27227
rect 7137 -27243 7964 -27241
rect 8085 -27243 8912 -27241
rect 9021 -27243 9848 -27241
rect 9952 -27242 10779 -27241
rect 10879 -27192 11894 -27131
rect 10879 -27227 11131 -27192
rect 11419 -27227 11894 -27192
rect 10879 -27243 11894 -27227
rect 12136 -27243 12147 -27001
rect 11883 -27254 12147 -27243
rect 5658 -27713 7357 -27669
rect 5658 -27747 5721 -27713
rect 5812 -27747 6161 -27713
rect 6252 -27747 6601 -27713
rect 6692 -27747 7357 -27713
rect 5658 -27759 7357 -27747
rect 5658 -27785 5872 -27759
rect 5558 -27817 5627 -27811
rect 5558 -28059 5577 -27886
rect 5611 -28059 5627 -27886
rect 5658 -27819 5664 -27785
rect 5743 -27789 5872 -27785
rect 6098 -27785 6312 -27759
rect 5743 -27819 5749 -27789
rect 5998 -27817 6067 -27811
rect 5658 -27977 5749 -27819
rect 5658 -28011 5664 -27977
rect 5743 -28011 5749 -27977
rect 5658 -28027 5749 -28011
rect 5781 -27881 5970 -27817
rect 5781 -27915 5787 -27881
rect 5864 -27915 5970 -27881
rect 4573 -28130 5520 -28064
rect 4427 -28374 5329 -28308
rect 1078 -29337 4860 -29278
rect 4919 -29337 4925 -29278
rect 5263 -29395 5329 -28374
rect 5454 -29177 5520 -28130
rect 5558 -28161 5627 -28059
rect 5781 -28073 5970 -27915
rect 5658 -28107 5787 -28073
rect 5864 -28107 5970 -28073
rect 5558 -28279 5628 -28161
rect 5658 -28235 5970 -28107
rect 5658 -28269 5670 -28235
rect 5846 -28269 5970 -28235
rect 5658 -28275 5858 -28269
rect 5558 -28313 5577 -28279
rect 5611 -28313 5628 -28279
rect 5558 -28330 5628 -28313
rect 5559 -28407 5628 -28330
rect 5558 -28466 5628 -28407
rect 5658 -28323 5858 -28316
rect 5658 -28357 5670 -28323
rect 5846 -28357 5858 -28323
rect 5886 -28330 5970 -28269
rect 5658 -28425 5858 -28357
rect 5658 -28459 5689 -28425
rect 5821 -28459 5858 -28425
rect 5658 -28466 5858 -28459
rect 5901 -28382 5970 -28330
rect 5559 -28582 5628 -28466
rect 5703 -28468 5823 -28466
rect 5703 -28520 5734 -28468
rect 5786 -28520 5823 -28468
rect 5901 -28472 5970 -28451
rect 5998 -28059 6017 -27886
rect 6051 -28059 6067 -27886
rect 6098 -27819 6104 -27785
rect 6183 -27789 6312 -27785
rect 6538 -27772 7357 -27759
rect 6538 -27785 6752 -27772
rect 6183 -27819 6189 -27789
rect 6438 -27817 6507 -27811
rect 6098 -27977 6189 -27819
rect 6098 -28011 6104 -27977
rect 6183 -28011 6189 -27977
rect 6098 -28027 6189 -28011
rect 6221 -27881 6410 -27817
rect 6221 -27915 6227 -27881
rect 6304 -27915 6410 -27881
rect 5998 -28279 6067 -28059
rect 6221 -28073 6410 -27915
rect 6098 -28107 6227 -28073
rect 6304 -28107 6410 -28073
rect 6098 -28235 6410 -28107
rect 6098 -28269 6110 -28235
rect 6286 -28269 6410 -28235
rect 6098 -28275 6298 -28269
rect 5998 -28313 6017 -28279
rect 6051 -28313 6067 -28279
rect 5703 -28551 5823 -28520
rect 5559 -28651 5901 -28582
rect 5559 -28663 5628 -28651
rect 5454 -29249 5520 -29243
rect 5263 -29461 5491 -29395
rect 5425 -33705 5491 -29461
rect 5832 -31244 5901 -28651
rect 5998 -28915 6067 -28313
rect 6098 -28323 6298 -28316
rect 6098 -28357 6110 -28323
rect 6286 -28357 6298 -28323
rect 6326 -28330 6410 -28269
rect 6098 -28425 6298 -28357
rect 6098 -28459 6129 -28425
rect 6261 -28459 6298 -28425
rect 6098 -28466 6172 -28459
rect 6143 -28501 6172 -28466
rect 6224 -28466 6298 -28459
rect 6341 -28384 6410 -28330
rect 6341 -28466 6410 -28453
rect 6438 -28059 6457 -27886
rect 6491 -28059 6507 -27886
rect 6538 -27819 6544 -27785
rect 6623 -27789 6752 -27785
rect 6623 -27819 6629 -27789
rect 6538 -27977 6629 -27819
rect 6538 -28011 6544 -27977
rect 6623 -28011 6629 -27977
rect 6538 -28027 6629 -28011
rect 6661 -27881 6850 -27817
rect 6661 -27915 6667 -27881
rect 6744 -27915 6850 -27881
rect 6438 -28279 6507 -28059
rect 6661 -28073 6850 -27915
rect 6538 -28107 6667 -28073
rect 6744 -28107 6850 -28073
rect 6538 -28235 6850 -28107
rect 6538 -28269 6550 -28235
rect 6726 -28269 6850 -28235
rect 6538 -28275 6738 -28269
rect 6438 -28313 6457 -28279
rect 6491 -28313 6507 -28279
rect 6224 -28501 6263 -28466
rect 6143 -28526 6263 -28501
rect 5992 -28921 6073 -28915
rect 5992 -28990 5998 -28921
rect 6067 -28924 6073 -28921
rect 6067 -28990 6085 -28924
rect 5992 -28996 6073 -28990
rect 5998 -31150 6067 -28996
rect 6438 -29056 6507 -28313
rect 6538 -28323 6738 -28316
rect 6538 -28357 6550 -28323
rect 6726 -28357 6738 -28323
rect 6766 -28330 6850 -28269
rect 6538 -28425 6738 -28357
rect 6781 -28375 6850 -28330
rect 7254 -28369 7357 -27772
rect 11860 -28369 12409 -28368
rect 12750 -28369 13092 -28368
rect 6538 -28459 6569 -28425
rect 6701 -28459 6738 -28425
rect 6538 -28466 6612 -28459
rect 6580 -28492 6612 -28466
rect 6664 -28466 6738 -28459
rect 6780 -28406 6850 -28375
rect 7137 -28370 7964 -28369
rect 8085 -28370 8912 -28369
rect 9021 -28370 9848 -28369
rect 9952 -28370 10779 -28369
rect 7137 -28385 10780 -28370
rect 6664 -28492 6700 -28466
rect 6580 -28535 6700 -28492
rect 6438 -29131 6507 -29125
rect 6780 -29018 6849 -28406
rect 7137 -28420 7389 -28385
rect 7677 -28420 8337 -28385
rect 8625 -28420 9273 -28385
rect 9561 -28420 10204 -28385
rect 10492 -28420 10780 -28385
rect 7137 -28481 10780 -28420
rect 10879 -28385 13092 -28369
rect 10879 -28420 11131 -28385
rect 11419 -28420 13092 -28385
rect 10879 -28481 13092 -28420
rect 7138 -28492 10780 -28481
rect 7138 -28602 7150 -28492
rect 7184 -28602 7342 -28492
rect 7376 -28602 7534 -28492
rect 7568 -28602 7726 -28492
rect 7760 -28602 7918 -28492
rect 7952 -28602 8098 -28492
rect 8132 -28602 8290 -28492
rect 8324 -28602 8482 -28492
rect 8516 -28602 8674 -28492
rect 8708 -28602 8866 -28492
rect 8900 -28602 9034 -28492
rect 9068 -28602 9226 -28492
rect 9260 -28602 9418 -28492
rect 9452 -28602 9610 -28492
rect 9644 -28602 9802 -28492
rect 9836 -28602 9965 -28492
rect 9999 -28602 10157 -28492
rect 10191 -28602 10349 -28492
rect 10383 -28602 10541 -28492
rect 10575 -28602 10733 -28492
rect 10767 -28602 10780 -28492
rect 7138 -28611 10780 -28602
rect 10880 -28492 13092 -28481
rect 10880 -28602 10892 -28492
rect 10926 -28602 11084 -28492
rect 11118 -28602 11276 -28492
rect 11310 -28602 11468 -28492
rect 11502 -28602 11660 -28492
rect 11694 -28602 13092 -28492
rect 10880 -28611 13092 -28602
rect 7138 -28680 8001 -28665
rect 7138 -28792 7245 -28680
rect 7280 -28792 7438 -28680
rect 7473 -28792 7630 -28680
rect 7665 -28792 7822 -28680
rect 7857 -28792 8001 -28680
rect 7138 -28799 8001 -28792
rect 8086 -28680 8949 -28665
rect 8086 -28792 8193 -28680
rect 8228 -28792 8386 -28680
rect 8421 -28792 8578 -28680
rect 8613 -28792 8770 -28680
rect 8805 -28792 8949 -28680
rect 8086 -28799 8949 -28792
rect 9022 -28680 9885 -28665
rect 9022 -28792 9129 -28680
rect 9164 -28792 9322 -28680
rect 9357 -28792 9514 -28680
rect 9549 -28792 9706 -28680
rect 9741 -28792 9885 -28680
rect 9022 -28799 9885 -28792
rect 9953 -28680 10816 -28665
rect 9953 -28792 10060 -28680
rect 10095 -28792 10253 -28680
rect 10288 -28792 10445 -28680
rect 10480 -28792 10637 -28680
rect 10672 -28792 10816 -28680
rect 9953 -28799 10816 -28792
rect 10880 -28680 11743 -28665
rect 10880 -28792 10987 -28680
rect 11022 -28792 11180 -28680
rect 11215 -28792 11372 -28680
rect 11407 -28792 11564 -28680
rect 11599 -28792 11743 -28680
rect 10880 -28799 11743 -28792
rect 7106 -28830 7158 -28829
rect 7102 -28835 7248 -28830
rect 7102 -28887 7106 -28835
rect 7158 -28846 7248 -28835
rect 7158 -28880 7198 -28846
rect 7232 -28880 7248 -28846
rect 7158 -28887 7248 -28880
rect 7102 -28896 7248 -28887
rect 7304 -28846 7441 -28830
rect 7304 -28880 7390 -28846
rect 7424 -28880 7441 -28846
rect 7304 -28896 7441 -28880
rect 7491 -28846 7632 -28831
rect 7491 -28880 7582 -28846
rect 7616 -28880 7632 -28846
rect 7304 -28924 7370 -28896
rect 7097 -28929 7370 -28924
rect 7097 -28981 7113 -28929
rect 7165 -28981 7370 -28929
rect 7491 -28897 7632 -28880
rect 7661 -28846 7825 -28830
rect 7661 -28880 7774 -28846
rect 7808 -28880 7825 -28846
rect 7661 -28896 7825 -28880
rect 7491 -28933 7557 -28897
rect 7594 -28898 7628 -28897
rect 7097 -28990 7370 -28981
rect 7409 -29018 7557 -28933
rect 6780 -29084 7327 -29018
rect 7393 -29084 7557 -29018
rect 6780 -31047 6849 -29084
rect 7661 -29112 7727 -28896
rect 7102 -29178 7727 -29112
rect 7106 -29379 7172 -29178
rect 7891 -29206 8001 -28799
rect 8050 -28836 8196 -28830
rect 8050 -28888 8069 -28836
rect 8122 -28846 8196 -28836
rect 8122 -28880 8146 -28846
rect 8180 -28880 8196 -28846
rect 8122 -28888 8196 -28880
rect 8050 -28896 8196 -28888
rect 8252 -28846 8389 -28830
rect 8252 -28880 8338 -28846
rect 8372 -28880 8389 -28846
rect 8252 -28896 8389 -28880
rect 8439 -28846 8580 -28831
rect 8439 -28880 8530 -28846
rect 8564 -28880 8580 -28846
rect 8252 -28924 8318 -28896
rect 8050 -28928 8318 -28924
rect 8050 -28980 8057 -28928
rect 8109 -28980 8318 -28928
rect 8439 -28897 8580 -28880
rect 8609 -28846 8773 -28830
rect 8609 -28880 8722 -28846
rect 8756 -28880 8773 -28846
rect 8609 -28896 8773 -28880
rect 8439 -28933 8505 -28897
rect 8542 -28898 8576 -28897
rect 8050 -28990 8318 -28980
rect 8357 -29011 8505 -28933
rect 8357 -29018 8424 -29011
rect 8050 -29063 8424 -29018
rect 8493 -29063 8505 -29011
rect 8050 -29084 8505 -29063
rect 8609 -29112 8675 -28896
rect 7106 -29451 7172 -29445
rect 7214 -29218 7413 -29206
rect 7214 -29230 7372 -29218
rect 7214 -29981 7298 -29230
rect 7333 -29981 7372 -29230
rect 7214 -30159 7227 -29981
rect 7406 -29994 7413 -29218
rect 7405 -30146 7413 -29994
rect 7750 -29218 8001 -29206
rect 7750 -29994 7756 -29218
rect 7790 -29221 8001 -29218
rect 8050 -29178 8675 -29112
rect 7790 -29636 8000 -29221
rect 8050 -29483 8116 -29178
rect 8839 -29206 8949 -28799
rect 8986 -28835 9132 -28830
rect 8986 -28887 9002 -28835
rect 9055 -28846 9132 -28835
rect 9055 -28880 9082 -28846
rect 9116 -28880 9132 -28846
rect 9055 -28887 9132 -28880
rect 8986 -28896 9132 -28887
rect 9188 -28846 9325 -28830
rect 9188 -28880 9274 -28846
rect 9308 -28880 9325 -28846
rect 9188 -28896 9325 -28880
rect 9375 -28846 9516 -28831
rect 9375 -28880 9466 -28846
rect 9500 -28880 9516 -28846
rect 9188 -28924 9254 -28896
rect 8986 -28933 9254 -28924
rect 9375 -28897 9516 -28880
rect 9545 -28846 9709 -28830
rect 9545 -28880 9658 -28846
rect 9692 -28880 9709 -28846
rect 9545 -28896 9709 -28880
rect 9375 -28933 9441 -28897
rect 9478 -28898 9512 -28897
rect 8986 -28985 9000 -28933
rect 9052 -28985 9254 -28933
rect 8986 -28990 9254 -28985
rect 9293 -29018 9441 -28933
rect 8986 -29024 9441 -29018
rect 8986 -29077 8989 -29024
rect 9042 -29077 9441 -29024
rect 8986 -29084 9441 -29077
rect 9545 -29112 9611 -28896
rect 8050 -29555 8116 -29549
rect 8162 -29218 8361 -29206
rect 8162 -29230 8320 -29218
rect 7790 -29702 7872 -29636
rect 7938 -29702 8000 -29636
rect 7790 -29994 8000 -29702
rect 7750 -30006 8000 -29994
rect 8162 -29981 8246 -29230
rect 8281 -29981 8320 -29230
rect 8354 -29994 8361 -29218
rect 7102 -30805 7168 -30799
rect 7102 -30962 7168 -30871
rect 7214 -30910 7298 -30159
rect 7333 -30910 7372 -30159
rect 7214 -30922 7372 -30910
rect 7406 -30922 7413 -30146
rect 7214 -30934 7413 -30922
rect 7750 -30146 8000 -30134
rect 7750 -30922 7756 -30146
rect 7790 -30429 8000 -30146
rect 7790 -30495 7853 -30429
rect 7919 -30495 8000 -30429
rect 7790 -30919 8000 -30495
rect 8340 -30146 8361 -29994
rect 8698 -29218 8949 -29206
rect 8698 -29994 8704 -29218
rect 8738 -29221 8949 -29218
rect 8986 -29177 9611 -29112
rect 8738 -29382 8948 -29221
rect 9052 -29178 9611 -29177
rect 9775 -29134 9885 -28799
rect 10706 -28830 10816 -28799
rect 9917 -28835 10063 -28830
rect 9917 -28887 9933 -28835
rect 9986 -28846 10063 -28835
rect 9986 -28880 10013 -28846
rect 10047 -28880 10063 -28846
rect 9986 -28887 10063 -28880
rect 9917 -28896 10063 -28887
rect 10119 -28846 10256 -28830
rect 10119 -28880 10205 -28846
rect 10239 -28880 10256 -28846
rect 10119 -28896 10256 -28880
rect 10306 -28846 10447 -28831
rect 10306 -28880 10397 -28846
rect 10431 -28880 10447 -28846
rect 10119 -28924 10185 -28896
rect 9917 -28933 10185 -28924
rect 10306 -28897 10447 -28880
rect 10476 -28846 10640 -28830
rect 10476 -28880 10589 -28846
rect 10623 -28880 10640 -28846
rect 10476 -28896 10640 -28880
rect 10706 -28846 10990 -28830
rect 10706 -28880 10940 -28846
rect 10974 -28880 10990 -28846
rect 10706 -28896 10990 -28880
rect 11046 -28846 11183 -28830
rect 11046 -28880 11132 -28846
rect 11166 -28880 11183 -28846
rect 11046 -28896 11183 -28880
rect 11233 -28846 11374 -28831
rect 11233 -28880 11324 -28846
rect 11358 -28880 11374 -28846
rect 10306 -28933 10372 -28897
rect 10409 -28898 10443 -28897
rect 9917 -28985 9935 -28933
rect 9987 -28985 10185 -28933
rect 9917 -28990 10185 -28985
rect 10224 -28980 10372 -28933
rect 10224 -29018 10262 -28980
rect 9917 -29049 10262 -29018
rect 10331 -29049 10372 -28980
rect 9917 -29084 10372 -29049
rect 10476 -29112 10542 -28896
rect 9775 -29200 9798 -29134
rect 9864 -29200 9885 -29134
rect 9775 -29206 9885 -29200
rect 8986 -29261 9052 -29243
rect 9098 -29218 9297 -29206
rect 9098 -29230 9256 -29218
rect 8738 -29448 8818 -29382
rect 8884 -29448 8948 -29382
rect 8738 -29994 8948 -29448
rect 8698 -30006 8948 -29994
rect 9098 -29981 9182 -29230
rect 9217 -29981 9256 -29230
rect 9290 -29994 9297 -29218
rect 8162 -30910 8246 -30159
rect 8281 -30910 8320 -30159
rect 7790 -30922 8001 -30919
rect 7750 -30934 8001 -30922
rect 7102 -31028 7727 -30962
rect 6774 -31116 6780 -31047
rect 6849 -31056 6855 -31047
rect 6849 -31116 7557 -31056
rect 6780 -31122 7557 -31116
rect 5998 -31214 6066 -31150
rect 5999 -31216 6066 -31214
rect 6132 -31216 7370 -31150
rect 7409 -31207 7557 -31122
rect 7304 -31244 7370 -31216
rect 7491 -31243 7557 -31207
rect 7594 -31243 7628 -31242
rect 5832 -31310 6941 -31244
rect 7007 -31260 7248 -31244
rect 7007 -31294 7198 -31260
rect 7232 -31294 7248 -31260
rect 7007 -31310 7248 -31294
rect 7304 -31260 7441 -31244
rect 7304 -31294 7390 -31260
rect 7424 -31294 7441 -31260
rect 7304 -31310 7441 -31294
rect 7491 -31260 7632 -31243
rect 7491 -31294 7582 -31260
rect 7616 -31294 7632 -31260
rect 7491 -31309 7632 -31294
rect 7661 -31244 7727 -31028
rect 7661 -31260 7825 -31244
rect 7661 -31294 7774 -31260
rect 7808 -31294 7825 -31260
rect 7661 -31310 7825 -31294
rect 5832 -31320 5901 -31310
rect 7891 -31341 8001 -30934
rect 8050 -30926 8116 -30920
rect 8162 -30922 8320 -30910
rect 8354 -30922 8361 -30146
rect 8162 -30934 8361 -30922
rect 8698 -30146 8948 -30134
rect 8698 -30922 8704 -30146
rect 8738 -30839 8948 -30146
rect 9276 -30146 9297 -29994
rect 9634 -29218 9885 -29206
rect 9634 -29994 9640 -29218
rect 9674 -29221 9885 -29218
rect 9917 -29178 10542 -29112
rect 9674 -29994 9884 -29221
rect 9917 -29273 9983 -29178
rect 10706 -29206 10816 -28896
rect 11046 -28924 11112 -28896
rect 10844 -28990 10860 -28924
rect 10926 -28990 11112 -28924
rect 11233 -28897 11374 -28880
rect 11403 -28846 11567 -28830
rect 11403 -28880 11516 -28846
rect 11550 -28880 11567 -28846
rect 11403 -28896 11567 -28880
rect 11233 -28933 11299 -28897
rect 11336 -28898 11370 -28897
rect 11151 -29018 11299 -28933
rect 10844 -29084 10858 -29018
rect 10924 -29084 11299 -29018
rect 11403 -29112 11469 -28896
rect 10844 -29178 10850 -29112
rect 10915 -29178 11469 -29112
rect 11633 -29206 11743 -28799
rect 9917 -29345 9983 -29339
rect 10029 -29218 10228 -29206
rect 10029 -29230 10187 -29218
rect 9634 -30006 9884 -29994
rect 10029 -29981 10113 -29230
rect 10148 -29981 10187 -29230
rect 10221 -29994 10228 -29218
rect 8738 -30905 8837 -30839
rect 8903 -30905 8948 -30839
rect 8738 -30919 8948 -30905
rect 8989 -30585 9055 -30579
rect 8738 -30922 8949 -30919
rect 8698 -30934 8949 -30922
rect 8116 -30992 8675 -30962
rect 8050 -31028 8675 -30992
rect 8050 -31063 8505 -31056
rect 8050 -31122 8401 -31063
rect 8357 -31127 8401 -31122
rect 8465 -31127 8505 -31063
rect 8050 -31159 8318 -31150
rect 8050 -31211 8079 -31159
rect 8131 -31211 8318 -31159
rect 8357 -31207 8505 -31127
rect 8050 -31216 8318 -31211
rect 8252 -31244 8318 -31216
rect 8439 -31243 8505 -31207
rect 8542 -31243 8576 -31242
rect 8050 -31253 8196 -31244
rect 8050 -31305 8063 -31253
rect 8128 -31260 8196 -31253
rect 8128 -31294 8146 -31260
rect 8180 -31294 8196 -31260
rect 8128 -31305 8196 -31294
rect 8050 -31310 8196 -31305
rect 8252 -31260 8389 -31244
rect 8252 -31294 8338 -31260
rect 8372 -31294 8389 -31260
rect 8252 -31310 8389 -31294
rect 8439 -31260 8580 -31243
rect 8439 -31294 8530 -31260
rect 8564 -31294 8580 -31260
rect 8439 -31309 8580 -31294
rect 8609 -31244 8675 -31028
rect 8609 -31260 8773 -31244
rect 8609 -31294 8722 -31260
rect 8756 -31294 8773 -31260
rect 8609 -31310 8773 -31294
rect 8839 -31341 8949 -30934
rect 8989 -30962 9055 -30651
rect 9098 -30910 9182 -30159
rect 9217 -30910 9256 -30159
rect 9098 -30922 9256 -30910
rect 9290 -30922 9297 -30146
rect 9098 -30934 9297 -30922
rect 9634 -30146 9884 -30134
rect 9634 -30922 9640 -30146
rect 9674 -30919 9884 -30146
rect 10206 -30145 10228 -29994
rect 10565 -29218 10816 -29206
rect 10565 -29994 10571 -29218
rect 10605 -29221 10816 -29218
rect 10956 -29218 11155 -29206
rect 10605 -29994 10815 -29221
rect 10565 -30006 10815 -29994
rect 10956 -29230 11114 -29218
rect 10956 -29981 11040 -29230
rect 11075 -29981 11114 -29230
rect 11148 -29994 11155 -29218
rect 9917 -30707 9983 -30701
rect 9674 -30922 9885 -30919
rect 9634 -30933 9885 -30922
rect 9634 -30934 9807 -30933
rect 8986 -31028 9611 -30962
rect 8986 -31122 8993 -31056
rect 9059 -31122 9441 -31056
rect 8986 -31216 9001 -31150
rect 9067 -31216 9254 -31150
rect 9293 -31207 9441 -31122
rect 9188 -31244 9254 -31216
rect 9375 -31243 9441 -31207
rect 9478 -31243 9512 -31242
rect 8986 -31253 9132 -31244
rect 8986 -31305 8992 -31253
rect 9057 -31260 9132 -31253
rect 9057 -31294 9082 -31260
rect 9116 -31294 9132 -31260
rect 9057 -31305 9132 -31294
rect 8986 -31310 9132 -31305
rect 9188 -31260 9325 -31244
rect 9188 -31294 9274 -31260
rect 9308 -31294 9325 -31260
rect 9188 -31310 9325 -31294
rect 9375 -31260 9516 -31243
rect 9375 -31294 9466 -31260
rect 9500 -31294 9516 -31260
rect 9375 -31309 9516 -31294
rect 9545 -31244 9611 -31028
rect 9775 -30997 9807 -30934
rect 9873 -30997 9885 -30933
rect 9545 -31260 9709 -31244
rect 9545 -31294 9658 -31260
rect 9692 -31294 9709 -31260
rect 9545 -31310 9709 -31294
rect 9775 -31341 9885 -30997
rect 9917 -30961 9983 -30773
rect 10029 -30909 10113 -30158
rect 10148 -30909 10187 -30158
rect 10029 -30921 10187 -30909
rect 10221 -30921 10228 -30145
rect 10029 -30933 10228 -30921
rect 10565 -30145 10815 -30133
rect 10565 -30921 10571 -30145
rect 10605 -30918 10815 -30145
rect 11134 -30146 11155 -29994
rect 11492 -29218 11743 -29206
rect 11492 -29994 11498 -29218
rect 11532 -29221 11743 -29218
rect 11860 -28835 13092 -28611
rect 11860 -29038 12189 -28835
rect 12410 -29038 13092 -28835
rect 11532 -29977 11742 -29221
rect 11860 -29536 13092 -29038
rect 11799 -29544 13092 -29536
rect 11799 -29595 11811 -29544
rect 12168 -29553 13092 -29544
rect 12168 -29595 12180 -29553
rect 11799 -29602 12180 -29595
rect 11860 -29640 11903 -29602
rect 12726 -29687 13092 -29553
rect 11875 -29699 12689 -29687
rect 12726 -29694 13137 -29687
rect 11875 -29789 11881 -29699
rect 11915 -29789 12073 -29699
rect 12107 -29789 12265 -29699
rect 12299 -29789 12457 -29699
rect 12491 -29789 12649 -29699
rect 12683 -29789 12689 -29699
rect 11875 -29801 12689 -29789
rect 12923 -29731 13137 -29694
rect 12923 -29765 12986 -29731
rect 13077 -29765 13137 -29731
rect 12923 -29803 13137 -29765
rect 11779 -29841 12209 -29829
rect 11779 -29931 11785 -29841
rect 11819 -29931 11977 -29841
rect 12011 -29931 12169 -29841
rect 12203 -29931 12209 -29841
rect 11779 -29943 12209 -29931
rect 12355 -29835 12827 -29829
rect 12355 -29841 12892 -29835
rect 12355 -29931 12361 -29841
rect 12395 -29931 12553 -29841
rect 12587 -29931 12745 -29841
rect 12779 -29851 12892 -29841
rect 12779 -29931 12842 -29851
rect 12355 -29943 12842 -29931
rect 11532 -29993 12263 -29977
rect 11532 -29994 12170 -29993
rect 11492 -30006 12170 -29994
rect 11737 -30027 12170 -30006
rect 12204 -30027 12263 -29993
rect 11737 -30043 12263 -30027
rect 12702 -30077 12842 -29943
rect 12876 -30077 12892 -29851
rect 12923 -29837 12929 -29803
rect 13008 -29807 13137 -29803
rect 13008 -29837 13014 -29807
rect 12923 -29995 13014 -29837
rect 12923 -30029 12929 -29995
rect 13008 -30029 13014 -29995
rect 12923 -30045 13014 -30029
rect 13046 -29899 13235 -29835
rect 13046 -29933 13052 -29899
rect 13129 -29933 13235 -29899
rect 13046 -30040 13235 -29933
rect 15447 -30040 15513 -19790
rect 15617 -19834 16719 -19818
rect 15617 -19868 16669 -19834
rect 16703 -19868 16719 -19834
rect 15617 -19884 16719 -19868
rect 11703 -30098 12363 -30082
rect 11703 -30132 12313 -30098
rect 12347 -30132 12363 -30098
rect 11703 -30134 12363 -30132
rect 10956 -30910 11040 -30159
rect 11075 -30910 11114 -30159
rect 10605 -30921 10816 -30918
rect 10565 -30933 10816 -30921
rect 9917 -31027 10542 -30961
rect 9917 -31063 10372 -31055
rect 9917 -31121 10264 -31063
rect 10224 -31123 10264 -31121
rect 10324 -31123 10372 -31063
rect 9917 -31215 9937 -31149
rect 10003 -31215 10185 -31149
rect 10224 -31206 10372 -31123
rect 10119 -31243 10185 -31215
rect 10306 -31242 10372 -31206
rect 10409 -31242 10443 -31241
rect 9917 -31253 10063 -31243
rect 9917 -31305 9951 -31253
rect 10016 -31259 10063 -31253
rect 10047 -31293 10063 -31259
rect 10016 -31305 10063 -31293
rect 9917 -31309 10063 -31305
rect 10119 -31259 10256 -31243
rect 10119 -31293 10205 -31259
rect 10239 -31293 10256 -31259
rect 10119 -31309 10256 -31293
rect 10306 -31259 10447 -31242
rect 10306 -31293 10397 -31259
rect 10431 -31293 10447 -31259
rect 10306 -31308 10447 -31293
rect 10476 -31243 10542 -31027
rect 10476 -31259 10640 -31243
rect 10476 -31293 10589 -31259
rect 10623 -31293 10640 -31259
rect 10476 -31309 10640 -31293
rect 10706 -31244 10816 -30933
rect 10956 -30922 11114 -30910
rect 11148 -30922 11155 -30146
rect 10956 -30934 11155 -30922
rect 11492 -30146 12363 -30134
rect 11492 -30922 11498 -30146
rect 11532 -30148 12363 -30146
rect 11532 -30179 11815 -30148
rect 11532 -30919 11742 -30179
rect 12259 -30182 12305 -30176
rect 12702 -30182 12892 -30077
rect 13046 -30091 15513 -30040
rect 12259 -30188 12892 -30182
rect 12259 -30364 12265 -30188
rect 12299 -30297 12892 -30188
rect 12923 -30125 13052 -30091
rect 13129 -30106 15513 -30091
rect 13129 -30125 13235 -30106
rect 12923 -30253 13235 -30125
rect 12923 -30287 12935 -30253
rect 13111 -30287 13235 -30253
rect 12923 -30293 13123 -30287
rect 12299 -30331 12842 -30297
rect 12876 -30331 12892 -30297
rect 12299 -30348 12892 -30331
rect 12923 -30341 13123 -30334
rect 12299 -30364 12827 -30348
rect 12259 -30376 12827 -30364
rect 12305 -30380 12827 -30376
rect 12923 -30375 12935 -30341
rect 13111 -30375 13123 -30341
rect 13151 -30348 13235 -30287
rect 12305 -30381 12825 -30380
rect 12305 -30382 12774 -30381
rect 12171 -30447 12394 -30440
rect 12171 -30495 12183 -30447
rect 12074 -30508 12183 -30495
rect 12382 -30495 12394 -30447
rect 12923 -30443 13123 -30375
rect 12923 -30477 12954 -30443
rect 13086 -30477 13123 -30443
rect 12921 -30484 13123 -30477
rect 12382 -30508 12473 -30495
rect 12074 -30611 12233 -30508
rect 12352 -30611 12473 -30508
rect 12921 -30533 13121 -30484
rect 12921 -30555 12960 -30533
rect 12074 -30685 12473 -30611
rect 12923 -30652 12960 -30555
rect 13079 -30555 13121 -30533
rect 13079 -30652 13113 -30555
rect 12923 -30710 13113 -30652
rect 11532 -30922 11743 -30919
rect 11492 -30934 11743 -30922
rect 10844 -31028 10850 -30962
rect 10916 -31028 11469 -30962
rect 10844 -31122 10888 -31056
rect 10954 -31122 11299 -31056
rect 10844 -31216 10859 -31150
rect 10925 -31216 11112 -31150
rect 11151 -31207 11299 -31122
rect 11046 -31244 11112 -31216
rect 11233 -31243 11299 -31207
rect 11336 -31243 11370 -31242
rect 10706 -31260 10990 -31244
rect 10706 -31294 10940 -31260
rect 10974 -31294 10990 -31260
rect 10706 -31310 10990 -31294
rect 11046 -31260 11183 -31244
rect 11046 -31294 11132 -31260
rect 11166 -31294 11183 -31260
rect 11046 -31310 11183 -31294
rect 11233 -31260 11374 -31243
rect 11233 -31294 11324 -31260
rect 11358 -31294 11374 -31260
rect 11233 -31309 11374 -31294
rect 11403 -31244 11469 -31028
rect 11403 -31260 11567 -31244
rect 11403 -31294 11516 -31260
rect 11550 -31294 11567 -31260
rect 11403 -31310 11567 -31294
rect 10706 -31340 10816 -31310
rect 7138 -31348 8001 -31341
rect 7138 -31460 7245 -31348
rect 7280 -31460 7438 -31348
rect 7473 -31460 7630 -31348
rect 7665 -31460 7822 -31348
rect 7857 -31460 8001 -31348
rect 7138 -31475 8001 -31460
rect 8086 -31348 8949 -31341
rect 8086 -31460 8193 -31348
rect 8228 -31460 8386 -31348
rect 8421 -31460 8578 -31348
rect 8613 -31460 8770 -31348
rect 8805 -31460 8949 -31348
rect 8086 -31475 8949 -31460
rect 9022 -31348 9885 -31341
rect 9022 -31460 9129 -31348
rect 9164 -31460 9322 -31348
rect 9357 -31460 9514 -31348
rect 9549 -31460 9706 -31348
rect 9741 -31460 9885 -31348
rect 9022 -31475 9885 -31460
rect 9953 -31347 10816 -31340
rect 11633 -31341 11743 -30934
rect 9953 -31459 10060 -31347
rect 10095 -31459 10253 -31347
rect 10288 -31459 10445 -31347
rect 10480 -31459 10637 -31347
rect 10672 -31459 10816 -31347
rect 9953 -31474 10816 -31459
rect 10880 -31348 11743 -31341
rect 10880 -31460 10987 -31348
rect 11022 -31460 11180 -31348
rect 11215 -31460 11372 -31348
rect 11407 -31460 11564 -31348
rect 11599 -31460 11743 -31348
rect 10880 -31475 11743 -31460
rect 7137 -31537 10779 -31528
rect 11883 -31529 12147 -31518
rect 7137 -31538 9965 -31537
rect 7137 -31648 7150 -31538
rect 7184 -31648 7342 -31538
rect 7376 -31648 7534 -31538
rect 7568 -31648 7726 -31538
rect 7760 -31648 7918 -31538
rect 7952 -31648 8098 -31538
rect 8132 -31648 8290 -31538
rect 8324 -31648 8482 -31538
rect 8516 -31648 8674 -31538
rect 8708 -31648 8866 -31538
rect 8900 -31648 9034 -31538
rect 9068 -31648 9226 -31538
rect 9260 -31648 9418 -31538
rect 9452 -31648 9610 -31538
rect 9644 -31648 9802 -31538
rect 9836 -31647 9965 -31538
rect 9999 -31647 10157 -31537
rect 10191 -31647 10349 -31537
rect 10383 -31647 10541 -31537
rect 10575 -31647 10733 -31537
rect 10767 -31647 10779 -31537
rect 9836 -31648 10779 -31647
rect 7137 -31719 10779 -31648
rect 10880 -31538 11894 -31529
rect 10880 -31648 10892 -31538
rect 10926 -31648 11084 -31538
rect 11118 -31648 11276 -31538
rect 11310 -31648 11468 -31538
rect 11502 -31648 11660 -31538
rect 11694 -31648 11894 -31538
rect 10880 -31659 11894 -31648
rect 7137 -31720 10204 -31719
rect 7137 -31755 7389 -31720
rect 7677 -31755 8337 -31720
rect 8625 -31755 9273 -31720
rect 9561 -31754 10204 -31720
rect 10492 -31754 10779 -31719
rect 9561 -31755 10779 -31754
rect 7137 -31769 10779 -31755
rect 7137 -31771 7964 -31769
rect 8085 -31771 8912 -31769
rect 9021 -31771 9848 -31769
rect 9952 -31770 10779 -31769
rect 10879 -31720 11894 -31659
rect 10879 -31755 11131 -31720
rect 11419 -31755 11894 -31720
rect 10879 -31771 11894 -31755
rect 12136 -31771 12147 -31529
rect 11883 -31782 12147 -31771
rect 5658 -32241 7357 -32197
rect 5658 -32275 5721 -32241
rect 5812 -32275 6161 -32241
rect 6252 -32275 6601 -32241
rect 6692 -32275 7357 -32241
rect 5658 -32287 7357 -32275
rect 5658 -32313 5872 -32287
rect 5558 -32345 5627 -32339
rect 5558 -32587 5577 -32414
rect 5611 -32587 5627 -32414
rect 5658 -32347 5664 -32313
rect 5743 -32317 5872 -32313
rect 6098 -32313 6312 -32287
rect 5743 -32347 5749 -32317
rect 5998 -32345 6067 -32339
rect 5658 -32505 5749 -32347
rect 5658 -32539 5664 -32505
rect 5743 -32539 5749 -32505
rect 5658 -32555 5749 -32539
rect 5781 -32409 5970 -32345
rect 5781 -32443 5787 -32409
rect 5864 -32443 5970 -32409
rect 5558 -32689 5627 -32587
rect 5781 -32601 5970 -32443
rect 5658 -32635 5787 -32601
rect 5864 -32635 5970 -32601
rect 5558 -32807 5628 -32689
rect 5658 -32763 5970 -32635
rect 5658 -32797 5670 -32763
rect 5846 -32797 5970 -32763
rect 5658 -32803 5858 -32797
rect 5558 -32841 5577 -32807
rect 5611 -32841 5628 -32807
rect 5558 -32858 5628 -32841
rect 5559 -32935 5628 -32858
rect 5558 -32994 5628 -32935
rect 5658 -32851 5858 -32844
rect 5658 -32885 5670 -32851
rect 5846 -32885 5858 -32851
rect 5886 -32858 5970 -32797
rect 5658 -32953 5858 -32885
rect 5658 -32987 5689 -32953
rect 5821 -32987 5858 -32953
rect 5658 -32994 5858 -32987
rect 5901 -32910 5970 -32858
rect 5559 -33110 5628 -32994
rect 5703 -32996 5823 -32994
rect 5703 -33048 5734 -32996
rect 5786 -33048 5823 -32996
rect 5901 -33000 5970 -32979
rect 5998 -32587 6017 -32414
rect 6051 -32587 6067 -32414
rect 6098 -32347 6104 -32313
rect 6183 -32317 6312 -32313
rect 6538 -32300 7357 -32287
rect 6538 -32313 6752 -32300
rect 6183 -32347 6189 -32317
rect 6438 -32345 6507 -32339
rect 6098 -32505 6189 -32347
rect 6098 -32539 6104 -32505
rect 6183 -32539 6189 -32505
rect 6098 -32555 6189 -32539
rect 6221 -32409 6410 -32345
rect 6221 -32443 6227 -32409
rect 6304 -32443 6410 -32409
rect 5998 -32807 6067 -32587
rect 6221 -32601 6410 -32443
rect 6098 -32635 6227 -32601
rect 6304 -32635 6410 -32601
rect 6098 -32763 6410 -32635
rect 6098 -32797 6110 -32763
rect 6286 -32797 6410 -32763
rect 6098 -32803 6298 -32797
rect 5998 -32841 6017 -32807
rect 6051 -32841 6067 -32807
rect 5703 -33079 5823 -33048
rect 5559 -33179 5901 -33110
rect 5559 -33191 5628 -33179
rect 5425 -33777 5491 -33771
rect 3663 -33801 3729 -33795
rect -413 -33867 3663 -33801
rect -11291 -34073 -11279 -34039
rect -11245 -34073 -11223 -34039
rect -11291 -34231 -11223 -34073
rect -11092 -34118 -11070 -33867
rect -11195 -34135 -11070 -34118
rect -11195 -34169 -11178 -34135
rect -11144 -34169 -11070 -34135
rect -11195 -34183 -11070 -34169
rect -11291 -34265 -11279 -34231
rect -11245 -34265 -11223 -34231
rect -11291 -34281 -11223 -34265
rect -11092 -34313 -11070 -34183
rect -11925 -34361 -11903 -34327
rect -11801 -34361 -11778 -34327
rect -11925 -34373 -11778 -34361
rect -12612 -34504 -11498 -34498
rect -12612 -34576 -12582 -34504
rect -12510 -34528 -11498 -34504
rect -12510 -34571 -11553 -34528
rect -11510 -34571 -11498 -34528
rect -12510 -34576 -11498 -34571
rect -12612 -34583 -11498 -34576
rect -11464 -34666 -11321 -34314
rect -11280 -34327 -11070 -34313
rect -11024 -34327 -11001 -33867
rect 3663 -33873 3729 -33867
rect -11280 -34361 -11264 -34327
rect -11158 -34361 -11001 -34327
rect -11280 -34368 -11001 -34361
rect -12612 -34670 -11321 -34666
rect -12746 -34671 -11321 -34670
rect -12746 -34760 -12726 -34671
rect -12637 -34758 -11321 -34671
rect -12637 -34760 -12476 -34758
rect 5832 -35772 5901 -33179
rect 5998 -33443 6067 -32841
rect 6098 -32851 6298 -32844
rect 6098 -32885 6110 -32851
rect 6286 -32885 6298 -32851
rect 6326 -32858 6410 -32797
rect 6098 -32953 6298 -32885
rect 6098 -32987 6129 -32953
rect 6261 -32987 6298 -32953
rect 6098 -32994 6172 -32987
rect 6143 -33029 6172 -32994
rect 6224 -32994 6298 -32987
rect 6341 -32912 6410 -32858
rect 6341 -32994 6410 -32981
rect 6438 -32587 6457 -32414
rect 6491 -32587 6507 -32414
rect 6538 -32347 6544 -32313
rect 6623 -32317 6752 -32313
rect 6623 -32347 6629 -32317
rect 6538 -32505 6629 -32347
rect 6538 -32539 6544 -32505
rect 6623 -32539 6629 -32505
rect 6538 -32555 6629 -32539
rect 6661 -32409 6850 -32345
rect 6661 -32443 6667 -32409
rect 6744 -32443 6850 -32409
rect 6438 -32807 6507 -32587
rect 6661 -32601 6850 -32443
rect 6538 -32635 6667 -32601
rect 6744 -32635 6850 -32601
rect 6538 -32763 6850 -32635
rect 6538 -32797 6550 -32763
rect 6726 -32797 6850 -32763
rect 6538 -32803 6738 -32797
rect 6438 -32841 6457 -32807
rect 6491 -32841 6507 -32807
rect 6224 -33029 6263 -32994
rect 6143 -33054 6263 -33029
rect 5992 -33449 6073 -33443
rect 5992 -33518 5998 -33449
rect 6067 -33452 6073 -33449
rect 6067 -33518 6085 -33452
rect 5992 -33524 6073 -33518
rect 5998 -35678 6067 -33524
rect 6438 -33584 6507 -32841
rect 6538 -32851 6738 -32844
rect 6538 -32885 6550 -32851
rect 6726 -32885 6738 -32851
rect 6766 -32858 6850 -32797
rect 6538 -32953 6738 -32885
rect 6781 -32903 6850 -32858
rect 7254 -32897 7357 -32300
rect 11860 -32897 12409 -32896
rect 12750 -32897 13092 -32896
rect 6538 -32987 6569 -32953
rect 6701 -32987 6738 -32953
rect 6538 -32994 6612 -32987
rect 6580 -33020 6612 -32994
rect 6664 -32994 6738 -32987
rect 6780 -32934 6850 -32903
rect 7137 -32898 7964 -32897
rect 8085 -32898 8912 -32897
rect 9021 -32898 9848 -32897
rect 9952 -32898 10779 -32897
rect 7137 -32913 10780 -32898
rect 6664 -33020 6700 -32994
rect 6580 -33063 6700 -33020
rect 6438 -33659 6507 -33653
rect 6780 -33546 6849 -32934
rect 7137 -32948 7389 -32913
rect 7677 -32948 8337 -32913
rect 8625 -32948 9273 -32913
rect 9561 -32948 10204 -32913
rect 10492 -32948 10780 -32913
rect 7137 -33009 10780 -32948
rect 10879 -32913 13092 -32897
rect 10879 -32948 11131 -32913
rect 11419 -32948 13092 -32913
rect 10879 -33009 13092 -32948
rect 7138 -33020 10780 -33009
rect 7138 -33130 7150 -33020
rect 7184 -33130 7342 -33020
rect 7376 -33130 7534 -33020
rect 7568 -33130 7726 -33020
rect 7760 -33130 7918 -33020
rect 7952 -33130 8098 -33020
rect 8132 -33130 8290 -33020
rect 8324 -33130 8482 -33020
rect 8516 -33130 8674 -33020
rect 8708 -33130 8866 -33020
rect 8900 -33130 9034 -33020
rect 9068 -33130 9226 -33020
rect 9260 -33130 9418 -33020
rect 9452 -33130 9610 -33020
rect 9644 -33130 9802 -33020
rect 9836 -33130 9965 -33020
rect 9999 -33130 10157 -33020
rect 10191 -33130 10349 -33020
rect 10383 -33130 10541 -33020
rect 10575 -33130 10733 -33020
rect 10767 -33130 10780 -33020
rect 7138 -33139 10780 -33130
rect 10880 -33020 13092 -33009
rect 10880 -33130 10892 -33020
rect 10926 -33130 11084 -33020
rect 11118 -33130 11276 -33020
rect 11310 -33130 11468 -33020
rect 11502 -33130 11660 -33020
rect 11694 -33130 13092 -33020
rect 10880 -33139 13092 -33130
rect 7138 -33208 8001 -33193
rect 7138 -33320 7245 -33208
rect 7280 -33320 7438 -33208
rect 7473 -33320 7630 -33208
rect 7665 -33320 7822 -33208
rect 7857 -33320 8001 -33208
rect 7138 -33327 8001 -33320
rect 8086 -33208 8949 -33193
rect 8086 -33320 8193 -33208
rect 8228 -33320 8386 -33208
rect 8421 -33320 8578 -33208
rect 8613 -33320 8770 -33208
rect 8805 -33320 8949 -33208
rect 8086 -33327 8949 -33320
rect 9022 -33208 9885 -33193
rect 9022 -33320 9129 -33208
rect 9164 -33320 9322 -33208
rect 9357 -33320 9514 -33208
rect 9549 -33320 9706 -33208
rect 9741 -33320 9885 -33208
rect 9022 -33327 9885 -33320
rect 9953 -33208 10816 -33193
rect 9953 -33320 10060 -33208
rect 10095 -33320 10253 -33208
rect 10288 -33320 10445 -33208
rect 10480 -33320 10637 -33208
rect 10672 -33320 10816 -33208
rect 9953 -33327 10816 -33320
rect 10880 -33208 11743 -33193
rect 10880 -33320 10987 -33208
rect 11022 -33320 11180 -33208
rect 11215 -33320 11372 -33208
rect 11407 -33320 11564 -33208
rect 11599 -33320 11743 -33208
rect 10880 -33327 11743 -33320
rect 7106 -33358 7158 -33357
rect 7102 -33363 7248 -33358
rect 7102 -33415 7106 -33363
rect 7158 -33374 7248 -33363
rect 7158 -33408 7198 -33374
rect 7232 -33408 7248 -33374
rect 7158 -33415 7248 -33408
rect 7102 -33424 7248 -33415
rect 7304 -33374 7441 -33358
rect 7304 -33408 7390 -33374
rect 7424 -33408 7441 -33374
rect 7304 -33424 7441 -33408
rect 7491 -33374 7632 -33359
rect 7491 -33408 7582 -33374
rect 7616 -33408 7632 -33374
rect 7304 -33452 7370 -33424
rect 7097 -33457 7370 -33452
rect 7097 -33509 7113 -33457
rect 7165 -33509 7370 -33457
rect 7491 -33425 7632 -33408
rect 7661 -33374 7825 -33358
rect 7661 -33408 7774 -33374
rect 7808 -33408 7825 -33374
rect 7661 -33424 7825 -33408
rect 7491 -33461 7557 -33425
rect 7594 -33426 7628 -33425
rect 7097 -33518 7370 -33509
rect 7409 -33546 7557 -33461
rect 6780 -33612 7327 -33546
rect 7393 -33612 7557 -33546
rect 6780 -35575 6849 -33612
rect 7661 -33640 7727 -33424
rect 7102 -33706 7727 -33640
rect 7106 -33907 7172 -33706
rect 7891 -33734 8001 -33327
rect 8050 -33364 8196 -33358
rect 8050 -33416 8069 -33364
rect 8122 -33374 8196 -33364
rect 8122 -33408 8146 -33374
rect 8180 -33408 8196 -33374
rect 8122 -33416 8196 -33408
rect 8050 -33424 8196 -33416
rect 8252 -33374 8389 -33358
rect 8252 -33408 8338 -33374
rect 8372 -33408 8389 -33374
rect 8252 -33424 8389 -33408
rect 8439 -33374 8580 -33359
rect 8439 -33408 8530 -33374
rect 8564 -33408 8580 -33374
rect 8252 -33452 8318 -33424
rect 8050 -33456 8318 -33452
rect 8050 -33508 8057 -33456
rect 8109 -33508 8318 -33456
rect 8439 -33425 8580 -33408
rect 8609 -33374 8773 -33358
rect 8609 -33408 8722 -33374
rect 8756 -33408 8773 -33374
rect 8609 -33424 8773 -33408
rect 8439 -33461 8505 -33425
rect 8542 -33426 8576 -33425
rect 8050 -33518 8318 -33508
rect 8357 -33539 8505 -33461
rect 8357 -33546 8424 -33539
rect 8050 -33591 8424 -33546
rect 8493 -33591 8505 -33539
rect 8050 -33612 8505 -33591
rect 8609 -33640 8675 -33424
rect 7106 -33979 7172 -33973
rect 7214 -33746 7413 -33734
rect 7214 -33758 7372 -33746
rect 7214 -34509 7298 -33758
rect 7333 -34509 7372 -33758
rect 7214 -34687 7227 -34509
rect 7406 -34522 7413 -33746
rect 7405 -34674 7413 -34522
rect 7750 -33746 8001 -33734
rect 7750 -34522 7756 -33746
rect 7790 -33749 8001 -33746
rect 8050 -33706 8675 -33640
rect 7790 -34164 8000 -33749
rect 8050 -34011 8116 -33706
rect 8839 -33734 8949 -33327
rect 8986 -33363 9132 -33358
rect 8986 -33415 9002 -33363
rect 9055 -33374 9132 -33363
rect 9055 -33408 9082 -33374
rect 9116 -33408 9132 -33374
rect 9055 -33415 9132 -33408
rect 8986 -33424 9132 -33415
rect 9188 -33374 9325 -33358
rect 9188 -33408 9274 -33374
rect 9308 -33408 9325 -33374
rect 9188 -33424 9325 -33408
rect 9375 -33374 9516 -33359
rect 9375 -33408 9466 -33374
rect 9500 -33408 9516 -33374
rect 9188 -33452 9254 -33424
rect 8986 -33461 9254 -33452
rect 9375 -33425 9516 -33408
rect 9545 -33374 9709 -33358
rect 9545 -33408 9658 -33374
rect 9692 -33408 9709 -33374
rect 9545 -33424 9709 -33408
rect 9375 -33461 9441 -33425
rect 9478 -33426 9512 -33425
rect 8986 -33513 9000 -33461
rect 9052 -33513 9254 -33461
rect 8986 -33518 9254 -33513
rect 9293 -33546 9441 -33461
rect 8986 -33552 9441 -33546
rect 8986 -33605 8989 -33552
rect 9042 -33605 9441 -33552
rect 8986 -33612 9441 -33605
rect 9545 -33640 9611 -33424
rect 8050 -34083 8116 -34077
rect 8162 -33746 8361 -33734
rect 8162 -33758 8320 -33746
rect 7790 -34230 7872 -34164
rect 7938 -34230 8000 -34164
rect 7790 -34522 8000 -34230
rect 7750 -34534 8000 -34522
rect 8162 -34509 8246 -33758
rect 8281 -34509 8320 -33758
rect 8354 -34522 8361 -33746
rect 7102 -35333 7168 -35327
rect 7102 -35490 7168 -35399
rect 7214 -35438 7298 -34687
rect 7333 -35438 7372 -34687
rect 7214 -35450 7372 -35438
rect 7406 -35450 7413 -34674
rect 7214 -35462 7413 -35450
rect 7750 -34674 8000 -34662
rect 7750 -35450 7756 -34674
rect 7790 -34957 8000 -34674
rect 7790 -35023 7853 -34957
rect 7919 -35023 8000 -34957
rect 7790 -35447 8000 -35023
rect 8340 -34674 8361 -34522
rect 8698 -33746 8949 -33734
rect 8698 -34522 8704 -33746
rect 8738 -33749 8949 -33746
rect 8986 -33705 9611 -33640
rect 8738 -33910 8948 -33749
rect 9052 -33706 9611 -33705
rect 9775 -33662 9885 -33327
rect 10706 -33358 10816 -33327
rect 9917 -33363 10063 -33358
rect 9917 -33415 9933 -33363
rect 9986 -33374 10063 -33363
rect 9986 -33408 10013 -33374
rect 10047 -33408 10063 -33374
rect 9986 -33415 10063 -33408
rect 9917 -33424 10063 -33415
rect 10119 -33374 10256 -33358
rect 10119 -33408 10205 -33374
rect 10239 -33408 10256 -33374
rect 10119 -33424 10256 -33408
rect 10306 -33374 10447 -33359
rect 10306 -33408 10397 -33374
rect 10431 -33408 10447 -33374
rect 10119 -33452 10185 -33424
rect 9917 -33461 10185 -33452
rect 10306 -33425 10447 -33408
rect 10476 -33374 10640 -33358
rect 10476 -33408 10589 -33374
rect 10623 -33408 10640 -33374
rect 10476 -33424 10640 -33408
rect 10706 -33374 10990 -33358
rect 10706 -33408 10940 -33374
rect 10974 -33408 10990 -33374
rect 10706 -33424 10990 -33408
rect 11046 -33374 11183 -33358
rect 11046 -33408 11132 -33374
rect 11166 -33408 11183 -33374
rect 11046 -33424 11183 -33408
rect 11233 -33374 11374 -33359
rect 11233 -33408 11324 -33374
rect 11358 -33408 11374 -33374
rect 10306 -33461 10372 -33425
rect 10409 -33426 10443 -33425
rect 9917 -33513 9935 -33461
rect 9987 -33513 10185 -33461
rect 9917 -33518 10185 -33513
rect 10224 -33508 10372 -33461
rect 10224 -33546 10262 -33508
rect 9917 -33577 10262 -33546
rect 10331 -33577 10372 -33508
rect 9917 -33612 10372 -33577
rect 10476 -33640 10542 -33424
rect 9775 -33728 9798 -33662
rect 9864 -33728 9885 -33662
rect 9775 -33734 9885 -33728
rect 8986 -33789 9052 -33771
rect 9098 -33746 9297 -33734
rect 9098 -33758 9256 -33746
rect 8738 -33976 8818 -33910
rect 8884 -33976 8948 -33910
rect 8738 -34522 8948 -33976
rect 8698 -34534 8948 -34522
rect 9098 -34509 9182 -33758
rect 9217 -34509 9256 -33758
rect 9290 -34522 9297 -33746
rect 8162 -35438 8246 -34687
rect 8281 -35438 8320 -34687
rect 7790 -35450 8001 -35447
rect 7750 -35462 8001 -35450
rect 7102 -35556 7727 -35490
rect 6774 -35644 6780 -35575
rect 6849 -35584 6855 -35575
rect 6849 -35644 7557 -35584
rect 6780 -35650 7557 -35644
rect 5998 -35742 6066 -35678
rect 5999 -35744 6066 -35742
rect 6132 -35744 7370 -35678
rect 7409 -35735 7557 -35650
rect 7304 -35772 7370 -35744
rect 7491 -35771 7557 -35735
rect 7594 -35771 7628 -35770
rect 5832 -35838 6941 -35772
rect 7007 -35788 7248 -35772
rect 7007 -35822 7198 -35788
rect 7232 -35822 7248 -35788
rect 7007 -35838 7248 -35822
rect 7304 -35788 7441 -35772
rect 7304 -35822 7390 -35788
rect 7424 -35822 7441 -35788
rect 7304 -35838 7441 -35822
rect 7491 -35788 7632 -35771
rect 7491 -35822 7582 -35788
rect 7616 -35822 7632 -35788
rect 7491 -35837 7632 -35822
rect 7661 -35772 7727 -35556
rect 7661 -35788 7825 -35772
rect 7661 -35822 7774 -35788
rect 7808 -35822 7825 -35788
rect 7661 -35838 7825 -35822
rect 5832 -35848 5901 -35838
rect 7891 -35869 8001 -35462
rect 8050 -35454 8116 -35448
rect 8162 -35450 8320 -35438
rect 8354 -35450 8361 -34674
rect 8162 -35462 8361 -35450
rect 8698 -34674 8948 -34662
rect 8698 -35450 8704 -34674
rect 8738 -35367 8948 -34674
rect 9276 -34674 9297 -34522
rect 9634 -33746 9885 -33734
rect 9634 -34522 9640 -33746
rect 9674 -33749 9885 -33746
rect 9917 -33706 10542 -33640
rect 9674 -34522 9884 -33749
rect 9917 -33801 9983 -33706
rect 10706 -33734 10816 -33424
rect 11046 -33452 11112 -33424
rect 10844 -33518 10860 -33452
rect 10926 -33518 11112 -33452
rect 11233 -33425 11374 -33408
rect 11403 -33374 11567 -33358
rect 11403 -33408 11516 -33374
rect 11550 -33408 11567 -33374
rect 11403 -33424 11567 -33408
rect 11233 -33461 11299 -33425
rect 11336 -33426 11370 -33425
rect 11151 -33546 11299 -33461
rect 10844 -33612 10858 -33546
rect 10924 -33612 11299 -33546
rect 11403 -33640 11469 -33424
rect 10844 -33706 10850 -33640
rect 10915 -33706 11469 -33640
rect 11633 -33734 11743 -33327
rect 9917 -33873 9983 -33867
rect 10029 -33746 10228 -33734
rect 10029 -33758 10187 -33746
rect 9634 -34534 9884 -34522
rect 10029 -34509 10113 -33758
rect 10148 -34509 10187 -33758
rect 10221 -34522 10228 -33746
rect 8738 -35433 8837 -35367
rect 8903 -35433 8948 -35367
rect 8738 -35447 8948 -35433
rect 8989 -35113 9055 -35107
rect 8738 -35450 8949 -35447
rect 8698 -35462 8949 -35450
rect 8116 -35520 8675 -35490
rect 8050 -35556 8675 -35520
rect 8050 -35591 8505 -35584
rect 8050 -35650 8401 -35591
rect 8357 -35655 8401 -35650
rect 8465 -35655 8505 -35591
rect 8050 -35687 8318 -35678
rect 8050 -35739 8079 -35687
rect 8131 -35739 8318 -35687
rect 8357 -35735 8505 -35655
rect 8050 -35744 8318 -35739
rect 8252 -35772 8318 -35744
rect 8439 -35771 8505 -35735
rect 8542 -35771 8576 -35770
rect 8050 -35781 8196 -35772
rect 8050 -35833 8063 -35781
rect 8128 -35788 8196 -35781
rect 8128 -35822 8146 -35788
rect 8180 -35822 8196 -35788
rect 8128 -35833 8196 -35822
rect 8050 -35838 8196 -35833
rect 8252 -35788 8389 -35772
rect 8252 -35822 8338 -35788
rect 8372 -35822 8389 -35788
rect 8252 -35838 8389 -35822
rect 8439 -35788 8580 -35771
rect 8439 -35822 8530 -35788
rect 8564 -35822 8580 -35788
rect 8439 -35837 8580 -35822
rect 8609 -35772 8675 -35556
rect 8609 -35788 8773 -35772
rect 8609 -35822 8722 -35788
rect 8756 -35822 8773 -35788
rect 8609 -35838 8773 -35822
rect 8839 -35869 8949 -35462
rect 8989 -35490 9055 -35179
rect 9098 -35438 9182 -34687
rect 9217 -35438 9256 -34687
rect 9098 -35450 9256 -35438
rect 9290 -35450 9297 -34674
rect 9098 -35462 9297 -35450
rect 9634 -34674 9884 -34662
rect 9634 -35450 9640 -34674
rect 9674 -35447 9884 -34674
rect 10206 -34673 10228 -34522
rect 10565 -33746 10816 -33734
rect 10565 -34522 10571 -33746
rect 10605 -33749 10816 -33746
rect 10956 -33746 11155 -33734
rect 10605 -34522 10815 -33749
rect 10565 -34534 10815 -34522
rect 10956 -33758 11114 -33746
rect 10956 -34509 11040 -33758
rect 11075 -34509 11114 -33758
rect 11148 -34522 11155 -33746
rect 9917 -35235 9983 -35229
rect 9674 -35450 9885 -35447
rect 9634 -35461 9885 -35450
rect 9634 -35462 9807 -35461
rect 8986 -35556 9611 -35490
rect 8986 -35650 8993 -35584
rect 9059 -35650 9441 -35584
rect 8986 -35744 9001 -35678
rect 9067 -35744 9254 -35678
rect 9293 -35735 9441 -35650
rect 9188 -35772 9254 -35744
rect 9375 -35771 9441 -35735
rect 9478 -35771 9512 -35770
rect 8986 -35781 9132 -35772
rect 8986 -35833 8992 -35781
rect 9057 -35788 9132 -35781
rect 9057 -35822 9082 -35788
rect 9116 -35822 9132 -35788
rect 9057 -35833 9132 -35822
rect 8986 -35838 9132 -35833
rect 9188 -35788 9325 -35772
rect 9188 -35822 9274 -35788
rect 9308 -35822 9325 -35788
rect 9188 -35838 9325 -35822
rect 9375 -35788 9516 -35771
rect 9375 -35822 9466 -35788
rect 9500 -35822 9516 -35788
rect 9375 -35837 9516 -35822
rect 9545 -35772 9611 -35556
rect 9775 -35525 9807 -35462
rect 9873 -35525 9885 -35461
rect 9545 -35788 9709 -35772
rect 9545 -35822 9658 -35788
rect 9692 -35822 9709 -35788
rect 9545 -35838 9709 -35822
rect 9775 -35869 9885 -35525
rect 9917 -35489 9983 -35301
rect 10029 -35437 10113 -34686
rect 10148 -35437 10187 -34686
rect 10029 -35449 10187 -35437
rect 10221 -35449 10228 -34673
rect 10029 -35461 10228 -35449
rect 10565 -34673 10815 -34661
rect 10565 -35449 10571 -34673
rect 10605 -35446 10815 -34673
rect 11134 -34674 11155 -34522
rect 11492 -33746 11743 -33734
rect 11492 -34522 11498 -33746
rect 11532 -33749 11743 -33746
rect 11860 -33363 13092 -33139
rect 11860 -33566 12189 -33363
rect 12410 -33566 13092 -33363
rect 11532 -34505 11742 -33749
rect 11860 -34064 13092 -33566
rect 11799 -34072 13092 -34064
rect 11799 -34123 11811 -34072
rect 12168 -34081 13092 -34072
rect 12168 -34123 12180 -34081
rect 11799 -34130 12180 -34123
rect 11860 -34168 11903 -34130
rect 12726 -34215 13092 -34081
rect 11875 -34227 12689 -34215
rect 12726 -34222 13137 -34215
rect 11875 -34317 11881 -34227
rect 11915 -34317 12073 -34227
rect 12107 -34317 12265 -34227
rect 12299 -34317 12457 -34227
rect 12491 -34317 12649 -34227
rect 12683 -34317 12689 -34227
rect 11875 -34329 12689 -34317
rect 12923 -34259 13137 -34222
rect 12923 -34293 12986 -34259
rect 13077 -34293 13137 -34259
rect 12923 -34331 13137 -34293
rect 11779 -34369 12209 -34357
rect 11779 -34459 11785 -34369
rect 11819 -34459 11977 -34369
rect 12011 -34459 12169 -34369
rect 12203 -34459 12209 -34369
rect 11779 -34471 12209 -34459
rect 12355 -34363 12827 -34357
rect 12355 -34369 12892 -34363
rect 12355 -34459 12361 -34369
rect 12395 -34459 12553 -34369
rect 12587 -34459 12745 -34369
rect 12779 -34379 12892 -34369
rect 12779 -34459 12842 -34379
rect 12355 -34471 12842 -34459
rect 11532 -34521 12263 -34505
rect 11532 -34522 12170 -34521
rect 11492 -34534 12170 -34522
rect 11737 -34555 12170 -34534
rect 12204 -34555 12263 -34521
rect 11737 -34571 12263 -34555
rect 12702 -34605 12842 -34471
rect 12876 -34605 12892 -34379
rect 12923 -34365 12929 -34331
rect 13008 -34335 13137 -34331
rect 13008 -34365 13014 -34335
rect 12923 -34523 13014 -34365
rect 12923 -34557 12929 -34523
rect 13008 -34557 13014 -34523
rect 12923 -34573 13014 -34557
rect 13046 -34427 13235 -34363
rect 13046 -34461 13052 -34427
rect 13129 -34461 13235 -34427
rect 13046 -34535 13235 -34461
rect 15619 -34535 15685 -19884
rect 16830 -19923 16967 -19607
rect 16249 -19935 16967 -19923
rect 16249 -20111 16255 -19935
rect 16289 -20111 16447 -19935
rect 16481 -20111 16967 -19935
rect 16249 -20123 16967 -20111
rect 16147 -20245 16221 -20177
rect 16480 -20245 16590 -20177
rect 16147 -20358 16211 -20245
rect 16541 -20358 16590 -20245
rect 16147 -20436 16221 -20358
rect 16480 -20436 16590 -20358
rect 11703 -34626 12363 -34610
rect 11703 -34660 12313 -34626
rect 12347 -34660 12363 -34626
rect 11703 -34662 12363 -34660
rect 10956 -35438 11040 -34687
rect 11075 -35438 11114 -34687
rect 10605 -35449 10816 -35446
rect 10565 -35461 10816 -35449
rect 9917 -35555 10542 -35489
rect 9917 -35591 10372 -35583
rect 9917 -35649 10264 -35591
rect 10224 -35651 10264 -35649
rect 10324 -35651 10372 -35591
rect 9917 -35743 9937 -35677
rect 10003 -35743 10185 -35677
rect 10224 -35734 10372 -35651
rect 10119 -35771 10185 -35743
rect 10306 -35770 10372 -35734
rect 10409 -35770 10443 -35769
rect 9917 -35781 10063 -35771
rect 9917 -35833 9951 -35781
rect 10016 -35787 10063 -35781
rect 10047 -35821 10063 -35787
rect 10016 -35833 10063 -35821
rect 9917 -35837 10063 -35833
rect 10119 -35787 10256 -35771
rect 10119 -35821 10205 -35787
rect 10239 -35821 10256 -35787
rect 10119 -35837 10256 -35821
rect 10306 -35787 10447 -35770
rect 10306 -35821 10397 -35787
rect 10431 -35821 10447 -35787
rect 10306 -35836 10447 -35821
rect 10476 -35771 10542 -35555
rect 10476 -35787 10640 -35771
rect 10476 -35821 10589 -35787
rect 10623 -35821 10640 -35787
rect 10476 -35837 10640 -35821
rect 10706 -35772 10816 -35461
rect 10956 -35450 11114 -35438
rect 11148 -35450 11155 -34674
rect 10956 -35462 11155 -35450
rect 11492 -34674 12363 -34662
rect 11492 -35450 11498 -34674
rect 11532 -34676 12363 -34674
rect 11532 -34707 11815 -34676
rect 11532 -35447 11742 -34707
rect 12259 -34710 12305 -34704
rect 12702 -34710 12892 -34605
rect 13046 -34601 15685 -34535
rect 13046 -34619 13235 -34601
rect 12259 -34716 12892 -34710
rect 12259 -34892 12265 -34716
rect 12299 -34825 12892 -34716
rect 12923 -34653 13052 -34619
rect 13129 -34653 13235 -34619
rect 12923 -34781 13235 -34653
rect 12923 -34815 12935 -34781
rect 13111 -34815 13235 -34781
rect 12923 -34821 13123 -34815
rect 12299 -34859 12842 -34825
rect 12876 -34859 12892 -34825
rect 12299 -34876 12892 -34859
rect 12923 -34869 13123 -34862
rect 12299 -34892 12827 -34876
rect 12259 -34904 12827 -34892
rect 12305 -34908 12827 -34904
rect 12923 -34903 12935 -34869
rect 13111 -34903 13123 -34869
rect 12305 -34909 12825 -34908
rect 12305 -34910 12774 -34909
rect 12171 -34975 12394 -34968
rect 12171 -35023 12183 -34975
rect 12074 -35036 12183 -35023
rect 12382 -35023 12394 -34975
rect 12923 -34971 13123 -34903
rect 12923 -35005 12954 -34971
rect 13086 -35005 13123 -34971
rect 12921 -35012 13123 -35005
rect 12382 -35036 12473 -35023
rect 12074 -35139 12233 -35036
rect 12352 -35139 12473 -35036
rect 12921 -35061 13121 -35012
rect 12921 -35083 12960 -35061
rect 12074 -35213 12473 -35139
rect 12923 -35180 12960 -35083
rect 13079 -35083 13121 -35061
rect 13079 -35180 13113 -35083
rect 12923 -35238 13113 -35180
rect 11532 -35450 11743 -35447
rect 11492 -35462 11743 -35450
rect 10844 -35556 10850 -35490
rect 10916 -35556 11469 -35490
rect 10844 -35650 10888 -35584
rect 10954 -35650 11299 -35584
rect 10844 -35744 10859 -35678
rect 10925 -35744 11112 -35678
rect 11151 -35735 11299 -35650
rect 11046 -35772 11112 -35744
rect 11233 -35771 11299 -35735
rect 11336 -35771 11370 -35770
rect 10706 -35788 10990 -35772
rect 10706 -35822 10940 -35788
rect 10974 -35822 10990 -35788
rect 10706 -35838 10990 -35822
rect 11046 -35788 11183 -35772
rect 11046 -35822 11132 -35788
rect 11166 -35822 11183 -35788
rect 11046 -35838 11183 -35822
rect 11233 -35788 11374 -35771
rect 11233 -35822 11324 -35788
rect 11358 -35822 11374 -35788
rect 11233 -35837 11374 -35822
rect 11403 -35772 11469 -35556
rect 11403 -35788 11567 -35772
rect 11403 -35822 11516 -35788
rect 11550 -35822 11567 -35788
rect 11403 -35838 11567 -35822
rect 10706 -35868 10816 -35838
rect 7138 -35876 8001 -35869
rect 7138 -35988 7245 -35876
rect 7280 -35988 7438 -35876
rect 7473 -35988 7630 -35876
rect 7665 -35988 7822 -35876
rect 7857 -35988 8001 -35876
rect 7138 -36003 8001 -35988
rect 8086 -35876 8949 -35869
rect 8086 -35988 8193 -35876
rect 8228 -35988 8386 -35876
rect 8421 -35988 8578 -35876
rect 8613 -35988 8770 -35876
rect 8805 -35988 8949 -35876
rect 8086 -36003 8949 -35988
rect 9022 -35876 9885 -35869
rect 9022 -35988 9129 -35876
rect 9164 -35988 9322 -35876
rect 9357 -35988 9514 -35876
rect 9549 -35988 9706 -35876
rect 9741 -35988 9885 -35876
rect 9022 -36003 9885 -35988
rect 9953 -35875 10816 -35868
rect 11633 -35869 11743 -35462
rect 13151 -35615 13235 -34815
rect 12913 -35634 13426 -35615
rect 12913 -35668 12930 -35634
rect 12964 -35668 13184 -35634
rect 13410 -35668 13426 -35634
rect 12913 -35684 13426 -35668
rect 9953 -35987 10060 -35875
rect 10095 -35987 10253 -35875
rect 10288 -35987 10445 -35875
rect 10480 -35987 10637 -35875
rect 10672 -35987 10816 -35875
rect 9953 -36002 10816 -35987
rect 10880 -35876 11743 -35869
rect 10880 -35988 10987 -35876
rect 11022 -35988 11180 -35876
rect 11215 -35988 11372 -35876
rect 11407 -35988 11564 -35876
rect 11599 -35988 11743 -35876
rect 12777 -35727 12927 -35715
rect 12777 -35746 12886 -35727
rect 12777 -35878 12784 -35746
rect 12818 -35878 12886 -35746
rect 12777 -35903 12886 -35878
rect 12920 -35903 12927 -35727
rect 12777 -35915 12927 -35903
rect 12968 -35727 13170 -35715
rect 12968 -35903 12974 -35727
rect 13008 -35838 13170 -35727
rect 13216 -35721 13574 -35715
rect 13216 -35800 13232 -35721
rect 13266 -35800 13424 -35721
rect 13458 -35778 13574 -35721
rect 13458 -35800 13496 -35778
rect 13216 -35806 13496 -35800
rect 13008 -35844 13426 -35838
rect 13008 -35903 13136 -35844
rect 12968 -35915 13136 -35903
rect 12777 -35955 12874 -35915
rect 12974 -35921 13136 -35915
rect 13170 -35921 13328 -35844
rect 13362 -35921 13426 -35844
rect 12974 -35943 13426 -35921
rect 10880 -36003 11743 -35988
rect 7137 -36065 10779 -36056
rect 11883 -36057 12147 -36046
rect 12543 -36052 12549 -35955
rect 12646 -36052 12874 -35955
rect 7137 -36066 9965 -36065
rect 7137 -36176 7150 -36066
rect 7184 -36176 7342 -36066
rect 7376 -36176 7534 -36066
rect 7568 -36176 7726 -36066
rect 7760 -36176 7918 -36066
rect 7952 -36176 8098 -36066
rect 8132 -36176 8290 -36066
rect 8324 -36176 8482 -36066
rect 8516 -36176 8674 -36066
rect 8708 -36176 8866 -36066
rect 8900 -36176 9034 -36066
rect 9068 -36176 9226 -36066
rect 9260 -36176 9418 -36066
rect 9452 -36176 9610 -36066
rect 9644 -36176 9802 -36066
rect 9836 -36175 9965 -36066
rect 9999 -36175 10157 -36065
rect 10191 -36175 10349 -36065
rect 10383 -36175 10541 -36065
rect 10575 -36175 10733 -36065
rect 10767 -36175 10779 -36065
rect 9836 -36176 10779 -36175
rect 7137 -36247 10779 -36176
rect 10880 -36066 11894 -36057
rect 10880 -36176 10892 -36066
rect 10926 -36176 11084 -36066
rect 11118 -36176 11276 -36066
rect 11310 -36176 11468 -36066
rect 11502 -36176 11660 -36066
rect 11694 -36176 11894 -36066
rect 10880 -36187 11894 -36176
rect 7137 -36248 10204 -36247
rect 7137 -36283 7389 -36248
rect 7677 -36283 8337 -36248
rect 8625 -36283 9273 -36248
rect 9561 -36282 10204 -36248
rect 10492 -36282 10779 -36247
rect 9561 -36283 10779 -36282
rect 7137 -36297 10779 -36283
rect 7137 -36299 7964 -36297
rect 8085 -36299 8912 -36297
rect 9021 -36299 9848 -36297
rect 9952 -36298 10779 -36297
rect 10879 -36248 11894 -36187
rect 10879 -36283 11131 -36248
rect 11419 -36283 11894 -36248
rect 10879 -36299 11894 -36283
rect 12136 -36299 12147 -36057
rect 12777 -36094 12874 -36052
rect 12913 -36013 13426 -35943
rect 12913 -36047 12930 -36013
rect 12964 -36047 13184 -36013
rect 13410 -36047 13426 -36013
rect 12913 -36063 13426 -36047
rect 13454 -35869 13496 -35806
rect 13530 -35869 13574 -35778
rect 13454 -35925 13574 -35869
rect 13454 -35959 13690 -35925
rect 13454 -36063 13558 -35959
rect 13662 -36063 13690 -35959
rect 13454 -36094 13690 -36063
rect 12777 -36106 12927 -36094
rect 12777 -36125 12886 -36106
rect 12777 -36257 12784 -36125
rect 12818 -36257 12886 -36125
rect 12777 -36282 12886 -36257
rect 12920 -36282 12927 -36106
rect 12777 -36294 12927 -36282
rect 12968 -36106 13170 -36094
rect 12968 -36282 12974 -36106
rect 13008 -36217 13170 -36106
rect 13216 -36095 13690 -36094
rect 13216 -36100 13574 -36095
rect 13216 -36179 13232 -36100
rect 13266 -36179 13424 -36100
rect 13458 -36157 13574 -36100
rect 13458 -36179 13496 -36157
rect 13216 -36185 13496 -36179
rect 13008 -36223 13426 -36217
rect 13008 -36282 13136 -36223
rect 12968 -36294 13136 -36282
rect 11883 -36310 12147 -36299
rect 12974 -36300 13136 -36294
rect 13170 -36300 13328 -36223
rect 13362 -36300 13426 -36223
rect 12974 -36322 13426 -36300
rect 13454 -36248 13496 -36185
rect 13530 -36248 13574 -36157
rect 13454 -36308 13574 -36248
rect 12913 -36406 13426 -36322
<< via1 >>
rect -21816 6725 -21727 6814
rect -27525 4452 -27436 4541
rect -24000 4445 -22878 4517
rect -22632 4418 -22560 4490
rect -25114 3839 -25005 3948
rect -22416 4366 -22230 4552
rect -15130 6556 -15022 6664
rect -19312 6376 -19240 6448
rect -18528 6279 -18439 6368
rect -24791 3409 -24197 3549
rect -20709 4445 -19587 4517
rect -21823 3876 -21714 3987
rect -16019 6124 -15947 6196
rect -15230 5884 -15141 5973
rect -19130 4372 -18949 4553
rect -21500 3409 -20906 3549
rect -17418 4445 -16296 4517
rect -18532 3887 -18423 3998
rect -12742 5681 -12670 5753
rect -11940 5537 -11851 5626
rect -15826 4378 -15648 4556
rect -18209 3409 -17615 3549
rect -14127 4445 -13005 4517
rect -15241 3891 -15132 4002
rect -12549 4387 -12374 4562
rect -9439 5385 -9367 5457
rect -8640 5227 -8551 5316
rect -6166 5269 -6096 5339
rect -14918 3409 -14324 3549
rect -10836 4445 -9714 4517
rect -11950 3880 -11841 3991
rect 1841 6169 2963 6241
rect 1565 5813 1674 5925
rect 3447 6169 4569 6241
rect 5151 6167 6273 6239
rect 4873 5815 4970 5924
rect 3195 5390 3247 5442
rect 4738 5472 4807 5541
rect -5351 4991 -5262 5080
rect -9267 4252 -9092 4429
rect -11627 3409 -11033 3549
rect -7546 4445 -6424 4517
rect -8660 3900 -8551 4009
rect -5978 4395 -5803 4570
rect 2301 4838 2361 4849
rect -2875 4746 -2803 4818
rect 2301 4792 2361 4838
rect 2301 4789 2361 4792
rect 3907 4838 3967 4849
rect 3907 4792 3967 4838
rect 3907 4789 3967 4792
rect 425 4612 497 4684
rect 4959 5087 5028 5230
rect 5611 4836 5671 4847
rect 5611 4790 5671 4836
rect 5611 4787 5671 4790
rect 7323 4787 7433 4802
rect 7323 4693 7433 4787
rect 7810 4785 7840 4802
rect 7840 4785 7919 4802
rect 7810 4693 7919 4785
rect -8337 3409 -7743 3549
rect -4255 4445 -3133 4517
rect -5369 3900 -5260 4009
rect -2683 4383 -2508 4558
rect -2058 4473 -1969 4562
rect -5046 3409 -4452 3549
rect -964 4445 158 4517
rect -2078 3883 -1969 3994
rect 602 4377 774 4549
rect 602 4060 774 4232
rect 2921 4209 2987 4275
rect 4885 4209 4951 4275
rect -1755 3409 -1161 3549
rect 5339 4011 5411 4083
rect 5558 3863 5627 3879
rect 5558 3810 5577 3863
rect 5577 3810 5611 3863
rect 5611 3810 5627 3863
rect -23398 3114 -23338 3125
rect -23398 3068 -23338 3114
rect -23398 3065 -23338 3068
rect -20107 3114 -20047 3125
rect -20107 3068 -20047 3114
rect -20107 3065 -20047 3068
rect -16816 3114 -16756 3125
rect -16816 3068 -16756 3114
rect -16816 3065 -16756 3068
rect -13525 3114 -13465 3125
rect -13525 3068 -13465 3114
rect -13525 3065 -13465 3068
rect -10234 3114 -10174 3125
rect -10234 3068 -10174 3114
rect -10234 3065 -10174 3068
rect -6944 3114 -6884 3125
rect -6944 3068 -6884 3114
rect -6944 3065 -6884 3068
rect -3653 3114 -3593 3125
rect -3653 3068 -3593 3114
rect -3653 3065 -3593 3068
rect -362 3114 -302 3125
rect -362 3068 -302 3114
rect -362 3065 -302 3068
rect -24670 2661 -23548 2733
rect -23111 2661 -21989 2733
rect -21379 2661 -20257 2733
rect -19820 2661 -18698 2733
rect -18088 2661 -16966 2733
rect -16529 2661 -15407 2733
rect -14797 2661 -13675 2733
rect -13238 2661 -12116 2733
rect -11506 2661 -10384 2733
rect -9947 2661 -8825 2733
rect -8216 2661 -7094 2733
rect -6657 2661 -5535 2733
rect -4925 2661 -3803 2733
rect -3366 2661 -2244 2733
rect -1634 2661 -512 2733
rect -75 2661 1047 2733
rect -24915 1830 -24874 1938
rect -24874 1830 -24825 1938
rect -24818 1597 -24742 1705
rect -23439 1790 -23364 1886
rect -23364 1790 -23291 1886
rect -23291 1790 -23289 1886
rect -23439 1789 -23289 1790
rect -21624 1830 -21583 1938
rect -21583 1830 -21534 1938
rect -23263 1601 -23147 1698
rect -24210 1330 -24150 1341
rect -24210 1284 -24150 1330
rect -24210 1281 -24150 1284
rect -22651 1330 -22591 1341
rect -22651 1284 -22591 1330
rect -21527 1597 -21451 1705
rect -20148 1790 -20073 1886
rect -20073 1790 -20000 1886
rect -20000 1790 -19998 1886
rect -20148 1789 -19998 1790
rect -18333 1830 -18292 1938
rect -18292 1830 -18243 1938
rect -19972 1601 -19856 1698
rect -21814 1321 -21723 1407
rect -20919 1330 -20859 1341
rect -22651 1281 -22591 1284
rect -20919 1284 -20859 1330
rect -20919 1281 -20859 1284
rect -19360 1330 -19300 1341
rect -19360 1284 -19300 1330
rect -18236 1597 -18160 1705
rect -16857 1790 -16782 1886
rect -16782 1790 -16709 1886
rect -16709 1790 -16707 1886
rect -16857 1789 -16707 1790
rect -15042 1830 -15001 1938
rect -15001 1830 -14952 1938
rect -16681 1601 -16565 1698
rect -18523 1321 -18432 1407
rect -17628 1330 -17568 1341
rect -19360 1281 -19300 1284
rect -17628 1284 -17568 1330
rect -17628 1281 -17568 1284
rect -16069 1330 -16009 1341
rect -16069 1284 -16009 1330
rect -14945 1597 -14869 1705
rect -13566 1790 -13491 1886
rect -13491 1790 -13418 1886
rect -13418 1790 -13416 1886
rect -13566 1789 -13416 1790
rect -11751 1830 -11710 1938
rect -11710 1830 -11661 1938
rect -13390 1601 -13274 1698
rect -15232 1321 -15141 1407
rect -14337 1330 -14277 1341
rect -16069 1281 -16009 1284
rect -14337 1284 -14277 1330
rect -14337 1281 -14277 1284
rect -12778 1330 -12718 1341
rect -12778 1284 -12718 1330
rect -11654 1597 -11578 1705
rect -10275 1790 -10200 1886
rect -10200 1790 -10127 1886
rect -10127 1790 -10125 1886
rect -10275 1789 -10125 1790
rect -8461 1830 -8420 1938
rect -8420 1830 -8371 1938
rect -10099 1601 -9983 1698
rect -11941 1321 -11850 1407
rect -11046 1330 -10986 1341
rect -12778 1281 -12718 1284
rect -11046 1284 -10986 1330
rect -11046 1281 -10986 1284
rect -9487 1330 -9427 1341
rect -9487 1284 -9427 1330
rect -8364 1597 -8288 1705
rect -6985 1790 -6910 1886
rect -6910 1790 -6837 1886
rect -6837 1790 -6835 1886
rect -6985 1789 -6835 1790
rect -5170 1830 -5129 1938
rect -5129 1830 -5080 1938
rect -6809 1601 -6693 1698
rect -8650 1321 -8559 1407
rect -7756 1330 -7696 1341
rect -9487 1281 -9427 1284
rect -7756 1284 -7696 1330
rect -7756 1281 -7696 1284
rect -6197 1330 -6137 1341
rect -6197 1284 -6137 1330
rect -5073 1597 -4997 1705
rect -3694 1790 -3619 1886
rect -3619 1790 -3546 1886
rect -3546 1790 -3544 1886
rect -3694 1789 -3544 1790
rect -1879 1830 -1838 1938
rect -1838 1830 -1789 1938
rect -3518 1601 -3402 1698
rect -5360 1321 -5269 1407
rect -4465 1330 -4405 1341
rect -6197 1281 -6137 1284
rect -4465 1284 -4405 1330
rect -4465 1281 -4405 1284
rect -2906 1330 -2846 1341
rect -2906 1284 -2846 1330
rect -1782 1597 -1706 1705
rect -403 1790 -328 1886
rect -328 1790 -255 1886
rect -255 1790 -253 1886
rect -403 1789 -253 1790
rect -227 1601 -111 1698
rect -2069 1321 -1978 1407
rect -1174 1330 -1114 1341
rect -2906 1281 -2846 1284
rect -1174 1284 -1114 1330
rect -1174 1281 -1114 1284
rect 385 1330 445 1341
rect 385 1284 445 1330
rect 1222 1321 1313 1407
rect 385 1281 445 1284
rect 5901 3245 5970 3314
rect 5734 3176 5786 3228
rect 5998 3863 6067 3879
rect 5998 3810 6017 3863
rect 6017 3810 6051 3863
rect 6051 3810 6067 3863
rect -23802 1123 -23703 1192
rect -23290 1130 -23219 1196
rect -20511 1123 -20412 1192
rect -19999 1130 -19928 1196
rect -17220 1123 -17121 1192
rect -16708 1130 -16637 1196
rect -13929 1123 -13830 1192
rect -13417 1130 -13346 1196
rect -10638 1123 -10539 1192
rect -10126 1130 -10055 1196
rect -7348 1123 -7249 1192
rect -6836 1130 -6765 1196
rect -4057 1123 -3958 1192
rect -3545 1130 -3474 1196
rect -766 1123 -667 1192
rect -254 1130 -183 1196
rect 1934 2453 2000 2519
rect -24412 988 -24156 1001
rect -24412 941 -24156 988
rect -24412 929 -24156 941
rect -23123 988 -22867 1001
rect -23123 941 -22891 988
rect -22891 941 -22867 988
rect -23123 929 -22867 941
rect -22406 988 -22150 1001
rect -22406 941 -22150 988
rect -22406 929 -22150 941
rect -21121 988 -20865 1001
rect -21121 941 -20865 988
rect -21121 929 -20865 941
rect -19832 988 -19576 1001
rect -19832 941 -19600 988
rect -19600 941 -19576 988
rect -19832 929 -19576 941
rect -19115 988 -18859 1001
rect -19115 941 -18859 988
rect -19115 929 -18859 941
rect -17830 988 -17574 1001
rect -17830 941 -17574 988
rect -17830 929 -17574 941
rect -16541 988 -16285 1001
rect -16541 941 -16309 988
rect -16309 941 -16285 988
rect -16541 929 -16285 941
rect -15824 988 -15568 1001
rect -15824 941 -15568 988
rect -15824 929 -15568 941
rect -14539 988 -14283 1001
rect -14539 941 -14283 988
rect -14539 929 -14283 941
rect -13250 988 -12994 1001
rect -13250 941 -13018 988
rect -13018 941 -12994 988
rect -13250 929 -12994 941
rect -12533 988 -12277 1001
rect -12533 941 -12277 988
rect -12533 929 -12277 941
rect -11248 988 -10992 1001
rect -11248 941 -10992 988
rect -11248 929 -10992 941
rect -9959 988 -9703 1001
rect -9959 941 -9727 988
rect -9727 941 -9703 988
rect -9959 929 -9703 941
rect -9242 988 -8986 1001
rect -9242 941 -8986 988
rect -9242 929 -8986 941
rect -7958 988 -7702 1001
rect -7958 941 -7702 988
rect -7958 929 -7702 941
rect -6669 988 -6413 1001
rect -6669 941 -6437 988
rect -6437 941 -6413 988
rect -6669 929 -6413 941
rect -5952 988 -5696 1001
rect -5952 941 -5696 988
rect -5952 929 -5696 941
rect -4667 988 -4411 1001
rect -4667 941 -4411 988
rect -4667 929 -4411 941
rect -3378 988 -3122 1001
rect -3378 941 -3146 988
rect -3146 941 -3122 988
rect -3378 929 -3122 941
rect -2661 988 -2405 1001
rect -2661 941 -2405 988
rect -2661 929 -2405 941
rect -1376 988 -1120 1001
rect -1376 941 -1120 988
rect -1376 929 -1120 941
rect -87 988 169 1001
rect -87 941 145 988
rect 145 941 169 988
rect -87 929 169 941
rect 630 988 886 1001
rect 630 941 886 988
rect 630 929 886 941
rect -24601 579 -24519 605
rect -24519 579 -24503 605
rect -24601 525 -24503 579
rect -24046 519 -23963 666
rect -24046 518 -23975 519
rect -23975 518 -23963 519
rect -23490 579 -23410 604
rect -23410 579 -23392 604
rect -23490 524 -23392 579
rect -24810 346 -24557 412
rect -22069 536 -21949 616
rect -23500 341 -23315 401
rect -21310 579 -21228 605
rect -21228 579 -21212 605
rect -21310 525 -21212 579
rect -22628 375 -22483 450
rect -24336 221 -24001 255
rect -24336 203 -24001 221
rect -20755 519 -20672 666
rect -20755 518 -20684 519
rect -20684 518 -20672 519
rect -20199 579 -20119 604
rect -20119 579 -20101 604
rect -20199 524 -20101 579
rect -21519 346 -21266 412
rect -23100 221 -23038 250
rect -23100 188 -23038 221
rect -18778 536 -18658 616
rect -20209 341 -20024 401
rect -18019 579 -17937 605
rect -17937 579 -17921 605
rect -18019 525 -17921 579
rect -19337 375 -19192 450
rect -22233 221 -22181 223
rect -22233 171 -22181 221
rect -21801 218 -21735 284
rect -25060 -214 -24969 -123
rect -21045 221 -20710 255
rect -21045 203 -20710 221
rect -17464 519 -17381 666
rect -17464 518 -17393 519
rect -17393 518 -17381 519
rect -16908 579 -16828 604
rect -16828 579 -16810 604
rect -16908 524 -16810 579
rect -18228 346 -17975 412
rect -19809 221 -19747 250
rect -19809 188 -19747 221
rect -15487 536 -15367 616
rect -16918 341 -16733 401
rect -14728 579 -14646 605
rect -14646 579 -14630 605
rect -14728 525 -14630 579
rect -16046 375 -15901 450
rect -18942 221 -18890 223
rect -18942 171 -18890 221
rect -18505 217 -18439 283
rect -17754 221 -17419 255
rect -17754 203 -17419 221
rect -14173 519 -14090 666
rect -14173 518 -14102 519
rect -14102 518 -14090 519
rect -13617 579 -13537 604
rect -13537 579 -13519 604
rect -13617 524 -13519 579
rect -14937 346 -14684 412
rect -16518 221 -16456 250
rect -16518 188 -16456 221
rect -12196 536 -12076 616
rect -13627 341 -13442 401
rect -11437 579 -11355 605
rect -11355 579 -11339 605
rect -11437 525 -11339 579
rect -12755 375 -12610 450
rect -15651 221 -15599 223
rect -15651 171 -15599 221
rect -15223 230 -15157 296
rect -14463 221 -14128 255
rect -14463 203 -14128 221
rect -10882 519 -10799 666
rect -10882 518 -10811 519
rect -10811 518 -10799 519
rect -10326 579 -10246 604
rect -10246 579 -10228 604
rect -10326 524 -10228 579
rect -11646 346 -11393 412
rect -13227 221 -13165 250
rect -13227 188 -13165 221
rect -8905 536 -8785 616
rect -10336 341 -10151 401
rect -8147 579 -8065 605
rect -8065 579 -8049 605
rect -8147 525 -8049 579
rect -9464 375 -9319 450
rect -12360 221 -12308 223
rect -11963 223 -11897 289
rect -12360 171 -12308 221
rect -11172 221 -10837 255
rect -11172 203 -10837 221
rect -7592 519 -7509 666
rect -7592 518 -7521 519
rect -7521 518 -7509 519
rect -7036 579 -6956 604
rect -6956 579 -6938 604
rect -7036 524 -6938 579
rect -8356 346 -8103 412
rect -9936 221 -9874 250
rect -9936 188 -9874 221
rect -5615 536 -5495 616
rect -7046 341 -6861 401
rect -4856 579 -4774 605
rect -4774 579 -4758 605
rect -4856 525 -4758 579
rect -6174 375 -6029 450
rect -9069 221 -9017 223
rect -9069 171 -9017 221
rect -8633 243 -8567 309
rect -7882 221 -7547 255
rect -7882 203 -7547 221
rect -4301 519 -4218 666
rect -4301 518 -4230 519
rect -4230 518 -4218 519
rect -3745 579 -3665 604
rect -3665 579 -3647 604
rect -3745 524 -3647 579
rect -5065 346 -4812 412
rect -6646 221 -6584 250
rect -6646 188 -6584 221
rect -2324 536 -2204 616
rect -3755 341 -3570 401
rect -1565 579 -1483 605
rect -1483 579 -1467 605
rect -1565 525 -1467 579
rect -2883 375 -2738 450
rect -5779 221 -5727 223
rect -5779 171 -5727 221
rect -5349 226 -5283 292
rect -4591 221 -4256 255
rect -4591 203 -4256 221
rect -1010 519 -927 666
rect -1010 518 -939 519
rect -939 518 -927 519
rect -454 579 -374 604
rect -374 579 -356 604
rect -454 524 -356 579
rect -1774 346 -1521 412
rect -3355 221 -3293 250
rect -3355 188 -3293 221
rect 967 536 1087 616
rect -464 341 -279 401
rect 408 375 553 450
rect -2488 221 -2436 223
rect -2488 171 -2436 221
rect -2061 195 -1995 261
rect -1300 221 -965 255
rect -1300 203 -965 221
rect -64 221 -2 250
rect -64 188 -2 221
rect 803 221 855 223
rect 803 171 855 221
rect 6172 3237 6224 3247
rect 6172 3195 6224 3237
rect 6341 3243 6410 3312
rect 6438 3863 6507 3879
rect 6438 3810 6457 3863
rect 6457 3810 6491 3863
rect 6491 3810 6507 3863
rect 5998 2706 6067 2775
rect 6612 3237 6664 3256
rect 6612 3204 6664 3237
rect 6438 2571 6507 2640
rect 7106 2809 7158 2861
rect 7113 2715 7165 2767
rect 7327 2612 7393 2678
rect 8069 2808 8122 2860
rect 8057 2716 8109 2768
rect 8424 2633 8493 2685
rect 7106 2251 7172 2317
rect 6966 2147 7032 2213
rect 7227 1702 7372 1715
rect 7372 1702 7405 1715
rect 7227 1550 7405 1702
rect 9002 2809 9055 2861
rect 9000 2711 9052 2763
rect 8989 2619 9042 2672
rect 8050 2147 8116 2213
rect 7872 1994 7938 2060
rect 8162 1702 8320 1715
rect 8320 1702 8340 1715
rect 7227 1537 7372 1550
rect 7372 1537 7405 1550
rect 6953 1045 7019 1111
rect 7102 825 7168 891
rect 7853 1201 7919 1267
rect 8162 1550 8340 1702
rect 8986 2453 9052 2519
rect 9933 2809 9986 2861
rect 9935 2711 9987 2763
rect 10262 2647 10331 2716
rect 9798 2496 9864 2562
rect 8818 2248 8884 2314
rect 9098 1702 9256 1715
rect 9256 1702 9276 1715
rect 8162 1537 8320 1550
rect 8320 1537 8340 1550
rect 6780 580 6849 649
rect 6066 480 6132 546
rect 6941 386 7007 452
rect 8050 704 8116 770
rect 9098 1550 9276 1702
rect 10860 2706 10926 2772
rect 10858 2612 10924 2678
rect 10850 2518 10915 2584
rect 9917 2357 9983 2423
rect 10029 1702 10187 1715
rect 10187 1702 10206 1715
rect 9098 1537 9256 1550
rect 9256 1537 9276 1550
rect 8837 791 8903 857
rect 8989 1045 9055 1111
rect 8401 569 8465 633
rect 8079 485 8131 537
rect 8063 391 8128 443
rect 10029 1551 10206 1702
rect 10956 1702 11114 1715
rect 11114 1702 11134 1715
rect 10029 1538 10187 1551
rect 10187 1538 10206 1551
rect 9917 923 9983 989
rect 8993 574 9059 640
rect 9001 480 9067 546
rect 8992 391 9057 443
rect 9807 699 9873 763
rect 10956 1550 11134 1702
rect 12189 2658 12410 2861
rect 10956 1537 11114 1550
rect 11114 1537 11134 1550
rect 10264 573 10324 633
rect 9937 481 10003 547
rect 9951 437 10016 443
rect 9951 403 10013 437
rect 10013 403 10016 437
rect 9951 391 10016 403
rect 12233 1188 12352 1204
rect 12233 1085 12352 1188
rect 12960 1044 13079 1163
rect 10850 668 10916 734
rect 10888 574 10954 640
rect 10859 480 10925 546
rect 248 -131 339 -40
rect 11894 -75 12136 167
rect 1625 -1375 1691 -1309
rect 3886 -1635 3970 -1551
rect -24410 -2347 -23856 -2327
rect -24410 -2419 -23856 -2347
rect -23605 -2247 -23436 -2225
rect -23605 -2281 -23565 -2247
rect -23565 -2281 -23474 -2247
rect -23474 -2281 -23436 -2247
rect -23605 -2304 -23436 -2281
rect -24410 -2467 -24401 -2419
rect -24401 -2467 -24243 -2419
rect -24243 -2467 -24209 -2419
rect -24209 -2467 -24051 -2419
rect -24051 -2467 -24017 -2419
rect -24017 -2467 -23859 -2419
rect -23859 -2467 -23856 -2419
rect -22373 -2347 -21819 -2327
rect -22373 -2419 -21819 -2347
rect -21585 -2247 -21416 -2225
rect -21585 -2281 -21545 -2247
rect -21545 -2281 -21454 -2247
rect -21454 -2281 -21416 -2247
rect -21585 -2304 -21416 -2281
rect -22373 -2467 -22364 -2419
rect -22364 -2467 -22206 -2419
rect -22206 -2467 -22172 -2419
rect -22172 -2467 -22014 -2419
rect -22014 -2467 -21980 -2419
rect -21980 -2467 -21822 -2419
rect -21822 -2467 -21819 -2419
rect -24635 -2791 -24492 -2648
rect -20643 -2347 -20089 -2327
rect -20643 -2419 -20089 -2347
rect -19844 -2247 -19675 -2225
rect -19844 -2281 -19804 -2247
rect -19804 -2281 -19713 -2247
rect -19713 -2281 -19675 -2247
rect -19844 -2304 -19675 -2281
rect -20643 -2467 -20634 -2419
rect -20634 -2467 -20476 -2419
rect -20476 -2467 -20442 -2419
rect -20442 -2467 -20284 -2419
rect -20284 -2467 -20250 -2419
rect -20250 -2467 -20092 -2419
rect -20092 -2467 -20089 -2419
rect -23601 -2891 -23452 -2878
rect -24550 -3165 -24428 -2987
rect -24184 -2995 -23844 -2983
rect -24184 -3033 -23844 -2995
rect -24184 -3057 -23851 -3033
rect -23851 -3057 -23844 -3033
rect -23601 -2959 -23452 -2891
rect -23601 -2974 -23597 -2959
rect -23597 -2974 -23465 -2959
rect -23465 -2974 -23452 -2959
rect -23253 -2866 -23121 -2747
rect -22731 -2767 -22413 -2674
rect -18883 -2347 -18329 -2327
rect -18883 -2419 -18329 -2347
rect -18065 -2247 -17896 -2225
rect -18065 -2281 -18025 -2247
rect -18025 -2281 -17934 -2247
rect -17934 -2281 -17896 -2247
rect -18065 -2304 -17896 -2281
rect -18883 -2467 -18874 -2419
rect -18874 -2467 -18716 -2419
rect -18716 -2467 -18682 -2419
rect -18682 -2467 -18524 -2419
rect -18524 -2467 -18490 -2419
rect -18490 -2467 -18332 -2419
rect -18332 -2467 -18329 -2419
rect -20889 -2772 -20682 -2675
rect -22594 -3080 -22431 -2852
rect -21581 -2891 -21432 -2878
rect -21293 -2859 -21209 -2775
rect -19043 -2780 -18894 -2673
rect -22147 -2995 -21807 -2983
rect -22147 -3033 -21807 -2995
rect -22147 -3057 -21814 -3033
rect -21814 -3057 -21807 -3033
rect -21581 -2959 -21432 -2891
rect -21581 -2974 -21577 -2959
rect -21577 -2974 -21445 -2959
rect -21445 -2974 -21432 -2959
rect -19840 -2891 -19691 -2878
rect -19555 -2864 -19471 -2780
rect -20417 -2995 -20077 -2983
rect -20417 -3033 -20077 -2995
rect -20917 -3165 -20741 -3042
rect -20417 -3057 -20084 -3033
rect -20084 -3057 -20077 -3033
rect -19840 -2959 -19691 -2891
rect -19840 -2974 -19836 -2959
rect -19836 -2974 -19704 -2959
rect -19704 -2974 -19691 -2959
rect -19241 -3087 -19043 -2934
rect -18061 -2891 -17912 -2878
rect -17693 -2852 -17579 -2696
rect -18657 -2995 -18317 -2983
rect -18657 -3033 -18317 -2995
rect -18657 -3057 -18324 -3033
rect -18324 -3057 -18317 -3033
rect -18061 -2959 -17912 -2891
rect -18061 -2974 -18057 -2959
rect -18057 -2974 -17925 -2959
rect -17925 -2974 -17912 -2959
rect -24807 -4337 -24618 -4064
rect -24359 -4159 -23805 -4139
rect -24359 -4231 -23805 -4159
rect -23561 -4059 -23392 -4037
rect -23561 -4093 -23521 -4059
rect -23521 -4093 -23430 -4059
rect -23430 -4093 -23392 -4059
rect -23561 -4116 -23392 -4093
rect -24359 -4279 -24350 -4231
rect -24350 -4279 -24192 -4231
rect -24192 -4279 -24158 -4231
rect -24158 -4279 -24000 -4231
rect -24000 -4279 -23966 -4231
rect -23966 -4279 -23808 -4231
rect -23808 -4279 -23805 -4231
rect -23557 -4703 -23408 -4690
rect -24133 -4807 -23793 -4795
rect -24133 -4845 -23793 -4807
rect -24133 -4869 -23800 -4845
rect -23800 -4869 -23793 -4845
rect -23557 -4771 -23408 -4703
rect -23557 -4786 -23553 -4771
rect -23553 -4786 -23421 -4771
rect -23421 -4786 -23408 -4771
rect -24615 -5133 -24479 -4997
rect -24359 -5451 -23805 -5431
rect -24359 -5523 -23805 -5451
rect -23563 -5351 -23394 -5329
rect -23563 -5385 -23523 -5351
rect -23523 -5385 -23432 -5351
rect -23432 -5385 -23394 -5351
rect -23563 -5408 -23394 -5385
rect -24359 -5571 -24350 -5523
rect -24350 -5571 -24192 -5523
rect -24192 -5571 -24158 -5523
rect -24158 -5571 -24000 -5523
rect -24000 -5571 -23966 -5523
rect -23966 -5571 -23808 -5523
rect -23808 -5571 -23805 -5523
rect -22623 -4159 -22069 -4139
rect -22623 -4231 -22069 -4159
rect -21823 -4059 -21654 -4037
rect -21823 -4093 -21783 -4059
rect -21783 -4093 -21692 -4059
rect -21692 -4093 -21654 -4059
rect -21823 -4116 -21654 -4093
rect -22623 -4279 -22614 -4231
rect -22614 -4279 -22456 -4231
rect -22456 -4279 -22422 -4231
rect -22422 -4279 -22264 -4231
rect -22264 -4279 -22230 -4231
rect -22230 -4279 -22072 -4231
rect -22072 -4279 -22069 -4231
rect -22836 -4594 -22690 -4481
rect -20603 -3899 -19481 -3827
rect -19044 -3899 -17922 -3827
rect -17744 -3858 -17655 -3763
rect -17312 -3899 -16190 -3827
rect -15753 -3899 -14631 -3827
rect -14460 -3946 -14361 -3762
rect -14021 -3899 -12899 -3827
rect -12462 -3899 -11340 -3827
rect -11165 -3905 -11074 -3761
rect -10730 -3899 -9608 -3827
rect -9171 -3899 -8049 -3827
rect -21819 -4703 -21670 -4690
rect -22397 -4807 -22057 -4795
rect -22397 -4845 -22057 -4807
rect -22397 -4869 -22064 -4845
rect -22064 -4869 -22057 -4845
rect -21819 -4771 -21670 -4703
rect -21819 -4786 -21815 -4771
rect -21815 -4786 -21683 -4771
rect -21683 -4786 -21670 -4771
rect -20848 -4730 -20807 -4622
rect -20807 -4730 -20758 -4622
rect -20751 -4963 -20675 -4855
rect -19372 -4770 -19297 -4674
rect -19297 -4770 -19224 -4674
rect -19224 -4770 -19222 -4674
rect -19372 -4771 -19222 -4770
rect -17557 -4730 -17516 -4622
rect -17516 -4730 -17467 -4622
rect -19196 -4959 -19080 -4862
rect -22868 -5133 -22732 -4997
rect -20143 -5230 -20083 -5219
rect -20143 -5276 -20083 -5230
rect -20143 -5279 -20083 -5276
rect -18584 -5230 -18524 -5219
rect -18584 -5276 -18524 -5230
rect -17460 -4963 -17384 -4855
rect -16081 -4770 -16006 -4674
rect -16006 -4770 -15933 -4674
rect -15933 -4770 -15931 -4674
rect -16081 -4771 -15931 -4770
rect -14266 -4730 -14225 -4622
rect -14225 -4730 -14176 -4622
rect -15905 -4959 -15789 -4862
rect -17747 -5239 -17656 -5153
rect -16852 -5230 -16792 -5219
rect -18584 -5279 -18524 -5276
rect -16852 -5276 -16792 -5230
rect -16852 -5279 -16792 -5276
rect -15293 -5230 -15233 -5219
rect -15293 -5276 -15233 -5230
rect -14169 -4963 -14093 -4855
rect -12790 -4770 -12715 -4674
rect -12715 -4770 -12642 -4674
rect -12642 -4770 -12640 -4674
rect -12790 -4771 -12640 -4770
rect -10975 -4730 -10934 -4622
rect -10934 -4730 -10885 -4622
rect -12614 -4959 -12498 -4862
rect -14456 -5239 -14365 -5153
rect -13561 -5230 -13501 -5219
rect -15293 -5279 -15233 -5276
rect -13561 -5276 -13501 -5230
rect -13561 -5279 -13501 -5276
rect -12002 -5230 -11942 -5219
rect -12002 -5276 -11942 -5230
rect -10878 -4963 -10802 -4855
rect -9499 -4770 -9424 -4674
rect -9424 -4770 -9351 -4674
rect -9351 -4770 -9349 -4674
rect -9499 -4771 -9349 -4770
rect -9323 -4959 -9207 -4862
rect -11165 -5239 -11074 -5153
rect -10270 -5230 -10210 -5219
rect -12002 -5279 -11942 -5276
rect -10270 -5276 -10210 -5230
rect -10270 -5279 -10210 -5276
rect -8711 -5230 -8651 -5219
rect -8711 -5276 -8651 -5230
rect -7874 -5239 -7783 -5153
rect -8711 -5279 -8651 -5276
rect -22623 -5451 -22069 -5431
rect -22623 -5523 -22069 -5451
rect -21829 -5351 -21660 -5329
rect -21829 -5385 -21789 -5351
rect -21789 -5385 -21698 -5351
rect -21698 -5385 -21660 -5351
rect -21829 -5408 -21660 -5385
rect -22623 -5571 -22614 -5523
rect -22614 -5571 -22456 -5523
rect -22456 -5571 -22422 -5523
rect -22422 -5571 -22264 -5523
rect -22264 -5571 -22230 -5523
rect -22230 -5571 -22072 -5523
rect -22072 -5571 -22069 -5523
rect -21003 -5435 -20885 -5333
rect -19735 -5437 -19636 -5368
rect -19223 -5430 -19152 -5364
rect -16444 -5437 -16345 -5368
rect -15932 -5430 -15861 -5364
rect -13153 -5437 -13054 -5368
rect -12641 -5430 -12570 -5364
rect -9862 -5437 -9763 -5368
rect -9350 -5430 -9279 -5364
rect -20345 -5572 -20089 -5559
rect -20345 -5619 -20089 -5572
rect -20345 -5631 -20089 -5619
rect -19056 -5572 -18800 -5559
rect -19056 -5619 -18824 -5572
rect -18824 -5619 -18800 -5572
rect -19056 -5631 -18800 -5619
rect -18339 -5572 -18083 -5559
rect -18339 -5619 -18083 -5572
rect -18339 -5631 -18083 -5619
rect -17054 -5572 -16798 -5559
rect -17054 -5619 -16798 -5572
rect -17054 -5631 -16798 -5619
rect -15765 -5572 -15509 -5559
rect -15765 -5619 -15533 -5572
rect -15533 -5619 -15509 -5572
rect -15765 -5631 -15509 -5619
rect -15048 -5572 -14792 -5559
rect -15048 -5619 -14792 -5572
rect -15048 -5631 -14792 -5619
rect -13763 -5572 -13507 -5559
rect -13763 -5619 -13507 -5572
rect -13763 -5631 -13507 -5619
rect -12474 -5572 -12218 -5559
rect -12474 -5619 -12242 -5572
rect -12242 -5619 -12218 -5572
rect -12474 -5631 -12218 -5619
rect -11757 -5572 -11501 -5559
rect -11757 -5619 -11501 -5572
rect -11757 -5631 -11501 -5619
rect -10472 -5572 -10216 -5559
rect -10472 -5619 -10216 -5572
rect -10472 -5631 -10216 -5619
rect -9183 -5572 -8927 -5559
rect -9183 -5619 -8951 -5572
rect -8951 -5619 -8927 -5572
rect -9183 -5631 -8927 -5619
rect -8466 -5572 -8210 -5559
rect -8466 -5619 -8210 -5572
rect -8466 -5631 -8210 -5619
rect -24612 -6247 -24466 -6049
rect -23559 -5995 -23410 -5982
rect -24133 -6099 -23793 -6087
rect -24133 -6137 -23793 -6099
rect -24133 -6161 -23800 -6137
rect -23800 -6161 -23793 -6137
rect -23559 -6063 -23410 -5995
rect -23559 -6078 -23555 -6063
rect -23555 -6078 -23423 -6063
rect -23423 -6078 -23410 -6063
rect -22884 -6046 -22652 -5936
rect -21560 -5922 -21347 -5731
rect -21825 -5995 -21676 -5982
rect -22397 -6099 -22057 -6087
rect -22397 -6137 -22057 -6099
rect -22397 -6161 -22064 -6137
rect -22064 -6161 -22057 -6137
rect -21825 -6063 -21676 -5995
rect -21825 -6078 -21821 -6063
rect -21821 -6078 -21689 -6063
rect -21689 -6078 -21676 -6063
rect -20534 -5981 -20452 -5955
rect -20452 -5981 -20436 -5955
rect -20534 -6035 -20436 -5981
rect -19979 -6041 -19896 -5894
rect -19979 -6042 -19908 -6041
rect -19908 -6042 -19896 -6041
rect -19423 -5981 -19343 -5956
rect -19343 -5981 -19325 -5956
rect -19423 -6036 -19325 -5981
rect -20743 -6214 -20490 -6148
rect -18002 -6024 -17882 -5944
rect -19433 -6219 -19248 -6159
rect -17243 -5981 -17161 -5955
rect -17161 -5981 -17145 -5955
rect -17243 -6035 -17145 -5981
rect -18561 -6185 -18416 -6110
rect -20269 -6339 -19934 -6305
rect -20269 -6357 -19934 -6339
rect -16688 -6041 -16605 -5894
rect -16688 -6042 -16617 -6041
rect -16617 -6042 -16605 -6041
rect -16132 -5981 -16052 -5956
rect -16052 -5981 -16034 -5956
rect -16132 -6036 -16034 -5981
rect -17452 -6214 -17199 -6148
rect -19033 -6339 -18971 -6310
rect -19033 -6372 -18971 -6339
rect -14711 -6024 -14591 -5944
rect -16142 -6219 -15957 -6159
rect -18166 -6339 -18114 -6337
rect -18166 -6389 -18114 -6339
rect -13952 -5981 -13870 -5955
rect -13870 -5981 -13854 -5955
rect -13952 -6035 -13854 -5981
rect -15270 -6185 -15125 -6110
rect -16978 -6339 -16643 -6305
rect -16978 -6357 -16643 -6339
rect -13397 -6041 -13314 -5894
rect -13397 -6042 -13326 -6041
rect -13326 -6042 -13314 -6041
rect -12841 -5981 -12761 -5956
rect -12761 -5981 -12743 -5956
rect -12841 -6036 -12743 -5981
rect -14161 -6214 -13908 -6148
rect -15742 -6339 -15680 -6310
rect -15742 -6372 -15680 -6339
rect -11420 -6024 -11300 -5944
rect -12851 -6219 -12666 -6159
rect -14875 -6339 -14823 -6337
rect -14875 -6389 -14823 -6339
rect -10661 -5981 -10579 -5955
rect -10579 -5981 -10563 -5955
rect -10661 -6035 -10563 -5981
rect -11979 -6185 -11834 -6110
rect -13687 -6339 -13352 -6305
rect -13687 -6357 -13352 -6339
rect -10106 -6041 -10023 -5894
rect -10106 -6042 -10035 -6041
rect -10035 -6042 -10023 -6041
rect -9550 -5981 -9470 -5956
rect -9470 -5981 -9452 -5956
rect -9550 -6036 -9452 -5981
rect -10870 -6214 -10617 -6148
rect -12451 -6339 -12389 -6310
rect -12451 -6372 -12389 -6339
rect -8129 -6024 -8009 -5944
rect -9560 -6219 -9375 -6159
rect -11584 -6339 -11532 -6337
rect -11584 -6389 -11532 -6339
rect -8688 -6185 -8543 -6110
rect -10396 -6339 -10061 -6305
rect -10396 -6357 -10061 -6339
rect -9160 -6339 -9098 -6310
rect -9160 -6372 -9098 -6339
rect -7873 -6291 -7807 -6225
rect -8293 -6339 -8241 -6337
rect -8293 -6389 -8241 -6339
rect -5439 -6599 -5373 -6533
rect -24359 -7424 -23805 -7404
rect -23562 -7324 -23393 -7302
rect -23562 -7358 -23521 -7324
rect -23521 -7358 -23430 -7324
rect -23430 -7358 -23393 -7324
rect -23562 -7381 -23393 -7358
rect -24359 -7496 -23805 -7424
rect -24359 -7544 -24350 -7496
rect -24350 -7544 -24192 -7496
rect -24192 -7544 -24158 -7496
rect -24158 -7544 -24000 -7496
rect -24000 -7544 -23966 -7496
rect -23966 -7544 -23808 -7496
rect -23808 -7544 -23805 -7496
rect -24611 -8015 -24368 -7911
rect -23558 -7968 -23409 -7955
rect -24133 -8072 -23793 -8060
rect -24133 -8110 -23793 -8072
rect -24133 -8134 -23800 -8110
rect -23800 -8134 -23793 -8110
rect -23558 -8036 -23409 -7968
rect -23558 -8051 -23553 -8036
rect -23553 -8051 -23421 -8036
rect -23421 -8051 -23409 -8036
rect -24359 -8716 -23805 -8696
rect -24359 -8788 -23805 -8716
rect -23560 -8616 -23391 -8594
rect -23560 -8650 -23520 -8616
rect -23520 -8650 -23429 -8616
rect -23429 -8650 -23391 -8616
rect -23560 -8673 -23391 -8650
rect -24359 -8836 -24350 -8788
rect -24350 -8836 -24192 -8788
rect -24192 -8836 -24158 -8788
rect -24158 -8836 -24000 -8788
rect -24000 -8836 -23966 -8788
rect -23966 -8836 -23808 -8788
rect -23808 -8836 -23805 -8788
rect -22622 -7424 -22068 -7404
rect -22622 -7496 -22068 -7424
rect -21827 -7324 -21658 -7302
rect -21827 -7358 -21787 -7324
rect -21787 -7358 -21696 -7324
rect -21696 -7358 -21658 -7324
rect -21827 -7381 -21658 -7358
rect -22622 -7544 -22613 -7496
rect -22613 -7544 -22455 -7496
rect -22455 -7544 -22421 -7496
rect -22421 -7544 -22263 -7496
rect -22263 -7544 -22229 -7496
rect -22229 -7544 -22071 -7496
rect -22071 -7544 -22068 -7496
rect -22808 -7856 -22688 -7749
rect -22857 -8015 -22628 -7907
rect -20603 -7164 -19481 -7092
rect -19044 -7164 -17922 -7092
rect -17744 -7123 -17655 -7028
rect -17312 -7164 -16190 -7092
rect -15753 -7164 -14631 -7092
rect -14460 -7211 -14361 -7027
rect -14021 -7164 -12899 -7092
rect -12462 -7164 -11340 -7092
rect -11165 -7170 -11074 -7026
rect -10730 -7164 -9608 -7092
rect -9171 -7164 -8049 -7092
rect -21823 -7968 -21674 -7955
rect -22396 -8072 -22056 -8060
rect -22396 -8110 -22056 -8072
rect -22396 -8134 -22063 -8110
rect -22063 -8134 -22056 -8110
rect -21823 -8036 -21674 -7968
rect -21823 -8051 -21819 -8036
rect -21819 -8051 -21687 -8036
rect -21687 -8051 -21674 -8036
rect -20848 -7995 -20807 -7887
rect -20807 -7995 -20758 -7887
rect -20751 -8228 -20675 -8120
rect -19372 -8035 -19297 -7939
rect -19297 -8035 -19224 -7939
rect -19224 -8035 -19222 -7939
rect -19372 -8036 -19222 -8035
rect -17557 -7995 -17516 -7887
rect -17516 -7995 -17467 -7887
rect -19196 -8224 -19080 -8127
rect -20143 -8495 -20083 -8484
rect -20143 -8541 -20083 -8495
rect -20143 -8544 -20083 -8541
rect -18584 -8495 -18524 -8484
rect -18584 -8541 -18524 -8495
rect -17460 -8228 -17384 -8120
rect -16081 -8035 -16006 -7939
rect -16006 -8035 -15933 -7939
rect -15933 -8035 -15931 -7939
rect -16081 -8036 -15931 -8035
rect -14266 -7995 -14225 -7887
rect -14225 -7995 -14176 -7887
rect -15905 -8224 -15789 -8127
rect -17747 -8504 -17656 -8418
rect -16852 -8495 -16792 -8484
rect -18584 -8544 -18524 -8541
rect -16852 -8541 -16792 -8495
rect -16852 -8544 -16792 -8541
rect -15293 -8495 -15233 -8484
rect -15293 -8541 -15233 -8495
rect -14169 -8228 -14093 -8120
rect -12790 -8035 -12715 -7939
rect -12715 -8035 -12642 -7939
rect -12642 -8035 -12640 -7939
rect -12790 -8036 -12640 -8035
rect -10975 -7995 -10934 -7887
rect -10934 -7995 -10885 -7887
rect -12614 -8224 -12498 -8127
rect -14456 -8504 -14365 -8418
rect -13561 -8495 -13501 -8484
rect -15293 -8544 -15233 -8541
rect -13561 -8541 -13501 -8495
rect -13561 -8544 -13501 -8541
rect -12002 -8495 -11942 -8484
rect -12002 -8541 -11942 -8495
rect -10878 -8228 -10802 -8120
rect -9499 -8035 -9424 -7939
rect -9424 -8035 -9351 -7939
rect -9351 -8035 -9349 -7939
rect -9499 -8036 -9349 -8035
rect -9323 -8224 -9207 -8127
rect -11165 -8504 -11074 -8418
rect -10270 -8495 -10210 -8484
rect -12002 -8544 -11942 -8541
rect -10270 -8541 -10210 -8495
rect -10270 -8544 -10210 -8541
rect -8711 -8495 -8651 -8484
rect -8711 -8541 -8651 -8495
rect -7874 -8504 -7783 -8418
rect -8711 -8544 -8651 -8541
rect -22623 -8716 -22069 -8696
rect -22623 -8788 -22069 -8716
rect -21823 -8616 -21654 -8594
rect -21823 -8650 -21783 -8616
rect -21783 -8650 -21692 -8616
rect -21692 -8650 -21654 -8616
rect -21823 -8673 -21654 -8650
rect -22623 -8836 -22614 -8788
rect -22614 -8836 -22456 -8788
rect -22456 -8836 -22422 -8788
rect -22422 -8836 -22264 -8788
rect -22264 -8836 -22230 -8788
rect -22230 -8836 -22072 -8788
rect -22072 -8836 -22069 -8788
rect -24601 -9146 -24445 -9039
rect -21003 -8700 -20885 -8598
rect -19735 -8702 -19636 -8633
rect -19223 -8695 -19152 -8629
rect -16444 -8702 -16345 -8633
rect -15932 -8695 -15861 -8629
rect -13153 -8702 -13054 -8633
rect -12641 -8695 -12570 -8629
rect -9862 -8702 -9763 -8633
rect -9350 -8695 -9279 -8629
rect -20345 -8837 -20089 -8824
rect -20345 -8884 -20089 -8837
rect -20345 -8896 -20089 -8884
rect -19056 -8837 -18800 -8824
rect -19056 -8884 -18824 -8837
rect -18824 -8884 -18800 -8837
rect -19056 -8896 -18800 -8884
rect -18339 -8837 -18083 -8824
rect -18339 -8884 -18083 -8837
rect -18339 -8896 -18083 -8884
rect -17054 -8837 -16798 -8824
rect -17054 -8884 -16798 -8837
rect -17054 -8896 -16798 -8884
rect -15765 -8837 -15509 -8824
rect -15765 -8884 -15533 -8837
rect -15533 -8884 -15509 -8837
rect -15765 -8896 -15509 -8884
rect -15048 -8837 -14792 -8824
rect -15048 -8884 -14792 -8837
rect -15048 -8896 -14792 -8884
rect -13763 -8837 -13507 -8824
rect -13763 -8884 -13507 -8837
rect -13763 -8896 -13507 -8884
rect -12474 -8837 -12218 -8824
rect -12474 -8884 -12242 -8837
rect -12242 -8884 -12218 -8837
rect -12474 -8896 -12218 -8884
rect -11757 -8837 -11501 -8824
rect -11757 -8884 -11501 -8837
rect -11757 -8896 -11501 -8884
rect -10472 -8837 -10216 -8824
rect -10472 -8884 -10216 -8837
rect -10472 -8896 -10216 -8884
rect -9183 -8837 -8927 -8824
rect -9183 -8884 -8951 -8837
rect -8951 -8884 -8927 -8837
rect -9183 -8896 -8927 -8884
rect -8466 -8837 -8210 -8824
rect -8466 -8884 -8210 -8837
rect -8466 -8896 -8210 -8884
rect -22885 -9148 -22683 -9037
rect -24612 -9512 -24466 -9314
rect -23556 -9260 -23407 -9247
rect -24133 -9364 -23793 -9352
rect -24133 -9402 -23793 -9364
rect -24133 -9426 -23800 -9402
rect -23800 -9426 -23793 -9402
rect -23556 -9328 -23407 -9260
rect -23556 -9343 -23552 -9328
rect -23552 -9343 -23420 -9328
rect -23420 -9343 -23407 -9328
rect -22891 -9303 -22686 -9211
rect -21573 -9193 -21351 -9019
rect -21819 -9260 -21670 -9247
rect -22397 -9364 -22057 -9352
rect -22397 -9402 -22057 -9364
rect -22397 -9426 -22064 -9402
rect -22064 -9426 -22057 -9402
rect -21819 -9328 -21670 -9260
rect -21819 -9343 -21815 -9328
rect -21815 -9343 -21683 -9328
rect -21683 -9343 -21670 -9328
rect -20534 -9246 -20452 -9220
rect -20452 -9246 -20436 -9220
rect -20534 -9300 -20436 -9246
rect -19979 -9306 -19896 -9159
rect -19979 -9307 -19908 -9306
rect -19908 -9307 -19896 -9306
rect -19423 -9246 -19343 -9221
rect -19343 -9246 -19325 -9221
rect -19423 -9301 -19325 -9246
rect -20743 -9479 -20490 -9413
rect -18002 -9289 -17882 -9209
rect -19433 -9484 -19248 -9424
rect -17243 -9246 -17161 -9220
rect -17161 -9246 -17145 -9220
rect -17243 -9300 -17145 -9246
rect -18561 -9450 -18416 -9375
rect -20269 -9604 -19934 -9570
rect -20269 -9622 -19934 -9604
rect -16688 -9306 -16605 -9159
rect -16688 -9307 -16617 -9306
rect -16617 -9307 -16605 -9306
rect -16132 -9246 -16052 -9221
rect -16052 -9246 -16034 -9221
rect -16132 -9301 -16034 -9246
rect -17452 -9479 -17199 -9413
rect -19033 -9604 -18971 -9575
rect -19033 -9637 -18971 -9604
rect -14711 -9289 -14591 -9209
rect -16142 -9484 -15957 -9424
rect -18166 -9604 -18114 -9602
rect -18166 -9654 -18114 -9604
rect -13952 -9246 -13870 -9220
rect -13870 -9246 -13854 -9220
rect -13952 -9300 -13854 -9246
rect -15270 -9450 -15125 -9375
rect -16978 -9604 -16643 -9570
rect -16978 -9622 -16643 -9604
rect -13397 -9306 -13314 -9159
rect -13397 -9307 -13326 -9306
rect -13326 -9307 -13314 -9306
rect -12841 -9246 -12761 -9221
rect -12761 -9246 -12743 -9221
rect -12841 -9301 -12743 -9246
rect -14161 -9479 -13908 -9413
rect -15742 -9604 -15680 -9575
rect -15742 -9637 -15680 -9604
rect -11420 -9289 -11300 -9209
rect -12851 -9484 -12666 -9424
rect -14875 -9604 -14823 -9602
rect -14875 -9654 -14823 -9604
rect -10661 -9246 -10579 -9220
rect -10579 -9246 -10563 -9220
rect -10661 -9300 -10563 -9246
rect -11979 -9450 -11834 -9375
rect -13687 -9604 -13352 -9570
rect -13687 -9622 -13352 -9604
rect -10106 -9306 -10023 -9159
rect -10106 -9307 -10035 -9306
rect -10035 -9307 -10023 -9306
rect -9550 -9246 -9470 -9221
rect -9470 -9246 -9452 -9221
rect -9550 -9301 -9452 -9246
rect -10870 -9479 -10617 -9413
rect -12451 -9604 -12389 -9575
rect -12451 -9637 -12389 -9604
rect -8129 -9289 -8009 -9209
rect -9560 -9484 -9375 -9424
rect -11584 -9604 -11532 -9602
rect -11584 -9654 -11532 -9604
rect -8688 -9450 -8543 -9375
rect -10396 -9604 -10061 -9570
rect -10396 -9622 -10061 -9604
rect -9160 -9604 -9098 -9575
rect -9160 -9637 -9098 -9604
rect -8293 -9604 -8241 -9602
rect -8293 -9654 -8241 -9604
rect -24359 -10688 -23805 -10668
rect -24359 -10760 -23805 -10688
rect -23560 -10588 -23391 -10566
rect -23560 -10622 -23520 -10588
rect -23520 -10622 -23429 -10588
rect -23429 -10622 -23391 -10588
rect -23560 -10645 -23391 -10622
rect -24359 -10808 -24350 -10760
rect -24350 -10808 -24192 -10760
rect -24192 -10808 -24158 -10760
rect -24158 -10808 -24000 -10760
rect -24000 -10808 -23966 -10760
rect -23966 -10808 -23808 -10760
rect -23808 -10808 -23805 -10760
rect -24837 -11059 -24748 -10970
rect -24563 -11278 -24335 -11187
rect -23556 -11232 -23407 -11219
rect -24133 -11336 -23793 -11324
rect -24133 -11374 -23793 -11336
rect -24133 -11398 -23800 -11374
rect -23800 -11398 -23793 -11374
rect -23556 -11300 -23407 -11232
rect -23556 -11315 -23552 -11300
rect -23552 -11315 -23420 -11300
rect -23420 -11315 -23407 -11300
rect -24359 -11980 -23805 -11960
rect -24359 -12052 -23805 -11980
rect -23560 -11880 -23391 -11858
rect -23560 -11914 -23520 -11880
rect -23520 -11914 -23429 -11880
rect -23429 -11914 -23391 -11880
rect -23560 -11937 -23391 -11914
rect -24359 -12100 -24350 -12052
rect -24350 -12100 -24192 -12052
rect -24192 -12100 -24158 -12052
rect -24158 -12100 -24000 -12052
rect -24000 -12100 -23966 -12052
rect -23966 -12100 -23808 -12052
rect -23808 -12100 -23805 -12052
rect -22622 -10688 -22068 -10668
rect -22622 -10760 -22068 -10688
rect -21827 -10588 -21658 -10566
rect -21827 -10622 -21787 -10588
rect -21787 -10622 -21696 -10588
rect -21696 -10622 -21658 -10588
rect -21827 -10645 -21658 -10622
rect -22622 -10808 -22613 -10760
rect -22613 -10808 -22455 -10760
rect -22455 -10808 -22421 -10760
rect -22421 -10808 -22263 -10760
rect -22263 -10808 -22229 -10760
rect -22229 -10808 -22071 -10760
rect -22071 -10808 -22068 -10760
rect -22832 -11113 -22650 -11019
rect -20603 -10428 -19481 -10356
rect -19044 -10428 -17922 -10356
rect -17744 -10387 -17655 -10292
rect -17312 -10428 -16190 -10356
rect -15753 -10428 -14631 -10356
rect -14460 -10475 -14361 -10291
rect -14021 -10428 -12899 -10356
rect -12462 -10428 -11340 -10356
rect -11165 -10434 -11074 -10290
rect -10730 -10428 -9608 -10356
rect -9171 -10428 -8049 -10356
rect -22848 -11275 -22644 -11179
rect -21823 -11232 -21674 -11219
rect -22396 -11336 -22056 -11324
rect -22396 -11374 -22056 -11336
rect -22396 -11398 -22063 -11374
rect -22063 -11398 -22056 -11374
rect -21823 -11300 -21674 -11232
rect -21823 -11315 -21819 -11300
rect -21819 -11315 -21687 -11300
rect -21687 -11315 -21674 -11300
rect -20848 -11259 -20807 -11151
rect -20807 -11259 -20758 -11151
rect -20751 -11492 -20675 -11384
rect -19372 -11299 -19297 -11203
rect -19297 -11299 -19224 -11203
rect -19224 -11299 -19222 -11203
rect -19372 -11300 -19222 -11299
rect -17557 -11259 -17516 -11151
rect -17516 -11259 -17467 -11151
rect -19196 -11488 -19080 -11391
rect -20143 -11759 -20083 -11748
rect -20143 -11805 -20083 -11759
rect -20143 -11808 -20083 -11805
rect -18584 -11759 -18524 -11748
rect -18584 -11805 -18524 -11759
rect -17460 -11492 -17384 -11384
rect -16081 -11299 -16006 -11203
rect -16006 -11299 -15933 -11203
rect -15933 -11299 -15931 -11203
rect -16081 -11300 -15931 -11299
rect -14266 -11259 -14225 -11151
rect -14225 -11259 -14176 -11151
rect -15905 -11488 -15789 -11391
rect -17747 -11768 -17656 -11682
rect -16852 -11759 -16792 -11748
rect -18584 -11808 -18524 -11805
rect -16852 -11805 -16792 -11759
rect -16852 -11808 -16792 -11805
rect -15293 -11759 -15233 -11748
rect -15293 -11805 -15233 -11759
rect -14169 -11492 -14093 -11384
rect -12790 -11299 -12715 -11203
rect -12715 -11299 -12642 -11203
rect -12642 -11299 -12640 -11203
rect -12790 -11300 -12640 -11299
rect -10975 -11259 -10934 -11151
rect -10934 -11259 -10885 -11151
rect -12614 -11488 -12498 -11391
rect -14456 -11768 -14365 -11682
rect -13561 -11759 -13501 -11748
rect -15293 -11808 -15233 -11805
rect -13561 -11805 -13501 -11759
rect -13561 -11808 -13501 -11805
rect -12002 -11759 -11942 -11748
rect -12002 -11805 -11942 -11759
rect -10878 -11492 -10802 -11384
rect -9499 -11299 -9424 -11203
rect -9424 -11299 -9351 -11203
rect -9351 -11299 -9349 -11203
rect -9499 -11300 -9349 -11299
rect -5043 -11227 -4977 -11161
rect -9323 -11488 -9207 -11391
rect -11165 -11768 -11074 -11682
rect -10270 -11759 -10210 -11748
rect -12002 -11808 -11942 -11805
rect -10270 -11805 -10210 -11759
rect -10270 -11808 -10210 -11805
rect -8711 -11759 -8651 -11748
rect -8711 -11805 -8651 -11759
rect -7874 -11768 -7783 -11682
rect -8711 -11808 -8651 -11805
rect -22622 -11980 -22068 -11960
rect -22622 -12052 -22068 -11980
rect -21831 -11880 -21662 -11858
rect -21831 -11914 -21791 -11880
rect -21791 -11914 -21700 -11880
rect -21700 -11914 -21662 -11880
rect -21831 -11937 -21662 -11914
rect -22622 -12100 -22613 -12052
rect -22613 -12100 -22455 -12052
rect -22455 -12100 -22421 -12052
rect -22421 -12100 -22263 -12052
rect -22263 -12100 -22229 -12052
rect -22229 -12100 -22071 -12052
rect -22071 -12100 -22068 -12052
rect -24570 -12400 -24353 -12313
rect -21003 -11964 -20885 -11862
rect -19735 -11966 -19636 -11897
rect -19223 -11959 -19152 -11893
rect -16444 -11966 -16345 -11897
rect -15932 -11959 -15861 -11893
rect -13153 -11966 -13054 -11897
rect -12641 -11959 -12570 -11893
rect -9862 -11966 -9763 -11897
rect -9350 -11959 -9279 -11893
rect -20345 -12101 -20089 -12088
rect -20345 -12148 -20089 -12101
rect -20345 -12160 -20089 -12148
rect -19056 -12101 -18800 -12088
rect -19056 -12148 -18824 -12101
rect -18824 -12148 -18800 -12101
rect -19056 -12160 -18800 -12148
rect -18339 -12101 -18083 -12088
rect -18339 -12148 -18083 -12101
rect -18339 -12160 -18083 -12148
rect -17054 -12101 -16798 -12088
rect -17054 -12148 -16798 -12101
rect -17054 -12160 -16798 -12148
rect -15765 -12101 -15509 -12088
rect -15765 -12148 -15533 -12101
rect -15533 -12148 -15509 -12101
rect -15765 -12160 -15509 -12148
rect -15048 -12101 -14792 -12088
rect -15048 -12148 -14792 -12101
rect -15048 -12160 -14792 -12148
rect -13763 -12101 -13507 -12088
rect -13763 -12148 -13507 -12101
rect -13763 -12160 -13507 -12148
rect -12474 -12101 -12218 -12088
rect -12474 -12148 -12242 -12101
rect -12242 -12148 -12218 -12101
rect -12474 -12160 -12218 -12148
rect -11757 -12101 -11501 -12088
rect -11757 -12148 -11501 -12101
rect -11757 -12160 -11501 -12148
rect -10472 -12101 -10216 -12088
rect -10472 -12148 -10216 -12101
rect -10472 -12160 -10216 -12148
rect -9183 -12101 -8927 -12088
rect -9183 -12148 -8951 -12101
rect -8951 -12148 -8927 -12101
rect -9183 -12160 -8927 -12148
rect -8466 -12101 -8210 -12088
rect -8466 -12148 -8210 -12101
rect -8466 -12160 -8210 -12148
rect -22868 -12408 -22670 -12316
rect -24612 -12776 -24466 -12578
rect -23556 -12524 -23407 -12511
rect -24133 -12628 -23793 -12616
rect -24133 -12666 -23793 -12628
rect -24133 -12690 -23800 -12666
rect -23800 -12690 -23793 -12666
rect -23556 -12592 -23407 -12524
rect -23556 -12607 -23552 -12592
rect -23552 -12607 -23420 -12592
rect -23420 -12607 -23407 -12592
rect -22730 -12560 -22611 -12472
rect -21554 -12462 -21355 -12276
rect -21827 -12524 -21678 -12511
rect -22396 -12628 -22056 -12616
rect -22396 -12666 -22056 -12628
rect -22396 -12690 -22063 -12666
rect -22063 -12690 -22056 -12666
rect -21827 -12592 -21678 -12524
rect -21827 -12607 -21823 -12592
rect -21823 -12607 -21691 -12592
rect -21691 -12607 -21678 -12592
rect -20534 -12510 -20452 -12484
rect -20452 -12510 -20436 -12484
rect -20534 -12564 -20436 -12510
rect -19979 -12570 -19896 -12423
rect -19979 -12571 -19908 -12570
rect -19908 -12571 -19896 -12570
rect -19423 -12510 -19343 -12485
rect -19343 -12510 -19325 -12485
rect -19423 -12565 -19325 -12510
rect -20743 -12743 -20490 -12677
rect -18002 -12553 -17882 -12473
rect -19433 -12748 -19248 -12688
rect -17243 -12510 -17161 -12484
rect -17161 -12510 -17145 -12484
rect -17243 -12564 -17145 -12510
rect -18561 -12714 -18416 -12639
rect -20269 -12868 -19934 -12834
rect -20269 -12886 -19934 -12868
rect -16688 -12570 -16605 -12423
rect -16688 -12571 -16617 -12570
rect -16617 -12571 -16605 -12570
rect -16132 -12510 -16052 -12485
rect -16052 -12510 -16034 -12485
rect -16132 -12565 -16034 -12510
rect -17452 -12743 -17199 -12677
rect -19033 -12868 -18971 -12839
rect -19033 -12901 -18971 -12868
rect -14711 -12553 -14591 -12473
rect -16142 -12748 -15957 -12688
rect -18166 -12868 -18114 -12866
rect -18166 -12918 -18114 -12868
rect -13952 -12510 -13870 -12484
rect -13870 -12510 -13854 -12484
rect -13952 -12564 -13854 -12510
rect -15270 -12714 -15125 -12639
rect -16978 -12868 -16643 -12834
rect -16978 -12886 -16643 -12868
rect -13397 -12570 -13314 -12423
rect -13397 -12571 -13326 -12570
rect -13326 -12571 -13314 -12570
rect -12841 -12510 -12761 -12485
rect -12761 -12510 -12743 -12485
rect -12841 -12565 -12743 -12510
rect -14161 -12743 -13908 -12677
rect -15742 -12868 -15680 -12839
rect -15742 -12901 -15680 -12868
rect -11420 -12553 -11300 -12473
rect -12851 -12748 -12666 -12688
rect -14875 -12868 -14823 -12866
rect -14875 -12918 -14823 -12868
rect -10661 -12510 -10579 -12484
rect -10579 -12510 -10563 -12484
rect -10661 -12564 -10563 -12510
rect -11979 -12714 -11834 -12639
rect -13687 -12868 -13352 -12834
rect -13687 -12886 -13352 -12868
rect -10106 -12570 -10023 -12423
rect -10106 -12571 -10035 -12570
rect -10035 -12571 -10023 -12570
rect -9550 -12510 -9470 -12485
rect -9470 -12510 -9452 -12485
rect -9550 -12565 -9452 -12510
rect -10870 -12743 -10617 -12677
rect -12451 -12868 -12389 -12839
rect -12451 -12901 -12389 -12868
rect -8129 -12553 -8009 -12473
rect -9560 -12748 -9375 -12688
rect -11584 -12868 -11532 -12866
rect -11584 -12918 -11532 -12868
rect -8688 -12714 -8543 -12639
rect -10396 -12868 -10061 -12834
rect -10396 -12886 -10061 -12868
rect -9160 -12868 -9098 -12839
rect -9160 -12901 -9098 -12868
rect -8293 -12868 -8241 -12866
rect -8293 -12918 -8241 -12868
rect -7799 -12909 -7688 -12798
rect -11151 -13445 -11085 -13379
rect -768 -12902 -684 -12818
rect -14443 -13643 -14377 -13577
rect -5286 -13312 -5233 -13259
rect -5814 -13492 -5730 -13408
rect -17730 -13759 -17671 -13700
rect -4626 -13818 -4542 -13734
rect -1201 -13750 -1117 -13666
rect -14808 -13976 -14756 -13924
rect -5370 -13928 -5318 -13876
rect -21025 -14541 -20959 -14475
rect -24839 -15290 -24743 -15194
rect -23421 -15176 -23320 -15075
rect -24916 -15658 -24844 -15586
rect -24903 -15828 -24812 -15739
rect -24835 -16464 -24739 -16368
rect -23378 -16372 -23277 -16271
rect -24908 -16842 -24836 -16770
rect -24925 -17012 -24836 -16923
rect -24829 -17696 -24733 -17600
rect -23369 -17584 -23268 -17483
rect -24921 -18054 -24851 -17984
rect -24917 -18217 -24824 -18128
rect -24815 -18810 -24719 -18714
rect -23361 -18725 -23260 -18624
rect -24870 -19175 -24798 -19103
rect -24889 -19345 -24796 -19256
rect -24815 -20004 -24719 -19908
rect -23338 -19897 -23237 -19796
rect -24936 -20363 -24864 -20291
rect -20399 -17986 -20347 -17934
rect -21929 -18169 -21877 -18117
rect -20643 -18174 -20554 -18085
rect -20414 -18486 -20356 -18434
rect -21935 -18678 -21883 -18626
rect -20650 -18667 -20561 -18578
rect -18072 -15355 -17998 -15281
rect -17966 -15658 -17894 -15586
rect -16905 -15382 -16853 -15330
rect -18123 -15827 -18034 -15738
rect -18084 -16757 -18010 -16683
rect -18082 -17052 -18010 -16980
rect -16906 -16789 -16852 -16735
rect -18089 -17202 -18000 -17113
rect -18088 -18143 -18014 -18069
rect -18065 -18455 -17995 -18385
rect -17036 -18219 -16984 -18167
rect -18099 -18604 -18010 -18515
rect -19377 -18771 -19311 -18705
rect -20399 -18966 -20347 -18914
rect -21935 -19161 -21883 -19109
rect -20651 -19153 -20562 -19064
rect -14708 -14140 -14656 -14088
rect -16338 -18040 -16286 -17988
rect -15052 -18045 -14963 -17956
rect -12473 -15345 -12401 -14223
rect -10855 -14108 -10779 -14032
rect -5963 -14065 -5881 -13983
rect -6954 -14194 -6902 -14142
rect -11081 -14885 -11070 -14825
rect -11070 -14885 -11024 -14825
rect -11024 -14885 -11021 -14825
rect -10850 -14386 -10795 -14331
rect -12724 -15658 -12652 -15586
rect -12555 -15837 -12456 -15738
rect -14612 -16016 -14560 -15964
rect -16344 -18549 -16292 -18497
rect -15059 -18538 -14970 -18449
rect -14496 -16238 -14444 -16186
rect -20404 -19466 -20352 -19414
rect -21935 -19683 -21883 -19631
rect -18086 -19549 -18012 -19475
rect -20655 -19660 -20566 -19571
rect -18016 -19685 -17953 -19622
rect -20324 -19946 -20272 -19894
rect -16921 -19674 -16869 -19622
rect -16344 -19032 -16292 -18980
rect -15060 -19024 -14971 -18935
rect -10307 -14826 -10252 -14771
rect -5026 -14370 -4910 -14254
rect -4004 -14347 -3907 -14250
rect -6834 -14542 -6782 -14490
rect -8490 -15481 -8438 -15429
rect -8676 -15568 -8604 -15496
rect -7204 -15486 -7115 -15397
rect -5008 -14566 -4936 -14494
rect -3899 -14557 -3833 -14491
rect -6664 -14922 -6612 -14870
rect -8496 -15990 -8444 -15938
rect -7211 -15979 -7122 -15890
rect -8554 -16224 -8482 -16152
rect -5020 -14991 -4916 -14887
rect -4004 -14980 -3907 -14883
rect -4966 -15378 -4894 -15306
rect -5020 -15810 -4916 -15706
rect -4004 -15799 -3907 -15702
rect -2304 -14167 -2200 -14063
rect -1288 -14171 -1191 -14074
rect -2288 -14566 -2216 -14494
rect -2304 -14986 -2200 -14882
rect -1288 -14990 -1191 -14893
rect -2264 -15378 -2192 -15306
rect -2304 -15805 -2200 -15701
rect -1288 -15809 -1191 -15712
rect -4995 -16195 -4925 -16125
rect -2285 -16195 -2215 -16125
rect -8496 -16473 -8444 -16421
rect -7212 -16465 -7123 -16376
rect -5020 -16629 -4916 -16525
rect -4004 -16618 -3907 -16521
rect -2304 -16624 -2200 -16520
rect -8551 -16754 -8482 -16685
rect -12471 -18161 -12399 -17039
rect -11079 -17701 -11068 -17641
rect -11068 -17701 -11022 -17641
rect -11022 -17701 -11019 -17641
rect -12666 -18468 -12594 -18396
rect -12633 -18662 -12544 -18573
rect -16344 -19554 -16292 -19502
rect -15064 -19531 -14975 -19442
rect -8496 -16995 -8444 -16943
rect -7216 -16972 -7127 -16883
rect -8549 -17274 -8480 -17205
rect -5397 -17243 -5307 -17154
rect -8493 -17464 -8441 -17412
rect -7215 -17447 -7126 -17358
rect -8554 -17684 -8485 -17615
rect -8491 -17921 -8439 -17869
rect -7210 -17899 -7121 -17810
rect -8554 -18166 -8485 -18097
rect -8489 -18386 -8437 -18334
rect -7210 -18341 -7121 -18252
rect -8554 -18636 -8485 -18567
rect -8485 -18867 -8433 -18815
rect -7216 -18822 -7127 -18733
rect -8584 -19170 -8512 -19098
rect -17986 -19978 -17915 -19907
rect -21932 -20152 -21880 -20100
rect -16341 -20023 -16289 -19971
rect -20654 -20135 -20565 -20046
rect -15063 -20006 -14974 -19917
rect -14808 -19918 -14756 -19866
rect -24902 -20533 -24811 -20444
rect -20399 -20406 -20347 -20354
rect -21930 -20609 -21878 -20557
rect -20649 -20587 -20560 -20498
rect -24815 -21200 -24719 -21104
rect -18572 -20866 -18520 -20814
rect -23329 -21095 -23228 -20994
rect -21928 -21074 -21876 -21022
rect -20649 -21029 -20560 -20940
rect -18090 -20943 -18016 -20869
rect -24924 -21569 -24852 -21497
rect -24913 -21739 -24823 -21650
rect -18053 -21237 -17992 -21176
rect -16339 -20480 -16287 -20428
rect -15058 -20458 -14969 -20369
rect -16916 -21075 -16854 -21013
rect -18692 -21346 -18640 -21294
rect -21924 -21555 -21872 -21503
rect -17968 -21404 -17904 -21340
rect -20655 -21510 -20566 -21421
rect -16337 -20945 -16285 -20893
rect -15058 -20900 -14969 -20811
rect -24805 -22508 -24709 -22412
rect -23332 -22389 -23231 -22288
rect -24890 -22870 -24818 -22798
rect -24913 -23040 -24819 -22951
rect -18088 -22347 -18014 -22273
rect -18061 -22666 -17995 -22600
rect -16726 -22047 -16662 -21983
rect -18071 -22834 -17982 -22745
rect -16333 -21426 -16281 -21374
rect -15064 -21381 -14975 -21292
rect -24825 -23814 -24729 -23718
rect -23372 -23705 -23271 -23604
rect -18090 -23749 -18016 -23675
rect -24926 -24180 -24854 -24108
rect -18042 -24058 -17970 -23986
rect -16688 -23445 -16610 -23367
rect -18063 -24220 -17974 -24131
rect -24907 -24350 -24813 -24261
rect -18084 -25129 -18010 -25055
rect -17956 -25422 -17884 -25350
rect -16688 -24849 -16614 -24775
rect -12471 -21118 -12399 -19996
rect -11079 -20658 -11068 -20598
rect -11068 -20658 -11022 -20598
rect -11022 -20658 -11019 -20598
rect -12609 -21437 -12539 -21367
rect -12628 -21616 -12539 -21527
rect -12750 -22150 -12698 -22098
rect -12872 -22336 -12820 -22284
rect -12471 -23697 -12399 -22575
rect -11079 -23237 -11068 -23177
rect -11068 -23237 -11022 -23177
rect -11022 -23237 -11019 -23177
rect -12676 -24014 -12613 -23951
rect -12685 -24163 -12614 -24092
rect -5586 -20474 -5534 -20422
rect -5702 -22456 -5650 -22404
rect -6032 -24414 -5980 -24362
rect -5854 -24410 -5802 -24358
rect -1288 -16628 -1191 -16531
rect 407 -15493 473 -15427
rect -5000 -17021 -4937 -16958
rect -5236 -17372 -5184 -17320
rect -5020 -17448 -4916 -17344
rect -4004 -17437 -3907 -17340
rect -4979 -17841 -4918 -17780
rect -5020 -18267 -4916 -18163
rect -4004 -18256 -3907 -18159
rect -5006 -18654 -4934 -18582
rect -5020 -19086 -4916 -18982
rect -4004 -19075 -3907 -18978
rect -5014 -19502 -4942 -19430
rect -5020 -19905 -4916 -19801
rect -4004 -19894 -3907 -19797
rect -5166 -20128 -5094 -20056
rect -5020 -20724 -4916 -20620
rect -4004 -20713 -3907 -20616
rect -3906 -21130 -3822 -21046
rect -5130 -21608 -5047 -21525
rect -6032 -25036 -5980 -24984
rect -13016 -25164 -12964 -25112
rect -17976 -25642 -17887 -25553
rect -12471 -26465 -12399 -25343
rect -10479 -25193 -10393 -25107
rect -11079 -26005 -11068 -25945
rect -11068 -26005 -11022 -25945
rect -11022 -26005 -11019 -25945
rect -12743 -26805 -12682 -26744
rect -12748 -26998 -12684 -26934
rect -10152 -25634 -10048 -25530
rect -12471 -29098 -12399 -27976
rect -11079 -28638 -11068 -28578
rect -11068 -28638 -11022 -28578
rect -11022 -28638 -11019 -28578
rect -12724 -29446 -12652 -29374
rect -12727 -29626 -12638 -29537
rect -12471 -31707 -12399 -30585
rect -11079 -31247 -11068 -31187
rect -11068 -31247 -11022 -31187
rect -11022 -31247 -11019 -31187
rect -12758 -31990 -12686 -31918
rect -12791 -32176 -12702 -32087
rect -9857 -33009 -9764 -32916
rect -12473 -34327 -12401 -33205
rect -5854 -25086 -5802 -25034
rect -5854 -25794 -5802 -25742
rect -6032 -33168 -5980 -33116
rect -2291 -17021 -2228 -16958
rect -2304 -17443 -2200 -17339
rect -1288 -17447 -1191 -17350
rect -2269 -17841 -2208 -17780
rect -2608 -18064 -2524 -17980
rect -2304 -18262 -2200 -18158
rect -1288 -18266 -1191 -18169
rect -2294 -18654 -2222 -18582
rect -2304 -19081 -2200 -18977
rect -1288 -19085 -1191 -18988
rect -2300 -19502 -2228 -19430
rect -2304 -19900 -2200 -19796
rect -2420 -20128 -2348 -20056
rect -413 -19683 -347 -19617
rect -1288 -19904 -1191 -19807
rect -2310 -20533 -2194 -20417
rect -1288 -20537 -1191 -20440
rect -2751 -21819 -2680 -21748
rect -2914 -22610 -2830 -22526
rect -3082 -25958 -2998 -25874
rect -3260 -33356 -3176 -33272
rect -698 -33578 -614 -33494
rect -11081 -33867 -11070 -33807
rect -11070 -33867 -11024 -33807
rect -11024 -33867 -11021 -33807
rect 816 -17896 900 -17812
rect 674 -21956 758 -21872
rect 490 -22780 574 -22696
rect 320 -26148 404 -26064
rect 1367 -20283 1433 -20217
rect 4164 -1686 4248 -1602
rect 4164 -13750 4248 -13666
rect 3886 -21130 3970 -21046
rect 1221 -21455 1287 -21389
rect 5558 -665 5627 -649
rect 5558 -718 5577 -665
rect 5577 -718 5611 -665
rect 5611 -718 5627 -665
rect 5901 -1283 5970 -1214
rect 5734 -1352 5786 -1300
rect 5998 -665 6067 -649
rect 5998 -718 6017 -665
rect 6017 -718 6051 -665
rect 6051 -718 6067 -665
rect 6172 -1291 6224 -1281
rect 6172 -1333 6224 -1291
rect 6341 -1285 6410 -1216
rect 6438 -665 6507 -649
rect 6438 -718 6457 -665
rect 6457 -718 6491 -665
rect 6491 -718 6507 -665
rect 5998 -1822 6067 -1753
rect 6612 -1291 6664 -1272
rect 6612 -1324 6664 -1291
rect 6438 -1957 6507 -1888
rect 7106 -1719 7158 -1667
rect 7113 -1813 7165 -1761
rect 7327 -1916 7393 -1850
rect 8069 -1720 8122 -1668
rect 8057 -1812 8109 -1760
rect 8424 -1895 8493 -1843
rect 7106 -2277 7172 -2211
rect 7227 -2826 7372 -2813
rect 7372 -2826 7405 -2813
rect 7227 -2978 7405 -2826
rect 9002 -1719 9055 -1667
rect 9000 -1817 9052 -1765
rect 8989 -1909 9042 -1856
rect 8050 -2381 8116 -2315
rect 7872 -2534 7938 -2468
rect 8162 -2826 8320 -2813
rect 8320 -2826 8340 -2813
rect 7227 -2991 7372 -2978
rect 7372 -2991 7405 -2978
rect 7102 -3703 7168 -3637
rect 7853 -3327 7919 -3261
rect 8162 -2978 8340 -2826
rect 8986 -2075 9052 -2009
rect 9933 -1719 9986 -1667
rect 9935 -1817 9987 -1765
rect 10262 -1881 10331 -1812
rect 9798 -2032 9864 -1966
rect 8818 -2280 8884 -2214
rect 9098 -2826 9256 -2813
rect 9256 -2826 9276 -2813
rect 8162 -2991 8320 -2978
rect 8320 -2991 8340 -2978
rect 6780 -3948 6849 -3879
rect 6066 -4048 6132 -3982
rect 6941 -4142 7007 -4076
rect 8050 -3824 8116 -3758
rect 9098 -2978 9276 -2826
rect 10860 -1822 10926 -1756
rect 10858 -1916 10924 -1850
rect 10850 -2010 10915 -1944
rect 9917 -2171 9983 -2105
rect 10029 -2826 10187 -2813
rect 10187 -2826 10206 -2813
rect 9098 -2991 9256 -2978
rect 9256 -2991 9276 -2978
rect 8837 -3737 8903 -3671
rect 8989 -3483 9055 -3417
rect 8401 -3959 8465 -3895
rect 8079 -4043 8131 -3991
rect 8063 -4137 8128 -4085
rect 10029 -2977 10206 -2826
rect 10956 -2826 11114 -2813
rect 11114 -2826 11134 -2813
rect 10029 -2990 10187 -2977
rect 10187 -2990 10206 -2977
rect 9917 -3605 9983 -3539
rect 8993 -3954 9059 -3888
rect 9001 -4048 9067 -3982
rect 8992 -4137 9057 -4085
rect 9807 -3829 9873 -3765
rect 10956 -2978 11134 -2826
rect 12189 -1870 12410 -1667
rect 10956 -2991 11114 -2978
rect 11114 -2991 11134 -2978
rect 10264 -3955 10324 -3895
rect 9937 -4047 10003 -3981
rect 9951 -4091 10016 -4085
rect 9951 -4125 10013 -4091
rect 10013 -4125 10016 -4091
rect 9951 -4137 10016 -4125
rect 12233 -3340 12352 -3324
rect 12233 -3443 12352 -3340
rect 12960 -3484 13079 -3365
rect 10850 -3860 10916 -3794
rect 10888 -3954 10954 -3888
rect 10859 -4048 10925 -3982
rect 11894 -4603 12136 -4361
rect 5558 -5093 5627 -5077
rect 5558 -5146 5577 -5093
rect 5577 -5146 5611 -5093
rect 5611 -5146 5627 -5093
rect 5901 -5711 5970 -5642
rect 5734 -5780 5786 -5728
rect 5998 -5093 6067 -5077
rect 5998 -5146 6017 -5093
rect 6017 -5146 6051 -5093
rect 6051 -5146 6067 -5093
rect 5419 -6503 5485 -6437
rect 6172 -5719 6224 -5709
rect 6172 -5761 6224 -5719
rect 6341 -5713 6410 -5644
rect 6438 -5093 6507 -5077
rect 6438 -5146 6457 -5093
rect 6457 -5146 6491 -5093
rect 6491 -5146 6507 -5093
rect 5998 -6250 6067 -6181
rect 6612 -5719 6664 -5700
rect 6612 -5752 6664 -5719
rect 6438 -6385 6507 -6316
rect 7106 -6147 7158 -6095
rect 7113 -6241 7165 -6189
rect 7327 -6344 7393 -6278
rect 8069 -6148 8122 -6096
rect 8057 -6240 8109 -6188
rect 8424 -6323 8493 -6271
rect 7106 -6705 7172 -6639
rect 7227 -7254 7372 -7241
rect 7372 -7254 7405 -7241
rect 7227 -7406 7405 -7254
rect 9002 -6147 9055 -6095
rect 9000 -6245 9052 -6193
rect 8989 -6337 9042 -6284
rect 8050 -6809 8116 -6743
rect 7872 -6962 7938 -6896
rect 8162 -7254 8320 -7241
rect 8320 -7254 8340 -7241
rect 7227 -7419 7372 -7406
rect 7372 -7419 7405 -7406
rect 7102 -8131 7168 -8065
rect 7853 -7755 7919 -7689
rect 8162 -7406 8340 -7254
rect 8986 -6503 9052 -6437
rect 9933 -6147 9986 -6095
rect 9935 -6245 9987 -6193
rect 10262 -6309 10331 -6240
rect 9798 -6460 9864 -6394
rect 8818 -6708 8884 -6642
rect 9098 -7254 9256 -7241
rect 9256 -7254 9276 -7241
rect 8162 -7419 8320 -7406
rect 8320 -7419 8340 -7406
rect 6780 -8376 6849 -8307
rect 6066 -8476 6132 -8410
rect 6941 -8570 7007 -8504
rect 8050 -8252 8116 -8186
rect 9098 -7406 9276 -7254
rect 10860 -6250 10926 -6184
rect 10858 -6344 10924 -6278
rect 10850 -6438 10915 -6372
rect 9917 -6599 9983 -6533
rect 10029 -7254 10187 -7241
rect 10187 -7254 10206 -7241
rect 9098 -7419 9256 -7406
rect 9256 -7419 9276 -7406
rect 8837 -8165 8903 -8099
rect 8989 -7911 9055 -7845
rect 8401 -8387 8465 -8323
rect 8079 -8471 8131 -8419
rect 8063 -8565 8128 -8513
rect 10029 -7405 10206 -7254
rect 10956 -7254 11114 -7241
rect 11114 -7254 11134 -7241
rect 10029 -7418 10187 -7405
rect 10187 -7418 10206 -7405
rect 9917 -8033 9983 -7967
rect 8993 -8382 9059 -8316
rect 9001 -8476 9067 -8410
rect 8992 -8565 9057 -8513
rect 9807 -8257 9873 -8193
rect 10956 -7406 11134 -7254
rect 12189 -6298 12410 -6095
rect 10956 -7419 11114 -7406
rect 11114 -7419 11134 -7406
rect 10264 -8383 10324 -8323
rect 9937 -8475 10003 -8409
rect 9951 -8519 10016 -8513
rect 9951 -8553 10013 -8519
rect 10013 -8553 10016 -8519
rect 9951 -8565 10016 -8553
rect 12233 -7768 12352 -7752
rect 12233 -7871 12352 -7768
rect 12960 -7912 13079 -7793
rect 10850 -8288 10916 -8222
rect 10888 -8382 10954 -8316
rect 10859 -8476 10925 -8410
rect 11894 -9031 12136 -8789
rect 5558 -9721 5627 -9705
rect 5558 -9774 5577 -9721
rect 5577 -9774 5611 -9721
rect 5611 -9774 5627 -9721
rect 5901 -10339 5970 -10270
rect 5734 -10408 5786 -10356
rect 5998 -9721 6067 -9705
rect 5998 -9774 6017 -9721
rect 6017 -9774 6051 -9721
rect 6051 -9774 6067 -9721
rect 5426 -11131 5492 -11065
rect 5354 -13118 5420 -13052
rect 6172 -10347 6224 -10337
rect 6172 -10389 6224 -10347
rect 6341 -10341 6410 -10272
rect 6438 -9721 6507 -9705
rect 6438 -9774 6457 -9721
rect 6457 -9774 6491 -9721
rect 6491 -9774 6507 -9721
rect 5998 -10878 6067 -10809
rect 6612 -10347 6664 -10328
rect 6612 -10380 6664 -10347
rect 6438 -11013 6507 -10944
rect 7106 -10775 7158 -10723
rect 7113 -10869 7165 -10817
rect 7327 -10972 7393 -10906
rect 8069 -10776 8122 -10724
rect 8057 -10868 8109 -10816
rect 8424 -10951 8493 -10899
rect 7106 -11333 7172 -11267
rect 7227 -11882 7372 -11869
rect 7372 -11882 7405 -11869
rect 7227 -12034 7405 -11882
rect 9002 -10775 9055 -10723
rect 9000 -10873 9052 -10821
rect 8989 -10965 9042 -10912
rect 8050 -11437 8116 -11371
rect 7872 -11590 7938 -11524
rect 8162 -11882 8320 -11869
rect 8320 -11882 8340 -11869
rect 7227 -12047 7372 -12034
rect 7372 -12047 7405 -12034
rect 7102 -12759 7168 -12693
rect 7853 -12383 7919 -12317
rect 8162 -12034 8340 -11882
rect 8986 -11131 9052 -11065
rect 9933 -10775 9986 -10723
rect 9935 -10873 9987 -10821
rect 10262 -10937 10331 -10868
rect 9798 -11088 9864 -11022
rect 8818 -11336 8884 -11270
rect 9098 -11882 9256 -11869
rect 9256 -11882 9276 -11869
rect 8162 -12047 8320 -12034
rect 8320 -12047 8340 -12034
rect 6780 -13004 6849 -12935
rect 6066 -13104 6132 -13038
rect 6941 -13198 7007 -13132
rect 8050 -12880 8116 -12814
rect 9098 -12034 9276 -11882
rect 10860 -10878 10926 -10812
rect 10858 -10972 10924 -10906
rect 10850 -11066 10915 -11000
rect 9917 -11227 9983 -11161
rect 10029 -11882 10187 -11869
rect 10187 -11882 10206 -11869
rect 9098 -12047 9256 -12034
rect 9256 -12047 9276 -12034
rect 8837 -12793 8903 -12727
rect 8989 -12539 9055 -12473
rect 8401 -13015 8465 -12951
rect 8079 -13099 8131 -13047
rect 8063 -13193 8128 -13141
rect 10029 -12033 10206 -11882
rect 10956 -11882 11114 -11869
rect 11114 -11882 11134 -11869
rect 10029 -12046 10187 -12033
rect 10187 -12046 10206 -12033
rect 9917 -12661 9983 -12595
rect 8993 -13010 9059 -12944
rect 9001 -13104 9067 -13038
rect 8992 -13193 9057 -13141
rect 9807 -12885 9873 -12821
rect 10956 -12034 11134 -11882
rect 12189 -10926 12410 -10723
rect 10956 -12047 11114 -12034
rect 11114 -12047 11134 -12034
rect 10264 -13011 10324 -12951
rect 9937 -13103 10003 -13037
rect 9951 -13147 10016 -13141
rect 9951 -13181 10013 -13147
rect 10013 -13181 10016 -13147
rect 9951 -13193 10016 -13181
rect 12233 -12396 12352 -12380
rect 12233 -12499 12352 -12396
rect 12960 -12540 13079 -12421
rect 10850 -12916 10916 -12850
rect 10888 -13010 10954 -12944
rect 10859 -13104 10925 -13038
rect 11894 -13659 12136 -13417
rect 5558 -14249 5627 -14233
rect 5558 -14302 5577 -14249
rect 5577 -14302 5611 -14249
rect 5611 -14302 5627 -14249
rect 5901 -14867 5970 -14798
rect 5734 -14936 5786 -14884
rect 5998 -14249 6067 -14233
rect 5998 -14302 6017 -14249
rect 6017 -14302 6051 -14249
rect 6051 -14302 6067 -14249
rect 5407 -17619 5473 -17552
rect 6172 -14875 6224 -14865
rect 6172 -14917 6224 -14875
rect 6341 -14869 6410 -14800
rect 6438 -14249 6507 -14233
rect 6438 -14302 6457 -14249
rect 6457 -14302 6491 -14249
rect 6491 -14302 6507 -14249
rect 5998 -15406 6067 -15337
rect 6612 -14875 6664 -14856
rect 6612 -14908 6664 -14875
rect 6438 -15541 6507 -15472
rect 7106 -15303 7158 -15251
rect 7113 -15397 7165 -15345
rect 7327 -15500 7393 -15434
rect 8069 -15304 8122 -15252
rect 8057 -15396 8109 -15344
rect 8424 -15479 8493 -15427
rect 7106 -15861 7172 -15795
rect 7227 -16410 7372 -16397
rect 7372 -16410 7405 -16397
rect 7227 -16562 7405 -16410
rect 9002 -15303 9055 -15251
rect 9000 -15401 9052 -15349
rect 8989 -15493 9042 -15440
rect 8050 -15965 8116 -15899
rect 7872 -16118 7938 -16052
rect 8162 -16410 8320 -16397
rect 8320 -16410 8340 -16397
rect 7227 -16575 7372 -16562
rect 7372 -16575 7405 -16562
rect 7102 -17287 7168 -17221
rect 7853 -16911 7919 -16845
rect 8162 -16562 8340 -16410
rect 8986 -15659 9052 -15593
rect 9933 -15303 9986 -15251
rect 9935 -15401 9987 -15349
rect 10262 -15465 10331 -15396
rect 9798 -15616 9864 -15550
rect 8818 -15864 8884 -15798
rect 9098 -16410 9256 -16397
rect 9256 -16410 9276 -16397
rect 8162 -16575 8320 -16562
rect 8320 -16575 8340 -16562
rect 6780 -17532 6849 -17463
rect 6066 -17632 6132 -17566
rect 6941 -17726 7007 -17660
rect 8050 -17408 8116 -17342
rect 9098 -16562 9276 -16410
rect 10860 -15406 10926 -15340
rect 10858 -15500 10924 -15434
rect 10850 -15594 10915 -15528
rect 9917 -15755 9983 -15689
rect 10029 -16410 10187 -16397
rect 10187 -16410 10206 -16397
rect 9098 -16575 9256 -16562
rect 9256 -16575 9276 -16562
rect 8837 -17321 8903 -17255
rect 8989 -17067 9055 -17001
rect 8401 -17543 8465 -17479
rect 8079 -17627 8131 -17575
rect 8063 -17721 8128 -17669
rect 10029 -16561 10206 -16410
rect 10956 -16410 11114 -16397
rect 11114 -16410 11134 -16397
rect 10029 -16574 10187 -16561
rect 10187 -16574 10206 -16561
rect 9917 -17189 9983 -17123
rect 8993 -17538 9059 -17472
rect 9001 -17632 9067 -17566
rect 8992 -17721 9057 -17669
rect 9807 -17413 9873 -17349
rect 10956 -16562 11134 -16410
rect 12189 -15454 12410 -15251
rect 10956 -16575 11114 -16562
rect 11114 -16575 11134 -16562
rect 10264 -17539 10324 -17479
rect 9937 -17631 10003 -17565
rect 9951 -17675 10016 -17669
rect 9951 -17709 10013 -17675
rect 10013 -17709 10016 -17675
rect 9951 -17721 10016 -17709
rect 12233 -16924 12352 -16908
rect 12233 -17027 12352 -16924
rect 12960 -17068 13079 -16949
rect 10850 -17444 10916 -17378
rect 10888 -17538 10954 -17472
rect 10859 -17632 10925 -17566
rect 16285 -16814 16543 -16737
rect 16285 -16927 16541 -16814
rect 16541 -16927 16543 -16814
rect 16285 -16995 16543 -16927
rect 4745 -21455 4811 -21389
rect 11894 -18187 12136 -17945
rect 15551 -18658 15695 -18514
rect 17526 -18154 17659 -18021
rect 5558 -18777 5627 -18761
rect 5558 -18830 5577 -18777
rect 5577 -18830 5611 -18777
rect 5611 -18830 5627 -18777
rect 5901 -19395 5970 -19326
rect 5734 -19464 5786 -19412
rect 5998 -18777 6067 -18761
rect 5998 -18830 6017 -18777
rect 6017 -18830 6051 -18777
rect 6051 -18830 6067 -18777
rect 6172 -19403 6224 -19393
rect 6172 -19445 6224 -19403
rect 6341 -19397 6410 -19328
rect 6438 -18777 6507 -18761
rect 6438 -18830 6457 -18777
rect 6457 -18830 6491 -18777
rect 6491 -18830 6507 -18777
rect 5998 -19934 6067 -19865
rect 6612 -19403 6664 -19384
rect 6612 -19436 6664 -19403
rect 6438 -20069 6507 -20000
rect 17977 -18940 18048 -18869
rect 7106 -19831 7158 -19779
rect 7113 -19925 7165 -19873
rect 7327 -20028 7393 -19962
rect 8069 -19832 8122 -19780
rect 8057 -19924 8109 -19872
rect 8424 -20007 8493 -19955
rect 7106 -20389 7172 -20323
rect 7227 -20938 7372 -20925
rect 7372 -20938 7405 -20925
rect 7227 -21090 7405 -20938
rect 9002 -19831 9055 -19779
rect 9000 -19929 9052 -19877
rect 8989 -20021 9042 -19968
rect 8050 -20493 8116 -20427
rect 7872 -20646 7938 -20580
rect 8162 -20938 8320 -20925
rect 8320 -20938 8340 -20925
rect 7227 -21103 7372 -21090
rect 7372 -21103 7405 -21090
rect 7102 -21815 7168 -21749
rect 7853 -21439 7919 -21373
rect 8162 -21090 8340 -20938
rect 8986 -20187 9052 -20121
rect 9933 -19831 9986 -19779
rect 9935 -19929 9987 -19877
rect 10262 -19993 10331 -19924
rect 9798 -20144 9864 -20078
rect 8818 -20392 8884 -20326
rect 9098 -20938 9256 -20925
rect 9256 -20938 9276 -20925
rect 8162 -21103 8320 -21090
rect 8320 -21103 8340 -21090
rect 6780 -22060 6849 -21991
rect 6066 -22160 6132 -22094
rect 6941 -22254 7007 -22188
rect 8050 -21936 8116 -21870
rect 9098 -21090 9276 -20938
rect 10860 -19934 10926 -19868
rect 10858 -20028 10924 -19962
rect 10850 -20122 10915 -20056
rect 9917 -20283 9983 -20217
rect 10029 -20938 10187 -20925
rect 10187 -20938 10206 -20925
rect 9098 -21103 9256 -21090
rect 9256 -21103 9276 -21090
rect 8837 -21849 8903 -21783
rect 8989 -21595 9055 -21529
rect 8401 -22071 8465 -22007
rect 8079 -22155 8131 -22103
rect 8063 -22249 8128 -22197
rect 10029 -21089 10206 -20938
rect 10956 -20938 11114 -20925
rect 11114 -20938 11134 -20925
rect 10029 -21102 10187 -21089
rect 10187 -21102 10206 -21089
rect 9917 -21717 9983 -21651
rect 8993 -22066 9059 -22000
rect 9001 -22160 9067 -22094
rect 8992 -22249 9057 -22197
rect 9807 -21941 9873 -21877
rect 10956 -21090 11134 -20938
rect 12189 -19982 12410 -19779
rect 10956 -21103 11114 -21090
rect 11114 -21103 11134 -21090
rect 10264 -22067 10324 -22007
rect 9937 -22159 10003 -22093
rect 9951 -22203 10016 -22197
rect 9951 -22237 10013 -22203
rect 10013 -22237 10016 -22203
rect 9951 -22249 10016 -22237
rect 12233 -21452 12352 -21436
rect 12233 -21555 12352 -21452
rect 12960 -21596 13079 -21477
rect 10850 -21972 10916 -21906
rect 10888 -22066 10954 -22000
rect 10859 -22160 10925 -22094
rect 11894 -22715 12136 -22473
rect 5558 -23305 5627 -23289
rect 5558 -23358 5577 -23305
rect 5577 -23358 5611 -23305
rect 5611 -23358 5627 -23305
rect 5901 -23923 5970 -23854
rect 5734 -23992 5786 -23940
rect 5998 -23305 6067 -23289
rect 5998 -23358 6017 -23305
rect 6017 -23358 6051 -23305
rect 6051 -23358 6067 -23305
rect 5732 -24715 5798 -24649
rect 5317 -24811 5383 -24745
rect 6172 -23931 6224 -23921
rect 6172 -23973 6224 -23931
rect 6341 -23925 6410 -23856
rect 6438 -23305 6507 -23289
rect 6438 -23358 6457 -23305
rect 6457 -23358 6491 -23305
rect 6491 -23358 6507 -23305
rect 5998 -24462 6067 -24393
rect 6612 -23931 6664 -23912
rect 6612 -23964 6664 -23931
rect 6438 -24597 6507 -24528
rect 7106 -24359 7158 -24307
rect 7113 -24453 7165 -24401
rect 7327 -24556 7393 -24490
rect 8069 -24360 8122 -24308
rect 8057 -24452 8109 -24400
rect 8424 -24535 8493 -24483
rect 7106 -24917 7172 -24851
rect 7227 -25466 7372 -25453
rect 7372 -25466 7405 -25453
rect 7227 -25618 7405 -25466
rect 9002 -24359 9055 -24307
rect 9000 -24457 9052 -24405
rect 8989 -24549 9042 -24496
rect 8050 -25021 8116 -24955
rect 7872 -25174 7938 -25108
rect 8162 -25466 8320 -25453
rect 8320 -25466 8340 -25453
rect 7227 -25631 7372 -25618
rect 7372 -25631 7405 -25618
rect 7102 -26343 7168 -26277
rect 7853 -25967 7919 -25901
rect 8162 -25618 8340 -25466
rect 8986 -24715 9052 -24649
rect 9933 -24359 9986 -24307
rect 9935 -24457 9987 -24405
rect 10262 -24521 10331 -24452
rect 9798 -24672 9864 -24606
rect 8818 -24920 8884 -24854
rect 9098 -25466 9256 -25453
rect 9256 -25466 9276 -25453
rect 8162 -25631 8320 -25618
rect 8320 -25631 8340 -25618
rect 6780 -26588 6849 -26519
rect 6066 -26688 6132 -26622
rect 6941 -26782 7007 -26716
rect 8050 -26464 8116 -26398
rect 9098 -25618 9276 -25466
rect 10860 -24462 10926 -24396
rect 10858 -24556 10924 -24490
rect 10850 -24650 10915 -24584
rect 9917 -24811 9983 -24745
rect 10029 -25466 10187 -25453
rect 10187 -25466 10206 -25453
rect 9098 -25631 9256 -25618
rect 9256 -25631 9276 -25618
rect 8837 -26377 8903 -26311
rect 8989 -26123 9055 -26057
rect 8401 -26599 8465 -26535
rect 8079 -26683 8131 -26631
rect 8063 -26777 8128 -26725
rect 10029 -25617 10206 -25466
rect 10956 -25466 11114 -25453
rect 11114 -25466 11134 -25453
rect 10029 -25630 10187 -25617
rect 10187 -25630 10206 -25617
rect 9917 -26245 9983 -26179
rect 8993 -26594 9059 -26528
rect 9001 -26688 9067 -26622
rect 8992 -26777 9057 -26725
rect 9807 -26469 9873 -26405
rect 10956 -25618 11134 -25466
rect 12189 -24510 12410 -24307
rect 10956 -25631 11114 -25618
rect 11114 -25631 11134 -25618
rect 10264 -26595 10324 -26535
rect 9937 -26687 10003 -26621
rect 9951 -26731 10016 -26725
rect 9951 -26765 10013 -26731
rect 10013 -26765 10016 -26731
rect 9951 -26777 10016 -26765
rect 12233 -25980 12352 -25964
rect 12233 -26083 12352 -25980
rect 12960 -26124 13079 -26005
rect 10850 -26500 10916 -26434
rect 10888 -26594 10954 -26528
rect 10859 -26688 10925 -26622
rect 11894 -27243 12136 -27001
rect 5558 -27833 5627 -27817
rect 5558 -27886 5577 -27833
rect 5577 -27886 5611 -27833
rect 5611 -27886 5627 -27833
rect 4860 -29337 4919 -29278
rect 5901 -28451 5970 -28382
rect 5734 -28520 5786 -28468
rect 5998 -27833 6067 -27817
rect 5998 -27886 6017 -27833
rect 6017 -27886 6051 -27833
rect 6051 -27886 6067 -27833
rect 5454 -29243 5520 -29177
rect 6172 -28459 6224 -28449
rect 6172 -28501 6224 -28459
rect 6341 -28453 6410 -28384
rect 6438 -27833 6507 -27817
rect 6438 -27886 6457 -27833
rect 6457 -27886 6491 -27833
rect 6491 -27886 6507 -27833
rect 5998 -28990 6067 -28921
rect 6612 -28459 6664 -28440
rect 6612 -28492 6664 -28459
rect 6438 -29125 6507 -29056
rect 7106 -28887 7158 -28835
rect 7113 -28981 7165 -28929
rect 7327 -29084 7393 -29018
rect 8069 -28888 8122 -28836
rect 8057 -28980 8109 -28928
rect 8424 -29063 8493 -29011
rect 7106 -29445 7172 -29379
rect 7227 -29994 7372 -29981
rect 7372 -29994 7405 -29981
rect 7227 -30146 7405 -29994
rect 9002 -28887 9055 -28835
rect 9000 -28985 9052 -28933
rect 8989 -29077 9042 -29024
rect 8050 -29549 8116 -29483
rect 7872 -29702 7938 -29636
rect 8162 -29994 8320 -29981
rect 8320 -29994 8340 -29981
rect 7227 -30159 7372 -30146
rect 7372 -30159 7405 -30146
rect 7102 -30871 7168 -30805
rect 7853 -30495 7919 -30429
rect 8162 -30146 8340 -29994
rect 8986 -29243 9052 -29177
rect 9933 -28887 9986 -28835
rect 9935 -28985 9987 -28933
rect 10262 -29049 10331 -28980
rect 9798 -29200 9864 -29134
rect 8818 -29448 8884 -29382
rect 9098 -29994 9256 -29981
rect 9256 -29994 9276 -29981
rect 8162 -30159 8320 -30146
rect 8320 -30159 8340 -30146
rect 6780 -31116 6849 -31047
rect 6066 -31216 6132 -31150
rect 6941 -31310 7007 -31244
rect 8050 -30992 8116 -30926
rect 9098 -30146 9276 -29994
rect 10860 -28990 10926 -28924
rect 10858 -29084 10924 -29018
rect 10850 -29178 10915 -29112
rect 9917 -29339 9983 -29273
rect 10029 -29994 10187 -29981
rect 10187 -29994 10206 -29981
rect 9098 -30159 9256 -30146
rect 9256 -30159 9276 -30146
rect 8837 -30905 8903 -30839
rect 8989 -30651 9055 -30585
rect 8401 -31127 8465 -31063
rect 8079 -31211 8131 -31159
rect 8063 -31305 8128 -31253
rect 10029 -30145 10206 -29994
rect 10956 -29994 11114 -29981
rect 11114 -29994 11134 -29981
rect 10029 -30158 10187 -30145
rect 10187 -30158 10206 -30145
rect 9917 -30773 9983 -30707
rect 8993 -31122 9059 -31056
rect 9001 -31216 9067 -31150
rect 8992 -31305 9057 -31253
rect 9807 -30997 9873 -30933
rect 10956 -30146 11134 -29994
rect 12189 -29038 12410 -28835
rect 10956 -30159 11114 -30146
rect 11114 -30159 11134 -30146
rect 10264 -31123 10324 -31063
rect 9937 -31215 10003 -31149
rect 9951 -31259 10016 -31253
rect 9951 -31293 10013 -31259
rect 10013 -31293 10016 -31259
rect 9951 -31305 10016 -31293
rect 12233 -30508 12352 -30492
rect 12233 -30611 12352 -30508
rect 12960 -30652 13079 -30533
rect 10850 -31028 10916 -30962
rect 10888 -31122 10954 -31056
rect 10859 -31216 10925 -31150
rect 11894 -31771 12136 -31529
rect 5558 -32361 5627 -32345
rect 5558 -32414 5577 -32361
rect 5577 -32414 5611 -32361
rect 5611 -32414 5627 -32361
rect 5901 -32979 5970 -32910
rect 5734 -33048 5786 -32996
rect 5998 -32361 6067 -32345
rect 5998 -32414 6017 -32361
rect 6017 -32414 6051 -32361
rect 6051 -32414 6067 -32361
rect 5425 -33771 5491 -33705
rect 3663 -33867 3729 -33801
rect -12582 -34576 -12510 -34504
rect -12726 -34760 -12637 -34671
rect 6172 -32987 6224 -32977
rect 6172 -33029 6224 -32987
rect 6341 -32981 6410 -32912
rect 6438 -32361 6507 -32345
rect 6438 -32414 6457 -32361
rect 6457 -32414 6491 -32361
rect 6491 -32414 6507 -32361
rect 5998 -33518 6067 -33449
rect 6612 -32987 6664 -32968
rect 6612 -33020 6664 -32987
rect 6438 -33653 6507 -33584
rect 7106 -33415 7158 -33363
rect 7113 -33509 7165 -33457
rect 7327 -33612 7393 -33546
rect 8069 -33416 8122 -33364
rect 8057 -33508 8109 -33456
rect 8424 -33591 8493 -33539
rect 7106 -33973 7172 -33907
rect 7227 -34522 7372 -34509
rect 7372 -34522 7405 -34509
rect 7227 -34674 7405 -34522
rect 9002 -33415 9055 -33363
rect 9000 -33513 9052 -33461
rect 8989 -33605 9042 -33552
rect 8050 -34077 8116 -34011
rect 7872 -34230 7938 -34164
rect 8162 -34522 8320 -34509
rect 8320 -34522 8340 -34509
rect 7227 -34687 7372 -34674
rect 7372 -34687 7405 -34674
rect 7102 -35399 7168 -35333
rect 7853 -35023 7919 -34957
rect 8162 -34674 8340 -34522
rect 8986 -33771 9052 -33705
rect 9933 -33415 9986 -33363
rect 9935 -33513 9987 -33461
rect 10262 -33577 10331 -33508
rect 9798 -33728 9864 -33662
rect 8818 -33976 8884 -33910
rect 9098 -34522 9256 -34509
rect 9256 -34522 9276 -34509
rect 8162 -34687 8320 -34674
rect 8320 -34687 8340 -34674
rect 6780 -35644 6849 -35575
rect 6066 -35744 6132 -35678
rect 6941 -35838 7007 -35772
rect 8050 -35520 8116 -35454
rect 9098 -34674 9276 -34522
rect 10860 -33518 10926 -33452
rect 10858 -33612 10924 -33546
rect 10850 -33706 10915 -33640
rect 9917 -33867 9983 -33801
rect 10029 -34522 10187 -34509
rect 10187 -34522 10206 -34509
rect 9098 -34687 9256 -34674
rect 9256 -34687 9276 -34674
rect 8837 -35433 8903 -35367
rect 8989 -35179 9055 -35113
rect 8401 -35655 8465 -35591
rect 8079 -35739 8131 -35687
rect 8063 -35833 8128 -35781
rect 10029 -34673 10206 -34522
rect 10956 -34522 11114 -34509
rect 11114 -34522 11134 -34509
rect 10029 -34686 10187 -34673
rect 10187 -34686 10206 -34673
rect 9917 -35301 9983 -35235
rect 8993 -35650 9059 -35584
rect 9001 -35744 9067 -35678
rect 8992 -35833 9057 -35781
rect 9807 -35525 9873 -35461
rect 10956 -34674 11134 -34522
rect 12189 -33566 12410 -33363
rect 16221 -20245 16480 -20177
rect 16221 -20358 16480 -20245
rect 16221 -20436 16480 -20358
rect 10956 -34687 11114 -34674
rect 11114 -34687 11134 -34674
rect 10264 -35651 10324 -35591
rect 9937 -35743 10003 -35677
rect 9951 -35787 10016 -35781
rect 9951 -35821 10013 -35787
rect 10013 -35821 10016 -35787
rect 9951 -35833 10016 -35821
rect 12233 -35036 12352 -35020
rect 12233 -35139 12352 -35036
rect 12960 -35180 13079 -35061
rect 10850 -35556 10916 -35490
rect 10888 -35650 10954 -35584
rect 10859 -35744 10925 -35678
rect 12549 -36052 12646 -35955
rect 11894 -36299 12136 -36057
rect 13558 -36063 13662 -35959
<< metal2 >>
rect -22627 7080 -22565 7084
rect -22632 7075 -22560 7080
rect -22632 7013 -22627 7075
rect -22565 7030 -22560 7075
rect -22565 7013 -21452 7030
rect -22632 6922 -21452 7013
rect -27531 4452 -27525 4541
rect -27436 4452 -27430 4541
rect -24042 4517 -22832 4545
rect -24042 4445 -24000 4517
rect -22878 4445 -22832 4517
rect -24042 4419 -22832 4445
rect -22632 4490 -22560 6922
rect -21560 6920 -21452 6922
rect -21816 6814 -21727 6820
rect -21560 6812 -17646 6920
rect -21816 6719 -21727 6725
rect -17754 6664 -17646 6812
rect -19307 6655 -19245 6659
rect -19312 6650 -19240 6655
rect -19312 6588 -19307 6650
rect -19245 6588 -19240 6650
rect -19312 6448 -19240 6588
rect -17754 6556 -15130 6664
rect -15022 6556 -15016 6664
rect -18524 6501 -18445 6505
rect -19312 6370 -19240 6376
rect -18528 6496 -18439 6501
rect -18528 6417 -18524 6496
rect -18445 6417 -18439 6496
rect -18528 6368 -18439 6417
rect -16019 6304 -15947 6309
rect -18528 6273 -18439 6279
rect -16023 6242 -16014 6304
rect -15952 6242 -15943 6304
rect -16019 6196 -15947 6242
rect 1795 6241 3005 6269
rect 1795 6169 1841 6241
rect 2963 6169 3005 6241
rect -15226 6155 -15147 6159
rect -16019 6118 -15947 6124
rect -15230 6150 -15141 6155
rect -15230 6071 -15226 6150
rect -15147 6071 -15141 6150
rect 1795 6143 3005 6169
rect 3401 6241 4611 6269
rect 3401 6169 3447 6241
rect 4569 6169 4611 6241
rect 3401 6143 4611 6169
rect 5105 6239 6315 6267
rect 5105 6167 5151 6239
rect 6273 6167 6315 6239
rect 5105 6141 6315 6167
rect -15230 5973 -15141 6071
rect -12737 5978 -12675 5982
rect -15230 5878 -15141 5884
rect -12742 5973 -12670 5978
rect -12742 5911 -12737 5973
rect -12675 5911 -12670 5973
rect -12742 5753 -12670 5911
rect 1559 5925 1679 5932
rect 1559 5813 1565 5925
rect 1674 5924 1679 5925
rect 1674 5815 4873 5924
rect 4970 5815 4976 5924
rect 1674 5813 1679 5815
rect 1559 5807 1679 5813
rect -11940 5784 -11851 5789
rect -11945 5705 -11936 5784
rect -11857 5705 -11848 5784
rect -12742 5675 -12670 5681
rect -11940 5626 -11851 5705
rect -9434 5613 -9372 5617
rect -11940 5531 -11851 5537
rect -9439 5608 -9367 5613
rect -9439 5546 -9434 5608
rect -9372 5546 -9367 5608
rect -9439 5457 -9367 5546
rect 4738 5541 4807 5547
rect -8636 5486 -8557 5490
rect -9439 5379 -9367 5385
rect -8640 5481 -8551 5486
rect -8640 5402 -8636 5481
rect -8557 5402 -8551 5481
rect -8640 5316 -8551 5402
rect 3195 5442 3247 5448
rect 3195 5384 3247 5390
rect -6173 5339 -6084 5346
rect -6173 5269 -6166 5339
rect -6096 5269 -6084 5339
rect -6173 5261 -6084 5269
rect -8640 5221 -8551 5227
rect -5363 5202 -5253 5215
rect -5363 5123 -5353 5202
rect -5268 5123 -5253 5202
rect -5363 5113 -5253 5123
rect -5351 5080 -5262 5113
rect -2870 5028 -2808 5032
rect -5351 4985 -5262 4991
rect -2875 5023 -2803 5028
rect -2875 4961 -2870 5023
rect -2808 4961 -2803 5023
rect -2875 4818 -2803 4961
rect -2054 4881 -1975 4885
rect -2875 4740 -2803 4746
rect -2058 4876 -1969 4881
rect -2058 4797 -2054 4876
rect -1975 4797 -1969 4876
rect -5978 4570 -5803 4576
rect -12549 4562 -12374 4568
rect -22632 4412 -22560 4418
rect -22416 4552 -22230 4558
rect -15826 4556 -15648 4562
rect -20751 4517 -19541 4545
rect -20751 4445 -20709 4517
rect -19587 4445 -19541 4517
rect -20751 4419 -19541 4445
rect -19136 4372 -19130 4553
rect -18949 4372 -18943 4553
rect -17460 4517 -16250 4545
rect -17460 4445 -17418 4517
rect -16296 4445 -16250 4517
rect -17460 4419 -16250 4445
rect -14169 4517 -12959 4545
rect -14169 4445 -14127 4517
rect -13005 4445 -12959 4517
rect -14169 4419 -12959 4445
rect -22416 4237 -22230 4366
rect -19130 4237 -18949 4372
rect -22416 4235 -18933 4237
rect -15826 4235 -15648 4378
rect -10878 4517 -9668 4545
rect -10878 4445 -10836 4517
rect -9714 4445 -9668 4517
rect -10878 4419 -9668 4445
rect -7588 4517 -6378 4545
rect -7588 4445 -7546 4517
rect -6424 4445 -6378 4517
rect -9273 4429 -9081 4436
rect -22416 4233 -15638 4235
rect -12549 4233 -12374 4387
rect -9273 4252 -9267 4429
rect -9092 4252 -9081 4429
rect -7588 4419 -6378 4445
rect -22416 4232 -12373 4233
rect -9273 4232 -9081 4252
rect -2691 4558 -2503 4564
rect -4297 4517 -3087 4545
rect -4297 4445 -4255 4517
rect -3133 4445 -3087 4517
rect -4297 4419 -3087 4445
rect -5978 4232 -5803 4395
rect -2691 4383 -2683 4558
rect -2508 4383 -2503 4558
rect -2058 4562 -1969 4797
rect 2290 4849 2372 4860
rect 2290 4789 2301 4849
rect 2361 4789 2372 4849
rect 2290 4778 2372 4789
rect 430 4726 492 4730
rect 425 4721 497 4726
rect 425 4684 430 4721
rect 492 4684 497 4721
rect 425 4606 497 4612
rect 602 4549 774 4555
rect -2058 4467 -1969 4473
rect -1006 4517 204 4545
rect -1006 4445 -964 4517
rect 158 4445 204 4517
rect -1006 4419 204 4445
rect -2691 4376 -2503 4383
rect -2683 4232 -2508 4376
rect 602 4232 774 4377
rect -22416 4060 602 4232
rect 774 4060 780 4232
rect 1625 4209 2921 4275
rect 2987 4209 2993 4275
rect -22416 4057 -2508 4060
rect -22416 4055 -12373 4057
rect -22416 4054 -15638 4055
rect 602 4054 774 4060
rect -22416 4051 -18933 4054
rect -8666 4009 -8545 4015
rect -25114 3948 -25005 4009
rect -25114 1718 -25005 3839
rect -21823 3987 -21714 4009
rect -18532 3998 -18423 4009
rect -15241 4002 -15132 4009
rect -18538 3887 -18532 3998
rect -18423 3887 -18417 3998
rect -24939 3549 -24166 3587
rect -24939 3409 -24791 3549
rect -24197 3409 -24166 3549
rect -24939 3378 -24166 3409
rect -24939 1961 -24825 3378
rect -23409 3125 -23327 3136
rect -23409 3065 -23398 3125
rect -23338 3065 -23327 3125
rect -23409 3054 -23327 3065
rect -24716 2733 -23506 2761
rect -24716 2661 -24670 2733
rect -23548 2661 -23506 2733
rect -24716 2635 -23506 2661
rect -23157 2733 -21947 2761
rect -23157 2661 -23111 2733
rect -21989 2661 -21947 2733
rect -23157 2635 -21947 2661
rect -24939 1938 -24536 1961
rect -24939 1830 -24915 1938
rect -24825 1830 -24536 1938
rect -24939 1808 -24536 1830
rect -24939 1807 -24825 1808
rect -25114 1717 -24757 1718
rect -25114 1705 -24728 1717
rect -25114 1605 -24818 1705
rect -24840 1597 -24818 1605
rect -24742 1597 -24728 1705
rect -24840 432 -24739 1597
rect -24632 632 -24536 1808
rect -23523 1886 -23251 1902
rect -23523 1789 -23439 1886
rect -23289 1789 -23251 1886
rect -23523 1754 -23251 1789
rect -24221 1341 -24139 1352
rect -24221 1281 -24210 1341
rect -24150 1281 -24139 1341
rect -24221 1270 -24139 1281
rect -23818 1192 -23687 1208
rect -23818 1123 -23802 1192
rect -23703 1123 -23687 1192
rect -24421 1001 -24147 1010
rect -24421 929 -24412 1001
rect -24156 929 -24147 1001
rect -24421 920 -24147 929
rect -24059 666 -23950 681
rect -24633 605 -24469 632
rect -24633 525 -24601 605
rect -24503 525 -24469 605
rect -24633 497 -24469 525
rect -24059 518 -24046 666
rect -23963 518 -23950 666
rect -24059 506 -23950 518
rect -24840 412 -24469 432
rect -24840 346 -24810 412
rect -24557 346 -24469 412
rect -24840 333 -24469 346
rect -24345 259 -23992 268
rect -24345 203 -24336 259
rect -24001 203 -23992 259
rect -24345 194 -23992 203
rect -23818 120 -23687 1123
rect -23523 627 -23427 1754
rect -23304 1698 -23098 1724
rect -23304 1601 -23263 1698
rect -23147 1601 -23098 1698
rect -21823 1718 -21714 3876
rect -21648 3549 -20875 3587
rect -21648 3409 -21500 3549
rect -20906 3409 -20875 3549
rect -21648 3378 -20875 3409
rect -21648 1961 -21534 3378
rect -20118 3125 -20036 3136
rect -20118 3065 -20107 3125
rect -20047 3065 -20036 3125
rect -20118 3054 -20036 3065
rect -21425 2733 -20215 2761
rect -21425 2661 -21379 2733
rect -20257 2661 -20215 2733
rect -21425 2635 -20215 2661
rect -19866 2733 -18656 2761
rect -19866 2661 -19820 2733
rect -18698 2661 -18656 2733
rect -19866 2635 -18656 2661
rect -21648 1938 -21245 1961
rect -21648 1830 -21624 1938
rect -21534 1830 -21245 1938
rect -21648 1808 -21245 1830
rect -21648 1807 -21534 1808
rect -21823 1717 -21466 1718
rect -21823 1705 -21437 1717
rect -21823 1605 -21527 1705
rect -23304 1581 -23098 1601
rect -21549 1597 -21527 1605
rect -21451 1597 -21437 1705
rect -23304 1196 -23209 1581
rect -21823 1407 -21714 1416
rect -22662 1341 -22580 1352
rect -22662 1281 -22651 1341
rect -22591 1281 -22580 1341
rect -22662 1270 -22580 1281
rect -21823 1321 -21814 1407
rect -21723 1321 -21714 1407
rect -23304 1130 -23290 1196
rect -23219 1130 -23209 1196
rect -23524 604 -23360 627
rect -23524 524 -23490 604
rect -23392 524 -23360 604
rect -23524 497 -23360 524
rect -23304 416 -23209 1130
rect -23132 1001 -22858 1010
rect -23132 929 -23123 1001
rect -22867 929 -22858 1001
rect -23132 920 -22858 929
rect -22415 1001 -22141 1010
rect -22415 929 -22406 1001
rect -22150 929 -22141 1001
rect -22415 920 -22141 929
rect -22114 616 -21936 667
rect -22114 536 -22069 616
rect -21949 536 -21936 616
rect -22114 519 -21936 536
rect -23524 401 -23209 416
rect -23524 341 -23500 401
rect -23315 341 -23209 401
rect -22640 450 -22465 461
rect -22640 375 -22628 450
rect -22483 375 -22465 450
rect -22640 363 -22465 375
rect -23524 331 -23209 341
rect -23111 250 -23027 262
rect -23111 188 -23100 250
rect -23038 188 -23027 250
rect -23111 177 -23027 188
rect -22246 225 -22168 236
rect -22246 169 -22235 225
rect -22179 169 -22168 225
rect -22246 158 -22168 169
rect -22114 120 -21994 519
rect -21823 284 -21714 1321
rect -21549 432 -21448 1597
rect -21341 632 -21245 1808
rect -20232 1886 -19960 1902
rect -20232 1789 -20148 1886
rect -19998 1789 -19960 1886
rect -20232 1754 -19960 1789
rect -20930 1341 -20848 1352
rect -20930 1281 -20919 1341
rect -20859 1281 -20848 1341
rect -20930 1270 -20848 1281
rect -20527 1192 -20396 1208
rect -20527 1123 -20511 1192
rect -20412 1123 -20396 1192
rect -21130 1001 -20856 1010
rect -21130 929 -21121 1001
rect -20865 929 -20856 1001
rect -21130 920 -20856 929
rect -20768 666 -20659 681
rect -21342 605 -21178 632
rect -21342 525 -21310 605
rect -21212 525 -21178 605
rect -21342 497 -21178 525
rect -20768 518 -20755 666
rect -20672 518 -20659 666
rect -20768 506 -20659 518
rect -21549 412 -21178 432
rect -21549 346 -21519 412
rect -21266 346 -21178 412
rect -21549 333 -21178 346
rect -21823 218 -21801 284
rect -21735 218 -21714 284
rect -21823 179 -21714 218
rect -21054 259 -20701 268
rect -21054 203 -21045 259
rect -20710 203 -20701 259
rect -21054 194 -20701 203
rect -23818 18 -21994 120
rect -20527 120 -20396 1123
rect -20232 627 -20136 1754
rect -20013 1698 -19807 1724
rect -20013 1601 -19972 1698
rect -19856 1601 -19807 1698
rect -18532 1718 -18423 3887
rect -18357 3549 -17584 3587
rect -18357 3409 -18209 3549
rect -17615 3409 -17584 3549
rect -18357 3378 -17584 3409
rect -18357 1961 -18243 3378
rect -16827 3125 -16745 3136
rect -16827 3065 -16816 3125
rect -16756 3065 -16745 3125
rect -16827 3054 -16745 3065
rect -18134 2733 -16924 2761
rect -18134 2661 -18088 2733
rect -16966 2661 -16924 2733
rect -18134 2635 -16924 2661
rect -16575 2733 -15365 2761
rect -16575 2661 -16529 2733
rect -15407 2661 -15365 2733
rect -16575 2635 -15365 2661
rect -18357 1938 -17954 1961
rect -18357 1830 -18333 1938
rect -18243 1830 -17954 1938
rect -18357 1808 -17954 1830
rect -18357 1807 -18243 1808
rect -18532 1717 -18175 1718
rect -18532 1705 -18146 1717
rect -18532 1605 -18236 1705
rect -20013 1581 -19807 1601
rect -18258 1597 -18236 1605
rect -18160 1597 -18146 1705
rect -20013 1196 -19918 1581
rect -18532 1407 -18423 1416
rect -19371 1341 -19289 1352
rect -19371 1281 -19360 1341
rect -19300 1281 -19289 1341
rect -19371 1270 -19289 1281
rect -18532 1321 -18523 1407
rect -18432 1321 -18423 1407
rect -20013 1130 -19999 1196
rect -19928 1130 -19918 1196
rect -20233 604 -20069 627
rect -20233 524 -20199 604
rect -20101 524 -20069 604
rect -20233 497 -20069 524
rect -20013 416 -19918 1130
rect -19841 1001 -19567 1010
rect -19841 929 -19832 1001
rect -19576 929 -19567 1001
rect -19841 920 -19567 929
rect -19124 1001 -18850 1010
rect -19124 929 -19115 1001
rect -18859 929 -18850 1001
rect -19124 920 -18850 929
rect -18823 616 -18645 667
rect -18823 536 -18778 616
rect -18658 536 -18645 616
rect -18823 519 -18645 536
rect -20233 401 -19918 416
rect -20233 341 -20209 401
rect -20024 341 -19918 401
rect -19349 450 -19174 461
rect -19349 375 -19337 450
rect -19192 375 -19174 450
rect -19349 363 -19174 375
rect -20233 331 -19918 341
rect -19820 250 -19736 262
rect -19820 188 -19809 250
rect -19747 188 -19736 250
rect -19820 177 -19736 188
rect -18955 225 -18877 236
rect -18955 169 -18944 225
rect -18888 169 -18877 225
rect -18955 158 -18877 169
rect -18823 120 -18703 519
rect -18532 283 -18423 1321
rect -18258 432 -18157 1597
rect -18050 632 -17954 1808
rect -16941 1886 -16669 1902
rect -16941 1789 -16857 1886
rect -16707 1789 -16669 1886
rect -16941 1754 -16669 1789
rect -17639 1341 -17557 1352
rect -17639 1281 -17628 1341
rect -17568 1281 -17557 1341
rect -17639 1270 -17557 1281
rect -17236 1192 -17105 1208
rect -17236 1123 -17220 1192
rect -17121 1123 -17105 1192
rect -17839 1001 -17565 1010
rect -17839 929 -17830 1001
rect -17574 929 -17565 1001
rect -17839 920 -17565 929
rect -17477 666 -17368 681
rect -18051 605 -17887 632
rect -18051 525 -18019 605
rect -17921 525 -17887 605
rect -18051 497 -17887 525
rect -17477 518 -17464 666
rect -17381 518 -17368 666
rect -17477 506 -17368 518
rect -18258 412 -17887 432
rect -18258 346 -18228 412
rect -17975 346 -17887 412
rect -18258 333 -17887 346
rect -18532 217 -18505 283
rect -18439 217 -18423 283
rect -18532 179 -18423 217
rect -17763 259 -17410 268
rect -17763 203 -17754 259
rect -17419 203 -17410 259
rect -17763 194 -17410 203
rect -20527 18 -18703 120
rect -17236 120 -17105 1123
rect -16941 627 -16845 1754
rect -16722 1698 -16516 1724
rect -16722 1601 -16681 1698
rect -16565 1601 -16516 1698
rect -15241 1718 -15132 3891
rect -11950 3991 -11841 4009
rect -8666 3900 -8660 4009
rect -8551 3900 -8545 4009
rect -8666 3894 -8545 3900
rect -5375 4009 -5254 4015
rect -5375 3900 -5369 4009
rect -5260 3900 -5254 4009
rect -5375 3894 -5254 3900
rect -2078 3994 -1969 4009
rect -15066 3549 -14293 3587
rect -15066 3409 -14918 3549
rect -14324 3409 -14293 3549
rect -15066 3378 -14293 3409
rect -15066 1961 -14952 3378
rect -13536 3125 -13454 3136
rect -13536 3065 -13525 3125
rect -13465 3065 -13454 3125
rect -13536 3054 -13454 3065
rect -14843 2733 -13633 2761
rect -14843 2661 -14797 2733
rect -13675 2661 -13633 2733
rect -14843 2635 -13633 2661
rect -13284 2733 -12074 2761
rect -13284 2661 -13238 2733
rect -12116 2661 -12074 2733
rect -13284 2635 -12074 2661
rect -15066 1938 -14663 1961
rect -15066 1830 -15042 1938
rect -14952 1830 -14663 1938
rect -15066 1808 -14663 1830
rect -15066 1807 -14952 1808
rect -15241 1717 -14884 1718
rect -15241 1705 -14855 1717
rect -15241 1605 -14945 1705
rect -16722 1581 -16516 1601
rect -14967 1597 -14945 1605
rect -14869 1597 -14855 1705
rect -16722 1196 -16627 1581
rect -15241 1407 -15132 1416
rect -16080 1341 -15998 1352
rect -16080 1281 -16069 1341
rect -16009 1281 -15998 1341
rect -16080 1270 -15998 1281
rect -15241 1321 -15232 1407
rect -15141 1321 -15132 1407
rect -16722 1130 -16708 1196
rect -16637 1130 -16627 1196
rect -16942 604 -16778 627
rect -16942 524 -16908 604
rect -16810 524 -16778 604
rect -16942 497 -16778 524
rect -16722 416 -16627 1130
rect -16550 1001 -16276 1010
rect -16550 929 -16541 1001
rect -16285 929 -16276 1001
rect -16550 920 -16276 929
rect -15833 1001 -15559 1010
rect -15833 929 -15824 1001
rect -15568 929 -15559 1001
rect -15833 920 -15559 929
rect -15532 616 -15354 667
rect -15532 536 -15487 616
rect -15367 536 -15354 616
rect -15532 519 -15354 536
rect -16942 401 -16627 416
rect -16942 341 -16918 401
rect -16733 341 -16627 401
rect -16058 450 -15883 461
rect -16058 375 -16046 450
rect -15901 375 -15883 450
rect -16058 363 -15883 375
rect -16942 331 -16627 341
rect -16529 250 -16445 262
rect -16529 188 -16518 250
rect -16456 188 -16445 250
rect -16529 177 -16445 188
rect -15664 225 -15586 236
rect -15664 169 -15653 225
rect -15597 169 -15586 225
rect -15664 158 -15586 169
rect -15532 120 -15412 519
rect -15241 296 -15132 1321
rect -14967 432 -14866 1597
rect -14759 632 -14663 1808
rect -13650 1886 -13378 1902
rect -13650 1789 -13566 1886
rect -13416 1789 -13378 1886
rect -13650 1754 -13378 1789
rect -14348 1341 -14266 1352
rect -14348 1281 -14337 1341
rect -14277 1281 -14266 1341
rect -14348 1270 -14266 1281
rect -13945 1192 -13814 1208
rect -13945 1123 -13929 1192
rect -13830 1123 -13814 1192
rect -14548 1001 -14274 1010
rect -14548 929 -14539 1001
rect -14283 929 -14274 1001
rect -14548 920 -14274 929
rect -14186 666 -14077 681
rect -14760 605 -14596 632
rect -14760 525 -14728 605
rect -14630 525 -14596 605
rect -14760 497 -14596 525
rect -14186 518 -14173 666
rect -14090 518 -14077 666
rect -14186 506 -14077 518
rect -14967 412 -14596 432
rect -14967 346 -14937 412
rect -14684 346 -14596 412
rect -14967 333 -14596 346
rect -15241 230 -15223 296
rect -15157 230 -15132 296
rect -15241 179 -15132 230
rect -14472 259 -14119 268
rect -14472 203 -14463 259
rect -14128 203 -14119 259
rect -14472 194 -14119 203
rect -17236 18 -15412 120
rect -13945 120 -13814 1123
rect -13650 627 -13554 1754
rect -13431 1698 -13225 1724
rect -13431 1601 -13390 1698
rect -13274 1601 -13225 1698
rect -11950 1718 -11841 3880
rect -11775 3549 -11002 3587
rect -11775 3409 -11627 3549
rect -11033 3409 -11002 3549
rect -11775 3378 -11002 3409
rect -11775 1961 -11661 3378
rect -10245 3125 -10163 3136
rect -10245 3065 -10234 3125
rect -10174 3065 -10163 3125
rect -10245 3054 -10163 3065
rect -11552 2733 -10342 2761
rect -11552 2661 -11506 2733
rect -10384 2661 -10342 2733
rect -11552 2635 -10342 2661
rect -9993 2733 -8783 2761
rect -9993 2661 -9947 2733
rect -8825 2661 -8783 2733
rect -9993 2635 -8783 2661
rect -11775 1938 -11372 1961
rect -11775 1830 -11751 1938
rect -11661 1830 -11372 1938
rect -11775 1808 -11372 1830
rect -11775 1807 -11661 1808
rect -11950 1717 -11593 1718
rect -11950 1705 -11564 1717
rect -11950 1605 -11654 1705
rect -13431 1581 -13225 1601
rect -11676 1597 -11654 1605
rect -11578 1597 -11564 1705
rect -13431 1196 -13336 1581
rect -11950 1407 -11841 1416
rect -12789 1341 -12707 1352
rect -12789 1281 -12778 1341
rect -12718 1281 -12707 1341
rect -12789 1270 -12707 1281
rect -11950 1321 -11941 1407
rect -11850 1321 -11841 1407
rect -13431 1130 -13417 1196
rect -13346 1130 -13336 1196
rect -13651 604 -13487 627
rect -13651 524 -13617 604
rect -13519 524 -13487 604
rect -13651 497 -13487 524
rect -13431 416 -13336 1130
rect -13259 1001 -12985 1010
rect -13259 929 -13250 1001
rect -12994 929 -12985 1001
rect -13259 920 -12985 929
rect -12542 1001 -12268 1010
rect -12542 929 -12533 1001
rect -12277 929 -12268 1001
rect -12542 920 -12268 929
rect -12241 616 -12063 667
rect -12241 536 -12196 616
rect -12076 536 -12063 616
rect -12241 519 -12063 536
rect -13651 401 -13336 416
rect -13651 341 -13627 401
rect -13442 341 -13336 401
rect -12767 450 -12592 461
rect -12767 375 -12755 450
rect -12610 375 -12592 450
rect -12767 363 -12592 375
rect -13651 331 -13336 341
rect -13238 250 -13154 262
rect -13238 188 -13227 250
rect -13165 188 -13154 250
rect -13238 177 -13154 188
rect -12373 225 -12295 236
rect -12373 169 -12362 225
rect -12306 169 -12295 225
rect -12373 158 -12295 169
rect -12241 120 -12121 519
rect -11950 295 -11841 1321
rect -11676 432 -11575 1597
rect -11468 632 -11372 1808
rect -10359 1886 -10087 1902
rect -10359 1789 -10275 1886
rect -10125 1789 -10087 1886
rect -10359 1754 -10087 1789
rect -11057 1341 -10975 1352
rect -11057 1281 -11046 1341
rect -10986 1281 -10975 1341
rect -11057 1270 -10975 1281
rect -10654 1192 -10523 1208
rect -10654 1123 -10638 1192
rect -10539 1123 -10523 1192
rect -11257 1001 -10983 1010
rect -11257 929 -11248 1001
rect -10992 929 -10983 1001
rect -11257 920 -10983 929
rect -10895 666 -10786 681
rect -11469 605 -11305 632
rect -11469 525 -11437 605
rect -11339 525 -11305 605
rect -11469 497 -11305 525
rect -10895 518 -10882 666
rect -10799 518 -10786 666
rect -10895 506 -10786 518
rect -11676 412 -11305 432
rect -11676 346 -11646 412
rect -11393 346 -11305 412
rect -11676 333 -11305 346
rect -11963 289 -11841 295
rect -11897 223 -11841 289
rect -11963 217 -11841 223
rect -11950 179 -11841 217
rect -11181 259 -10828 268
rect -11181 203 -11172 259
rect -10837 203 -10828 259
rect -11181 194 -10828 203
rect -13945 18 -12121 120
rect -10654 120 -10523 1123
rect -10359 627 -10263 1754
rect -10140 1698 -9934 1724
rect -10140 1601 -10099 1698
rect -9983 1601 -9934 1698
rect -8660 1718 -8551 3894
rect -8485 3549 -7712 3587
rect -8485 3409 -8337 3549
rect -7743 3409 -7712 3549
rect -8485 3378 -7712 3409
rect -8485 1961 -8371 3378
rect -6955 3125 -6873 3136
rect -6955 3065 -6944 3125
rect -6884 3065 -6873 3125
rect -6955 3054 -6873 3065
rect -8262 2733 -7052 2761
rect -8262 2661 -8216 2733
rect -7094 2661 -7052 2733
rect -8262 2635 -7052 2661
rect -6703 2733 -5493 2761
rect -6703 2661 -6657 2733
rect -5535 2661 -5493 2733
rect -6703 2635 -5493 2661
rect -8485 1938 -8082 1961
rect -8485 1830 -8461 1938
rect -8371 1830 -8082 1938
rect -8485 1808 -8082 1830
rect -8485 1807 -8371 1808
rect -8660 1717 -8303 1718
rect -8660 1705 -8274 1717
rect -8660 1605 -8364 1705
rect -10140 1581 -9934 1601
rect -8386 1597 -8364 1605
rect -8288 1597 -8274 1705
rect -10140 1196 -10045 1581
rect -8659 1407 -8550 1416
rect -9498 1341 -9416 1352
rect -9498 1281 -9487 1341
rect -9427 1281 -9416 1341
rect -9498 1270 -9416 1281
rect -8659 1321 -8650 1407
rect -8559 1321 -8550 1407
rect -10140 1130 -10126 1196
rect -10055 1130 -10045 1196
rect -10360 604 -10196 627
rect -10360 524 -10326 604
rect -10228 524 -10196 604
rect -10360 497 -10196 524
rect -10140 416 -10045 1130
rect -9968 1001 -9694 1010
rect -9968 929 -9959 1001
rect -9703 929 -9694 1001
rect -9968 920 -9694 929
rect -9251 1001 -8977 1010
rect -9251 929 -9242 1001
rect -8986 929 -8977 1001
rect -9251 920 -8977 929
rect -8950 616 -8772 667
rect -8950 536 -8905 616
rect -8785 536 -8772 616
rect -8950 519 -8772 536
rect -10360 401 -10045 416
rect -10360 341 -10336 401
rect -10151 341 -10045 401
rect -9476 450 -9301 461
rect -9476 375 -9464 450
rect -9319 375 -9301 450
rect -9476 363 -9301 375
rect -10360 331 -10045 341
rect -9947 250 -9863 262
rect -9947 188 -9936 250
rect -9874 188 -9863 250
rect -9947 177 -9863 188
rect -9082 225 -9004 236
rect -9082 169 -9071 225
rect -9015 169 -9004 225
rect -9082 158 -9004 169
rect -8950 120 -8830 519
rect -8659 309 -8550 1321
rect -8386 432 -8285 1597
rect -8178 632 -8082 1808
rect -7069 1886 -6797 1902
rect -7069 1789 -6985 1886
rect -6835 1789 -6797 1886
rect -7069 1754 -6797 1789
rect -7767 1341 -7685 1352
rect -7767 1281 -7756 1341
rect -7696 1281 -7685 1341
rect -7767 1270 -7685 1281
rect -7364 1192 -7233 1208
rect -7364 1123 -7348 1192
rect -7249 1123 -7233 1192
rect -7967 1001 -7693 1010
rect -7967 929 -7958 1001
rect -7702 929 -7693 1001
rect -7967 920 -7693 929
rect -7605 666 -7496 681
rect -8179 605 -8015 632
rect -8179 525 -8147 605
rect -8049 525 -8015 605
rect -8179 497 -8015 525
rect -7605 518 -7592 666
rect -7509 518 -7496 666
rect -7605 506 -7496 518
rect -8386 412 -8015 432
rect -8386 346 -8356 412
rect -8103 346 -8015 412
rect -8386 333 -8015 346
rect -8659 243 -8633 309
rect -8567 243 -8550 309
rect -8659 179 -8550 243
rect -7891 259 -7538 268
rect -7891 203 -7882 259
rect -7547 203 -7538 259
rect -7891 194 -7538 203
rect -10654 18 -8830 120
rect -7364 120 -7233 1123
rect -7069 627 -6973 1754
rect -6850 1698 -6644 1724
rect -6850 1601 -6809 1698
rect -6693 1601 -6644 1698
rect -5369 1718 -5260 3894
rect -5194 3549 -4421 3587
rect -5194 3409 -5046 3549
rect -4452 3409 -4421 3549
rect -5194 3378 -4421 3409
rect -5194 1961 -5080 3378
rect -3664 3125 -3582 3136
rect -3664 3065 -3653 3125
rect -3593 3065 -3582 3125
rect -3664 3054 -3582 3065
rect -4971 2733 -3761 2761
rect -4971 2661 -4925 2733
rect -3803 2661 -3761 2733
rect -4971 2635 -3761 2661
rect -3412 2733 -2202 2761
rect -3412 2661 -3366 2733
rect -2244 2661 -2202 2733
rect -3412 2635 -2202 2661
rect -5194 1938 -4791 1961
rect -5194 1830 -5170 1938
rect -5080 1830 -4791 1938
rect -5194 1808 -4791 1830
rect -5194 1807 -5080 1808
rect -5369 1717 -5012 1718
rect -5369 1705 -4983 1717
rect -5369 1605 -5073 1705
rect -6850 1581 -6644 1601
rect -5095 1597 -5073 1605
rect -4997 1597 -4983 1705
rect -6850 1196 -6755 1581
rect -5369 1407 -5260 1416
rect -6208 1341 -6126 1352
rect -6208 1281 -6197 1341
rect -6137 1281 -6126 1341
rect -6208 1270 -6126 1281
rect -5369 1321 -5360 1407
rect -5269 1321 -5260 1407
rect -6850 1130 -6836 1196
rect -6765 1130 -6755 1196
rect -7070 604 -6906 627
rect -7070 524 -7036 604
rect -6938 524 -6906 604
rect -7070 497 -6906 524
rect -6850 416 -6755 1130
rect -6678 1001 -6404 1010
rect -6678 929 -6669 1001
rect -6413 929 -6404 1001
rect -6678 920 -6404 929
rect -5961 1001 -5687 1010
rect -5961 929 -5952 1001
rect -5696 929 -5687 1001
rect -5961 920 -5687 929
rect -5660 616 -5482 667
rect -5660 536 -5615 616
rect -5495 536 -5482 616
rect -5660 519 -5482 536
rect -7070 401 -6755 416
rect -7070 341 -7046 401
rect -6861 341 -6755 401
rect -6186 450 -6011 461
rect -6186 375 -6174 450
rect -6029 375 -6011 450
rect -6186 363 -6011 375
rect -7070 331 -6755 341
rect -6657 250 -6573 262
rect -6657 188 -6646 250
rect -6584 188 -6573 250
rect -6657 177 -6573 188
rect -5792 225 -5714 236
rect -5792 169 -5781 225
rect -5725 169 -5714 225
rect -5792 158 -5714 169
rect -5660 120 -5540 519
rect -5369 292 -5260 1321
rect -5095 432 -4994 1597
rect -4887 632 -4791 1808
rect -3778 1886 -3506 1902
rect -3778 1789 -3694 1886
rect -3544 1789 -3506 1886
rect -3778 1754 -3506 1789
rect -4476 1341 -4394 1352
rect -4476 1281 -4465 1341
rect -4405 1281 -4394 1341
rect -4476 1270 -4394 1281
rect -4073 1192 -3942 1208
rect -4073 1123 -4057 1192
rect -3958 1123 -3942 1192
rect -4676 1001 -4402 1010
rect -4676 929 -4667 1001
rect -4411 929 -4402 1001
rect -4676 920 -4402 929
rect -4314 666 -4205 681
rect -4888 605 -4724 632
rect -4888 525 -4856 605
rect -4758 525 -4724 605
rect -4888 497 -4724 525
rect -4314 518 -4301 666
rect -4218 518 -4205 666
rect -4314 506 -4205 518
rect -5095 412 -4724 432
rect -5095 346 -5065 412
rect -4812 346 -4724 412
rect -5095 333 -4724 346
rect -5369 226 -5349 292
rect -5283 226 -5260 292
rect -5369 179 -5260 226
rect -4600 259 -4247 268
rect -4600 203 -4591 259
rect -4256 203 -4247 259
rect -4600 194 -4247 203
rect -7364 18 -5540 120
rect -4073 120 -3942 1123
rect -3778 627 -3682 1754
rect -3559 1698 -3353 1724
rect -3559 1601 -3518 1698
rect -3402 1601 -3353 1698
rect -2078 1718 -1969 3883
rect -1903 3549 -1130 3587
rect -1903 3409 -1755 3549
rect -1161 3409 -1130 3549
rect -1903 3378 -1130 3409
rect -1903 1961 -1789 3378
rect -373 3125 -291 3136
rect -373 3065 -362 3125
rect -302 3065 -291 3125
rect -373 3054 -291 3065
rect -1680 2733 -470 2761
rect -1680 2661 -1634 2733
rect -512 2661 -470 2733
rect -1680 2635 -470 2661
rect -121 2733 1089 2761
rect -121 2661 -75 2733
rect 1047 2661 1089 2733
rect -121 2635 1089 2661
rect -1903 1938 -1500 1961
rect -1903 1830 -1879 1938
rect -1789 1830 -1500 1938
rect -1903 1808 -1500 1830
rect -1903 1807 -1789 1808
rect -2078 1717 -1721 1718
rect -2078 1705 -1692 1717
rect -2078 1605 -1782 1705
rect -3559 1581 -3353 1601
rect -1804 1597 -1782 1605
rect -1706 1597 -1692 1705
rect -3559 1196 -3464 1581
rect -2078 1407 -1969 1416
rect -2917 1341 -2835 1352
rect -2917 1281 -2906 1341
rect -2846 1281 -2835 1341
rect -2917 1270 -2835 1281
rect -2078 1321 -2069 1407
rect -1978 1321 -1969 1407
rect -3559 1130 -3545 1196
rect -3474 1130 -3464 1196
rect -3779 604 -3615 627
rect -3779 524 -3745 604
rect -3647 524 -3615 604
rect -3779 497 -3615 524
rect -3559 416 -3464 1130
rect -3387 1001 -3113 1010
rect -3387 929 -3378 1001
rect -3122 929 -3113 1001
rect -3387 920 -3113 929
rect -2670 1001 -2396 1010
rect -2670 929 -2661 1001
rect -2405 929 -2396 1001
rect -2670 920 -2396 929
rect -2369 616 -2191 667
rect -2369 536 -2324 616
rect -2204 536 -2191 616
rect -2369 519 -2191 536
rect -3779 401 -3464 416
rect -3779 341 -3755 401
rect -3570 341 -3464 401
rect -2895 450 -2720 461
rect -2895 375 -2883 450
rect -2738 375 -2720 450
rect -2895 363 -2720 375
rect -3779 331 -3464 341
rect -3366 250 -3282 262
rect -3366 188 -3355 250
rect -3293 188 -3282 250
rect -3366 177 -3282 188
rect -2501 225 -2423 236
rect -2501 169 -2490 225
rect -2434 169 -2423 225
rect -2501 158 -2423 169
rect -2369 120 -2249 519
rect -2078 261 -1969 1321
rect -1804 432 -1703 1597
rect -1596 632 -1500 1808
rect -487 1886 -215 1902
rect -487 1789 -403 1886
rect -253 1789 -215 1886
rect -487 1754 -215 1789
rect -1185 1341 -1103 1352
rect -1185 1281 -1174 1341
rect -1114 1281 -1103 1341
rect -1185 1270 -1103 1281
rect -782 1192 -651 1208
rect -782 1123 -766 1192
rect -667 1123 -651 1192
rect -1385 1001 -1111 1010
rect -1385 929 -1376 1001
rect -1120 929 -1111 1001
rect -1385 920 -1111 929
rect -1023 666 -914 681
rect -1597 605 -1433 632
rect -1597 525 -1565 605
rect -1467 525 -1433 605
rect -1597 497 -1433 525
rect -1023 518 -1010 666
rect -927 518 -914 666
rect -1023 506 -914 518
rect -1804 412 -1433 432
rect -1804 346 -1774 412
rect -1521 346 -1433 412
rect -1804 333 -1433 346
rect -2078 195 -2061 261
rect -1995 195 -1969 261
rect -2078 179 -1969 195
rect -1309 259 -956 268
rect -1309 203 -1300 259
rect -965 203 -956 259
rect -1309 194 -956 203
rect -4073 18 -2249 120
rect -782 120 -651 1123
rect -487 627 -391 1754
rect -268 1698 -62 1724
rect -268 1601 -227 1698
rect -111 1601 -62 1698
rect -268 1581 -62 1601
rect -268 1196 -173 1581
rect 1213 1407 1322 1416
rect 374 1341 456 1352
rect 374 1281 385 1341
rect 445 1281 456 1341
rect 374 1270 456 1281
rect 1213 1321 1222 1407
rect 1313 1321 1322 1407
rect -268 1130 -254 1196
rect -183 1130 -173 1196
rect -488 604 -324 627
rect -488 524 -454 604
rect -356 524 -324 604
rect -488 497 -324 524
rect -268 416 -173 1130
rect -96 1001 178 1010
rect -96 929 -87 1001
rect 169 929 178 1001
rect -96 920 178 929
rect 621 1001 895 1010
rect 621 929 630 1001
rect 886 929 895 1001
rect 621 920 895 929
rect 922 616 1100 667
rect 922 536 967 616
rect 1087 536 1100 616
rect 922 519 1100 536
rect -488 401 -173 416
rect -488 341 -464 401
rect -279 341 -173 401
rect 396 450 571 461
rect 396 375 408 450
rect 553 375 571 450
rect 396 363 571 375
rect -488 331 -173 341
rect -75 250 9 262
rect -75 188 -64 250
rect -2 188 9 250
rect -75 177 9 188
rect 790 225 868 236
rect 790 169 801 225
rect 857 169 868 225
rect 790 158 868 169
rect 922 120 1042 519
rect 1213 179 1322 1321
rect -782 18 1042 120
rect -25060 -123 -24969 -117
rect 242 -123 248 -40
rect -24969 -131 248 -123
rect 339 -131 345 -40
rect -24969 -214 339 -131
rect -25060 -220 -24969 -214
rect -24635 -2113 -18960 -1976
rect 1225 -2009 1291 179
rect 1625 -1298 1691 4209
rect 3198 4128 3243 5384
rect 4738 5193 4807 5472
rect 4959 5230 5028 5236
rect 4738 5124 4959 5193
rect 4885 5087 4959 5124
rect 4885 5081 5028 5087
rect 4885 5060 4978 5081
rect 3896 4849 3978 4860
rect 3896 4789 3907 4849
rect 3967 4789 3978 4849
rect 3896 4778 3978 4789
rect 4885 4275 4951 5060
rect 5583 4847 5692 4879
rect 5583 4787 5611 4847
rect 5671 4802 5692 4847
rect 7313 4802 7444 4812
rect 5671 4787 7323 4802
rect 5583 4693 7323 4787
rect 7433 4693 7810 4802
rect 7919 4693 7925 4802
rect 7313 4683 7444 4693
rect 4879 4209 4885 4275
rect 4951 4209 4957 4275
rect 3198 4083 5411 4128
rect 5558 4099 5627 4128
rect 5333 4011 5339 4083
rect 5411 4011 5417 4083
rect 5339 3863 5411 4011
rect 5558 3879 5627 4029
rect 5998 4099 6067 4128
rect 6438 4081 6507 4128
rect 5998 3879 6067 4029
rect 6436 4022 6445 4081
rect 6504 4022 6513 4081
rect 6438 3879 6507 4022
rect 5552 3810 5558 3879
rect 5627 3810 5633 3879
rect 5992 3810 5998 3879
rect 6067 3810 6073 3879
rect 6432 3810 6438 3879
rect 6507 3810 6513 3879
rect 5901 3425 7113 3494
rect 5901 3314 5970 3425
rect 5703 3230 5823 3258
rect 5901 3239 5970 3245
rect 6158 3249 6236 3259
rect 5703 3174 5732 3230
rect 5788 3174 5823 3230
rect 6158 3193 6170 3249
rect 6226 3193 6236 3249
rect 6335 3243 6341 3312
rect 6410 3243 6416 3312
rect 6580 3258 6700 3274
rect 6158 3178 6236 3193
rect 5703 3145 5823 3174
rect 6341 3033 6410 3243
rect 6580 3202 6610 3258
rect 6666 3202 6700 3258
rect 6580 3161 6700 3202
rect 6299 2974 6410 3033
rect 6299 2875 6367 2974
rect 6295 2817 6304 2875
rect 6362 2817 6371 2875
rect 7044 2870 7113 3425
rect 7044 2861 10140 2870
rect 6299 2812 6367 2817
rect 7044 2809 7106 2861
rect 7158 2860 9002 2861
rect 7158 2809 8069 2860
rect 7044 2808 8069 2809
rect 8122 2809 9002 2860
rect 9055 2809 9933 2861
rect 9986 2809 10140 2861
rect 8122 2808 10140 2809
rect 7044 2801 10140 2808
rect 12187 2869 12431 2880
rect 12187 2861 12198 2869
rect 5992 2775 6073 2781
rect 5992 2706 5998 2775
rect 6067 2770 6073 2775
rect 6067 2768 8115 2770
rect 6067 2767 8057 2768
rect 6067 2715 7113 2767
rect 7165 2716 8057 2767
rect 8109 2716 8115 2768
rect 7165 2715 8115 2716
rect 6067 2711 8115 2715
rect 8182 2720 8914 2773
rect 9929 2767 10000 2769
rect 6067 2706 6073 2711
rect 5992 2700 6073 2706
rect 7321 2678 7393 2683
rect 8182 2678 8248 2720
rect 6429 2640 6516 2649
rect 6429 2571 6438 2640
rect 6507 2571 6516 2640
rect 7321 2612 7327 2678
rect 7393 2612 8248 2678
rect 8424 2685 8493 2691
rect 8861 2672 8914 2720
rect 8989 2709 8998 2765
rect 9054 2709 9063 2765
rect 9923 2711 9935 2767
rect 9991 2711 10000 2767
rect 10256 2716 10336 2722
rect 9929 2705 9993 2711
rect 8541 2640 8600 2644
rect 8493 2635 8605 2640
rect 8493 2633 8541 2635
rect 7321 2606 7393 2612
rect 8424 2576 8541 2633
rect 8600 2576 8605 2635
rect 8861 2619 8989 2672
rect 9042 2619 9048 2672
rect 10256 2647 10262 2716
rect 10331 2647 10336 2716
rect 10256 2640 10336 2647
rect 10405 2706 10860 2772
rect 10926 2706 10932 2772
rect 8424 2571 8605 2576
rect 6429 2562 6516 2571
rect 8541 2567 8600 2571
rect 10405 2562 10471 2706
rect 1934 2519 2000 2525
rect 2000 2453 8986 2519
rect 9052 2453 9058 2519
rect 9792 2496 9798 2562
rect 9864 2496 10471 2562
rect 10536 2612 10858 2678
rect 10924 2612 10930 2678
rect 12187 2658 12189 2861
rect 12187 2647 12198 2658
rect 12420 2647 12441 2869
rect 12187 2636 12431 2647
rect 1934 2447 2000 2453
rect 5732 2357 9917 2423
rect 9983 2357 9989 2423
rect 6576 2317 6642 2357
rect 5732 2251 7106 2317
rect 7172 2251 7178 2317
rect 10536 2314 10602 2612
rect 6576 2215 6642 2251
rect 8812 2248 8818 2314
rect 8884 2248 10602 2314
rect 10659 2518 10850 2584
rect 10915 2518 10921 2584
rect 6576 2213 6683 2215
rect 5732 2147 6966 2213
rect 7032 2147 8050 2213
rect 8116 2147 8122 2213
rect 6617 1111 6683 2147
rect 10659 2060 10725 2518
rect 7866 1994 7872 2060
rect 7938 1994 10725 2060
rect 7156 1715 11207 1787
rect 7156 1537 7227 1715
rect 7405 1537 8162 1715
rect 8340 1537 9098 1715
rect 9276 1538 10029 1715
rect 10206 1538 10956 1715
rect 9276 1537 10956 1538
rect 11134 1537 11207 1715
rect 7156 1466 11207 1537
rect 12414 1296 12821 1408
rect 12128 1292 12821 1296
rect 7847 1201 7853 1267
rect 7919 1201 10121 1267
rect 5732 1045 6953 1111
rect 7019 1045 8989 1111
rect 9055 1045 9061 1111
rect 6617 989 6683 1045
rect 10055 989 10121 1201
rect 12128 1266 13042 1292
rect 12128 1204 13186 1266
rect 12128 1085 12233 1204
rect 12352 1163 13186 1204
rect 12352 1085 12960 1163
rect 12128 1044 12960 1085
rect 13079 1044 13186 1163
rect 5732 923 9917 989
rect 9983 923 9989 989
rect 10055 923 10704 989
rect 12128 979 13186 1044
rect 3886 825 7102 891
rect 7168 825 7174 891
rect 1618 -1309 1704 -1298
rect 1618 -1375 1625 -1309
rect 1691 -1375 1704 -1309
rect 1618 -1380 1704 -1375
rect 3886 -1551 3970 825
rect 8831 791 8837 857
rect 8903 791 10588 857
rect 4166 733 8050 770
rect 4164 704 8050 733
rect 8116 704 8122 770
rect 3880 -1635 3886 -1551
rect 3970 -1635 3976 -1551
rect 4164 -1602 4248 704
rect 9801 699 9807 763
rect 9873 699 10453 763
rect 8396 668 8470 674
rect 6780 649 6849 655
rect 6849 596 8206 635
rect 8396 633 8405 668
rect 8461 633 8470 668
rect 8396 604 8401 633
rect 6780 574 6849 580
rect 6066 546 6132 552
rect 6132 537 8139 546
rect 6132 485 8079 537
rect 8131 485 8139 537
rect 8167 527 8206 596
rect 8465 604 8470 633
rect 8615 574 8993 640
rect 9059 574 9065 640
rect 10264 633 10324 639
rect 10257 575 10264 631
rect 10324 575 10331 631
rect 8401 563 8465 569
rect 8616 527 8655 574
rect 10264 567 10324 573
rect 8167 488 8655 527
rect 6132 480 8139 485
rect 8992 480 9001 546
rect 9067 480 9076 546
rect 9931 481 9937 547
rect 10003 481 10012 547
rect 10387 546 10453 699
rect 10522 640 10588 791
rect 10638 734 10704 923
rect 12467 820 13186 979
rect 12796 787 13186 820
rect 10638 668 10850 734
rect 10916 668 10922 734
rect 10522 574 10888 640
rect 10954 574 10963 640
rect 10387 480 10859 546
rect 10925 480 10931 546
rect 6066 474 6132 480
rect 6934 386 6941 452
rect 7007 443 10062 452
rect 7007 391 8063 443
rect 8128 391 8992 443
rect 9057 391 9951 443
rect 10016 391 10062 443
rect 7007 386 10062 391
rect 6941 380 7007 386
rect 11883 167 12147 178
rect 11883 -75 11894 167
rect 12136 -75 12147 167
rect 11883 -86 12147 -75
rect 5558 -450 5627 -400
rect 5998 -424 6067 -400
rect 5554 -509 5563 -450
rect 5622 -509 5631 -450
rect 5994 -483 6003 -424
rect 6062 -483 6071 -424
rect 6438 -455 6507 -400
rect 5558 -649 5627 -509
rect 5998 -649 6067 -483
rect 6434 -514 6443 -455
rect 6502 -514 6511 -455
rect 6438 -649 6507 -514
rect 5552 -718 5558 -649
rect 5627 -718 5633 -649
rect 5992 -718 5998 -649
rect 6067 -718 6073 -649
rect 6432 -718 6438 -649
rect 6507 -718 6513 -649
rect 5901 -1103 7113 -1034
rect 5901 -1214 5970 -1103
rect 5703 -1298 5823 -1270
rect 5901 -1289 5970 -1283
rect 6158 -1279 6236 -1269
rect 5703 -1354 5732 -1298
rect 5788 -1354 5823 -1298
rect 6158 -1335 6170 -1279
rect 6226 -1335 6236 -1279
rect 6335 -1285 6341 -1216
rect 6410 -1285 6416 -1216
rect 6580 -1270 6700 -1254
rect 6158 -1350 6236 -1335
rect 5703 -1383 5823 -1354
rect 6341 -1495 6410 -1285
rect 6580 -1326 6610 -1270
rect 6666 -1326 6700 -1270
rect 6580 -1367 6700 -1326
rect 6299 -1554 6410 -1495
rect 4158 -1686 4164 -1602
rect 4248 -1686 4254 -1602
rect 6299 -1653 6367 -1554
rect 6295 -1711 6304 -1653
rect 6362 -1711 6371 -1653
rect 7044 -1658 7113 -1103
rect 7044 -1667 10140 -1658
rect 6299 -1716 6367 -1711
rect 7044 -1719 7106 -1667
rect 7158 -1668 9002 -1667
rect 7158 -1719 8069 -1668
rect 7044 -1720 8069 -1719
rect 8122 -1719 9002 -1668
rect 9055 -1719 9933 -1667
rect 9986 -1719 10140 -1667
rect 8122 -1720 10140 -1719
rect 7044 -1727 10140 -1720
rect 12187 -1659 12431 -1648
rect 12187 -1667 12198 -1659
rect 5992 -1753 6073 -1747
rect 5992 -1822 5998 -1753
rect 6067 -1758 6073 -1753
rect 6067 -1760 8115 -1758
rect 6067 -1761 8057 -1760
rect 6067 -1813 7113 -1761
rect 7165 -1812 8057 -1761
rect 8109 -1812 8115 -1760
rect 7165 -1813 8115 -1812
rect 6067 -1817 8115 -1813
rect 8182 -1808 8914 -1755
rect 9929 -1761 10000 -1759
rect 6067 -1822 6073 -1817
rect 5992 -1828 6073 -1822
rect 7321 -1850 7393 -1845
rect 8182 -1850 8248 -1808
rect 6429 -1888 6516 -1879
rect 6429 -1957 6438 -1888
rect 6507 -1957 6516 -1888
rect 7321 -1916 7327 -1850
rect 7393 -1916 8248 -1850
rect 8424 -1843 8493 -1837
rect 8861 -1856 8914 -1808
rect 8989 -1819 8998 -1763
rect 9054 -1819 9063 -1763
rect 9923 -1817 9935 -1761
rect 9991 -1817 10000 -1761
rect 10256 -1812 10336 -1806
rect 9929 -1823 9993 -1817
rect 8541 -1888 8600 -1884
rect 8493 -1893 8605 -1888
rect 8493 -1895 8541 -1893
rect 7321 -1922 7393 -1916
rect 8424 -1952 8541 -1895
rect 8600 -1952 8605 -1893
rect 8861 -1909 8989 -1856
rect 9042 -1909 9048 -1856
rect 10256 -1881 10262 -1812
rect 10331 -1881 10336 -1812
rect 10256 -1888 10336 -1881
rect 10405 -1822 10860 -1756
rect 10926 -1822 10932 -1756
rect 8424 -1957 8605 -1952
rect 6429 -1966 6516 -1957
rect 8541 -1961 8600 -1957
rect 10405 -1966 10471 -1822
rect 1225 -2075 8986 -2009
rect 9052 -2075 9058 -2009
rect 9792 -2032 9798 -1966
rect 9864 -2032 10471 -1966
rect 10536 -1916 10858 -1850
rect 10924 -1916 10930 -1850
rect 12187 -1870 12189 -1667
rect 12187 -1881 12198 -1870
rect 12420 -1881 12441 -1659
rect 12187 -1892 12431 -1881
rect -25216 -2524 -25155 -2520
rect -24635 -2524 -24492 -2113
rect -23628 -2225 -23414 -2203
rect -24448 -2327 -23814 -2293
rect -23628 -2304 -23605 -2225
rect -23436 -2304 -23414 -2225
rect -23628 -2323 -23414 -2304
rect -24448 -2467 -24410 -2327
rect -23856 -2467 -23814 -2327
rect -24448 -2506 -23814 -2467
rect -25220 -2529 -24492 -2524
rect -25220 -2591 -25216 -2529
rect -25155 -2591 -24492 -2529
rect -25220 -2595 -24492 -2591
rect -25216 -2600 -25155 -2595
rect -24635 -2648 -24492 -2595
rect -22793 -2655 -22650 -2113
rect -21608 -2225 -21394 -2203
rect -22411 -2327 -21777 -2293
rect -21608 -2304 -21585 -2225
rect -21416 -2304 -21394 -2225
rect -21608 -2323 -21394 -2304
rect -22411 -2467 -22373 -2327
rect -21819 -2467 -21777 -2327
rect -22411 -2506 -21777 -2467
rect -20952 -2652 -20809 -2113
rect -19867 -2225 -19653 -2203
rect -20681 -2327 -20047 -2293
rect -19867 -2304 -19844 -2225
rect -19675 -2304 -19653 -2225
rect -19867 -2323 -19653 -2304
rect -20681 -2467 -20643 -2327
rect -20089 -2467 -20047 -2327
rect -20681 -2506 -20047 -2467
rect -22793 -2674 -22379 -2655
rect -24635 -2797 -24492 -2791
rect -23295 -2720 -23221 -2716
rect -23295 -2747 -23074 -2720
rect -23628 -2878 -23428 -2850
rect -24603 -2987 -24394 -2940
rect -24603 -3165 -24550 -2987
rect -24428 -3165 -24394 -2987
rect -24213 -2983 -23813 -2955
rect -24213 -3057 -24184 -2983
rect -23844 -3057 -23813 -2983
rect -23628 -2974 -23601 -2878
rect -23452 -2974 -23428 -2878
rect -23295 -2866 -23253 -2747
rect -23121 -2866 -23074 -2747
rect -22793 -2767 -22731 -2674
rect -22413 -2767 -22379 -2674
rect -20952 -2675 -20644 -2652
rect -22793 -2791 -22379 -2767
rect -21319 -2720 -21288 -2716
rect -21319 -2775 -21179 -2720
rect -23295 -2907 -23074 -2866
rect -23628 -3000 -23428 -2974
rect -24213 -3078 -23813 -3057
rect -24603 -3194 -24394 -3165
rect -23260 -3504 -23074 -2907
rect -22627 -2852 -22400 -2819
rect -22627 -3080 -22594 -2852
rect -22431 -3080 -22400 -2852
rect -21608 -2878 -21408 -2850
rect -22176 -2983 -21776 -2955
rect -22176 -3057 -22147 -2983
rect -21807 -3057 -21776 -2983
rect -21608 -2974 -21581 -2878
rect -21432 -2974 -21408 -2878
rect -21608 -3000 -21408 -2974
rect -21319 -2859 -21293 -2775
rect -21209 -2859 -21179 -2775
rect -20952 -2772 -20889 -2675
rect -20682 -2772 -20644 -2675
rect -19111 -2653 -18968 -2113
rect -8187 -2171 9917 -2105
rect 9983 -2171 9989 -2105
rect -18088 -2225 -17874 -2203
rect -18921 -2327 -18287 -2293
rect -18088 -2304 -18065 -2225
rect -17896 -2304 -17874 -2225
rect -18088 -2323 -17874 -2304
rect -18921 -2467 -18883 -2327
rect -18329 -2467 -18287 -2327
rect -18921 -2506 -18287 -2467
rect -19111 -2673 -18806 -2653
rect -20952 -2792 -20644 -2772
rect -19567 -2721 -19528 -2716
rect -19567 -2780 -19444 -2721
rect -22176 -3078 -21776 -3057
rect -22627 -3113 -22400 -3080
rect -21319 -3398 -21179 -2859
rect -19867 -2878 -19667 -2850
rect -20446 -2983 -20046 -2955
rect -20944 -3042 -20726 -3021
rect -20944 -3165 -20917 -3042
rect -20741 -3165 -20726 -3042
rect -20446 -3057 -20417 -2983
rect -20077 -3057 -20046 -2983
rect -19867 -2974 -19840 -2878
rect -19691 -2974 -19667 -2878
rect -19567 -2864 -19555 -2780
rect -19471 -2864 -19444 -2780
rect -19111 -2780 -19043 -2673
rect -18894 -2780 -18806 -2673
rect -19111 -2792 -18806 -2780
rect -17726 -2696 -17436 -2677
rect -19567 -2904 -19444 -2864
rect -19867 -3000 -19667 -2974
rect -20446 -3078 -20046 -3057
rect -20944 -3186 -20726 -3165
rect -19539 -3246 -19444 -2904
rect -18088 -2878 -17888 -2850
rect -17726 -2852 -17693 -2696
rect -17579 -2852 -17436 -2696
rect -17726 -2864 -17436 -2852
rect -19292 -2934 -19012 -2908
rect -19292 -3087 -19241 -2934
rect -19043 -3087 -19012 -2934
rect -18686 -2983 -18286 -2955
rect -18686 -3057 -18657 -2983
rect -18317 -3057 -18286 -2983
rect -18088 -2974 -18061 -2878
rect -17912 -2974 -17888 -2878
rect -18088 -3000 -17888 -2974
rect -18686 -3078 -18286 -3057
rect -17591 -3045 -17436 -2864
rect -8187 -3045 -8121 -2171
rect 5732 -2226 7106 -2211
rect -6334 -2274 7106 -2226
rect -19292 -3115 -19012 -3087
rect -17591 -3167 -7885 -3045
rect -17586 -3195 -7885 -3167
rect -19539 -3247 -10885 -3246
rect -19539 -3355 -10874 -3247
rect -22329 -3504 -22012 -3495
rect -23260 -3565 -22012 -3504
rect -21329 -3509 -14165 -3398
rect -23260 -3617 -17462 -3565
rect -22329 -3678 -17462 -3617
rect -22329 -3687 -22012 -3678
rect -22913 -3714 -22744 -3704
rect -22913 -3742 -22451 -3714
rect -22913 -3848 -22600 -3742
rect -22476 -3848 -22451 -3742
rect -22913 -3877 -22451 -3848
rect -24861 -4064 -24578 -3997
rect -24861 -4337 -24807 -4064
rect -24618 -4337 -24578 -4064
rect -23584 -4037 -23370 -4015
rect -24397 -4139 -23763 -4105
rect -23584 -4116 -23561 -4037
rect -23392 -4116 -23370 -4037
rect -23584 -4135 -23370 -4116
rect -24397 -4279 -24359 -4139
rect -23805 -4279 -23763 -4139
rect -24397 -4318 -23763 -4279
rect -24861 -4379 -24578 -4337
rect -22913 -4468 -22744 -3877
rect -21846 -4037 -21632 -4015
rect -22661 -4139 -22027 -4105
rect -21846 -4116 -21823 -4037
rect -21654 -4116 -21632 -4037
rect -21846 -4135 -21632 -4116
rect -22661 -4279 -22623 -4139
rect -22069 -4279 -22027 -4139
rect -22661 -4318 -22027 -4279
rect -23210 -4469 -22736 -4468
rect -23210 -4480 -22655 -4469
rect -23210 -4594 -23195 -4480
rect -23064 -4481 -22655 -4480
rect -23064 -4594 -22836 -4481
rect -22690 -4594 -22655 -4481
rect -23210 -4603 -22655 -4594
rect -23584 -4690 -23384 -4662
rect -24162 -4795 -23762 -4767
rect -24162 -4869 -24133 -4795
rect -23793 -4869 -23762 -4795
rect -23584 -4786 -23557 -4690
rect -23408 -4786 -23384 -4690
rect -21846 -4690 -21646 -4662
rect -23584 -4812 -23384 -4786
rect -22426 -4795 -22026 -4767
rect -24162 -4890 -23762 -4869
rect -22426 -4869 -22397 -4795
rect -22057 -4869 -22026 -4795
rect -21846 -4786 -21819 -4690
rect -21670 -4786 -21646 -4690
rect -21047 -4756 -20938 -3746
rect -20872 -4599 -20758 -3746
rect -17756 -3763 -17647 -3746
rect -20649 -3827 -19439 -3799
rect -20649 -3899 -20603 -3827
rect -19481 -3899 -19439 -3827
rect -20649 -3925 -19439 -3899
rect -19090 -3827 -17880 -3799
rect -19090 -3899 -19044 -3827
rect -17922 -3899 -17880 -3827
rect -19090 -3925 -17880 -3899
rect -17756 -3858 -17744 -3763
rect -17655 -3858 -17647 -3763
rect -17586 -3823 -17463 -3678
rect -14465 -3762 -14356 -3746
rect -20872 -4622 -20469 -4599
rect -20872 -4730 -20848 -4622
rect -20758 -4730 -20469 -4622
rect -20872 -4752 -20469 -4730
rect -20872 -4753 -20758 -4752
rect -21356 -4763 -20938 -4756
rect -21846 -4812 -21646 -4786
rect -22426 -4890 -22026 -4869
rect -21395 -4842 -20938 -4763
rect -21395 -4843 -20690 -4842
rect -21395 -4855 -20661 -4843
rect -21395 -4896 -20751 -4855
rect -24622 -4997 -24472 -4989
rect -25512 -5030 -25432 -5026
rect -25060 -5030 -24615 -4997
rect -25512 -5035 -24615 -5030
rect -25512 -5097 -25504 -5035
rect -25442 -5097 -24615 -5035
rect -25512 -5102 -24615 -5097
rect -25512 -5106 -25432 -5102
rect -25060 -5133 -24615 -5102
rect -24479 -5133 -22868 -4997
rect -22732 -5133 -22726 -4997
rect -24622 -5141 -24472 -5133
rect -23586 -5329 -23372 -5307
rect -24397 -5431 -23763 -5397
rect -23586 -5408 -23563 -5329
rect -23394 -5408 -23372 -5329
rect -21852 -5329 -21638 -5307
rect -23586 -5427 -23372 -5408
rect -24397 -5571 -24359 -5431
rect -23805 -5571 -23763 -5431
rect -24397 -5610 -23763 -5571
rect -22661 -5431 -22027 -5397
rect -21852 -5408 -21829 -5329
rect -21660 -5408 -21638 -5329
rect -21852 -5427 -21638 -5408
rect -22661 -5571 -22623 -5431
rect -22069 -5571 -22027 -5431
rect -22661 -5610 -22027 -5571
rect -21562 -5705 -21477 -5703
rect -21395 -5705 -21304 -4896
rect -21047 -4955 -20751 -4896
rect -20773 -4963 -20751 -4955
rect -20675 -4963 -20661 -4855
rect -21610 -5731 -21304 -5705
rect -21610 -5922 -21560 -5731
rect -21347 -5922 -21304 -5731
rect -22912 -5936 -22624 -5924
rect -23586 -5982 -23386 -5954
rect -24637 -6049 -24439 -6020
rect -24637 -6247 -24612 -6049
rect -24466 -6247 -24439 -6049
rect -24162 -6087 -23762 -6059
rect -24162 -6161 -24133 -6087
rect -23793 -6161 -23762 -6087
rect -23586 -6078 -23559 -5982
rect -23410 -6078 -23386 -5982
rect -23586 -6104 -23386 -6078
rect -22912 -6046 -22884 -5936
rect -22652 -6046 -22624 -5936
rect -24162 -6182 -23762 -6161
rect -24637 -6262 -24439 -6247
rect -22912 -6441 -22862 -6046
rect -22773 -6059 -22624 -6046
rect -21852 -5982 -21652 -5954
rect -21610 -5968 -21304 -5922
rect -21039 -5333 -20854 -5317
rect -21039 -5435 -21003 -5333
rect -20885 -5435 -20854 -5333
rect -22773 -6339 -22736 -6059
rect -22426 -6087 -22026 -6059
rect -22426 -6161 -22397 -6087
rect -22057 -6161 -22026 -6087
rect -21852 -6078 -21825 -5982
rect -21676 -6078 -21652 -5982
rect -21852 -6104 -21652 -6078
rect -22426 -6182 -22026 -6161
rect -22773 -6441 -22737 -6339
rect -22912 -6485 -22737 -6441
rect -21039 -6427 -20854 -5435
rect -20773 -6128 -20672 -4963
rect -20565 -5928 -20469 -4752
rect -19456 -4674 -19184 -4658
rect -19456 -4771 -19372 -4674
rect -19222 -4771 -19184 -4674
rect -19456 -4806 -19184 -4771
rect -20154 -5219 -20072 -5208
rect -20154 -5279 -20143 -5219
rect -20083 -5279 -20072 -5219
rect -20154 -5290 -20072 -5279
rect -19751 -5368 -19620 -5352
rect -19751 -5437 -19735 -5368
rect -19636 -5437 -19620 -5368
rect -20354 -5559 -20080 -5550
rect -20354 -5631 -20345 -5559
rect -20089 -5631 -20080 -5559
rect -20354 -5640 -20080 -5631
rect -19992 -5894 -19883 -5879
rect -20566 -5955 -20402 -5928
rect -20566 -6035 -20534 -5955
rect -20436 -6035 -20402 -5955
rect -20566 -6063 -20402 -6035
rect -19992 -6042 -19979 -5894
rect -19896 -6042 -19883 -5894
rect -19992 -6054 -19883 -6042
rect -20773 -6148 -20402 -6128
rect -20773 -6214 -20743 -6148
rect -20490 -6214 -20402 -6148
rect -20773 -6227 -20402 -6214
rect -20278 -6301 -19925 -6292
rect -20278 -6357 -20269 -6301
rect -19934 -6357 -19925 -6301
rect -20278 -6366 -19925 -6357
rect -21039 -6431 -20757 -6427
rect -21039 -6521 -20729 -6431
rect -21034 -6632 -20729 -6521
rect -19751 -6440 -19620 -5437
rect -19456 -5933 -19360 -4806
rect -19237 -4862 -19031 -4836
rect -19237 -4959 -19196 -4862
rect -19080 -4959 -19031 -4862
rect -17756 -4842 -17647 -3858
rect -17581 -4599 -17467 -3823
rect -17358 -3827 -16148 -3799
rect -17358 -3899 -17312 -3827
rect -16190 -3899 -16148 -3827
rect -17358 -3925 -16148 -3899
rect -15799 -3827 -14589 -3799
rect -15799 -3899 -15753 -3827
rect -14631 -3899 -14589 -3827
rect -15799 -3925 -14589 -3899
rect -14465 -3946 -14460 -3762
rect -14361 -3946 -14356 -3762
rect -14294 -3855 -14166 -3509
rect -11174 -3761 -11065 -3746
rect -14067 -3827 -12857 -3799
rect -17581 -4622 -17178 -4599
rect -17581 -4730 -17557 -4622
rect -17467 -4730 -17178 -4622
rect -17581 -4752 -17178 -4730
rect -17581 -4753 -17467 -4752
rect -17756 -4843 -17399 -4842
rect -17756 -4855 -17370 -4843
rect -17756 -4955 -17460 -4855
rect -19237 -4979 -19031 -4959
rect -17482 -4963 -17460 -4955
rect -17384 -4963 -17370 -4855
rect -19237 -5364 -19142 -4979
rect -17756 -5153 -17647 -5144
rect -18595 -5219 -18513 -5208
rect -18595 -5279 -18584 -5219
rect -18524 -5279 -18513 -5219
rect -18595 -5290 -18513 -5279
rect -17756 -5239 -17747 -5153
rect -17656 -5239 -17647 -5153
rect -19237 -5430 -19223 -5364
rect -19152 -5430 -19142 -5364
rect -19457 -5956 -19293 -5933
rect -19457 -6036 -19423 -5956
rect -19325 -6036 -19293 -5956
rect -19457 -6063 -19293 -6036
rect -19237 -6144 -19142 -5430
rect -19065 -5559 -18791 -5550
rect -19065 -5631 -19056 -5559
rect -18800 -5631 -18791 -5559
rect -19065 -5640 -18791 -5631
rect -18348 -5559 -18074 -5550
rect -18348 -5631 -18339 -5559
rect -18083 -5631 -18074 -5559
rect -18348 -5640 -18074 -5631
rect -18047 -5944 -17869 -5893
rect -18047 -6024 -18002 -5944
rect -17882 -6024 -17869 -5944
rect -18047 -6041 -17869 -6024
rect -19457 -6159 -19142 -6144
rect -19457 -6219 -19433 -6159
rect -19248 -6219 -19142 -6159
rect -18573 -6110 -18398 -6099
rect -18573 -6185 -18561 -6110
rect -18416 -6185 -18398 -6110
rect -18573 -6197 -18398 -6185
rect -19457 -6229 -19142 -6219
rect -19044 -6310 -18960 -6298
rect -19044 -6372 -19033 -6310
rect -18971 -6372 -18960 -6310
rect -19044 -6383 -18960 -6372
rect -18179 -6335 -18101 -6324
rect -18179 -6391 -18168 -6335
rect -18112 -6391 -18101 -6335
rect -18179 -6402 -18101 -6391
rect -18047 -6440 -17927 -6041
rect -17756 -6359 -17647 -5239
rect -17482 -6128 -17381 -4963
rect -17274 -5928 -17178 -4752
rect -16165 -4674 -15893 -4658
rect -16165 -4771 -16081 -4674
rect -15931 -4771 -15893 -4674
rect -16165 -4806 -15893 -4771
rect -16863 -5219 -16781 -5208
rect -16863 -5279 -16852 -5219
rect -16792 -5279 -16781 -5219
rect -16863 -5290 -16781 -5279
rect -16460 -5368 -16329 -5352
rect -16460 -5437 -16444 -5368
rect -16345 -5437 -16329 -5368
rect -17063 -5559 -16789 -5550
rect -17063 -5631 -17054 -5559
rect -16798 -5631 -16789 -5559
rect -17063 -5640 -16789 -5631
rect -16701 -5894 -16592 -5879
rect -17275 -5955 -17111 -5928
rect -17275 -6035 -17243 -5955
rect -17145 -6035 -17111 -5955
rect -17275 -6063 -17111 -6035
rect -16701 -6042 -16688 -5894
rect -16605 -6042 -16592 -5894
rect -16701 -6054 -16592 -6042
rect -17482 -6148 -17111 -6128
rect -17482 -6214 -17452 -6148
rect -17199 -6214 -17111 -6148
rect -17482 -6227 -17111 -6214
rect -16987 -6301 -16634 -6292
rect -16987 -6357 -16978 -6301
rect -16643 -6357 -16634 -6301
rect -19751 -6542 -17927 -6440
rect -17769 -6444 -17637 -6359
rect -16987 -6366 -16634 -6357
rect -16460 -6440 -16329 -5437
rect -16165 -5933 -16069 -4806
rect -15946 -4862 -15740 -4836
rect -15946 -4959 -15905 -4862
rect -15789 -4959 -15740 -4862
rect -14465 -4842 -14356 -3946
rect -14290 -4599 -14176 -3855
rect -14067 -3899 -14021 -3827
rect -12899 -3899 -12857 -3827
rect -14067 -3925 -12857 -3899
rect -12508 -3827 -11298 -3799
rect -12508 -3899 -12462 -3827
rect -11340 -3899 -11298 -3827
rect -12508 -3925 -11298 -3899
rect -11174 -3905 -11165 -3761
rect -11074 -3905 -11065 -3761
rect -11016 -3843 -10874 -3355
rect -10776 -3827 -9566 -3799
rect -14290 -4622 -13887 -4599
rect -14290 -4730 -14266 -4622
rect -14176 -4730 -13887 -4622
rect -14290 -4752 -13887 -4730
rect -14290 -4753 -14176 -4752
rect -14465 -4843 -14108 -4842
rect -14465 -4855 -14079 -4843
rect -14465 -4955 -14169 -4855
rect -15946 -4979 -15740 -4959
rect -14191 -4963 -14169 -4955
rect -14093 -4963 -14079 -4855
rect -15946 -5364 -15851 -4979
rect -14465 -5153 -14356 -5144
rect -15304 -5219 -15222 -5208
rect -15304 -5279 -15293 -5219
rect -15233 -5279 -15222 -5219
rect -15304 -5290 -15222 -5279
rect -14465 -5239 -14456 -5153
rect -14365 -5239 -14356 -5153
rect -15946 -5430 -15932 -5364
rect -15861 -5430 -15851 -5364
rect -16166 -5956 -16002 -5933
rect -16166 -6036 -16132 -5956
rect -16034 -6036 -16002 -5956
rect -16166 -6063 -16002 -6036
rect -15946 -6144 -15851 -5430
rect -15774 -5559 -15500 -5550
rect -15774 -5631 -15765 -5559
rect -15509 -5631 -15500 -5559
rect -15774 -5640 -15500 -5631
rect -15057 -5559 -14783 -5550
rect -15057 -5631 -15048 -5559
rect -14792 -5631 -14783 -5559
rect -15057 -5640 -14783 -5631
rect -14756 -5944 -14578 -5893
rect -14756 -6024 -14711 -5944
rect -14591 -6024 -14578 -5944
rect -14756 -6041 -14578 -6024
rect -16166 -6159 -15851 -6144
rect -16166 -6219 -16142 -6159
rect -15957 -6219 -15851 -6159
rect -15282 -6110 -15107 -6099
rect -15282 -6185 -15270 -6110
rect -15125 -6185 -15107 -6110
rect -15282 -6197 -15107 -6185
rect -16166 -6229 -15851 -6219
rect -15753 -6310 -15669 -6298
rect -15753 -6372 -15742 -6310
rect -15680 -6372 -15669 -6310
rect -15753 -6383 -15669 -6372
rect -14888 -6335 -14810 -6324
rect -14888 -6391 -14877 -6335
rect -14821 -6391 -14810 -6335
rect -14888 -6402 -14810 -6391
rect -14756 -6440 -14636 -6041
rect -14465 -6314 -14356 -5239
rect -14191 -6128 -14090 -4963
rect -13983 -5928 -13887 -4752
rect -12874 -4674 -12602 -4658
rect -12874 -4771 -12790 -4674
rect -12640 -4771 -12602 -4674
rect -12874 -4806 -12602 -4771
rect -13572 -5219 -13490 -5208
rect -13572 -5279 -13561 -5219
rect -13501 -5279 -13490 -5219
rect -13572 -5290 -13490 -5279
rect -13169 -5368 -13038 -5352
rect -13169 -5437 -13153 -5368
rect -13054 -5437 -13038 -5368
rect -13772 -5559 -13498 -5550
rect -13772 -5631 -13763 -5559
rect -13507 -5631 -13498 -5559
rect -13772 -5640 -13498 -5631
rect -13410 -5894 -13301 -5879
rect -13984 -5955 -13820 -5928
rect -13984 -6035 -13952 -5955
rect -13854 -6035 -13820 -5955
rect -13984 -6063 -13820 -6035
rect -13410 -6042 -13397 -5894
rect -13314 -6042 -13301 -5894
rect -13410 -6054 -13301 -6042
rect -14191 -6148 -13820 -6128
rect -14191 -6214 -14161 -6148
rect -13908 -6214 -13820 -6148
rect -14191 -6227 -13820 -6214
rect -13696 -6301 -13343 -6292
rect -14470 -6418 -14163 -6314
rect -13696 -6357 -13687 -6301
rect -13352 -6357 -13343 -6301
rect -13696 -6366 -13343 -6357
rect -17769 -6574 -17406 -6444
rect -16460 -6542 -14636 -6440
rect -17702 -6575 -17406 -6574
rect -24648 -6678 -21343 -6658
rect -24648 -6684 -21515 -6678
rect -25655 -6746 -25576 -6742
rect -24648 -6746 -24619 -6684
rect -25659 -6751 -24619 -6746
rect -25659 -6832 -25655 -6751
rect -25576 -6824 -24619 -6751
rect -24490 -6818 -21515 -6684
rect -21386 -6818 -21343 -6678
rect -24490 -6824 -21343 -6818
rect -25576 -6832 -21343 -6824
rect -25659 -6835 -21343 -6832
rect -25655 -6841 -25576 -6835
rect -24648 -6845 -21343 -6835
rect -23585 -7302 -23371 -7280
rect -24397 -7404 -23763 -7370
rect -23585 -7381 -23562 -7302
rect -23393 -7381 -23371 -7302
rect -21850 -7302 -21636 -7280
rect -23585 -7400 -23371 -7381
rect -24397 -7544 -24359 -7404
rect -23805 -7544 -23763 -7404
rect -24397 -7583 -23763 -7544
rect -22660 -7404 -22026 -7370
rect -21850 -7381 -21827 -7302
rect -21658 -7381 -21636 -7302
rect -21850 -7400 -21636 -7381
rect -22660 -7544 -22622 -7404
rect -22068 -7544 -22026 -7404
rect -22660 -7583 -22026 -7544
rect -23210 -7743 -22667 -7733
rect -23210 -7857 -23198 -7743
rect -23067 -7745 -22667 -7743
rect -23064 -7749 -22667 -7745
rect -23064 -7856 -22808 -7749
rect -22688 -7856 -22667 -7749
rect -23210 -7859 -23195 -7857
rect -23064 -7859 -22667 -7856
rect -23210 -7868 -22667 -7859
rect -24632 -7911 -24342 -7897
rect -24632 -8015 -24611 -7911
rect -24368 -8015 -24342 -7911
rect -22910 -7907 -22614 -7897
rect -24632 -8033 -24342 -8015
rect -23585 -7955 -23385 -7927
rect -24632 -8292 -24456 -8033
rect -24162 -8060 -23762 -8032
rect -24162 -8134 -24133 -8060
rect -23793 -8134 -23762 -8060
rect -23585 -8051 -23558 -7955
rect -23409 -8051 -23385 -7955
rect -23585 -8077 -23385 -8051
rect -22910 -8015 -22857 -7907
rect -22628 -8015 -22614 -7907
rect -22910 -8038 -22614 -8015
rect -21850 -7955 -21650 -7927
rect -24162 -8155 -23762 -8134
rect -22910 -8292 -22734 -8038
rect -22425 -8060 -22025 -8032
rect -22425 -8134 -22396 -8060
rect -22056 -8134 -22025 -8060
rect -21850 -8051 -21823 -7955
rect -21674 -8051 -21650 -7955
rect -21047 -8021 -20938 -7011
rect -20873 -7053 -20729 -6632
rect -17756 -7028 -17647 -7011
rect -20872 -7864 -20758 -7053
rect -20649 -7092 -19439 -7064
rect -20649 -7164 -20603 -7092
rect -19481 -7164 -19439 -7092
rect -20649 -7190 -19439 -7164
rect -19090 -7092 -17880 -7064
rect -19090 -7164 -19044 -7092
rect -17922 -7164 -17880 -7092
rect -19090 -7190 -17880 -7164
rect -17756 -7123 -17744 -7028
rect -17655 -7123 -17647 -7028
rect -17592 -7079 -17408 -6575
rect -14289 -7011 -14166 -6418
rect -13169 -6440 -13038 -5437
rect -12874 -5933 -12778 -4806
rect -12655 -4862 -12449 -4836
rect -12655 -4959 -12614 -4862
rect -12498 -4959 -12449 -4862
rect -11174 -4842 -11065 -3905
rect -10999 -4599 -10885 -3843
rect -10776 -3899 -10730 -3827
rect -9608 -3899 -9566 -3827
rect -10776 -3925 -9566 -3899
rect -9217 -3827 -8007 -3799
rect -9217 -3899 -9171 -3827
rect -8049 -3899 -8007 -3827
rect -9217 -3925 -8007 -3899
rect -10999 -4622 -10596 -4599
rect -10999 -4730 -10975 -4622
rect -10885 -4730 -10596 -4622
rect -10999 -4752 -10596 -4730
rect -10999 -4753 -10885 -4752
rect -11174 -4843 -10817 -4842
rect -11174 -4855 -10788 -4843
rect -11174 -4955 -10878 -4855
rect -12655 -4979 -12449 -4959
rect -10900 -4963 -10878 -4955
rect -10802 -4963 -10788 -4855
rect -12655 -5364 -12560 -4979
rect -11174 -5153 -11065 -5144
rect -12013 -5219 -11931 -5208
rect -12013 -5279 -12002 -5219
rect -11942 -5279 -11931 -5219
rect -12013 -5290 -11931 -5279
rect -11174 -5239 -11165 -5153
rect -11074 -5239 -11065 -5153
rect -12655 -5430 -12641 -5364
rect -12570 -5430 -12560 -5364
rect -12875 -5956 -12711 -5933
rect -12875 -6036 -12841 -5956
rect -12743 -6036 -12711 -5956
rect -12875 -6063 -12711 -6036
rect -12655 -6144 -12560 -5430
rect -12483 -5559 -12209 -5550
rect -12483 -5631 -12474 -5559
rect -12218 -5631 -12209 -5559
rect -12483 -5640 -12209 -5631
rect -11766 -5559 -11492 -5550
rect -11766 -5631 -11757 -5559
rect -11501 -5631 -11492 -5559
rect -11766 -5640 -11492 -5631
rect -11465 -5944 -11287 -5893
rect -11465 -6024 -11420 -5944
rect -11300 -6024 -11287 -5944
rect -11465 -6041 -11287 -6024
rect -12875 -6159 -12560 -6144
rect -12875 -6219 -12851 -6159
rect -12666 -6219 -12560 -6159
rect -11991 -6110 -11816 -6099
rect -11991 -6185 -11979 -6110
rect -11834 -6185 -11816 -6110
rect -11991 -6197 -11816 -6185
rect -12875 -6229 -12560 -6219
rect -12462 -6310 -12378 -6298
rect -12462 -6372 -12451 -6310
rect -12389 -6372 -12378 -6310
rect -12462 -6383 -12378 -6372
rect -11597 -6335 -11519 -6324
rect -11597 -6391 -11586 -6335
rect -11530 -6391 -11519 -6335
rect -11597 -6402 -11519 -6391
rect -11465 -6440 -11345 -6041
rect -13169 -6542 -11345 -6440
rect -11174 -6332 -11065 -5239
rect -10900 -6128 -10799 -4963
rect -10692 -5928 -10596 -4752
rect -9583 -4674 -9311 -4658
rect -9583 -4771 -9499 -4674
rect -9349 -4771 -9311 -4674
rect -9583 -4806 -9311 -4771
rect -10281 -5219 -10199 -5208
rect -10281 -5279 -10270 -5219
rect -10210 -5279 -10199 -5219
rect -10281 -5290 -10199 -5279
rect -9878 -5368 -9747 -5352
rect -9878 -5437 -9862 -5368
rect -9763 -5437 -9747 -5368
rect -10481 -5559 -10207 -5550
rect -10481 -5631 -10472 -5559
rect -10216 -5631 -10207 -5559
rect -10481 -5640 -10207 -5631
rect -10119 -5894 -10010 -5879
rect -10693 -5955 -10529 -5928
rect -10693 -6035 -10661 -5955
rect -10563 -6035 -10529 -5955
rect -10693 -6063 -10529 -6035
rect -10119 -6042 -10106 -5894
rect -10023 -6042 -10010 -5894
rect -10119 -6054 -10010 -6042
rect -10900 -6148 -10529 -6128
rect -10900 -6214 -10870 -6148
rect -10617 -6214 -10529 -6148
rect -10900 -6227 -10529 -6214
rect -10405 -6301 -10052 -6292
rect -11174 -6472 -11047 -6332
rect -10405 -6357 -10396 -6301
rect -10061 -6357 -10052 -6301
rect -10405 -6366 -10052 -6357
rect -9878 -6440 -9747 -5437
rect -9583 -5933 -9487 -4806
rect -9364 -4862 -9158 -4836
rect -9364 -4959 -9323 -4862
rect -9207 -4959 -9158 -4862
rect -9364 -4979 -9158 -4959
rect -9364 -5364 -9269 -4979
rect -7883 -5153 -7774 -5144
rect -8722 -5219 -8640 -5208
rect -8722 -5279 -8711 -5219
rect -8651 -5279 -8640 -5219
rect -8722 -5290 -8640 -5279
rect -7883 -5239 -7874 -5153
rect -7783 -5239 -7774 -5153
rect -9364 -5430 -9350 -5364
rect -9279 -5430 -9269 -5364
rect -9584 -5956 -9420 -5933
rect -9584 -6036 -9550 -5956
rect -9452 -6036 -9420 -5956
rect -9584 -6063 -9420 -6036
rect -9364 -6144 -9269 -5430
rect -9192 -5559 -8918 -5550
rect -9192 -5631 -9183 -5559
rect -8927 -5631 -8918 -5559
rect -9192 -5640 -8918 -5631
rect -8475 -5559 -8201 -5550
rect -8475 -5631 -8466 -5559
rect -8210 -5631 -8201 -5559
rect -8475 -5640 -8201 -5631
rect -8174 -5944 -7996 -5893
rect -8174 -6024 -8129 -5944
rect -8009 -6024 -7996 -5944
rect -8174 -6041 -7996 -6024
rect -9584 -6159 -9269 -6144
rect -9584 -6219 -9560 -6159
rect -9375 -6219 -9269 -6159
rect -8700 -6110 -8525 -6099
rect -8700 -6185 -8688 -6110
rect -8543 -6185 -8525 -6110
rect -8700 -6197 -8525 -6185
rect -9584 -6229 -9269 -6219
rect -9171 -6310 -9087 -6298
rect -9171 -6372 -9160 -6310
rect -9098 -6372 -9087 -6310
rect -9171 -6383 -9087 -6372
rect -8306 -6335 -8228 -6324
rect -8306 -6391 -8295 -6335
rect -8239 -6391 -8228 -6335
rect -8306 -6402 -8228 -6391
rect -8174 -6440 -8054 -6041
rect -7883 -6175 -7774 -5239
rect -7890 -6225 -7762 -6175
rect -7890 -6291 -7873 -6225
rect -7807 -6269 -7762 -6225
rect -7807 -6291 -7688 -6269
rect -7890 -6367 -7688 -6291
rect -7888 -6380 -7688 -6367
rect -7883 -6381 -7774 -6380
rect -11004 -6472 -10876 -6471
rect -11179 -6628 -10876 -6472
rect -9878 -6542 -8054 -6440
rect -11174 -6629 -11047 -6628
rect -14465 -7027 -14356 -7011
rect -20872 -7887 -20469 -7864
rect -20872 -7995 -20848 -7887
rect -20758 -7995 -20469 -7887
rect -20872 -8017 -20469 -7995
rect -20872 -8018 -20758 -8017
rect -21356 -8028 -20938 -8021
rect -21850 -8077 -21650 -8051
rect -22425 -8155 -22025 -8134
rect -21395 -8107 -20938 -8028
rect -21395 -8108 -20690 -8107
rect -21395 -8120 -20661 -8108
rect -25809 -8297 -25749 -8293
rect -24634 -8297 -22734 -8292
rect -25814 -8302 -22734 -8297
rect -25814 -8362 -25809 -8302
rect -25749 -8362 -22734 -8302
rect -25814 -8367 -22734 -8362
rect -25809 -8371 -25749 -8367
rect -24634 -8427 -22734 -8367
rect -24632 -9025 -24456 -8427
rect -23583 -8594 -23369 -8572
rect -24397 -8696 -23763 -8662
rect -23583 -8673 -23560 -8594
rect -23391 -8673 -23369 -8594
rect -23583 -8692 -23369 -8673
rect -24397 -8836 -24359 -8696
rect -23805 -8836 -23763 -8696
rect -24397 -8875 -23763 -8836
rect -22910 -9025 -22734 -8427
rect -21395 -8161 -20751 -8120
rect -21846 -8594 -21632 -8572
rect -22661 -8696 -22027 -8662
rect -21846 -8673 -21823 -8594
rect -21654 -8673 -21632 -8594
rect -21846 -8692 -21632 -8673
rect -22661 -8836 -22623 -8696
rect -22069 -8836 -22027 -8696
rect -22661 -8875 -22027 -8836
rect -21562 -8970 -21477 -8968
rect -21395 -8970 -21304 -8161
rect -21047 -8220 -20751 -8161
rect -20773 -8228 -20751 -8220
rect -20675 -8228 -20661 -8120
rect -21610 -9019 -21304 -8970
rect -24632 -9039 -24432 -9025
rect -24632 -9146 -24601 -9039
rect -24445 -9146 -24432 -9039
rect -24632 -9160 -24432 -9146
rect -22910 -9026 -22688 -9025
rect -22910 -9037 -22658 -9026
rect -22910 -9148 -22885 -9037
rect -22683 -9148 -22658 -9037
rect -22910 -9160 -22658 -9148
rect -22913 -9211 -22653 -9189
rect -23583 -9247 -23383 -9219
rect -24637 -9314 -24439 -9285
rect -24637 -9512 -24612 -9314
rect -24466 -9512 -24439 -9314
rect -24162 -9352 -23762 -9324
rect -24162 -9426 -24133 -9352
rect -23793 -9426 -23762 -9352
rect -23583 -9343 -23556 -9247
rect -23407 -9343 -23383 -9247
rect -22913 -9303 -22891 -9211
rect -22686 -9303 -22653 -9211
rect -21610 -9193 -21573 -9019
rect -21351 -9193 -21304 -9019
rect -22913 -9325 -22866 -9303
rect -23583 -9369 -23383 -9343
rect -24162 -9447 -23762 -9426
rect -24637 -9527 -24439 -9512
rect -22911 -9685 -22866 -9325
rect -22773 -9325 -22653 -9303
rect -21846 -9247 -21646 -9219
rect -21610 -9233 -21304 -9193
rect -21039 -8598 -20854 -8582
rect -21039 -8700 -21003 -8598
rect -20885 -8700 -20854 -8598
rect -22773 -9604 -22736 -9325
rect -22426 -9352 -22026 -9324
rect -22426 -9426 -22397 -9352
rect -22057 -9426 -22026 -9352
rect -21846 -9343 -21819 -9247
rect -21670 -9343 -21646 -9247
rect -21846 -9369 -21646 -9343
rect -22426 -9447 -22026 -9426
rect -22911 -9706 -22862 -9685
rect -22773 -9706 -22737 -9604
rect -22911 -9750 -22737 -9706
rect -21039 -9726 -20854 -8700
rect -20773 -9393 -20672 -8228
rect -20565 -9193 -20469 -8017
rect -19456 -7939 -19184 -7923
rect -19456 -8036 -19372 -7939
rect -19222 -8036 -19184 -7939
rect -19456 -8071 -19184 -8036
rect -20154 -8484 -20072 -8473
rect -20154 -8544 -20143 -8484
rect -20083 -8544 -20072 -8484
rect -20154 -8555 -20072 -8544
rect -19751 -8633 -19620 -8617
rect -19751 -8702 -19735 -8633
rect -19636 -8702 -19620 -8633
rect -20354 -8824 -20080 -8815
rect -20354 -8896 -20345 -8824
rect -20089 -8896 -20080 -8824
rect -20354 -8905 -20080 -8896
rect -19992 -9159 -19883 -9144
rect -20566 -9220 -20402 -9193
rect -20566 -9300 -20534 -9220
rect -20436 -9300 -20402 -9220
rect -20566 -9328 -20402 -9300
rect -19992 -9307 -19979 -9159
rect -19896 -9307 -19883 -9159
rect -19992 -9319 -19883 -9307
rect -20773 -9413 -20402 -9393
rect -20773 -9479 -20743 -9413
rect -20490 -9479 -20402 -9413
rect -20773 -9492 -20402 -9479
rect -20278 -9566 -19925 -9557
rect -20278 -9622 -20269 -9566
rect -19934 -9622 -19925 -9566
rect -20278 -9631 -19925 -9622
rect -19751 -9705 -19620 -8702
rect -19456 -9198 -19360 -8071
rect -19237 -8127 -19031 -8101
rect -19237 -8224 -19196 -8127
rect -19080 -8224 -19031 -8127
rect -17756 -8107 -17647 -7123
rect -17581 -7864 -17467 -7079
rect -17358 -7092 -16148 -7064
rect -17358 -7164 -17312 -7092
rect -16190 -7164 -16148 -7092
rect -17358 -7190 -16148 -7164
rect -15799 -7092 -14589 -7064
rect -15799 -7164 -15753 -7092
rect -14631 -7164 -14589 -7092
rect -15799 -7190 -14589 -7164
rect -14465 -7211 -14460 -7027
rect -14361 -7211 -14356 -7027
rect -17581 -7887 -17178 -7864
rect -17581 -7995 -17557 -7887
rect -17467 -7995 -17178 -7887
rect -17581 -8017 -17178 -7995
rect -17581 -8018 -17467 -8017
rect -17756 -8108 -17399 -8107
rect -17756 -8120 -17370 -8108
rect -17756 -8220 -17460 -8120
rect -19237 -8244 -19031 -8224
rect -17482 -8228 -17460 -8220
rect -17384 -8228 -17370 -8120
rect -19237 -8629 -19142 -8244
rect -17756 -8418 -17647 -8409
rect -18595 -8484 -18513 -8473
rect -18595 -8544 -18584 -8484
rect -18524 -8544 -18513 -8484
rect -18595 -8555 -18513 -8544
rect -17756 -8504 -17747 -8418
rect -17656 -8504 -17647 -8418
rect -19237 -8695 -19223 -8629
rect -19152 -8695 -19142 -8629
rect -19457 -9221 -19293 -9198
rect -19457 -9301 -19423 -9221
rect -19325 -9301 -19293 -9221
rect -19457 -9328 -19293 -9301
rect -19237 -9409 -19142 -8695
rect -19065 -8824 -18791 -8815
rect -19065 -8896 -19056 -8824
rect -18800 -8896 -18791 -8824
rect -19065 -8905 -18791 -8896
rect -18348 -8824 -18074 -8815
rect -18348 -8896 -18339 -8824
rect -18083 -8896 -18074 -8824
rect -18348 -8905 -18074 -8896
rect -18047 -9209 -17869 -9158
rect -18047 -9289 -18002 -9209
rect -17882 -9289 -17869 -9209
rect -18047 -9306 -17869 -9289
rect -19457 -9424 -19142 -9409
rect -19457 -9484 -19433 -9424
rect -19248 -9484 -19142 -9424
rect -18573 -9375 -18398 -9364
rect -18573 -9450 -18561 -9375
rect -18416 -9450 -18398 -9375
rect -18573 -9462 -18398 -9450
rect -19457 -9494 -19142 -9484
rect -19044 -9575 -18960 -9563
rect -19044 -9637 -19033 -9575
rect -18971 -9637 -18960 -9575
rect -19044 -9648 -18960 -9637
rect -18179 -9600 -18101 -9589
rect -18179 -9656 -18168 -9600
rect -18112 -9656 -18101 -9600
rect -18179 -9667 -18101 -9656
rect -18047 -9705 -17927 -9306
rect -17756 -9606 -17647 -8504
rect -17482 -9393 -17381 -8228
rect -17274 -9193 -17178 -8017
rect -16165 -7939 -15893 -7923
rect -16165 -8036 -16081 -7939
rect -15931 -8036 -15893 -7939
rect -16165 -8071 -15893 -8036
rect -16863 -8484 -16781 -8473
rect -16863 -8544 -16852 -8484
rect -16792 -8544 -16781 -8484
rect -16863 -8555 -16781 -8544
rect -16460 -8633 -16329 -8617
rect -16460 -8702 -16444 -8633
rect -16345 -8702 -16329 -8633
rect -17063 -8824 -16789 -8815
rect -17063 -8896 -17054 -8824
rect -16798 -8896 -16789 -8824
rect -17063 -8905 -16789 -8896
rect -16701 -9159 -16592 -9144
rect -17275 -9220 -17111 -9193
rect -17275 -9300 -17243 -9220
rect -17145 -9300 -17111 -9220
rect -17275 -9328 -17111 -9300
rect -16701 -9307 -16688 -9159
rect -16605 -9307 -16592 -9159
rect -16701 -9319 -16592 -9307
rect -17482 -9413 -17111 -9393
rect -17482 -9479 -17452 -9413
rect -17199 -9479 -17111 -9413
rect -17482 -9492 -17111 -9479
rect -16987 -9566 -16634 -9557
rect -21055 -9852 -20730 -9726
rect -19751 -9807 -17927 -9705
rect -17763 -9728 -17429 -9606
rect -16987 -9622 -16978 -9566
rect -16643 -9622 -16634 -9566
rect -16987 -9631 -16634 -9622
rect -16460 -9705 -16329 -8702
rect -16165 -9198 -16069 -8071
rect -15946 -8127 -15740 -8101
rect -15946 -8224 -15905 -8127
rect -15789 -8224 -15740 -8127
rect -14465 -8107 -14356 -7211
rect -14290 -7094 -14166 -7011
rect -11174 -7026 -11065 -7011
rect -14067 -7092 -12857 -7064
rect -14290 -7864 -14176 -7094
rect -14067 -7164 -14021 -7092
rect -12899 -7164 -12857 -7092
rect -14067 -7190 -12857 -7164
rect -12508 -7092 -11298 -7064
rect -12508 -7164 -12462 -7092
rect -11340 -7164 -11298 -7092
rect -12508 -7190 -11298 -7164
rect -11174 -7170 -11165 -7026
rect -11074 -7170 -11065 -7026
rect -11004 -7070 -10876 -6628
rect -14290 -7887 -13887 -7864
rect -14290 -7995 -14266 -7887
rect -14176 -7995 -13887 -7887
rect -14290 -8017 -13887 -7995
rect -14290 -8018 -14176 -8017
rect -14465 -8108 -14108 -8107
rect -14465 -8120 -14079 -8108
rect -14465 -8220 -14169 -8120
rect -15946 -8244 -15740 -8224
rect -14191 -8228 -14169 -8220
rect -14093 -8228 -14079 -8120
rect -15946 -8629 -15851 -8244
rect -14465 -8418 -14356 -8409
rect -15304 -8484 -15222 -8473
rect -15304 -8544 -15293 -8484
rect -15233 -8544 -15222 -8484
rect -15304 -8555 -15222 -8544
rect -14465 -8504 -14456 -8418
rect -14365 -8504 -14356 -8418
rect -15946 -8695 -15932 -8629
rect -15861 -8695 -15851 -8629
rect -16166 -9221 -16002 -9198
rect -16166 -9301 -16132 -9221
rect -16034 -9301 -16002 -9221
rect -16166 -9328 -16002 -9301
rect -15946 -9409 -15851 -8695
rect -15774 -8824 -15500 -8815
rect -15774 -8896 -15765 -8824
rect -15509 -8896 -15500 -8824
rect -15774 -8905 -15500 -8896
rect -15057 -8824 -14783 -8815
rect -15057 -8896 -15048 -8824
rect -14792 -8896 -14783 -8824
rect -15057 -8905 -14783 -8896
rect -14756 -9209 -14578 -9158
rect -14756 -9289 -14711 -9209
rect -14591 -9289 -14578 -9209
rect -14756 -9306 -14578 -9289
rect -16166 -9424 -15851 -9409
rect -16166 -9484 -16142 -9424
rect -15957 -9484 -15851 -9424
rect -15282 -9375 -15107 -9364
rect -15282 -9450 -15270 -9375
rect -15125 -9450 -15107 -9375
rect -15282 -9462 -15107 -9450
rect -16166 -9494 -15851 -9484
rect -15753 -9575 -15669 -9563
rect -15753 -9637 -15742 -9575
rect -15680 -9637 -15669 -9575
rect -15753 -9648 -15669 -9637
rect -14888 -9600 -14810 -9589
rect -14888 -9656 -14877 -9600
rect -14821 -9656 -14810 -9600
rect -14888 -9667 -14810 -9656
rect -14756 -9705 -14636 -9306
rect -14465 -9618 -14356 -8504
rect -14191 -9393 -14090 -8228
rect -13983 -9193 -13887 -8017
rect -12874 -7939 -12602 -7923
rect -12874 -8036 -12790 -7939
rect -12640 -8036 -12602 -7939
rect -12874 -8071 -12602 -8036
rect -13572 -8484 -13490 -8473
rect -13572 -8544 -13561 -8484
rect -13501 -8544 -13490 -8484
rect -13572 -8555 -13490 -8544
rect -13169 -8633 -13038 -8617
rect -13169 -8702 -13153 -8633
rect -13054 -8702 -13038 -8633
rect -13772 -8824 -13498 -8815
rect -13772 -8896 -13763 -8824
rect -13507 -8896 -13498 -8824
rect -13772 -8905 -13498 -8896
rect -13410 -9159 -13301 -9144
rect -13984 -9220 -13820 -9193
rect -13984 -9300 -13952 -9220
rect -13854 -9300 -13820 -9220
rect -13984 -9328 -13820 -9300
rect -13410 -9307 -13397 -9159
rect -13314 -9307 -13301 -9159
rect -13410 -9319 -13301 -9307
rect -14191 -9413 -13820 -9393
rect -14191 -9479 -14161 -9413
rect -13908 -9479 -13820 -9413
rect -14191 -9492 -13820 -9479
rect -13696 -9566 -13343 -9557
rect -25990 -10155 -25880 -10146
rect -25305 -10155 -23050 -10101
rect -25990 -10160 -23050 -10155
rect -25990 -10241 -25978 -10160
rect -25899 -10236 -23050 -10160
rect -25899 -10241 -25048 -10236
rect -25990 -10244 -25048 -10241
rect -25990 -10252 -25880 -10244
rect -23583 -10566 -23369 -10544
rect -24397 -10668 -23763 -10634
rect -23583 -10645 -23560 -10566
rect -23391 -10645 -23369 -10566
rect -23583 -10664 -23369 -10645
rect -24397 -10808 -24359 -10668
rect -23805 -10808 -23763 -10668
rect -24397 -10847 -23763 -10808
rect -25369 -10976 -24837 -10970
rect -25374 -11055 -25365 -10976
rect -25286 -11055 -24837 -10976
rect -25369 -11059 -24837 -11055
rect -24748 -11059 -24742 -10970
rect -23185 -10997 -23050 -10236
rect -21850 -10566 -21636 -10544
rect -22660 -10668 -22026 -10634
rect -21850 -10645 -21827 -10566
rect -21658 -10645 -21636 -10566
rect -21850 -10664 -21636 -10645
rect -22660 -10808 -22622 -10668
rect -22068 -10808 -22026 -10668
rect -22660 -10847 -22026 -10808
rect -23210 -11007 -22577 -10997
rect -23210 -11121 -23198 -11007
rect -23061 -11019 -22577 -11007
rect -23061 -11113 -22832 -11019
rect -22650 -11113 -22577 -11019
rect -23061 -11121 -22577 -11113
rect -23210 -11123 -23195 -11121
rect -23064 -11123 -22577 -11121
rect -23210 -11132 -22577 -11123
rect -24632 -11187 -24269 -11161
rect -24632 -11278 -24563 -11187
rect -24335 -11278 -24269 -11187
rect -22910 -11179 -22591 -11161
rect -24632 -11297 -24269 -11278
rect -23583 -11219 -23383 -11191
rect -24632 -11556 -24456 -11297
rect -24162 -11324 -23762 -11296
rect -24162 -11398 -24133 -11324
rect -23793 -11398 -23762 -11324
rect -23583 -11315 -23556 -11219
rect -23407 -11315 -23383 -11219
rect -23583 -11341 -23383 -11315
rect -22910 -11275 -22848 -11179
rect -22644 -11275 -22591 -11179
rect -22910 -11297 -22591 -11275
rect -21850 -11219 -21650 -11191
rect -24162 -11419 -23762 -11398
rect -22910 -11556 -22734 -11297
rect -22425 -11324 -22025 -11296
rect -22425 -11398 -22396 -11324
rect -22056 -11398 -22025 -11324
rect -21850 -11315 -21823 -11219
rect -21674 -11315 -21650 -11219
rect -21047 -11285 -20938 -10275
rect -20875 -10373 -20745 -9852
rect -17756 -10292 -17647 -10275
rect -20649 -10356 -19439 -10328
rect -20872 -11128 -20758 -10373
rect -20649 -10428 -20603 -10356
rect -19481 -10428 -19439 -10356
rect -20649 -10454 -19439 -10428
rect -19090 -10356 -17880 -10328
rect -19090 -10428 -19044 -10356
rect -17922 -10428 -17880 -10356
rect -19090 -10454 -17880 -10428
rect -17756 -10387 -17744 -10292
rect -17655 -10387 -17647 -10292
rect -20872 -11151 -20469 -11128
rect -20872 -11259 -20848 -11151
rect -20758 -11259 -20469 -11151
rect -20872 -11281 -20469 -11259
rect -20872 -11282 -20758 -11281
rect -21356 -11292 -20938 -11285
rect -21850 -11341 -21650 -11315
rect -22425 -11419 -22025 -11398
rect -21395 -11371 -20938 -11292
rect -21395 -11372 -20690 -11371
rect -21395 -11384 -20661 -11372
rect -26164 -11586 -26102 -11582
rect -24634 -11586 -22734 -11556
rect -26169 -11591 -22734 -11586
rect -26169 -11653 -26164 -11591
rect -26102 -11653 -22734 -11591
rect -26169 -11658 -22734 -11653
rect -26164 -11662 -26102 -11658
rect -24634 -11691 -22734 -11658
rect -24632 -12289 -24456 -11691
rect -23583 -11858 -23369 -11836
rect -24397 -11960 -23763 -11926
rect -23583 -11937 -23560 -11858
rect -23391 -11937 -23369 -11858
rect -23583 -11956 -23369 -11937
rect -24397 -12100 -24359 -11960
rect -23805 -12100 -23763 -11960
rect -24397 -12139 -23763 -12100
rect -22910 -12289 -22734 -11691
rect -21395 -11425 -20751 -11384
rect -21854 -11858 -21640 -11836
rect -22660 -11960 -22026 -11926
rect -21854 -11937 -21831 -11858
rect -21662 -11937 -21640 -11858
rect -21854 -11956 -21640 -11937
rect -22660 -12100 -22622 -11960
rect -22068 -12100 -22026 -11960
rect -22660 -12139 -22026 -12100
rect -21562 -12234 -21477 -12232
rect -21395 -12234 -21304 -11425
rect -21047 -11484 -20751 -11425
rect -20773 -11492 -20751 -11484
rect -20675 -11492 -20661 -11384
rect -21610 -12276 -21304 -12234
rect -24632 -12313 -24325 -12289
rect -24632 -12400 -24570 -12313
rect -24353 -12400 -24325 -12313
rect -24632 -12424 -24325 -12400
rect -22910 -12316 -22637 -12289
rect -22910 -12408 -22868 -12316
rect -22670 -12408 -22637 -12316
rect -22910 -12424 -22637 -12408
rect -22911 -12460 -22572 -12454
rect -22912 -12472 -22572 -12460
rect -23583 -12511 -23383 -12483
rect -24637 -12578 -24439 -12549
rect -24637 -12776 -24612 -12578
rect -24466 -12776 -24439 -12578
rect -24162 -12616 -23762 -12588
rect -24162 -12690 -24133 -12616
rect -23793 -12690 -23762 -12616
rect -23583 -12607 -23556 -12511
rect -23407 -12607 -23383 -12511
rect -23583 -12633 -23383 -12607
rect -22912 -12503 -22730 -12472
rect -22912 -12518 -22866 -12503
rect -24162 -12711 -23762 -12690
rect -24637 -12791 -24439 -12776
rect -22912 -12964 -22869 -12518
rect -22777 -12524 -22730 -12503
rect -22773 -12560 -22730 -12524
rect -22611 -12560 -22572 -12472
rect -21610 -12462 -21554 -12276
rect -21355 -12462 -21304 -12276
rect -22773 -12589 -22572 -12560
rect -21854 -12511 -21654 -12483
rect -21610 -12497 -21304 -12462
rect -21039 -11862 -20854 -11846
rect -21039 -11964 -21003 -11862
rect -20885 -11964 -20854 -11862
rect -22773 -12868 -22736 -12589
rect -22425 -12616 -22025 -12588
rect -22425 -12690 -22396 -12616
rect -22056 -12690 -22025 -12616
rect -21854 -12607 -21827 -12511
rect -21678 -12607 -21654 -12511
rect -21854 -12633 -21654 -12607
rect -22425 -12711 -22025 -12690
rect -22912 -12970 -22862 -12964
rect -22773 -12970 -22737 -12868
rect -22912 -13014 -22737 -12970
rect -22912 -13016 -22744 -13014
rect -26340 -13054 -22744 -13016
rect -21039 -13050 -20854 -11964
rect -20773 -12657 -20672 -11492
rect -20565 -12457 -20469 -11281
rect -19456 -11203 -19184 -11187
rect -19456 -11300 -19372 -11203
rect -19222 -11300 -19184 -11203
rect -19456 -11335 -19184 -11300
rect -20154 -11748 -20072 -11737
rect -20154 -11808 -20143 -11748
rect -20083 -11808 -20072 -11748
rect -20154 -11819 -20072 -11808
rect -19751 -11897 -19620 -11881
rect -19751 -11966 -19735 -11897
rect -19636 -11966 -19620 -11897
rect -20354 -12088 -20080 -12079
rect -20354 -12160 -20345 -12088
rect -20089 -12160 -20080 -12088
rect -20354 -12169 -20080 -12160
rect -19992 -12423 -19883 -12408
rect -20566 -12484 -20402 -12457
rect -20566 -12564 -20534 -12484
rect -20436 -12564 -20402 -12484
rect -20566 -12592 -20402 -12564
rect -19992 -12571 -19979 -12423
rect -19896 -12571 -19883 -12423
rect -19992 -12583 -19883 -12571
rect -20773 -12677 -20402 -12657
rect -20773 -12743 -20743 -12677
rect -20490 -12743 -20402 -12677
rect -20773 -12756 -20402 -12743
rect -20278 -12830 -19925 -12821
rect -20278 -12886 -20269 -12830
rect -19934 -12886 -19925 -12830
rect -20278 -12895 -19925 -12886
rect -19751 -12969 -19620 -11966
rect -19456 -12462 -19360 -11335
rect -19237 -11391 -19031 -11365
rect -19237 -11488 -19196 -11391
rect -19080 -11488 -19031 -11391
rect -17756 -11371 -17647 -10387
rect -17588 -10392 -17452 -9728
rect -16460 -9807 -14636 -9705
rect -14474 -9763 -14158 -9618
rect -13696 -9622 -13687 -9566
rect -13352 -9622 -13343 -9566
rect -13696 -9631 -13343 -9622
rect -13169 -9705 -13038 -8702
rect -12874 -9198 -12778 -8071
rect -12655 -8127 -12449 -8101
rect -12655 -8224 -12614 -8127
rect -12498 -8224 -12449 -8127
rect -11174 -8107 -11065 -7170
rect -10999 -7864 -10885 -7070
rect -10776 -7092 -9566 -7064
rect -10776 -7164 -10730 -7092
rect -9608 -7164 -9566 -7092
rect -10776 -7190 -9566 -7164
rect -9217 -7092 -8007 -7064
rect -9217 -7164 -9171 -7092
rect -8049 -7164 -8007 -7092
rect -9217 -7190 -8007 -7164
rect -10999 -7887 -10596 -7864
rect -10999 -7995 -10975 -7887
rect -10885 -7995 -10596 -7887
rect -10999 -8017 -10596 -7995
rect -10999 -8018 -10885 -8017
rect -11174 -8108 -10817 -8107
rect -11174 -8120 -10788 -8108
rect -11174 -8220 -10878 -8120
rect -12655 -8244 -12449 -8224
rect -10900 -8228 -10878 -8220
rect -10802 -8228 -10788 -8120
rect -12655 -8629 -12560 -8244
rect -11174 -8418 -11065 -8409
rect -12013 -8484 -11931 -8473
rect -12013 -8544 -12002 -8484
rect -11942 -8544 -11931 -8484
rect -12013 -8555 -11931 -8544
rect -11174 -8504 -11165 -8418
rect -11074 -8504 -11065 -8418
rect -12655 -8695 -12641 -8629
rect -12570 -8695 -12560 -8629
rect -12875 -9221 -12711 -9198
rect -12875 -9301 -12841 -9221
rect -12743 -9301 -12711 -9221
rect -12875 -9328 -12711 -9301
rect -12655 -9409 -12560 -8695
rect -12483 -8824 -12209 -8815
rect -12483 -8896 -12474 -8824
rect -12218 -8896 -12209 -8824
rect -12483 -8905 -12209 -8896
rect -11766 -8824 -11492 -8815
rect -11766 -8896 -11757 -8824
rect -11501 -8896 -11492 -8824
rect -11766 -8905 -11492 -8896
rect -11465 -9209 -11287 -9158
rect -11465 -9289 -11420 -9209
rect -11300 -9289 -11287 -9209
rect -11465 -9306 -11287 -9289
rect -12875 -9424 -12560 -9409
rect -12875 -9484 -12851 -9424
rect -12666 -9484 -12560 -9424
rect -11991 -9375 -11816 -9364
rect -11991 -9450 -11979 -9375
rect -11834 -9450 -11816 -9375
rect -11991 -9462 -11816 -9450
rect -12875 -9494 -12560 -9484
rect -12462 -9575 -12378 -9563
rect -12462 -9637 -12451 -9575
rect -12389 -9637 -12378 -9575
rect -12462 -9648 -12378 -9637
rect -11597 -9600 -11519 -9589
rect -11597 -9656 -11586 -9600
rect -11530 -9656 -11519 -9600
rect -11597 -9667 -11519 -9656
rect -11465 -9705 -11345 -9306
rect -11174 -9600 -11065 -8504
rect -10900 -9393 -10799 -8228
rect -10692 -9193 -10596 -8017
rect -9583 -7939 -9311 -7923
rect -9583 -8036 -9499 -7939
rect -9349 -8036 -9311 -7939
rect -9583 -8071 -9311 -8036
rect -10281 -8484 -10199 -8473
rect -10281 -8544 -10270 -8484
rect -10210 -8544 -10199 -8484
rect -10281 -8555 -10199 -8544
rect -9878 -8633 -9747 -8617
rect -9878 -8702 -9862 -8633
rect -9763 -8702 -9747 -8633
rect -10481 -8824 -10207 -8815
rect -10481 -8896 -10472 -8824
rect -10216 -8896 -10207 -8824
rect -10481 -8905 -10207 -8896
rect -10119 -9159 -10010 -9144
rect -10693 -9220 -10529 -9193
rect -10693 -9300 -10661 -9220
rect -10563 -9300 -10529 -9220
rect -10693 -9328 -10529 -9300
rect -10119 -9307 -10106 -9159
rect -10023 -9307 -10010 -9159
rect -10119 -9319 -10010 -9307
rect -10900 -9413 -10529 -9393
rect -10900 -9479 -10870 -9413
rect -10617 -9479 -10529 -9413
rect -10900 -9492 -10529 -9479
rect -10405 -9566 -10052 -9557
rect -11174 -9646 -10879 -9600
rect -10405 -9622 -10396 -9566
rect -10061 -9622 -10052 -9566
rect -10405 -9631 -10052 -9622
rect -14465 -10291 -14356 -10275
rect -17358 -10356 -16148 -10328
rect -17581 -11128 -17467 -10392
rect -17358 -10428 -17312 -10356
rect -16190 -10428 -16148 -10356
rect -17358 -10454 -16148 -10428
rect -15799 -10356 -14589 -10328
rect -15799 -10428 -15753 -10356
rect -14631 -10428 -14589 -10356
rect -15799 -10454 -14589 -10428
rect -14465 -10475 -14460 -10291
rect -14361 -10475 -14356 -10291
rect -14300 -10420 -14170 -9763
rect -13169 -9807 -11345 -9705
rect -11170 -9736 -10879 -9646
rect -9878 -9705 -9747 -8702
rect -9583 -9198 -9487 -8071
rect -9364 -8127 -9158 -8101
rect -9364 -8224 -9323 -8127
rect -9207 -8224 -9158 -8127
rect -9364 -8244 -9158 -8224
rect -9364 -8629 -9269 -8244
rect -7883 -8418 -7774 -8409
rect -8722 -8484 -8640 -8473
rect -8722 -8544 -8711 -8484
rect -8651 -8544 -8640 -8484
rect -8722 -8555 -8640 -8544
rect -7883 -8504 -7874 -8418
rect -7783 -8504 -7774 -8418
rect -9364 -8695 -9350 -8629
rect -9279 -8695 -9269 -8629
rect -9584 -9221 -9420 -9198
rect -9584 -9301 -9550 -9221
rect -9452 -9301 -9420 -9221
rect -9584 -9328 -9420 -9301
rect -9364 -9409 -9269 -8695
rect -9192 -8824 -8918 -8815
rect -9192 -8896 -9183 -8824
rect -8927 -8896 -8918 -8824
rect -9192 -8905 -8918 -8896
rect -8475 -8824 -8201 -8815
rect -8475 -8896 -8466 -8824
rect -8210 -8896 -8201 -8824
rect -8475 -8905 -8201 -8896
rect -8174 -9209 -7996 -9158
rect -8174 -9289 -8129 -9209
rect -8009 -9289 -7996 -9209
rect -8174 -9306 -7996 -9289
rect -9584 -9424 -9269 -9409
rect -9584 -9484 -9560 -9424
rect -9375 -9484 -9269 -9424
rect -8700 -9375 -8525 -9364
rect -8700 -9450 -8688 -9375
rect -8543 -9450 -8525 -9375
rect -8700 -9462 -8525 -9450
rect -9584 -9494 -9269 -9484
rect -9171 -9575 -9087 -9563
rect -9171 -9637 -9160 -9575
rect -9098 -9637 -9087 -9575
rect -9171 -9648 -9087 -9637
rect -8306 -9600 -8228 -9589
rect -8306 -9656 -8295 -9600
rect -8239 -9656 -8228 -9600
rect -8306 -9667 -8228 -9656
rect -8174 -9705 -8054 -9306
rect -7883 -9527 -7774 -8504
rect -7888 -9534 -7756 -9527
rect -7888 -9645 -7688 -9534
rect -7883 -9646 -7774 -9645
rect -11174 -10290 -11065 -10275
rect -14067 -10356 -12857 -10328
rect -17581 -11151 -17178 -11128
rect -17581 -11259 -17557 -11151
rect -17467 -11259 -17178 -11151
rect -17581 -11281 -17178 -11259
rect -17581 -11282 -17467 -11281
rect -17756 -11372 -17399 -11371
rect -17756 -11384 -17370 -11372
rect -17756 -11484 -17460 -11384
rect -19237 -11508 -19031 -11488
rect -17482 -11492 -17460 -11484
rect -17384 -11492 -17370 -11384
rect -19237 -11893 -19142 -11508
rect -17756 -11682 -17647 -11673
rect -18595 -11748 -18513 -11737
rect -18595 -11808 -18584 -11748
rect -18524 -11808 -18513 -11748
rect -18595 -11819 -18513 -11808
rect -17756 -11768 -17747 -11682
rect -17656 -11768 -17647 -11682
rect -19237 -11959 -19223 -11893
rect -19152 -11959 -19142 -11893
rect -19457 -12485 -19293 -12462
rect -19457 -12565 -19423 -12485
rect -19325 -12565 -19293 -12485
rect -19457 -12592 -19293 -12565
rect -19237 -12673 -19142 -11959
rect -19065 -12088 -18791 -12079
rect -19065 -12160 -19056 -12088
rect -18800 -12160 -18791 -12088
rect -19065 -12169 -18791 -12160
rect -18348 -12088 -18074 -12079
rect -18348 -12160 -18339 -12088
rect -18083 -12160 -18074 -12088
rect -18348 -12169 -18074 -12160
rect -18047 -12473 -17869 -12422
rect -18047 -12553 -18002 -12473
rect -17882 -12553 -17869 -12473
rect -18047 -12570 -17869 -12553
rect -19457 -12688 -19142 -12673
rect -19457 -12748 -19433 -12688
rect -19248 -12748 -19142 -12688
rect -18573 -12639 -18398 -12628
rect -18573 -12714 -18561 -12639
rect -18416 -12714 -18398 -12639
rect -18573 -12726 -18398 -12714
rect -19457 -12758 -19142 -12748
rect -19044 -12839 -18960 -12827
rect -19044 -12901 -19033 -12839
rect -18971 -12901 -18960 -12839
rect -19044 -12912 -18960 -12901
rect -18179 -12864 -18101 -12853
rect -18179 -12920 -18168 -12864
rect -18112 -12920 -18101 -12864
rect -18179 -12931 -18101 -12920
rect -18047 -12969 -17927 -12570
rect -17756 -12910 -17647 -11768
rect -17482 -12657 -17381 -11492
rect -17274 -12457 -17178 -11281
rect -16165 -11203 -15893 -11187
rect -16165 -11300 -16081 -11203
rect -15931 -11300 -15893 -11203
rect -16165 -11335 -15893 -11300
rect -16863 -11748 -16781 -11737
rect -16863 -11808 -16852 -11748
rect -16792 -11808 -16781 -11748
rect -16863 -11819 -16781 -11808
rect -16460 -11897 -16329 -11881
rect -16460 -11966 -16444 -11897
rect -16345 -11966 -16329 -11897
rect -17063 -12088 -16789 -12079
rect -17063 -12160 -17054 -12088
rect -16798 -12160 -16789 -12088
rect -17063 -12169 -16789 -12160
rect -16701 -12423 -16592 -12408
rect -17275 -12484 -17111 -12457
rect -17275 -12564 -17243 -12484
rect -17145 -12564 -17111 -12484
rect -17275 -12592 -17111 -12564
rect -16701 -12571 -16688 -12423
rect -16605 -12571 -16592 -12423
rect -16701 -12583 -16592 -12571
rect -17482 -12677 -17111 -12657
rect -17482 -12743 -17452 -12677
rect -17199 -12743 -17111 -12677
rect -17482 -12756 -17111 -12743
rect -16987 -12830 -16634 -12821
rect -16987 -12886 -16978 -12830
rect -16643 -12886 -16634 -12830
rect -16987 -12895 -16634 -12886
rect -26340 -13063 -22742 -13054
rect -26340 -13144 -26327 -13063
rect -26248 -13144 -22742 -13063
rect -26340 -13184 -22742 -13144
rect -21025 -14475 -20959 -13050
rect -19751 -13071 -17927 -12969
rect -17730 -13700 -17671 -12910
rect -16460 -12969 -16329 -11966
rect -16165 -12462 -16069 -11335
rect -15946 -11391 -15740 -11365
rect -15946 -11488 -15905 -11391
rect -15789 -11488 -15740 -11391
rect -14465 -11371 -14356 -10475
rect -14290 -11128 -14176 -10420
rect -14067 -10428 -14021 -10356
rect -12899 -10428 -12857 -10356
rect -14067 -10454 -12857 -10428
rect -12508 -10356 -11298 -10328
rect -12508 -10428 -12462 -10356
rect -11340 -10428 -11298 -10356
rect -12508 -10454 -11298 -10428
rect -11174 -10434 -11165 -10290
rect -11074 -10434 -11065 -10290
rect -11004 -10392 -10880 -9736
rect -9878 -9807 -8054 -9705
rect -10776 -10356 -9566 -10328
rect -14290 -11151 -13887 -11128
rect -14290 -11259 -14266 -11151
rect -14176 -11259 -13887 -11151
rect -14290 -11281 -13887 -11259
rect -14290 -11282 -14176 -11281
rect -14465 -11372 -14108 -11371
rect -14465 -11384 -14079 -11372
rect -14465 -11484 -14169 -11384
rect -15946 -11508 -15740 -11488
rect -14191 -11492 -14169 -11484
rect -14093 -11492 -14079 -11384
rect -15946 -11893 -15851 -11508
rect -14465 -11682 -14356 -11673
rect -15304 -11748 -15222 -11737
rect -15304 -11808 -15293 -11748
rect -15233 -11808 -15222 -11748
rect -15304 -11819 -15222 -11808
rect -14465 -11768 -14456 -11682
rect -14365 -11768 -14356 -11682
rect -15946 -11959 -15932 -11893
rect -15861 -11959 -15851 -11893
rect -16166 -12485 -16002 -12462
rect -16166 -12565 -16132 -12485
rect -16034 -12565 -16002 -12485
rect -16166 -12592 -16002 -12565
rect -15946 -12673 -15851 -11959
rect -15774 -12088 -15500 -12079
rect -15774 -12160 -15765 -12088
rect -15509 -12160 -15500 -12088
rect -15774 -12169 -15500 -12160
rect -15057 -12088 -14783 -12079
rect -15057 -12160 -15048 -12088
rect -14792 -12160 -14783 -12088
rect -15057 -12169 -14783 -12160
rect -14756 -12473 -14578 -12422
rect -14756 -12553 -14711 -12473
rect -14591 -12553 -14578 -12473
rect -14756 -12570 -14578 -12553
rect -16166 -12688 -15851 -12673
rect -16166 -12748 -16142 -12688
rect -15957 -12748 -15851 -12688
rect -15282 -12639 -15107 -12628
rect -15282 -12714 -15270 -12639
rect -15125 -12714 -15107 -12639
rect -15282 -12726 -15107 -12714
rect -16166 -12758 -15851 -12748
rect -15753 -12839 -15669 -12827
rect -15753 -12901 -15742 -12839
rect -15680 -12901 -15669 -12839
rect -15753 -12912 -15669 -12901
rect -14888 -12864 -14810 -12853
rect -14888 -12920 -14877 -12864
rect -14821 -12920 -14810 -12864
rect -14888 -12931 -14810 -12920
rect -14756 -12969 -14636 -12570
rect -14465 -12910 -14356 -11768
rect -14191 -12657 -14090 -11492
rect -13983 -12457 -13887 -11281
rect -12874 -11203 -12602 -11187
rect -12874 -11300 -12790 -11203
rect -12640 -11300 -12602 -11203
rect -12874 -11335 -12602 -11300
rect -13572 -11748 -13490 -11737
rect -13572 -11808 -13561 -11748
rect -13501 -11808 -13490 -11748
rect -13572 -11819 -13490 -11808
rect -13169 -11897 -13038 -11881
rect -13169 -11966 -13153 -11897
rect -13054 -11966 -13038 -11897
rect -13772 -12088 -13498 -12079
rect -13772 -12160 -13763 -12088
rect -13507 -12160 -13498 -12088
rect -13772 -12169 -13498 -12160
rect -13410 -12423 -13301 -12408
rect -13984 -12484 -13820 -12457
rect -13984 -12564 -13952 -12484
rect -13854 -12564 -13820 -12484
rect -13984 -12592 -13820 -12564
rect -13410 -12571 -13397 -12423
rect -13314 -12571 -13301 -12423
rect -13410 -12583 -13301 -12571
rect -14191 -12677 -13820 -12657
rect -14191 -12743 -14161 -12677
rect -13908 -12743 -13820 -12677
rect -14191 -12756 -13820 -12743
rect -13696 -12830 -13343 -12821
rect -13696 -12886 -13687 -12830
rect -13352 -12886 -13343 -12830
rect -13696 -12895 -13343 -12886
rect -16460 -13071 -14636 -12969
rect -14443 -13577 -14377 -12910
rect -13169 -12969 -13038 -11966
rect -12874 -12462 -12778 -11335
rect -12655 -11391 -12449 -11365
rect -12655 -11488 -12614 -11391
rect -12498 -11488 -12449 -11391
rect -11174 -11371 -11065 -10434
rect -10999 -11128 -10885 -10392
rect -10776 -10428 -10730 -10356
rect -9608 -10428 -9566 -10356
rect -10776 -10454 -9566 -10428
rect -9217 -10356 -8007 -10328
rect -9217 -10428 -9171 -10356
rect -8049 -10428 -8007 -10356
rect -9217 -10454 -8007 -10428
rect -10999 -11151 -10596 -11128
rect -10999 -11259 -10975 -11151
rect -10885 -11259 -10596 -11151
rect -10999 -11281 -10596 -11259
rect -10999 -11282 -10885 -11281
rect -11174 -11372 -10817 -11371
rect -11174 -11384 -10788 -11372
rect -11174 -11484 -10878 -11384
rect -12655 -11508 -12449 -11488
rect -10900 -11492 -10878 -11484
rect -10802 -11492 -10788 -11384
rect -12655 -11893 -12560 -11508
rect -11174 -11682 -11065 -11673
rect -12013 -11748 -11931 -11737
rect -12013 -11808 -12002 -11748
rect -11942 -11808 -11931 -11748
rect -12013 -11819 -11931 -11808
rect -11174 -11768 -11165 -11682
rect -11074 -11768 -11065 -11682
rect -12655 -11959 -12641 -11893
rect -12570 -11959 -12560 -11893
rect -12875 -12485 -12711 -12462
rect -12875 -12565 -12841 -12485
rect -12743 -12565 -12711 -12485
rect -12875 -12592 -12711 -12565
rect -12655 -12673 -12560 -11959
rect -12483 -12088 -12209 -12079
rect -12483 -12160 -12474 -12088
rect -12218 -12160 -12209 -12088
rect -12483 -12169 -12209 -12160
rect -11766 -12088 -11492 -12079
rect -11766 -12160 -11757 -12088
rect -11501 -12160 -11492 -12088
rect -11766 -12169 -11492 -12160
rect -11465 -12473 -11287 -12422
rect -11465 -12553 -11420 -12473
rect -11300 -12553 -11287 -12473
rect -11465 -12570 -11287 -12553
rect -12875 -12688 -12560 -12673
rect -12875 -12748 -12851 -12688
rect -12666 -12748 -12560 -12688
rect -11991 -12639 -11816 -12628
rect -11991 -12714 -11979 -12639
rect -11834 -12714 -11816 -12639
rect -11991 -12726 -11816 -12714
rect -12875 -12758 -12560 -12748
rect -12462 -12839 -12378 -12827
rect -12462 -12901 -12451 -12839
rect -12389 -12901 -12378 -12839
rect -12462 -12912 -12378 -12901
rect -11597 -12864 -11519 -12853
rect -11597 -12920 -11586 -12864
rect -11530 -12920 -11519 -12864
rect -11597 -12931 -11519 -12920
rect -11465 -12969 -11345 -12570
rect -11174 -12910 -11065 -11768
rect -10900 -12657 -10799 -11492
rect -10692 -12457 -10596 -11281
rect -9583 -11203 -9311 -11187
rect -9583 -11300 -9499 -11203
rect -9349 -11300 -9311 -11203
rect -9583 -11335 -9311 -11300
rect -10281 -11748 -10199 -11737
rect -10281 -11808 -10270 -11748
rect -10210 -11808 -10199 -11748
rect -10281 -11819 -10199 -11808
rect -9878 -11897 -9747 -11881
rect -9878 -11966 -9862 -11897
rect -9763 -11966 -9747 -11897
rect -10481 -12088 -10207 -12079
rect -10481 -12160 -10472 -12088
rect -10216 -12160 -10207 -12088
rect -10481 -12169 -10207 -12160
rect -10119 -12423 -10010 -12408
rect -10693 -12484 -10529 -12457
rect -10693 -12564 -10661 -12484
rect -10563 -12564 -10529 -12484
rect -10693 -12592 -10529 -12564
rect -10119 -12571 -10106 -12423
rect -10023 -12571 -10010 -12423
rect -10119 -12583 -10010 -12571
rect -10900 -12677 -10529 -12657
rect -10900 -12743 -10870 -12677
rect -10617 -12743 -10529 -12677
rect -10900 -12756 -10529 -12743
rect -10405 -12830 -10052 -12821
rect -10405 -12886 -10396 -12830
rect -10061 -12886 -10052 -12830
rect -10405 -12895 -10052 -12886
rect -13169 -13071 -11345 -12969
rect -11151 -13379 -11085 -12910
rect -9878 -12969 -9747 -11966
rect -9583 -12462 -9487 -11335
rect -9364 -11391 -9158 -11365
rect -9364 -11488 -9323 -11391
rect -9207 -11488 -9158 -11391
rect -9364 -11508 -9158 -11488
rect -9364 -11893 -9269 -11508
rect -7883 -11682 -7774 -11673
rect -8722 -11748 -8640 -11737
rect -8722 -11808 -8711 -11748
rect -8651 -11808 -8640 -11748
rect -8722 -11819 -8640 -11808
rect -7883 -11768 -7874 -11682
rect -7783 -11768 -7774 -11682
rect -9364 -11959 -9350 -11893
rect -9279 -11959 -9269 -11893
rect -9584 -12485 -9420 -12462
rect -9584 -12565 -9550 -12485
rect -9452 -12565 -9420 -12485
rect -9584 -12592 -9420 -12565
rect -9364 -12673 -9269 -11959
rect -9192 -12088 -8918 -12079
rect -9192 -12160 -9183 -12088
rect -8927 -12160 -8918 -12088
rect -9192 -12169 -8918 -12160
rect -8475 -12088 -8201 -12079
rect -8475 -12160 -8466 -12088
rect -8210 -12160 -8201 -12088
rect -8475 -12169 -8201 -12160
rect -8174 -12473 -7996 -12422
rect -8174 -12553 -8129 -12473
rect -8009 -12553 -7996 -12473
rect -8174 -12570 -7996 -12553
rect -9584 -12688 -9269 -12673
rect -9584 -12748 -9560 -12688
rect -9375 -12748 -9269 -12688
rect -8700 -12639 -8525 -12628
rect -8700 -12714 -8688 -12639
rect -8543 -12714 -8525 -12639
rect -8700 -12726 -8525 -12714
rect -9584 -12758 -9269 -12748
rect -9171 -12839 -9087 -12827
rect -9171 -12901 -9160 -12839
rect -9098 -12901 -9087 -12839
rect -9171 -12912 -9087 -12901
rect -8306 -12864 -8228 -12853
rect -8306 -12920 -8295 -12864
rect -8239 -12920 -8228 -12864
rect -8306 -12931 -8228 -12920
rect -8174 -12969 -8054 -12570
rect -7883 -12791 -7774 -11768
rect -7888 -12798 -7756 -12791
rect -7888 -12909 -7799 -12798
rect -7688 -12909 -7682 -12798
rect -7883 -12910 -7774 -12909
rect -9878 -13071 -8054 -12969
rect -11151 -13451 -11085 -13445
rect -14443 -13649 -14377 -13643
rect -17730 -13765 -17671 -13759
rect -6334 -13840 -6286 -2274
rect 5732 -2277 7106 -2274
rect 7172 -2277 7178 -2211
rect 10536 -2214 10602 -1916
rect 8812 -2280 8818 -2214
rect 8884 -2280 10602 -2214
rect 10659 -2010 10850 -1944
rect 10915 -2010 10921 -1944
rect 5732 -2328 8050 -2315
rect -20148 -13888 -6286 -13840
rect -6254 -2376 8050 -2328
rect -21031 -14541 -21025 -14475
rect -20959 -14541 -20953 -14475
rect -23433 -15075 -23310 -15063
rect -23433 -15176 -23421 -15075
rect -23320 -15176 -23310 -15075
rect -24849 -15194 -24733 -15184
rect -23433 -15191 -23310 -15176
rect -24849 -15290 -24839 -15194
rect -24743 -15290 -24733 -15194
rect -24849 -15300 -24733 -15290
rect -24936 -15658 -24916 -15586
rect -24844 -15658 -24820 -15586
rect -24936 -15739 -24800 -15738
rect -24936 -15828 -24903 -15739
rect -24812 -15828 -24800 -15739
rect -23390 -16271 -23267 -16259
rect -24845 -16368 -24729 -16358
rect -24845 -16464 -24835 -16368
rect -24739 -16464 -24729 -16368
rect -23390 -16372 -23378 -16271
rect -23277 -16372 -23267 -16271
rect -23390 -16387 -23267 -16372
rect -24845 -16474 -24729 -16464
rect -24920 -16842 -24908 -16770
rect -24836 -16842 -24820 -16770
rect -24925 -16923 -24836 -16917
rect -24836 -17012 -24827 -16923
rect -24925 -17018 -24836 -17012
rect -23381 -17483 -23258 -17471
rect -23381 -17584 -23369 -17483
rect -23268 -17584 -23258 -17483
rect -24839 -17600 -24723 -17590
rect -23381 -17599 -23258 -17584
rect -24839 -17696 -24829 -17600
rect -24733 -17696 -24723 -17600
rect -24839 -17706 -24723 -17696
rect -20399 -17934 -20347 -17928
rect -24921 -17982 -24851 -17978
rect -24934 -17984 -24834 -17982
rect -24934 -18054 -24921 -17984
rect -24851 -18054 -24834 -17984
rect -20148 -17936 -20100 -13888
rect -14808 -13920 -14756 -13918
rect -6254 -13920 -6206 -2376
rect 5732 -2381 8050 -2376
rect 8116 -2381 8122 -2315
rect 10659 -2468 10725 -2010
rect 7866 -2534 7872 -2468
rect 7938 -2534 10725 -2468
rect 7156 -2813 11207 -2741
rect 7156 -2991 7227 -2813
rect 7405 -2991 8162 -2813
rect 8340 -2991 9098 -2813
rect 9276 -2990 10029 -2813
rect 10206 -2990 10956 -2813
rect 9276 -2991 10956 -2990
rect 11134 -2991 11207 -2813
rect 7156 -3062 11207 -2991
rect 12414 -3232 12821 -3120
rect 12128 -3236 12821 -3232
rect 7847 -3327 7853 -3261
rect 7919 -3327 10121 -3261
rect 5732 -3426 8989 -3417
rect -14808 -13924 -6206 -13920
rect -20347 -17984 -20100 -17936
rect -20070 -13988 -14888 -13940
rect -14756 -13968 -6206 -13924
rect -6160 -3483 8989 -3426
rect 9055 -3483 9061 -3417
rect -6160 -3486 6238 -3483
rect -14808 -13982 -14756 -13976
rect -20399 -17992 -20347 -17986
rect -24921 -18060 -24851 -18054
rect -20643 -18080 -20554 -18079
rect -20654 -18085 -20543 -18080
rect -21944 -18113 -21862 -18102
rect -24936 -18128 -24806 -18126
rect -24936 -18217 -24917 -18128
rect -24824 -18217 -24806 -18128
rect -21944 -18173 -21933 -18113
rect -21873 -18173 -21862 -18113
rect -21944 -18184 -21862 -18173
rect -20654 -18174 -20643 -18085
rect -20554 -18174 -20543 -18085
rect -20654 -18179 -20543 -18174
rect -20643 -18180 -20554 -18179
rect -24936 -18218 -24806 -18217
rect -20408 -18434 -20356 -18428
rect -20420 -18486 -20414 -18434
rect -20070 -18436 -20022 -13988
rect -14936 -14010 -14888 -13988
rect -20356 -18484 -20022 -18436
rect -19958 -14084 -14970 -14036
rect -14936 -14058 -10918 -14010
rect -6160 -14032 -6100 -3486
rect -6062 -3539 5820 -3536
rect 10055 -3539 10121 -3327
rect 12128 -3262 13042 -3236
rect 12128 -3324 13186 -3262
rect 12128 -3443 12233 -3324
rect 12352 -3365 13186 -3324
rect 12352 -3443 12960 -3365
rect 12128 -3484 12960 -3443
rect 13079 -3484 13186 -3365
rect -6062 -3584 9917 -3539
rect -20408 -18492 -20356 -18486
rect -20650 -18573 -20561 -18572
rect -20661 -18578 -20550 -18573
rect -23373 -18624 -23250 -18612
rect -24825 -18714 -24709 -18704
rect -24825 -18810 -24815 -18714
rect -24719 -18810 -24709 -18714
rect -23373 -18725 -23361 -18624
rect -23260 -18725 -23250 -18624
rect -21950 -18622 -21868 -18611
rect -21950 -18682 -21939 -18622
rect -21879 -18682 -21868 -18622
rect -20661 -18667 -20650 -18578
rect -20561 -18667 -20550 -18578
rect -20661 -18672 -20550 -18667
rect -20650 -18673 -20561 -18672
rect -21950 -18693 -21868 -18682
rect -23373 -18740 -23250 -18725
rect -24825 -18820 -24709 -18810
rect -20406 -18914 -20340 -18908
rect -20406 -18966 -20399 -18914
rect -20347 -18916 -20340 -18914
rect -19958 -18916 -19910 -14084
rect -15018 -14170 -14970 -14084
rect -14714 -14140 -14708 -14088
rect -14656 -14090 -14650 -14088
rect -14656 -14138 -11022 -14090
rect -14656 -14140 -14650 -14138
rect -15018 -14218 -12652 -14170
rect -18084 -15281 -17986 -15269
rect -18084 -15355 -18072 -15281
rect -17998 -15355 -17986 -15281
rect -18084 -15367 -17986 -15355
rect -16924 -15326 -16836 -15311
rect -16924 -15386 -16909 -15326
rect -16849 -15386 -16836 -15326
rect -16924 -15401 -16836 -15386
rect -12700 -15454 -12652 -14218
rect -12501 -14223 -12375 -14181
rect -12501 -15345 -12473 -14223
rect -12401 -15345 -12375 -14223
rect -11070 -14250 -11022 -14138
rect -10966 -14152 -10918 -14058
rect -10861 -14108 -10855 -14032
rect -10779 -14108 -6092 -14032
rect -6062 -14136 -6014 -3584
rect 5732 -3605 9917 -3584
rect 9983 -3605 9989 -3539
rect 10055 -3605 10704 -3539
rect 12128 -3549 13186 -3484
rect -5959 -3703 7102 -3637
rect 7168 -3703 7174 -3637
rect -5959 -3793 -5893 -3703
rect 8831 -3737 8837 -3671
rect 8903 -3737 10588 -3671
rect -5963 -13983 -5881 -3793
rect -5799 -3824 8050 -3758
rect 8116 -3824 8122 -3758
rect -5799 -4072 -5733 -3824
rect 9801 -3829 9807 -3765
rect 9873 -3829 10453 -3765
rect 8396 -3860 8470 -3854
rect 6780 -3879 6849 -3873
rect 6849 -3932 8206 -3893
rect 8396 -3895 8405 -3860
rect 8461 -3895 8470 -3860
rect 8396 -3924 8401 -3895
rect 6780 -3954 6849 -3948
rect 6066 -3982 6132 -3976
rect 6132 -3991 8139 -3982
rect 6132 -4043 8079 -3991
rect 8131 -4043 8139 -3991
rect 8167 -4001 8206 -3932
rect 8465 -3924 8470 -3895
rect 8615 -3954 8993 -3888
rect 9059 -3954 9065 -3888
rect 10264 -3895 10324 -3889
rect 10257 -3953 10264 -3897
rect 10324 -3953 10331 -3897
rect 8401 -3965 8465 -3959
rect 8616 -4001 8655 -3954
rect 10264 -3961 10324 -3955
rect 8167 -4040 8655 -4001
rect 6132 -4048 8139 -4043
rect 8992 -4048 9001 -3982
rect 9067 -4048 9076 -3982
rect 9931 -4047 9937 -3981
rect 10003 -4047 10012 -3981
rect 10387 -3982 10453 -3829
rect 10522 -3888 10588 -3737
rect 10638 -3794 10704 -3605
rect 12467 -3708 13186 -3549
rect 12796 -3741 13186 -3708
rect 10638 -3860 10850 -3794
rect 10916 -3860 10922 -3794
rect 10522 -3954 10888 -3888
rect 10954 -3954 10963 -3888
rect 10387 -4048 10859 -3982
rect 10925 -4048 10931 -3982
rect 6066 -4054 6132 -4048
rect -5814 -13408 -5730 -4072
rect 6934 -4142 6941 -4076
rect 7007 -4085 10062 -4076
rect 7007 -4137 8063 -4085
rect 8128 -4137 8992 -4085
rect 9057 -4137 9951 -4085
rect 10016 -4137 10062 -4085
rect 7007 -4142 10062 -4137
rect 6941 -4148 7007 -4142
rect 11883 -4361 12147 -4350
rect 11883 -4603 11894 -4361
rect 12136 -4603 12147 -4361
rect 11883 -4614 12147 -4603
rect 5558 -4860 5627 -4828
rect 5554 -4919 5563 -4860
rect 5622 -4919 5631 -4860
rect 5998 -4880 6067 -4828
rect 5558 -5077 5627 -4919
rect 5994 -4939 6003 -4880
rect 6062 -4939 6071 -4880
rect 6438 -4889 6507 -4828
rect 5998 -5077 6067 -4939
rect 6433 -4948 6442 -4889
rect 6501 -4948 6510 -4889
rect 6438 -5077 6507 -4948
rect 5552 -5146 5558 -5077
rect 5627 -5146 5633 -5077
rect 5992 -5146 5998 -5077
rect 6067 -5146 6073 -5077
rect 6432 -5146 6438 -5077
rect 6507 -5146 6513 -5077
rect 5901 -5531 7113 -5462
rect 5901 -5642 5970 -5531
rect 5703 -5726 5823 -5698
rect 5901 -5717 5970 -5711
rect 6158 -5707 6236 -5697
rect 5703 -5782 5732 -5726
rect 5788 -5782 5823 -5726
rect 6158 -5763 6170 -5707
rect 6226 -5763 6236 -5707
rect 6335 -5713 6341 -5644
rect 6410 -5713 6416 -5644
rect 6580 -5698 6700 -5682
rect 6158 -5778 6236 -5763
rect 5703 -5811 5823 -5782
rect 6341 -5923 6410 -5713
rect 6580 -5754 6610 -5698
rect 6666 -5754 6700 -5698
rect 6580 -5795 6700 -5754
rect 6299 -5982 6410 -5923
rect 6299 -6081 6367 -5982
rect 6295 -6139 6304 -6081
rect 6362 -6139 6371 -6081
rect 7044 -6086 7113 -5531
rect 7044 -6095 10140 -6086
rect 6299 -6144 6367 -6139
rect 7044 -6147 7106 -6095
rect 7158 -6096 9002 -6095
rect 7158 -6147 8069 -6096
rect 7044 -6148 8069 -6147
rect 8122 -6147 9002 -6096
rect 9055 -6147 9933 -6095
rect 9986 -6147 10140 -6095
rect 8122 -6148 10140 -6147
rect 7044 -6155 10140 -6148
rect 12187 -6087 12431 -6076
rect 12187 -6095 12198 -6087
rect 5992 -6181 6073 -6175
rect 5992 -6250 5998 -6181
rect 6067 -6186 6073 -6181
rect 6067 -6188 8115 -6186
rect 6067 -6189 8057 -6188
rect 6067 -6241 7113 -6189
rect 7165 -6240 8057 -6189
rect 8109 -6240 8115 -6188
rect 7165 -6241 8115 -6240
rect 6067 -6245 8115 -6241
rect 8182 -6236 8914 -6183
rect 9929 -6189 10000 -6187
rect 6067 -6250 6073 -6245
rect 5992 -6256 6073 -6250
rect 7321 -6278 7393 -6273
rect 8182 -6278 8248 -6236
rect 6429 -6316 6516 -6307
rect 6429 -6385 6438 -6316
rect 6507 -6385 6516 -6316
rect 7321 -6344 7327 -6278
rect 7393 -6344 8248 -6278
rect 8424 -6271 8493 -6265
rect 8861 -6284 8914 -6236
rect 8989 -6247 8998 -6191
rect 9054 -6247 9063 -6191
rect 9923 -6245 9935 -6189
rect 9991 -6245 10000 -6189
rect 10256 -6240 10336 -6234
rect 9929 -6251 9993 -6245
rect 8541 -6316 8600 -6312
rect 8493 -6321 8605 -6316
rect 8493 -6323 8541 -6321
rect 7321 -6350 7393 -6344
rect 8424 -6380 8541 -6323
rect 8600 -6380 8605 -6321
rect 8861 -6337 8989 -6284
rect 9042 -6337 9048 -6284
rect 10256 -6309 10262 -6240
rect 10331 -6309 10336 -6240
rect 10256 -6316 10336 -6309
rect 10405 -6250 10860 -6184
rect 10926 -6250 10932 -6184
rect 8424 -6385 8605 -6380
rect 6429 -6394 6516 -6385
rect 8541 -6389 8600 -6385
rect 10405 -6394 10471 -6250
rect 5419 -6432 5485 -6431
rect 5412 -6437 5485 -6432
rect 5412 -6503 5419 -6437
rect 5485 -6503 8986 -6437
rect 9052 -6503 9058 -6437
rect 9792 -6460 9798 -6394
rect 9864 -6460 10471 -6394
rect 10536 -6344 10858 -6278
rect 10924 -6344 10930 -6278
rect 12187 -6298 12189 -6095
rect 12187 -6309 12198 -6298
rect 12420 -6309 12441 -6087
rect 12187 -6320 12431 -6309
rect 5412 -6504 5485 -6503
rect -5445 -6599 -5439 -6533
rect -5373 -6599 9917 -6533
rect 9983 -6599 9989 -6533
rect -5694 -6639 -5646 -6638
rect -5694 -6705 7106 -6639
rect 7172 -6705 7178 -6639
rect 10536 -6642 10602 -6344
rect -5820 -13492 -5814 -13408
rect -5730 -13492 -5724 -13408
rect -5963 -14071 -5881 -14065
rect -6958 -14142 -6014 -14136
rect -10966 -14200 -7014 -14152
rect -6960 -14194 -6954 -14142
rect -6902 -14184 -6014 -14142
rect -6902 -14194 -6896 -14184
rect -7062 -14232 -7014 -14200
rect -5694 -14232 -5646 -6705
rect 8812 -6708 8818 -6642
rect 8884 -6708 10602 -6642
rect 10659 -6438 10850 -6372
rect 10915 -6438 10921 -6372
rect -5615 -6766 8050 -6743
rect -11070 -14298 -7108 -14250
rect -7062 -14280 -5646 -14232
rect -5616 -6809 8050 -6766
rect 8116 -6809 8122 -6743
rect -7156 -14314 -7108 -14298
rect -5616 -14314 -5568 -6809
rect 10659 -6896 10725 -6438
rect 7866 -6962 7872 -6896
rect 7938 -6962 10725 -6896
rect 7156 -7241 11207 -7169
rect 7156 -7419 7227 -7241
rect 7405 -7419 8162 -7241
rect 8340 -7419 9098 -7241
rect 9276 -7418 10029 -7241
rect 10206 -7418 10956 -7241
rect 9276 -7419 10956 -7418
rect 11134 -7419 11207 -7241
rect 7156 -7490 11207 -7419
rect 12414 -7660 12821 -7548
rect 12128 -7664 12821 -7660
rect 7847 -7755 7853 -7689
rect 7919 -7755 10121 -7689
rect -5507 -7847 8989 -7845
rect -10856 -14386 -10850 -14331
rect -10795 -14386 -7187 -14331
rect -7156 -14362 -5568 -14314
rect -5536 -7911 8989 -7847
rect 9055 -7911 9061 -7845
rect -7242 -14402 -7187 -14386
rect -5536 -14402 -5481 -7911
rect 10055 -7967 10121 -7755
rect 12128 -7690 13042 -7664
rect 12128 -7752 13186 -7690
rect 12128 -7871 12233 -7752
rect 12352 -7793 13186 -7752
rect 12352 -7871 12960 -7793
rect 12128 -7912 12960 -7871
rect 13079 -7912 13186 -7793
rect -5451 -8033 9917 -7967
rect 9983 -8033 9989 -7967
rect 10055 -8033 10704 -7967
rect 12128 -7977 13186 -7912
rect -12501 -15391 -12375 -15345
rect -12114 -14474 -7308 -14426
rect -7242 -14457 -5481 -14402
rect -12114 -15454 -12066 -14474
rect -7356 -14586 -7308 -14474
rect -5450 -14490 -5398 -8033
rect -5367 -8131 7102 -8065
rect 7168 -8131 7174 -8065
rect -5366 -13870 -5322 -8131
rect 8831 -8165 8837 -8099
rect 8903 -8165 10588 -8099
rect -5286 -8186 -5233 -8180
rect -5286 -8252 8050 -8186
rect 8116 -8252 8122 -8186
rect -5286 -13259 -5233 -8252
rect 9801 -8257 9807 -8193
rect 9873 -8257 10453 -8193
rect 8396 -8288 8470 -8282
rect 6780 -8307 6849 -8301
rect 6849 -8360 8206 -8321
rect 8396 -8323 8405 -8288
rect 8461 -8323 8470 -8288
rect 8396 -8352 8401 -8323
rect 6780 -8382 6849 -8376
rect 6066 -8410 6132 -8404
rect 6132 -8419 8139 -8410
rect 6132 -8471 8079 -8419
rect 8131 -8471 8139 -8419
rect 8167 -8429 8206 -8360
rect 8465 -8352 8470 -8323
rect 8615 -8382 8993 -8316
rect 9059 -8382 9065 -8316
rect 10264 -8323 10324 -8317
rect 10257 -8381 10264 -8325
rect 10324 -8381 10331 -8325
rect 8401 -8393 8465 -8387
rect 8616 -8429 8655 -8382
rect 10264 -8389 10324 -8383
rect 8167 -8468 8655 -8429
rect 6132 -8476 8139 -8471
rect 8992 -8476 9001 -8410
rect 9067 -8476 9076 -8410
rect 9931 -8475 9937 -8409
rect 10003 -8475 10012 -8409
rect 10387 -8410 10453 -8257
rect 10522 -8316 10588 -8165
rect 10638 -8222 10704 -8033
rect 12467 -8136 13186 -7977
rect 12796 -8169 13186 -8136
rect 10638 -8288 10850 -8222
rect 10916 -8288 10922 -8222
rect 10522 -8382 10888 -8316
rect 10954 -8382 10963 -8316
rect 10387 -8476 10859 -8410
rect 10925 -8476 10931 -8410
rect 6066 -8482 6132 -8476
rect 6934 -8570 6941 -8504
rect 7007 -8513 10062 -8504
rect 7007 -8565 8063 -8513
rect 8128 -8565 8992 -8513
rect 9057 -8565 9951 -8513
rect 10016 -8565 10062 -8513
rect 7007 -8570 10062 -8565
rect 6941 -8576 7007 -8570
rect 11883 -8789 12147 -8778
rect 11883 -9031 11894 -8789
rect 12136 -9031 12147 -8789
rect 11883 -9042 12147 -9031
rect 5558 -9523 5627 -9456
rect 5554 -9582 5563 -9523
rect 5622 -9582 5631 -9523
rect 5998 -9528 6067 -9456
rect 6438 -9514 6507 -9456
rect 5558 -9705 5627 -9582
rect 5994 -9587 6003 -9528
rect 6062 -9587 6071 -9528
rect 6436 -9573 6445 -9514
rect 6504 -9573 6513 -9514
rect 5998 -9705 6067 -9587
rect 6438 -9705 6507 -9573
rect 5552 -9774 5558 -9705
rect 5627 -9774 5633 -9705
rect 5992 -9774 5998 -9705
rect 6067 -9774 6073 -9705
rect 6432 -9774 6438 -9705
rect 6507 -9774 6513 -9705
rect 5901 -10159 7113 -10090
rect 5901 -10270 5970 -10159
rect 5703 -10354 5823 -10326
rect 5901 -10345 5970 -10339
rect 6158 -10335 6236 -10325
rect 5703 -10410 5732 -10354
rect 5788 -10410 5823 -10354
rect 6158 -10391 6170 -10335
rect 6226 -10391 6236 -10335
rect 6335 -10341 6341 -10272
rect 6410 -10341 6416 -10272
rect 6580 -10326 6700 -10310
rect 6158 -10406 6236 -10391
rect 5703 -10439 5823 -10410
rect 6341 -10551 6410 -10341
rect 6580 -10382 6610 -10326
rect 6666 -10382 6700 -10326
rect 6580 -10423 6700 -10382
rect 6299 -10610 6410 -10551
rect 6299 -10709 6367 -10610
rect 6295 -10767 6304 -10709
rect 6362 -10767 6371 -10709
rect 7044 -10714 7113 -10159
rect 7044 -10723 10140 -10714
rect 6299 -10772 6367 -10767
rect 7044 -10775 7106 -10723
rect 7158 -10724 9002 -10723
rect 7158 -10775 8069 -10724
rect 7044 -10776 8069 -10775
rect 8122 -10775 9002 -10724
rect 9055 -10775 9933 -10723
rect 9986 -10775 10140 -10723
rect 8122 -10776 10140 -10775
rect 7044 -10783 10140 -10776
rect 12187 -10715 12431 -10704
rect 12187 -10723 12198 -10715
rect 5992 -10809 6073 -10803
rect 5992 -10878 5998 -10809
rect 6067 -10814 6073 -10809
rect 6067 -10816 8115 -10814
rect 6067 -10817 8057 -10816
rect 6067 -10869 7113 -10817
rect 7165 -10868 8057 -10817
rect 8109 -10868 8115 -10816
rect 7165 -10869 8115 -10868
rect 6067 -10873 8115 -10869
rect 8182 -10864 8914 -10811
rect 9929 -10817 10000 -10815
rect 6067 -10878 6073 -10873
rect 5992 -10884 6073 -10878
rect 7321 -10906 7393 -10901
rect 8182 -10906 8248 -10864
rect 6429 -10944 6516 -10935
rect 6429 -11013 6438 -10944
rect 6507 -11013 6516 -10944
rect 7321 -10972 7327 -10906
rect 7393 -10972 8248 -10906
rect 8424 -10899 8493 -10893
rect 8861 -10912 8914 -10864
rect 8989 -10875 8998 -10819
rect 9054 -10875 9063 -10819
rect 9923 -10873 9935 -10817
rect 9991 -10873 10000 -10817
rect 10256 -10868 10336 -10862
rect 9929 -10879 9993 -10873
rect 8541 -10944 8600 -10940
rect 8493 -10949 8605 -10944
rect 8493 -10951 8541 -10949
rect 7321 -10978 7393 -10972
rect 8424 -11008 8541 -10951
rect 8600 -11008 8605 -10949
rect 8861 -10965 8989 -10912
rect 9042 -10965 9048 -10912
rect 10256 -10937 10262 -10868
rect 10331 -10937 10336 -10868
rect 10256 -10944 10336 -10937
rect 10405 -10878 10860 -10812
rect 10926 -10878 10932 -10812
rect 8424 -11013 8605 -11008
rect 6429 -11022 6516 -11013
rect 8541 -11017 8600 -11013
rect 10405 -11022 10471 -10878
rect 5420 -11131 5426 -11065
rect 5492 -11131 8986 -11065
rect 9052 -11131 9058 -11065
rect 9792 -11088 9798 -11022
rect 9864 -11088 10471 -11022
rect 10536 -10972 10858 -10906
rect 10924 -10972 10930 -10906
rect 12187 -10926 12189 -10723
rect 12187 -10937 12198 -10926
rect 12420 -10937 12441 -10715
rect 12187 -10948 12431 -10937
rect -5049 -11227 -5043 -11161
rect -4977 -11227 9917 -11161
rect 9983 -11227 9989 -11161
rect -5195 -11276 7106 -11267
rect -5286 -13318 -5233 -13312
rect -5200 -11333 7106 -11276
rect 7172 -11333 7178 -11267
rect 10536 -11270 10602 -10972
rect -5200 -13382 -5152 -11333
rect 8812 -11336 8818 -11270
rect 8884 -11336 10602 -11270
rect 10659 -11066 10850 -11000
rect 10915 -11066 10921 -11000
rect -5115 -11379 8050 -11371
rect -5284 -13430 -5152 -13382
rect -5116 -11437 8050 -11379
rect 8116 -11437 8122 -11371
rect -5370 -13876 -5318 -13870
rect -5370 -13934 -5318 -13928
rect -5284 -13988 -5236 -13430
rect -5116 -13469 -5061 -11437
rect 10659 -11524 10725 -11066
rect 7866 -11590 7872 -11524
rect 7938 -11590 10725 -11524
rect 7156 -11869 11207 -11797
rect 7156 -12047 7227 -11869
rect 7405 -12047 8162 -11869
rect 8340 -12047 9098 -11869
rect 9276 -12046 10029 -11869
rect 10206 -12046 10956 -11869
rect 9276 -12047 10956 -12046
rect 11134 -12047 11207 -11869
rect 7156 -12118 11207 -12047
rect 12414 -12288 12821 -12176
rect 12128 -12292 12821 -12288
rect 7847 -12383 7853 -12317
rect 7919 -12383 10121 -12317
rect -6840 -14542 -6834 -14490
rect -6782 -14542 -5398 -14490
rect -5368 -14036 -5236 -13988
rect -5196 -13524 -5061 -13469
rect -5022 -12473 -4974 -12472
rect -5022 -12539 8989 -12473
rect 9055 -12539 9061 -12473
rect -5368 -14586 -5320 -14036
rect -5196 -14083 -5141 -13524
rect -5022 -13566 -4974 -12539
rect -7356 -14634 -5320 -14586
rect -5284 -14138 -5141 -14083
rect -5108 -13614 -4974 -13566
rect -4796 -12595 -4748 -12592
rect 10055 -12595 10121 -12383
rect 12128 -12318 13042 -12292
rect 12128 -12380 13186 -12318
rect 12128 -12499 12233 -12380
rect 12352 -12421 13186 -12380
rect 12352 -12499 12960 -12421
rect 12128 -12540 12960 -12499
rect 13079 -12540 13186 -12421
rect -4796 -12661 9917 -12595
rect 9983 -12661 9989 -12595
rect 10055 -12661 10704 -12595
rect 12128 -12605 13186 -12540
rect -5284 -14685 -5229 -14138
rect -5108 -14180 -5060 -13614
rect -10150 -14690 -5229 -14685
rect -10606 -14738 -5229 -14690
rect -11092 -14825 -11010 -14814
rect -11092 -14885 -11081 -14825
rect -11021 -14885 -11010 -14825
rect -11092 -14896 -11010 -14885
rect -12700 -15502 -12066 -15454
rect -17978 -15586 -17880 -15576
rect -17978 -15658 -17966 -15586
rect -17894 -15658 -17880 -15586
rect -17978 -15666 -17880 -15658
rect -12734 -15586 -12608 -15552
rect -12734 -15658 -12724 -15586
rect -12652 -15658 -12608 -15586
rect -12734 -15672 -12608 -15658
rect -18130 -15738 -18026 -15730
rect -18130 -15827 -18123 -15738
rect -18034 -15827 -18026 -15738
rect -18130 -15836 -18026 -15827
rect -12566 -15738 -12440 -15728
rect -12566 -15837 -12555 -15738
rect -12456 -15837 -12440 -15738
rect -12566 -15848 -12440 -15837
rect -14612 -15964 -14560 -15958
rect -10606 -15966 -10558 -14738
rect -10150 -14740 -5229 -14738
rect -5194 -14228 -5060 -14180
rect -10313 -14826 -10307 -14771
rect -10252 -14778 -6429 -14771
rect -5194 -14778 -5146 -14228
rect -5026 -14254 -4910 -14248
rect -5026 -14376 -4910 -14370
rect -5020 -14494 -4926 -14484
rect -5020 -14566 -5008 -14494
rect -4936 -14566 -4926 -14494
rect -5020 -14576 -4926 -14566
rect -4796 -14726 -4748 -12661
rect -4633 -12759 7102 -12693
rect 7168 -12759 7174 -12693
rect -4626 -13734 -4542 -12759
rect 8831 -12793 8837 -12727
rect 8903 -12793 10588 -12727
rect 5732 -12818 8050 -12814
rect -774 -12902 -768 -12818
rect -684 -12880 8050 -12818
rect 8116 -12880 8122 -12814
rect -684 -12902 5792 -12880
rect 9801 -12885 9807 -12821
rect 9873 -12885 10453 -12821
rect 8396 -12916 8470 -12910
rect 6780 -12935 6849 -12929
rect 6849 -12988 8206 -12949
rect 8396 -12951 8405 -12916
rect 8461 -12951 8470 -12916
rect 8396 -12980 8401 -12951
rect 6780 -13010 6849 -13004
rect 6066 -13038 6132 -13032
rect 5354 -13052 5420 -13046
rect 6132 -13047 8139 -13038
rect 6132 -13099 8079 -13047
rect 8131 -13099 8139 -13047
rect 8167 -13057 8206 -12988
rect 8465 -12980 8470 -12951
rect 8615 -13010 8993 -12944
rect 9059 -13010 9065 -12944
rect 10264 -12951 10324 -12945
rect 10257 -13009 10264 -12953
rect 10324 -13009 10331 -12953
rect 8401 -13021 8465 -13015
rect 8616 -13057 8655 -13010
rect 10264 -13017 10324 -13011
rect 8167 -13096 8655 -13057
rect 6132 -13104 8139 -13099
rect 8992 -13104 9001 -13038
rect 9067 -13104 9076 -13038
rect 9931 -13103 9937 -13037
rect 10003 -13103 10012 -13037
rect 10387 -13038 10453 -12885
rect 10522 -12944 10588 -12793
rect 10638 -12850 10704 -12661
rect 12467 -12764 13186 -12605
rect 12796 -12797 13186 -12764
rect 10638 -12916 10850 -12850
rect 10916 -12916 10922 -12850
rect 10522 -13010 10888 -12944
rect 10954 -13010 10963 -12944
rect 10387 -13104 10859 -13038
rect 10925 -13104 10931 -13038
rect 6066 -13110 6132 -13104
rect 4164 -13666 4248 -13660
rect -1207 -13750 -1201 -13666
rect -1117 -13750 4164 -13666
rect 4164 -13756 4248 -13750
rect -4626 -13824 -4542 -13818
rect -2304 -14063 -2200 -14054
rect -2304 -14176 -2200 -14167
rect -1288 -14074 -1191 -14065
rect -1288 -14180 -1191 -14171
rect -4004 -14250 -3907 -14241
rect -4004 -14356 -3907 -14347
rect -3912 -14491 -3812 -14472
rect -3912 -14557 -3899 -14491
rect -3833 -14557 -3812 -14491
rect -3912 -14574 -3812 -14557
rect -2296 -14494 -2202 -14482
rect -2296 -14566 -2288 -14494
rect -2216 -14566 -2202 -14494
rect -2296 -14574 -2202 -14566
rect -10252 -14826 -5146 -14778
rect -5110 -14774 -4748 -14726
rect -6674 -14870 -6600 -14860
rect -6674 -14922 -6664 -14870
rect -6612 -14872 -6600 -14870
rect -5110 -14872 -5062 -14774
rect -6612 -14920 -5062 -14872
rect -5020 -14887 -4916 -14878
rect -6612 -14922 -6600 -14920
rect -6674 -14930 -6600 -14922
rect -4004 -14883 -3907 -14874
rect -4004 -14989 -3907 -14980
rect -2304 -14882 -2200 -14873
rect -5020 -15000 -4916 -14991
rect -2304 -14995 -2200 -14986
rect -1288 -14893 -1191 -14884
rect -1288 -14999 -1191 -14990
rect -4974 -15306 -4880 -15294
rect -7204 -15392 -7115 -15391
rect -7215 -15397 -7104 -15392
rect -8505 -15425 -8423 -15414
rect -8505 -15485 -8494 -15425
rect -8434 -15485 -8423 -15425
rect -8690 -15496 -8594 -15486
rect -8505 -15496 -8423 -15485
rect -7215 -15486 -7204 -15397
rect -7115 -15486 -7104 -15397
rect -7215 -15491 -7104 -15486
rect -7204 -15492 -7115 -15491
rect -8690 -15568 -8676 -15496
rect -8604 -15568 -8594 -15496
rect -8690 -15588 -8594 -15568
rect -6114 -15533 -6066 -15372
rect -4974 -15378 -4966 -15306
rect -4894 -15378 -4880 -15306
rect -4974 -15386 -4880 -15378
rect -2276 -15306 -2182 -15296
rect -2276 -15378 -2264 -15306
rect -2192 -15378 -2182 -15306
rect -2276 -15388 -2182 -15378
rect 401 -15493 407 -15427
rect 473 -15493 4595 -15427
rect -6114 -15599 4429 -15533
rect -6114 -15644 -6066 -15599
rect -14560 -16014 -10558 -15966
rect -10500 -15692 -6066 -15644
rect -14612 -16022 -14560 -16016
rect -10500 -16086 -10452 -15692
rect -5020 -15706 -4916 -15697
rect -20347 -18964 -19910 -18916
rect -19848 -16134 -10452 -16086
rect -10410 -15772 -5990 -15724
rect -20347 -18966 -20340 -18964
rect -20406 -18972 -20340 -18966
rect -20651 -19059 -20562 -19058
rect -20662 -19064 -20551 -19059
rect -24870 -19102 -24798 -19097
rect -24892 -19103 -24778 -19102
rect -24892 -19175 -24870 -19103
rect -24798 -19175 -24778 -19103
rect -24892 -19176 -24778 -19175
rect -21950 -19105 -21868 -19094
rect -21950 -19165 -21939 -19105
rect -21879 -19165 -21868 -19105
rect -20662 -19153 -20651 -19064
rect -20562 -19153 -20551 -19064
rect -20662 -19158 -20551 -19153
rect -20651 -19159 -20562 -19158
rect -21950 -19176 -21868 -19165
rect -24870 -19181 -24798 -19176
rect -24916 -19345 -24889 -19256
rect -24796 -19345 -24780 -19256
rect -24916 -19346 -24780 -19345
rect -20404 -19414 -20352 -19408
rect -19848 -19416 -19800 -16134
rect -14502 -16238 -14496 -16186
rect -14444 -16188 -14438 -16186
rect -10410 -16188 -10362 -15772
rect -7211 -15885 -7122 -15884
rect -7222 -15890 -7111 -15885
rect -8511 -15934 -8429 -15923
rect -8511 -15994 -8500 -15934
rect -8440 -15994 -8429 -15934
rect -7222 -15979 -7211 -15890
rect -7122 -15979 -7111 -15890
rect -6038 -15930 -5990 -15772
rect -4004 -15702 -3907 -15693
rect -4004 -15808 -3907 -15799
rect -2304 -15701 -2200 -15692
rect -5020 -15819 -4916 -15810
rect -2304 -15814 -2200 -15805
rect -1288 -15712 -1191 -15703
rect -1288 -15818 -1191 -15809
rect 4363 -15795 4429 -15599
rect 4529 -15689 4595 -15493
rect 5354 -15593 5420 -13118
rect 6934 -13198 6941 -13132
rect 7007 -13141 10062 -13132
rect 7007 -13193 8063 -13141
rect 8128 -13193 8992 -13141
rect 9057 -13193 9951 -13141
rect 10016 -13193 10062 -13141
rect 7007 -13198 10062 -13193
rect 6941 -13204 7007 -13198
rect 11883 -13417 12147 -13406
rect 11883 -13659 11894 -13417
rect 12136 -13659 12147 -13417
rect 11883 -13670 12147 -13659
rect 5558 -14050 5627 -13984
rect 5998 -14034 6067 -13984
rect 6438 -14017 6507 -13984
rect 5554 -14109 5563 -14050
rect 5622 -14109 5631 -14050
rect 5994 -14093 6003 -14034
rect 6062 -14093 6071 -14034
rect 6433 -14076 6442 -14017
rect 6501 -14076 6510 -14017
rect 5558 -14233 5627 -14109
rect 5998 -14233 6067 -14093
rect 6438 -14233 6507 -14076
rect 5552 -14302 5558 -14233
rect 5627 -14302 5633 -14233
rect 5992 -14302 5998 -14233
rect 6067 -14302 6073 -14233
rect 6432 -14302 6438 -14233
rect 6507 -14302 6513 -14233
rect 5901 -14687 7113 -14618
rect 5901 -14798 5970 -14687
rect 5703 -14882 5823 -14854
rect 5901 -14873 5970 -14867
rect 6158 -14863 6236 -14853
rect 5703 -14938 5732 -14882
rect 5788 -14938 5823 -14882
rect 6158 -14919 6170 -14863
rect 6226 -14919 6236 -14863
rect 6335 -14869 6341 -14800
rect 6410 -14869 6416 -14800
rect 6580 -14854 6700 -14838
rect 6158 -14934 6236 -14919
rect 5703 -14967 5823 -14938
rect 6341 -15079 6410 -14869
rect 6580 -14910 6610 -14854
rect 6666 -14910 6700 -14854
rect 6580 -14951 6700 -14910
rect 6299 -15138 6410 -15079
rect 6299 -15237 6367 -15138
rect 6295 -15295 6304 -15237
rect 6362 -15295 6371 -15237
rect 7044 -15242 7113 -14687
rect 7044 -15251 10140 -15242
rect 6299 -15300 6367 -15295
rect 7044 -15303 7106 -15251
rect 7158 -15252 9002 -15251
rect 7158 -15303 8069 -15252
rect 7044 -15304 8069 -15303
rect 8122 -15303 9002 -15252
rect 9055 -15303 9933 -15251
rect 9986 -15303 10140 -15251
rect 8122 -15304 10140 -15303
rect 7044 -15311 10140 -15304
rect 12187 -15243 12431 -15232
rect 12187 -15251 12198 -15243
rect 5992 -15337 6073 -15331
rect 5992 -15406 5998 -15337
rect 6067 -15342 6073 -15337
rect 6067 -15344 8115 -15342
rect 6067 -15345 8057 -15344
rect 6067 -15397 7113 -15345
rect 7165 -15396 8057 -15345
rect 8109 -15396 8115 -15344
rect 7165 -15397 8115 -15396
rect 6067 -15401 8115 -15397
rect 8182 -15392 8914 -15339
rect 9929 -15345 10000 -15343
rect 6067 -15406 6073 -15401
rect 5992 -15412 6073 -15406
rect 7321 -15434 7393 -15429
rect 8182 -15434 8248 -15392
rect 6429 -15472 6516 -15463
rect 6429 -15541 6438 -15472
rect 6507 -15541 6516 -15472
rect 7321 -15500 7327 -15434
rect 7393 -15500 8248 -15434
rect 8424 -15427 8493 -15421
rect 8861 -15440 8914 -15392
rect 8989 -15403 8998 -15347
rect 9054 -15403 9063 -15347
rect 9923 -15401 9935 -15345
rect 9991 -15401 10000 -15345
rect 10256 -15396 10336 -15390
rect 9929 -15407 9993 -15401
rect 8541 -15472 8600 -15468
rect 8493 -15477 8605 -15472
rect 8493 -15479 8541 -15477
rect 7321 -15506 7393 -15500
rect 8424 -15536 8541 -15479
rect 8600 -15536 8605 -15477
rect 8861 -15493 8989 -15440
rect 9042 -15493 9048 -15440
rect 10256 -15465 10262 -15396
rect 10331 -15465 10336 -15396
rect 10256 -15472 10336 -15465
rect 10405 -15406 10860 -15340
rect 10926 -15406 10932 -15340
rect 8424 -15541 8605 -15536
rect 6429 -15550 6516 -15541
rect 8541 -15545 8600 -15541
rect 10405 -15550 10471 -15406
rect 5354 -15659 8986 -15593
rect 9052 -15659 9058 -15593
rect 9792 -15616 9798 -15550
rect 9864 -15616 10471 -15550
rect 10536 -15500 10858 -15434
rect 10924 -15500 10930 -15434
rect 12187 -15454 12189 -15251
rect 12187 -15465 12198 -15454
rect 12420 -15465 12441 -15243
rect 12187 -15476 12431 -15465
rect 4529 -15755 9917 -15689
rect 9983 -15755 9989 -15689
rect 4363 -15861 7106 -15795
rect 7172 -15861 7178 -15795
rect 10536 -15798 10602 -15500
rect 8812 -15864 8818 -15798
rect 8884 -15864 10602 -15798
rect 10659 -15594 10850 -15528
rect 10915 -15594 10921 -15528
rect 5732 -15920 8050 -15899
rect -6038 -15952 -3582 -15930
rect 4366 -15952 8050 -15920
rect -6038 -15965 8050 -15952
rect 8116 -15965 8122 -15899
rect -6038 -15968 5918 -15965
rect -6038 -15978 4414 -15968
rect -7222 -15984 -7111 -15979
rect -7211 -15985 -7122 -15984
rect -8511 -16005 -8429 -15994
rect -3647 -16000 4414 -15978
rect 10659 -16052 10725 -15594
rect -5002 -16125 -4908 -16110
rect -14444 -16236 -10362 -16188
rect -8570 -16152 -8470 -16140
rect -8570 -16224 -8554 -16152
rect -8482 -16224 -8470 -16152
rect -5002 -16195 -4995 -16125
rect -4925 -16195 -4908 -16125
rect -5002 -16202 -4908 -16195
rect -2294 -16125 -2200 -16114
rect 7866 -16118 7872 -16052
rect 7938 -16118 10725 -16052
rect -2294 -16195 -2285 -16125
rect -2215 -16195 -2200 -16125
rect -2294 -16206 -2200 -16195
rect -8570 -16236 -8470 -16224
rect -14444 -16238 -14438 -16236
rect -7212 -16371 -7123 -16370
rect -7223 -16376 -7112 -16371
rect -8511 -16417 -8429 -16406
rect -8511 -16477 -8500 -16417
rect -8440 -16477 -8429 -16417
rect -7223 -16465 -7212 -16376
rect -7123 -16465 -7112 -16376
rect -7223 -16470 -7112 -16465
rect 7156 -16397 11207 -16325
rect -7212 -16471 -7123 -16470
rect -8511 -16488 -8429 -16477
rect -5020 -16525 -4916 -16516
rect -4004 -16521 -3907 -16512
rect -4004 -16627 -3907 -16618
rect -2304 -16520 -2200 -16511
rect -5020 -16638 -4916 -16629
rect -2304 -16633 -2200 -16624
rect -1288 -16531 -1191 -16522
rect -1288 -16637 -1191 -16628
rect 7156 -16575 7227 -16397
rect 7405 -16575 8162 -16397
rect 8340 -16575 9098 -16397
rect 9276 -16574 10029 -16397
rect 10206 -16574 10956 -16397
rect 9276 -16575 10956 -16574
rect 11134 -16575 11207 -16397
rect 7156 -16646 11207 -16575
rect -18096 -16683 -17998 -16671
rect -18096 -16757 -18084 -16683
rect -18010 -16757 -17998 -16683
rect -8566 -16685 -8470 -16670
rect -18096 -16769 -17998 -16757
rect -16924 -16732 -16834 -16717
rect -16924 -16792 -16909 -16732
rect -16849 -16792 -16834 -16732
rect -8566 -16754 -8551 -16685
rect -8482 -16754 -8470 -16685
rect -8566 -16768 -8470 -16754
rect -16924 -16807 -16834 -16792
rect 12414 -16816 12821 -16704
rect 12128 -16820 12821 -16816
rect 16250 -16737 16588 -16694
rect -7216 -16878 -7127 -16877
rect -7227 -16883 -7116 -16878
rect -8511 -16939 -8429 -16928
rect -18077 -16980 -18015 -16976
rect -18088 -17052 -18082 -16980
rect -18010 -17052 -18004 -16980
rect -12499 -17039 -12373 -16997
rect -8511 -16999 -8500 -16939
rect -8440 -16999 -8429 -16939
rect -7227 -16972 -7216 -16883
rect -7127 -16972 -7116 -16883
rect 7847 -16911 7853 -16845
rect 7919 -16911 10121 -16845
rect -7227 -16977 -7116 -16972
rect -5010 -16958 -4916 -16940
rect -7216 -16978 -7127 -16977
rect -8511 -17010 -8429 -16999
rect -5010 -17021 -5000 -16958
rect -4937 -17021 -4916 -16958
rect -5010 -17032 -4916 -17021
rect -2298 -16958 -2204 -16938
rect -2298 -17021 -2291 -16958
rect -2228 -17021 -2204 -16958
rect -2298 -17030 -2204 -17021
rect 1537 -17001 5798 -16982
rect -18077 -17056 -18015 -17052
rect -18096 -17113 -17992 -17102
rect -18096 -17202 -18089 -17113
rect -18000 -17202 -17992 -17113
rect -18096 -17208 -17992 -17202
rect -15052 -17951 -14963 -17950
rect -15063 -17956 -14952 -17951
rect -16353 -17984 -16271 -17973
rect -16353 -18044 -16342 -17984
rect -16282 -18044 -16271 -17984
rect -16353 -18055 -16271 -18044
rect -15063 -18045 -15052 -17956
rect -14963 -18045 -14952 -17956
rect -15063 -18050 -14952 -18045
rect -15052 -18051 -14963 -18050
rect -18100 -18069 -18002 -18057
rect -18100 -18143 -18088 -18069
rect -18014 -18143 -18002 -18069
rect -18100 -18155 -18002 -18143
rect -17054 -18163 -16968 -18151
rect -17054 -18223 -17040 -18163
rect -16980 -18223 -16968 -18163
rect -12499 -18161 -12471 -17039
rect -12399 -18161 -12373 -17039
rect 1537 -17067 8989 -17001
rect 9055 -17067 9061 -17001
rect -5407 -17154 -5288 -17149
rect 1537 -17154 1622 -17067
rect 10055 -17123 10121 -16911
rect 12128 -16846 13042 -16820
rect 12128 -16908 13186 -16846
rect 12128 -17027 12233 -16908
rect 12352 -16949 13186 -16908
rect 12352 -17027 12960 -16949
rect 12128 -17068 12960 -17027
rect 13079 -17068 13186 -16949
rect 16250 -16995 16285 -16737
rect 16543 -16995 16588 -16737
rect 16250 -17028 16588 -16995
rect 5732 -17130 9917 -17123
rect -8560 -17205 -8464 -17188
rect -8560 -17274 -8549 -17205
rect -8480 -17274 -8464 -17205
rect -5414 -17243 -5397 -17154
rect -5307 -17243 1624 -17154
rect 1680 -17178 9917 -17130
rect -5407 -17252 -5288 -17243
rect -8560 -17286 -8464 -17274
rect -7215 -17353 -7126 -17352
rect -7226 -17358 -7115 -17353
rect -8508 -17408 -8426 -17397
rect -8508 -17468 -8497 -17408
rect -8437 -17468 -8426 -17408
rect -7226 -17447 -7215 -17358
rect -7126 -17447 -7115 -17358
rect -5242 -17372 -5236 -17320
rect -5184 -17372 -5178 -17320
rect -5020 -17344 -4916 -17335
rect -7226 -17452 -7115 -17447
rect -7215 -17453 -7126 -17452
rect -8508 -17479 -8426 -17468
rect -5234 -17548 -5186 -17372
rect -4004 -17340 -3907 -17331
rect -4004 -17446 -3907 -17437
rect -2304 -17339 -2200 -17330
rect -5020 -17457 -4916 -17448
rect -2304 -17452 -2200 -17443
rect -1288 -17350 -1191 -17341
rect -1288 -17456 -1191 -17447
rect 1680 -17548 1728 -17178
rect 5732 -17189 9917 -17178
rect 9983 -17189 9989 -17123
rect 10055 -17189 10704 -17123
rect 12128 -17133 13186 -17068
rect 1799 -17224 7102 -17221
rect -5234 -17596 1728 -17548
rect 1794 -17287 7102 -17224
rect 7168 -17287 7174 -17221
rect -8570 -17615 -8474 -17598
rect -11090 -17641 -11008 -17630
rect -11090 -17701 -11079 -17641
rect -11019 -17701 -11008 -17641
rect -8570 -17684 -8554 -17615
rect -8485 -17684 -8474 -17615
rect 1794 -17648 1878 -17287
rect 8831 -17321 8837 -17255
rect 8903 -17321 10588 -17255
rect 1941 -17408 8050 -17342
rect 8116 -17408 8122 -17342
rect -8570 -17696 -8474 -17684
rect -11090 -17712 -11008 -17701
rect -926 -17732 1878 -17648
rect -4988 -17780 -4894 -17758
rect -7210 -17805 -7121 -17804
rect -7221 -17810 -7110 -17805
rect -8506 -17865 -8424 -17854
rect -8506 -17925 -8495 -17865
rect -8435 -17925 -8424 -17865
rect -7221 -17899 -7210 -17810
rect -7121 -17899 -7110 -17810
rect -4988 -17841 -4979 -17780
rect -4918 -17841 -4894 -17780
rect -4988 -17850 -4894 -17841
rect -2280 -17780 -2186 -17760
rect -2280 -17841 -2269 -17780
rect -2208 -17841 -2186 -17780
rect -2280 -17852 -2186 -17841
rect -7221 -17904 -7110 -17899
rect -7210 -17905 -7121 -17904
rect -8506 -17936 -8424 -17925
rect -926 -17980 -842 -17732
rect 1942 -17812 2026 -17408
rect 9801 -17413 9807 -17349
rect 9873 -17413 10453 -17349
rect 8396 -17444 8470 -17438
rect 6780 -17463 6849 -17457
rect 6849 -17516 8206 -17477
rect 8396 -17479 8405 -17444
rect 8461 -17479 8470 -17444
rect 8396 -17508 8401 -17479
rect 6780 -17538 6849 -17532
rect 810 -17896 816 -17812
rect 900 -17896 2026 -17812
rect 5407 -17552 5473 -17546
rect -2614 -18064 -2608 -17980
rect -2524 -18064 -842 -17980
rect -12499 -18207 -12373 -18161
rect -8568 -18097 -8472 -18080
rect -8568 -18166 -8554 -18097
rect -8485 -18166 -8472 -18097
rect -8568 -18178 -8472 -18166
rect -5020 -18163 -4916 -18154
rect -17054 -18237 -16968 -18223
rect -7210 -18247 -7121 -18246
rect -7221 -18252 -7110 -18247
rect -8504 -18330 -8422 -18319
rect -18060 -18385 -18000 -18381
rect -18071 -18455 -18065 -18385
rect -17995 -18455 -17989 -18385
rect -8504 -18390 -8493 -18330
rect -8433 -18390 -8422 -18330
rect -7221 -18341 -7210 -18252
rect -7121 -18341 -7110 -18252
rect -4004 -18159 -3907 -18150
rect -4004 -18265 -3907 -18256
rect -2304 -18158 -2200 -18149
rect -5020 -18276 -4916 -18267
rect -2304 -18271 -2200 -18262
rect -1288 -18169 -1191 -18160
rect -1288 -18275 -1191 -18266
rect -7221 -18346 -7110 -18341
rect -7210 -18347 -7121 -18346
rect -12661 -18396 -12599 -18392
rect -15059 -18444 -14970 -18443
rect -15070 -18449 -14959 -18444
rect -18060 -18459 -18000 -18455
rect -16359 -18493 -16277 -18482
rect -18094 -18515 -18015 -18511
rect -18105 -18604 -18099 -18515
rect -18010 -18604 -18004 -18515
rect -16359 -18553 -16348 -18493
rect -16288 -18553 -16277 -18493
rect -15070 -18538 -15059 -18449
rect -14970 -18538 -14959 -18449
rect -12672 -18468 -12666 -18396
rect -12594 -18468 -12588 -18396
rect -8504 -18401 -8422 -18390
rect -12661 -18472 -12599 -18468
rect -15070 -18543 -14959 -18538
rect -15059 -18544 -14970 -18543
rect -16359 -18564 -16277 -18553
rect -8564 -18567 -8468 -18548
rect -12628 -18573 -12549 -18569
rect -18094 -18608 -18015 -18604
rect -12639 -18662 -12633 -18573
rect -12544 -18662 -12538 -18573
rect -8564 -18636 -8554 -18567
rect -8485 -18636 -8468 -18567
rect -8564 -18646 -8468 -18636
rect -5014 -18582 -4920 -18572
rect -5014 -18654 -5006 -18582
rect -4934 -18654 -4920 -18582
rect -12628 -18666 -12549 -18662
rect -5014 -18664 -4920 -18654
rect -2302 -18582 -2208 -18572
rect -2302 -18654 -2294 -18582
rect -2222 -18654 -2208 -18582
rect -2302 -18664 -2208 -18654
rect -19377 -18705 -19311 -18699
rect -19311 -18771 -14471 -18705
rect -19377 -18777 -19311 -18771
rect -15060 -18930 -14971 -18929
rect -15071 -18935 -14960 -18930
rect -16359 -18976 -16277 -18965
rect -16359 -19036 -16348 -18976
rect -16288 -19036 -16277 -18976
rect -15071 -19024 -15060 -18935
rect -14971 -19024 -14960 -18935
rect -15071 -19029 -14960 -19024
rect -15060 -19030 -14971 -19029
rect -16359 -19047 -16277 -19036
rect -20352 -19464 -19800 -19416
rect -15064 -19437 -14975 -19436
rect -15075 -19442 -14964 -19437
rect -20404 -19472 -20352 -19466
rect -18098 -19475 -18000 -19463
rect -18098 -19549 -18086 -19475
rect -18012 -19549 -18000 -19475
rect -18098 -19561 -18000 -19549
rect -16359 -19498 -16277 -19487
rect -16359 -19558 -16348 -19498
rect -16288 -19558 -16277 -19498
rect -15075 -19531 -15064 -19442
rect -14975 -19531 -14964 -19442
rect -15075 -19536 -14964 -19531
rect -15064 -19537 -14975 -19536
rect -20655 -19566 -20566 -19565
rect -20666 -19571 -20555 -19566
rect -16359 -19569 -16277 -19558
rect -21950 -19627 -21868 -19616
rect -21950 -19687 -21939 -19627
rect -21879 -19687 -21868 -19627
rect -20666 -19660 -20655 -19571
rect -20566 -19660 -20555 -19571
rect -20666 -19665 -20555 -19660
rect -18024 -19622 -17942 -19614
rect -20655 -19666 -20566 -19665
rect -21950 -19698 -21868 -19687
rect -18024 -19685 -18016 -19622
rect -17953 -19685 -17942 -19622
rect -18024 -19692 -17942 -19685
rect -16934 -19618 -16854 -19609
rect -16934 -19678 -16925 -19618
rect -16865 -19678 -16854 -19618
rect -16934 -19689 -16854 -19678
rect -14537 -19617 -14471 -18771
rect -7216 -18733 -7127 -18724
rect -8500 -18811 -8418 -18800
rect -8500 -18871 -8489 -18811
rect -8429 -18871 -8418 -18811
rect -7216 -18831 -7127 -18822
rect -8500 -18882 -8418 -18871
rect -5020 -18982 -4916 -18973
rect -4004 -18978 -3907 -18969
rect -4004 -19084 -3907 -19075
rect -2304 -18977 -2200 -18968
rect -8584 -19098 -8512 -19092
rect -5020 -19095 -4916 -19086
rect -2304 -19090 -2200 -19081
rect -1288 -18988 -1191 -18979
rect -1288 -19094 -1191 -19085
rect -8584 -19176 -8512 -19170
rect -5026 -19430 -4932 -19420
rect -5026 -19502 -5014 -19430
rect -4942 -19502 -4932 -19430
rect -5026 -19512 -4932 -19502
rect -2308 -19430 -2214 -19420
rect -2308 -19502 -2300 -19430
rect -2228 -19502 -2214 -19430
rect -2308 -19512 -2214 -19502
rect -14537 -19683 -413 -19617
rect -347 -19683 -341 -19617
rect -20317 -19762 -10635 -19753
rect -23350 -19796 -23227 -19784
rect -23350 -19897 -23338 -19796
rect -23237 -19897 -23227 -19796
rect -20322 -19819 -10635 -19762
rect -20322 -19894 -20274 -19819
rect -14808 -19866 -14756 -19860
rect -24825 -19908 -24709 -19898
rect -24825 -20004 -24815 -19908
rect -24719 -20004 -24709 -19908
rect -23350 -19912 -23227 -19897
rect -20330 -19946 -20324 -19894
rect -20272 -19946 -20266 -19894
rect -17994 -19907 -17906 -19898
rect -17994 -19978 -17986 -19907
rect -17915 -19978 -17906 -19907
rect -15063 -19912 -14974 -19911
rect -15074 -19917 -14963 -19912
rect -17994 -19986 -17906 -19978
rect -16356 -19967 -16274 -19956
rect -24825 -20014 -24709 -20004
rect -16356 -20027 -16345 -19967
rect -16285 -20027 -16274 -19967
rect -15074 -20006 -15063 -19917
rect -14974 -20006 -14963 -19917
rect -14756 -19916 -10766 -19868
rect -14808 -19924 -14756 -19918
rect -15074 -20011 -14963 -20006
rect -12499 -19996 -12373 -19954
rect -15063 -20012 -14974 -20011
rect -16356 -20038 -16274 -20027
rect -20654 -20041 -20565 -20040
rect -20665 -20046 -20554 -20041
rect -21947 -20096 -21865 -20085
rect -21947 -20156 -21936 -20096
rect -21876 -20156 -21865 -20096
rect -20665 -20135 -20654 -20046
rect -20565 -20135 -20554 -20046
rect -20665 -20140 -20554 -20135
rect -20654 -20141 -20565 -20140
rect -21947 -20167 -21865 -20156
rect -24956 -20291 -24844 -20290
rect -24956 -20363 -24936 -20291
rect -24864 -20363 -24844 -20291
rect -24956 -20364 -24844 -20363
rect -20399 -20354 -20347 -20348
rect -20347 -20360 -18426 -20356
rect -20347 -20404 -18421 -20360
rect -15058 -20364 -14969 -20363
rect -20399 -20412 -20347 -20406
rect -24940 -20444 -24792 -20436
rect -24940 -20533 -24902 -20444
rect -24811 -20533 -24792 -20444
rect -20649 -20493 -20560 -20492
rect -24940 -20534 -24792 -20533
rect -20660 -20498 -20549 -20493
rect -21945 -20553 -21863 -20542
rect -21945 -20613 -21934 -20553
rect -21874 -20613 -21863 -20553
rect -20660 -20587 -20649 -20498
rect -20560 -20587 -20549 -20498
rect -20660 -20592 -20549 -20587
rect -20649 -20593 -20560 -20592
rect -21945 -20624 -21863 -20613
rect -18572 -20814 -18520 -20808
rect -18572 -20872 -18520 -20866
rect -20649 -20935 -20560 -20934
rect -20660 -20940 -20549 -20935
rect -23341 -20994 -23218 -20982
rect -24825 -21104 -24709 -21094
rect -24825 -21200 -24815 -21104
rect -24719 -21200 -24709 -21104
rect -23341 -21095 -23329 -20994
rect -23228 -21095 -23218 -20994
rect -21943 -21018 -21861 -21007
rect -21943 -21078 -21932 -21018
rect -21872 -21078 -21861 -21018
rect -20660 -21029 -20649 -20940
rect -20560 -21029 -20549 -20940
rect -20660 -21034 -20549 -21029
rect -20649 -21035 -20560 -21034
rect -21943 -21089 -21861 -21078
rect -23341 -21110 -23218 -21095
rect -24825 -21210 -24709 -21200
rect -18698 -21346 -18692 -21294
rect -18640 -21346 -18634 -21294
rect -20655 -21421 -20566 -21412
rect -24936 -21497 -24812 -21464
rect -24936 -21569 -24924 -21497
rect -24852 -21569 -24812 -21497
rect -24936 -21574 -24812 -21569
rect -21939 -21499 -21857 -21488
rect -21939 -21559 -21928 -21499
rect -21868 -21559 -21857 -21499
rect -20655 -21519 -20566 -21510
rect -21939 -21570 -21857 -21559
rect -24936 -21650 -24812 -21638
rect -24936 -21739 -24913 -21650
rect -24823 -21739 -24812 -21650
rect -24936 -21748 -24812 -21739
rect -18690 -21784 -18642 -21346
rect -18570 -21672 -18522 -20872
rect -18466 -21596 -18421 -20404
rect -15069 -20369 -14958 -20364
rect -16354 -20424 -16272 -20413
rect -16354 -20484 -16343 -20424
rect -16283 -20484 -16272 -20424
rect -15069 -20458 -15058 -20369
rect -14969 -20458 -14958 -20369
rect -15069 -20463 -14958 -20458
rect -15058 -20464 -14969 -20463
rect -16354 -20495 -16272 -20484
rect -15058 -20806 -14969 -20805
rect -15069 -20811 -14958 -20806
rect -18102 -20869 -18004 -20857
rect -18102 -20943 -18090 -20869
rect -18016 -20943 -18004 -20869
rect -18102 -20955 -18004 -20943
rect -16352 -20889 -16270 -20878
rect -16352 -20949 -16341 -20889
rect -16281 -20949 -16270 -20889
rect -15069 -20900 -15058 -20811
rect -14969 -20900 -14958 -20811
rect -15069 -20905 -14958 -20900
rect -15058 -20906 -14969 -20905
rect -16352 -20960 -16270 -20949
rect -16930 -21013 -16836 -20995
rect -16930 -21075 -16916 -21013
rect -16854 -21075 -16836 -21013
rect -16930 -21091 -16836 -21075
rect -12499 -21118 -12471 -19996
rect -12399 -21118 -12373 -19996
rect -10814 -20290 -10766 -19916
rect -10701 -20195 -10635 -19819
rect -5020 -19801 -4916 -19792
rect -4004 -19797 -3907 -19788
rect -4004 -19903 -3907 -19894
rect -2304 -19796 -2200 -19787
rect -5020 -19914 -4916 -19905
rect -2304 -19909 -2200 -19900
rect -1288 -19807 -1191 -19798
rect -1288 -19913 -1191 -19904
rect -5174 -20056 -5074 -20044
rect -5174 -20128 -5166 -20056
rect -5094 -20128 -5074 -20056
rect -2420 -20056 -2348 -20050
rect -2424 -20123 -2420 -20061
rect -2348 -20123 -2344 -20061
rect 5407 -20121 5473 -17619
rect 6066 -17566 6132 -17560
rect 6132 -17575 8139 -17566
rect 6132 -17627 8079 -17575
rect 8131 -17627 8139 -17575
rect 8167 -17585 8206 -17516
rect 8465 -17508 8470 -17479
rect 8615 -17538 8993 -17472
rect 9059 -17538 9065 -17472
rect 10264 -17479 10324 -17473
rect 10257 -17537 10264 -17481
rect 10324 -17537 10331 -17481
rect 8401 -17549 8465 -17543
rect 8616 -17585 8655 -17538
rect 10264 -17545 10324 -17539
rect 8167 -17624 8655 -17585
rect 6132 -17632 8139 -17627
rect 8992 -17632 9001 -17566
rect 9067 -17632 9076 -17566
rect 9931 -17631 9937 -17565
rect 10003 -17631 10012 -17565
rect 10387 -17566 10453 -17413
rect 10522 -17472 10588 -17321
rect 10638 -17378 10704 -17189
rect 12467 -17292 13186 -17133
rect 12796 -17325 13186 -17292
rect 10638 -17444 10850 -17378
rect 10916 -17444 10922 -17378
rect 10522 -17538 10888 -17472
rect 10954 -17538 10963 -17472
rect 10387 -17632 10859 -17566
rect 10925 -17632 10931 -17566
rect 6066 -17638 6132 -17632
rect 6934 -17726 6941 -17660
rect 7007 -17669 10062 -17660
rect 7007 -17721 8063 -17669
rect 8128 -17721 8992 -17669
rect 9057 -17721 9951 -17669
rect 10016 -17721 10062 -17669
rect 7007 -17726 10062 -17721
rect 6941 -17732 7007 -17726
rect 11883 -17945 12147 -17934
rect 11883 -18187 11894 -17945
rect 12136 -18187 12147 -17945
rect 17515 -18021 17672 -18008
rect 17515 -18154 17526 -18021
rect 17659 -18154 17672 -18021
rect 17515 -18165 17672 -18154
rect 11883 -18198 12147 -18187
rect 5558 -18556 5627 -18512
rect 5554 -18615 5563 -18556
rect 5622 -18615 5631 -18556
rect 5998 -18574 6067 -18512
rect 6438 -18567 6507 -18512
rect 15538 -18514 15708 -18501
rect 5558 -18761 5627 -18615
rect 5994 -18633 6003 -18574
rect 6062 -18633 6071 -18574
rect 6431 -18626 6440 -18567
rect 6499 -18626 6508 -18567
rect 5998 -18761 6067 -18633
rect 6438 -18761 6507 -18626
rect 15538 -18658 15551 -18514
rect 15695 -18658 15708 -18514
rect 15538 -18671 15708 -18658
rect 5552 -18830 5558 -18761
rect 5627 -18830 5633 -18761
rect 5992 -18830 5998 -18761
rect 6067 -18830 6073 -18761
rect 6432 -18830 6438 -18761
rect 6507 -18830 6513 -18761
rect 17966 -18869 18059 -18858
rect 17966 -18940 17977 -18869
rect 18048 -18940 18059 -18869
rect 17966 -18951 18059 -18940
rect 5901 -19215 7113 -19146
rect 5901 -19326 5970 -19215
rect 5703 -19410 5823 -19382
rect 5901 -19401 5970 -19395
rect 6158 -19391 6236 -19381
rect 5703 -19466 5732 -19410
rect 5788 -19466 5823 -19410
rect 6158 -19447 6170 -19391
rect 6226 -19447 6236 -19391
rect 6335 -19397 6341 -19328
rect 6410 -19397 6416 -19328
rect 6580 -19382 6700 -19366
rect 6158 -19462 6236 -19447
rect 5703 -19495 5823 -19466
rect 6341 -19607 6410 -19397
rect 6580 -19438 6610 -19382
rect 6666 -19438 6700 -19382
rect 6580 -19479 6700 -19438
rect 6299 -19666 6410 -19607
rect 6299 -19765 6367 -19666
rect 6295 -19823 6304 -19765
rect 6362 -19823 6371 -19765
rect 7044 -19770 7113 -19215
rect 7044 -19779 10140 -19770
rect 6299 -19828 6367 -19823
rect 7044 -19831 7106 -19779
rect 7158 -19780 9002 -19779
rect 7158 -19831 8069 -19780
rect 7044 -19832 8069 -19831
rect 8122 -19831 9002 -19780
rect 9055 -19831 9933 -19779
rect 9986 -19831 10140 -19779
rect 8122 -19832 10140 -19831
rect 7044 -19839 10140 -19832
rect 12187 -19771 12431 -19760
rect 12187 -19779 12198 -19771
rect 5992 -19865 6073 -19859
rect 5992 -19934 5998 -19865
rect 6067 -19870 6073 -19865
rect 6067 -19872 8115 -19870
rect 6067 -19873 8057 -19872
rect 6067 -19925 7113 -19873
rect 7165 -19924 8057 -19873
rect 8109 -19924 8115 -19872
rect 7165 -19925 8115 -19924
rect 6067 -19929 8115 -19925
rect 8182 -19920 8914 -19867
rect 9929 -19873 10000 -19871
rect 6067 -19934 6073 -19929
rect 5992 -19940 6073 -19934
rect 7321 -19962 7393 -19957
rect 8182 -19962 8248 -19920
rect 6429 -20000 6516 -19991
rect 6429 -20069 6438 -20000
rect 6507 -20069 6516 -20000
rect 7321 -20028 7327 -19962
rect 7393 -20028 8248 -19962
rect 8424 -19955 8493 -19949
rect 8861 -19968 8914 -19920
rect 8989 -19931 8998 -19875
rect 9054 -19931 9063 -19875
rect 9923 -19929 9935 -19873
rect 9991 -19929 10000 -19873
rect 10256 -19924 10336 -19918
rect 9929 -19935 9993 -19929
rect 8541 -20000 8600 -19996
rect 8493 -20005 8605 -20000
rect 8493 -20007 8541 -20005
rect 7321 -20034 7393 -20028
rect 8424 -20064 8541 -20007
rect 8600 -20064 8605 -20005
rect 8861 -20021 8989 -19968
rect 9042 -20021 9048 -19968
rect 10256 -19993 10262 -19924
rect 10331 -19993 10336 -19924
rect 10256 -20000 10336 -19993
rect 10405 -19934 10860 -19868
rect 10926 -19934 10932 -19868
rect 8424 -20069 8605 -20064
rect 6429 -20078 6516 -20069
rect 8541 -20073 8600 -20069
rect 10405 -20078 10471 -19934
rect -5174 -20134 -5074 -20128
rect -2420 -20134 -2348 -20128
rect 5407 -20187 8986 -20121
rect 9052 -20187 9058 -20121
rect 9792 -20144 9798 -20078
rect 9864 -20144 10471 -20078
rect 10536 -20028 10858 -19962
rect 10924 -20028 10930 -19962
rect 12187 -19982 12189 -19779
rect 12187 -19993 12198 -19982
rect 12420 -19993 12441 -19771
rect 12187 -20004 12431 -19993
rect -10701 -20261 -337 -20195
rect -10814 -20338 -446 -20290
rect -5586 -20422 -5534 -20416
rect -5586 -20480 -5534 -20474
rect -2310 -20417 -2194 -20411
rect -11090 -20598 -11008 -20587
rect -11090 -20658 -11079 -20598
rect -11019 -20658 -11008 -20598
rect -11090 -20669 -11008 -20658
rect -12499 -21164 -12373 -21118
rect -18051 -21176 -17995 -21170
rect -18059 -21237 -18053 -21176
rect -17992 -21237 -17986 -21176
rect -18051 -21244 -17995 -21237
rect -15064 -21292 -14975 -21283
rect -17974 -21340 -17886 -21322
rect -17974 -21404 -17968 -21340
rect -17904 -21404 -17886 -21340
rect -17974 -21410 -17886 -21404
rect -16348 -21370 -16266 -21359
rect -16348 -21430 -16337 -21370
rect -16277 -21430 -16266 -21370
rect -15064 -21390 -14975 -21381
rect -12618 -21367 -12524 -21354
rect -16348 -21441 -16266 -21430
rect -12618 -21437 -12609 -21367
rect -12539 -21437 -12524 -21367
rect -12618 -21448 -12524 -21437
rect -12640 -21527 -12518 -21518
rect -18466 -21641 -16235 -21596
rect -12640 -21616 -12628 -21527
rect -12539 -21616 -12518 -21527
rect -12640 -21624 -12518 -21616
rect -18570 -21720 -16310 -21672
rect -18690 -21832 -16420 -21784
rect -16738 -21983 -16646 -21969
rect -16738 -22047 -16726 -21983
rect -16662 -22047 -16646 -21983
rect -16738 -22061 -16646 -22047
rect -16468 -22230 -16420 -21832
rect -16358 -22116 -16310 -21720
rect -16280 -22020 -16235 -21641
rect -5584 -21664 -5536 -20480
rect -494 -20430 -446 -20338
rect -403 -20323 -337 -20261
rect 1361 -20283 1367 -20217
rect 1433 -20283 9917 -20217
rect 9983 -20283 9989 -20217
rect -403 -20389 7106 -20323
rect 7172 -20389 7178 -20323
rect 10536 -20326 10602 -20028
rect 8812 -20392 8818 -20326
rect 8884 -20392 10602 -20326
rect 10659 -20122 10850 -20056
rect 10915 -20122 10921 -20056
rect 5732 -20430 8050 -20427
rect -2310 -20539 -2194 -20533
rect -1288 -20440 -1191 -20431
rect -494 -20478 8050 -20430
rect 5732 -20493 8050 -20478
rect 8116 -20493 8122 -20427
rect -1288 -20546 -1191 -20537
rect 10659 -20580 10725 -20122
rect 16196 -20177 16516 -20147
rect 16196 -20436 16221 -20177
rect 16480 -20436 16516 -20177
rect 16196 -20467 16516 -20436
rect -5020 -20620 -4916 -20611
rect -4004 -20616 -3907 -20607
rect 7866 -20646 7872 -20580
rect 7938 -20646 10725 -20580
rect -4004 -20722 -3907 -20713
rect -5020 -20733 -4916 -20724
rect 7156 -20925 11207 -20853
rect 3886 -21046 3970 -21040
rect -3912 -21130 -3906 -21046
rect -3822 -21130 3886 -21046
rect 3886 -21136 3970 -21130
rect 7156 -21103 7227 -20925
rect 7405 -21103 8162 -20925
rect 8340 -21103 9098 -20925
rect 9276 -21102 10029 -20925
rect 10206 -21102 10956 -20925
rect 9276 -21103 10956 -21102
rect 11134 -21103 11207 -20925
rect 7156 -21174 11207 -21103
rect 12414 -21344 12821 -21232
rect 12128 -21348 12821 -21344
rect 1221 -21389 1287 -21383
rect 1287 -21455 4745 -21389
rect 4811 -21455 4817 -21389
rect 7847 -21439 7853 -21373
rect 7919 -21439 10121 -21373
rect 1221 -21461 1287 -21455
rect -5136 -21608 -5130 -21525
rect -5047 -21529 6237 -21525
rect -5047 -21595 8989 -21529
rect 9055 -21595 9061 -21529
rect -5047 -21608 6237 -21595
rect 10055 -21651 10121 -21439
rect 12128 -21374 13042 -21348
rect 12128 -21436 13186 -21374
rect 12128 -21555 12233 -21436
rect 12352 -21477 13186 -21436
rect 12352 -21555 12960 -21477
rect 12128 -21596 12960 -21555
rect 13079 -21596 13186 -21477
rect 5732 -21664 9917 -21651
rect -5584 -21712 9917 -21664
rect 5732 -21717 9917 -21712
rect 9983 -21717 9989 -21651
rect 10055 -21717 10704 -21651
rect 12128 -21661 13186 -21596
rect -2757 -21819 -2751 -21748
rect -2680 -21749 6679 -21748
rect -2680 -21815 7102 -21749
rect 7168 -21815 7174 -21749
rect -2680 -21819 6679 -21815
rect 8831 -21849 8837 -21783
rect 8903 -21849 10588 -21783
rect 5732 -21872 8050 -21870
rect 668 -21956 674 -21872
rect 758 -21936 8050 -21872
rect 8116 -21936 8122 -21870
rect 758 -21956 5966 -21936
rect 9801 -21941 9807 -21877
rect 9873 -21941 10453 -21877
rect 8396 -21972 8470 -21966
rect 6780 -21991 6849 -21985
rect -16280 -22065 5277 -22020
rect -16358 -22164 -12790 -22116
rect -12756 -22150 -12750 -22098
rect -12698 -22100 -12692 -22098
rect -12698 -22148 5166 -22100
rect -12698 -22150 -12692 -22148
rect -12838 -22182 -12790 -22164
rect -12838 -22230 -10534 -22182
rect -18100 -22273 -18002 -22261
rect -23344 -22288 -23221 -22276
rect -23344 -22389 -23332 -22288
rect -23231 -22389 -23221 -22288
rect -18100 -22347 -18088 -22273
rect -18014 -22347 -18002 -22273
rect -16468 -22278 -12972 -22230
rect -18100 -22359 -18002 -22347
rect -24815 -22412 -24699 -22402
rect -23344 -22404 -23221 -22389
rect -13020 -22400 -12972 -22278
rect -12872 -22284 -12820 -22278
rect -12820 -22334 -10620 -22286
rect -12872 -22342 -12820 -22336
rect -24815 -22508 -24805 -22412
rect -24709 -22508 -24699 -22412
rect -13020 -22448 -10720 -22400
rect -24815 -22518 -24699 -22508
rect -12499 -22575 -12373 -22533
rect -18074 -22600 -17972 -22582
rect -18074 -22666 -18061 -22600
rect -17995 -22666 -17972 -22600
rect -18074 -22678 -17972 -22666
rect -18080 -22745 -17952 -22724
rect -24900 -22798 -24806 -22786
rect -24900 -22870 -24890 -22798
rect -24818 -22870 -24806 -22798
rect -18080 -22834 -18071 -22745
rect -17982 -22834 -17952 -22745
rect -18080 -22846 -17952 -22834
rect -24900 -22882 -24806 -22870
rect -24926 -22951 -24808 -22942
rect -24926 -23040 -24913 -22951
rect -24819 -23040 -24808 -22951
rect -24926 -23052 -24808 -23040
rect -16706 -23367 -16596 -23349
rect -16706 -23445 -16688 -23367
rect -16610 -23445 -16596 -23367
rect -16706 -23459 -16596 -23445
rect -23384 -23604 -23261 -23592
rect -23384 -23705 -23372 -23604
rect -23271 -23705 -23261 -23604
rect -24835 -23718 -24719 -23708
rect -24835 -23814 -24825 -23718
rect -24729 -23814 -24719 -23718
rect -23384 -23720 -23261 -23705
rect -18102 -23675 -18004 -23663
rect -18102 -23749 -18090 -23675
rect -18016 -23749 -18004 -23675
rect -12499 -23697 -12471 -22575
rect -12399 -23697 -12373 -22575
rect -11090 -23177 -11008 -23166
rect -11090 -23237 -11079 -23177
rect -11019 -23237 -11008 -23177
rect -11090 -23248 -11008 -23237
rect -12499 -23743 -12373 -23697
rect -18102 -23761 -18004 -23749
rect -24835 -23824 -24719 -23814
rect -12688 -23951 -12602 -23946
rect -12688 -23952 -12676 -23951
rect -18050 -23986 -17962 -23978
rect -18050 -24058 -18042 -23986
rect -17970 -24058 -17962 -23986
rect -12736 -24014 -12676 -23952
rect -12613 -23952 -12602 -23951
rect -12613 -24014 -12578 -23952
rect -12736 -24016 -12578 -24014
rect -18050 -24066 -17962 -24058
rect -12738 -24092 -12574 -24076
rect -24938 -24108 -24848 -24102
rect -24938 -24180 -24926 -24108
rect -24854 -24180 -24848 -24108
rect -24938 -24186 -24848 -24180
rect -18084 -24131 -17958 -24102
rect -18084 -24220 -18063 -24131
rect -17974 -24220 -17958 -24131
rect -12738 -24163 -12685 -24092
rect -12614 -24163 -12574 -24092
rect -12738 -24164 -12574 -24163
rect -18084 -24246 -17958 -24220
rect -24920 -24261 -24800 -24250
rect -24920 -24350 -24907 -24261
rect -24813 -24350 -24800 -24261
rect -24920 -24362 -24800 -24350
rect -16704 -24775 -16598 -24759
rect -16704 -24849 -16688 -24775
rect -16614 -24849 -16598 -24775
rect -16704 -24865 -16598 -24849
rect -18096 -25055 -17998 -25043
rect -18096 -25129 -18084 -25055
rect -18010 -25129 -17998 -25055
rect -18096 -25141 -17998 -25129
rect -13022 -25164 -13016 -25112
rect -12964 -25114 -12958 -25112
rect -12964 -25162 -10844 -25114
rect -12964 -25164 -12958 -25162
rect -12499 -25343 -12373 -25301
rect -17964 -25350 -17878 -25344
rect -17964 -25422 -17956 -25350
rect -17884 -25422 -17878 -25350
rect -17964 -25428 -17878 -25422
rect -17982 -25553 -17878 -25480
rect -17982 -25642 -17976 -25553
rect -17887 -25642 -17878 -25553
rect -17982 -25650 -17878 -25642
rect -12499 -26465 -12471 -25343
rect -12399 -26465 -12373 -25343
rect -10892 -25824 -10844 -25162
rect -10768 -25724 -10720 -22448
rect -10668 -25368 -10620 -22334
rect -10582 -25242 -10534 -22230
rect -10479 -22299 5069 -22213
rect -10479 -25098 -10393 -22299
rect -5708 -22456 -5702 -22404
rect -5650 -22406 -5644 -22404
rect -5650 -22454 4942 -22406
rect -5650 -22456 -5644 -22454
rect -2920 -22610 -2914 -22526
rect -2830 -22529 4836 -22526
rect -2830 -22610 4849 -22529
rect 490 -22696 574 -22690
rect 574 -22705 4656 -22696
rect 574 -22780 4717 -22705
rect 490 -22786 574 -22780
rect -5854 -24358 -5802 -24352
rect -6038 -24414 -6032 -24362
rect -5980 -24414 -5974 -24362
rect -6030 -24978 -5982 -24414
rect -5854 -24416 -5802 -24410
rect -6032 -24984 -5980 -24978
rect -5852 -25028 -5804 -24416
rect -6032 -25042 -5980 -25036
rect -5854 -25034 -5802 -25028
rect -5854 -25092 -5802 -25086
rect -10490 -25107 -10366 -25098
rect -10490 -25193 -10479 -25107
rect -10393 -25193 -10366 -25107
rect -10490 -25206 -10366 -25193
rect -10582 -25290 4462 -25242
rect -10668 -25416 4354 -25368
rect -10158 -25634 -10152 -25530
rect -10048 -25634 4226 -25530
rect -10768 -25772 -5970 -25724
rect -10892 -25872 -6064 -25824
rect -11090 -25945 -11008 -25934
rect -11090 -26005 -11079 -25945
rect -11019 -26005 -11008 -25945
rect -11090 -26016 -11008 -26005
rect -12499 -26511 -12373 -26465
rect -6112 -26420 -6064 -25872
rect -6018 -26332 -5970 -25772
rect -5854 -25742 -5802 -25736
rect -5802 -25792 4004 -25744
rect -5854 -25800 -5802 -25794
rect -3088 -25958 -3082 -25874
rect -2998 -25958 3902 -25874
rect 314 -26148 320 -26064
rect 404 -26148 3740 -26064
rect -6018 -26380 3558 -26332
rect -6112 -26468 3472 -26420
rect -12770 -26744 -12612 -26742
rect -12770 -26805 -12743 -26744
rect -12682 -26805 -12612 -26744
rect -12770 -26806 -12612 -26805
rect -12794 -26998 -12748 -26934
rect -12684 -26998 -12636 -26934
rect -12499 -27976 -12373 -27934
rect -12499 -29098 -12471 -27976
rect -12399 -29098 -12373 -27976
rect -11090 -28578 -11008 -28567
rect -11090 -28638 -11079 -28578
rect -11019 -28638 -11008 -28578
rect -11090 -28649 -11008 -28638
rect -12499 -29144 -12373 -29098
rect -12758 -29446 -12724 -29374
rect -12652 -29446 -12598 -29374
rect -12772 -29537 -12586 -29520
rect -12772 -29626 -12727 -29537
rect -12638 -29626 -12586 -29537
rect -12499 -30585 -12373 -30543
rect -12499 -31707 -12471 -30585
rect -12399 -31707 -12373 -30585
rect -11090 -31187 -11008 -31176
rect -11090 -31247 -11079 -31187
rect -11019 -31247 -11008 -31187
rect -11090 -31258 -11008 -31247
rect -12499 -31753 -12373 -31707
rect -12834 -31918 -12670 -31900
rect -12834 -31990 -12758 -31918
rect -12686 -31990 -12670 -31918
rect -12838 -32087 -12674 -32086
rect -12838 -32176 -12791 -32087
rect -12702 -32176 -12674 -32087
rect -9857 -32916 -9764 -32910
rect -9764 -33009 3112 -32916
rect -9857 -33015 -9764 -33009
rect -12501 -33205 -12375 -33163
rect -6038 -33168 -6032 -33116
rect -5980 -33118 -5974 -33116
rect -5980 -33166 2846 -33118
rect -5980 -33168 -5974 -33166
rect -12501 -34327 -12473 -33205
rect -12401 -34327 -12375 -33205
rect -3266 -33356 -3260 -33272
rect -3176 -33356 2696 -33272
rect -704 -33578 -698 -33494
rect -614 -33578 2428 -33494
rect -11092 -33807 -11010 -33796
rect -11092 -33867 -11081 -33807
rect -11021 -33867 -11010 -33807
rect -11092 -33878 -11010 -33867
rect -12501 -34373 -12375 -34327
rect -12582 -34504 -12510 -34498
rect -12582 -34582 -12510 -34576
rect -12746 -34671 -12582 -34670
rect -12746 -34760 -12726 -34671
rect -12637 -34760 -12582 -34671
rect 2344 -35454 2428 -33578
rect 2612 -35333 2696 -33356
rect 2798 -35235 2846 -33166
rect 3025 -35113 3091 -33009
rect 3424 -34011 3472 -26468
rect 3510 -33907 3558 -26380
rect 3656 -30926 3740 -26148
rect 3818 -30805 3902 -25958
rect 3956 -30722 4004 -25792
rect 4122 -30562 4226 -25634
rect 4306 -29500 4354 -25416
rect 4414 -29390 4462 -25290
rect 4651 -26398 4717 -22780
rect 4783 -26277 4849 -22610
rect 4894 -26179 4942 -22454
rect 4983 -26057 5069 -22299
rect 5118 -24962 5166 -22148
rect 5232 -24861 5277 -22065
rect 6849 -22044 8206 -22005
rect 8396 -22007 8405 -21972
rect 8461 -22007 8470 -21972
rect 8396 -22036 8401 -22007
rect 6780 -22066 6849 -22060
rect 6066 -22094 6132 -22088
rect 6132 -22103 8139 -22094
rect 6132 -22155 8079 -22103
rect 8131 -22155 8139 -22103
rect 8167 -22113 8206 -22044
rect 8465 -22036 8470 -22007
rect 8615 -22066 8993 -22000
rect 9059 -22066 9065 -22000
rect 10264 -22007 10324 -22001
rect 10257 -22065 10264 -22009
rect 10324 -22065 10331 -22009
rect 8401 -22077 8465 -22071
rect 8616 -22113 8655 -22066
rect 10264 -22073 10324 -22067
rect 8167 -22152 8655 -22113
rect 6132 -22160 8139 -22155
rect 8992 -22160 9001 -22094
rect 9067 -22160 9076 -22094
rect 9931 -22159 9937 -22093
rect 10003 -22159 10012 -22093
rect 10387 -22094 10453 -21941
rect 10522 -22000 10588 -21849
rect 10638 -21906 10704 -21717
rect 12467 -21820 13186 -21661
rect 12796 -21853 13186 -21820
rect 10638 -21972 10850 -21906
rect 10916 -21972 10922 -21906
rect 10522 -22066 10888 -22000
rect 10954 -22066 10963 -22000
rect 10387 -22160 10859 -22094
rect 10925 -22160 10931 -22094
rect 6066 -22166 6132 -22160
rect 6934 -22254 6941 -22188
rect 7007 -22197 10062 -22188
rect 7007 -22249 8063 -22197
rect 8128 -22249 8992 -22197
rect 9057 -22249 9951 -22197
rect 10016 -22249 10062 -22197
rect 7007 -22254 10062 -22249
rect 6941 -22260 7007 -22254
rect 11883 -22473 12147 -22462
rect 11883 -22715 11894 -22473
rect 12136 -22715 12147 -22473
rect 11883 -22726 12147 -22715
rect 5558 -23100 5627 -23040
rect 5998 -23090 6067 -23040
rect 6438 -23065 6507 -23040
rect 5554 -23159 5563 -23100
rect 5622 -23159 5631 -23100
rect 5994 -23149 6003 -23090
rect 6062 -23149 6071 -23090
rect 6438 -23124 6448 -23065
rect 6507 -23124 6516 -23065
rect 5558 -23289 5627 -23159
rect 5998 -23289 6067 -23149
rect 6438 -23289 6507 -23124
rect 5552 -23358 5558 -23289
rect 5627 -23358 5633 -23289
rect 5992 -23358 5998 -23289
rect 6067 -23358 6073 -23289
rect 6432 -23358 6438 -23289
rect 6507 -23358 6513 -23289
rect 5901 -23743 7113 -23674
rect 5901 -23854 5970 -23743
rect 5703 -23938 5823 -23910
rect 5901 -23929 5970 -23923
rect 6158 -23919 6236 -23909
rect 5703 -23994 5732 -23938
rect 5788 -23994 5823 -23938
rect 6158 -23975 6170 -23919
rect 6226 -23975 6236 -23919
rect 6335 -23925 6341 -23856
rect 6410 -23925 6416 -23856
rect 6580 -23910 6700 -23894
rect 6158 -23990 6236 -23975
rect 5703 -24023 5823 -23994
rect 6341 -24135 6410 -23925
rect 6580 -23966 6610 -23910
rect 6666 -23966 6700 -23910
rect 6580 -24007 6700 -23966
rect 6299 -24194 6410 -24135
rect 6299 -24293 6367 -24194
rect 6295 -24351 6304 -24293
rect 6362 -24351 6371 -24293
rect 7044 -24298 7113 -23743
rect 7044 -24307 10140 -24298
rect 6299 -24356 6367 -24351
rect 7044 -24359 7106 -24307
rect 7158 -24308 9002 -24307
rect 7158 -24359 8069 -24308
rect 7044 -24360 8069 -24359
rect 8122 -24359 9002 -24308
rect 9055 -24359 9933 -24307
rect 9986 -24359 10140 -24307
rect 8122 -24360 10140 -24359
rect 7044 -24367 10140 -24360
rect 12187 -24299 12431 -24288
rect 12187 -24307 12198 -24299
rect 5992 -24393 6073 -24387
rect 5992 -24462 5998 -24393
rect 6067 -24398 6073 -24393
rect 6067 -24400 8115 -24398
rect 6067 -24401 8057 -24400
rect 6067 -24453 7113 -24401
rect 7165 -24452 8057 -24401
rect 8109 -24452 8115 -24400
rect 7165 -24453 8115 -24452
rect 6067 -24457 8115 -24453
rect 8182 -24448 8914 -24395
rect 9929 -24401 10000 -24399
rect 6067 -24462 6073 -24457
rect 5992 -24468 6073 -24462
rect 7321 -24490 7393 -24485
rect 8182 -24490 8248 -24448
rect 6429 -24528 6516 -24519
rect 6429 -24597 6438 -24528
rect 6507 -24597 6516 -24528
rect 7321 -24556 7327 -24490
rect 7393 -24556 8248 -24490
rect 8424 -24483 8493 -24477
rect 8861 -24496 8914 -24448
rect 8989 -24459 8998 -24403
rect 9054 -24459 9063 -24403
rect 9923 -24457 9935 -24401
rect 9991 -24457 10000 -24401
rect 10256 -24452 10336 -24446
rect 9929 -24463 9993 -24457
rect 8541 -24528 8600 -24524
rect 8493 -24533 8605 -24528
rect 8493 -24535 8541 -24533
rect 7321 -24562 7393 -24556
rect 8424 -24592 8541 -24535
rect 8600 -24592 8605 -24533
rect 8861 -24549 8989 -24496
rect 9042 -24549 9048 -24496
rect 10256 -24521 10262 -24452
rect 10331 -24521 10336 -24452
rect 10256 -24528 10336 -24521
rect 10405 -24462 10860 -24396
rect 10926 -24462 10932 -24396
rect 8424 -24597 8605 -24592
rect 6429 -24606 6516 -24597
rect 8541 -24601 8600 -24597
rect 10405 -24606 10471 -24462
rect 5726 -24715 5732 -24649
rect 5798 -24715 8986 -24649
rect 9052 -24715 9058 -24649
rect 9792 -24672 9798 -24606
rect 9864 -24672 10471 -24606
rect 10536 -24556 10858 -24490
rect 10924 -24556 10930 -24490
rect 12187 -24510 12189 -24307
rect 12187 -24521 12198 -24510
rect 12420 -24521 12441 -24299
rect 12187 -24532 12431 -24521
rect 5311 -24811 5317 -24745
rect 5383 -24811 9917 -24745
rect 9983 -24811 9989 -24745
rect 5732 -24861 7106 -24851
rect 5232 -24906 7106 -24861
rect 5732 -24917 7106 -24906
rect 7172 -24917 7178 -24851
rect 10536 -24854 10602 -24556
rect 8812 -24920 8818 -24854
rect 8884 -24920 10602 -24854
rect 10659 -24650 10850 -24584
rect 10915 -24650 10921 -24584
rect 5732 -24962 8050 -24955
rect 5118 -25010 8050 -24962
rect 5732 -25021 8050 -25010
rect 8116 -25021 8122 -24955
rect 10659 -25108 10725 -24650
rect 7866 -25174 7872 -25108
rect 7938 -25174 10725 -25108
rect 7156 -25453 11207 -25381
rect 7156 -25631 7227 -25453
rect 7405 -25631 8162 -25453
rect 8340 -25631 9098 -25453
rect 9276 -25630 10029 -25453
rect 10206 -25630 10956 -25453
rect 9276 -25631 10956 -25630
rect 11134 -25631 11207 -25453
rect 7156 -25702 11207 -25631
rect 12414 -25872 12821 -25760
rect 12128 -25876 12821 -25872
rect 7847 -25967 7853 -25901
rect 7919 -25967 10121 -25901
rect 4983 -26123 8989 -26057
rect 9055 -26123 9061 -26057
rect 10055 -26179 10121 -25967
rect 12128 -25902 13042 -25876
rect 12128 -25964 13186 -25902
rect 12128 -26083 12233 -25964
rect 12352 -26005 13186 -25964
rect 12352 -26083 12960 -26005
rect 12128 -26124 12960 -26083
rect 13079 -26124 13186 -26005
rect 4894 -26228 9917 -26179
rect 4899 -26245 9917 -26228
rect 9983 -26245 9989 -26179
rect 10055 -26245 10704 -26179
rect 12128 -26189 13186 -26124
rect 4783 -26343 7102 -26277
rect 7168 -26343 7174 -26277
rect 8831 -26377 8837 -26311
rect 8903 -26377 10588 -26311
rect 4651 -26464 8050 -26398
rect 8116 -26464 8122 -26398
rect 9801 -26469 9807 -26405
rect 9873 -26469 10453 -26405
rect 8396 -26500 8470 -26494
rect 6780 -26519 6849 -26513
rect 6849 -26572 8206 -26533
rect 8396 -26535 8405 -26500
rect 8461 -26535 8470 -26500
rect 8396 -26564 8401 -26535
rect 6780 -26594 6849 -26588
rect 6066 -26622 6132 -26616
rect 6132 -26631 8139 -26622
rect 6132 -26683 8079 -26631
rect 8131 -26683 8139 -26631
rect 8167 -26641 8206 -26572
rect 8465 -26564 8470 -26535
rect 8615 -26594 8993 -26528
rect 9059 -26594 9065 -26528
rect 10264 -26535 10324 -26529
rect 10257 -26593 10264 -26537
rect 10324 -26593 10331 -26537
rect 8401 -26605 8465 -26599
rect 8616 -26641 8655 -26594
rect 10264 -26601 10324 -26595
rect 8167 -26680 8655 -26641
rect 6132 -26688 8139 -26683
rect 8992 -26688 9001 -26622
rect 9067 -26688 9076 -26622
rect 9931 -26687 9937 -26621
rect 10003 -26687 10012 -26621
rect 10387 -26622 10453 -26469
rect 10522 -26528 10588 -26377
rect 10638 -26434 10704 -26245
rect 12467 -26348 13186 -26189
rect 12796 -26381 13186 -26348
rect 10638 -26500 10850 -26434
rect 10916 -26500 10922 -26434
rect 10522 -26594 10888 -26528
rect 10954 -26594 10963 -26528
rect 10387 -26688 10859 -26622
rect 10925 -26688 10931 -26622
rect 6066 -26694 6132 -26688
rect 6934 -26782 6941 -26716
rect 7007 -26725 10062 -26716
rect 7007 -26777 8063 -26725
rect 8128 -26777 8992 -26725
rect 9057 -26777 9951 -26725
rect 10016 -26777 10062 -26725
rect 7007 -26782 10062 -26777
rect 6941 -26788 7007 -26782
rect 11883 -27001 12147 -26990
rect 11883 -27243 11894 -27001
rect 12136 -27243 12147 -27001
rect 11883 -27254 12147 -27243
rect 5558 -27640 5627 -27568
rect 5998 -27635 6067 -27568
rect 6438 -27581 6507 -27568
rect 5554 -27699 5563 -27640
rect 5622 -27699 5631 -27640
rect 5994 -27694 6003 -27635
rect 6062 -27694 6071 -27635
rect 6429 -27640 6438 -27581
rect 6497 -27640 6507 -27581
rect 5558 -27817 5627 -27699
rect 5998 -27817 6067 -27694
rect 6438 -27817 6507 -27640
rect 5552 -27886 5558 -27817
rect 5627 -27886 5633 -27817
rect 5992 -27886 5998 -27817
rect 6067 -27886 6073 -27817
rect 6432 -27886 6438 -27817
rect 6507 -27886 6513 -27817
rect 5901 -28271 7113 -28202
rect 5901 -28382 5970 -28271
rect 5703 -28466 5823 -28438
rect 5901 -28457 5970 -28451
rect 6158 -28447 6236 -28437
rect 5703 -28522 5732 -28466
rect 5788 -28522 5823 -28466
rect 6158 -28503 6170 -28447
rect 6226 -28503 6236 -28447
rect 6335 -28453 6341 -28384
rect 6410 -28453 6416 -28384
rect 6580 -28438 6700 -28422
rect 6158 -28518 6236 -28503
rect 5703 -28551 5823 -28522
rect 6341 -28663 6410 -28453
rect 6580 -28494 6610 -28438
rect 6666 -28494 6700 -28438
rect 6580 -28535 6700 -28494
rect 6299 -28722 6410 -28663
rect 6299 -28821 6367 -28722
rect 6295 -28879 6304 -28821
rect 6362 -28879 6371 -28821
rect 7044 -28826 7113 -28271
rect 7044 -28835 10140 -28826
rect 6299 -28884 6367 -28879
rect 7044 -28887 7106 -28835
rect 7158 -28836 9002 -28835
rect 7158 -28887 8069 -28836
rect 7044 -28888 8069 -28887
rect 8122 -28887 9002 -28836
rect 9055 -28887 9933 -28835
rect 9986 -28887 10140 -28835
rect 8122 -28888 10140 -28887
rect 7044 -28895 10140 -28888
rect 12187 -28827 12431 -28816
rect 12187 -28835 12198 -28827
rect 5992 -28921 6073 -28915
rect 5992 -28990 5998 -28921
rect 6067 -28926 6073 -28921
rect 6067 -28928 8115 -28926
rect 6067 -28929 8057 -28928
rect 6067 -28981 7113 -28929
rect 7165 -28980 8057 -28929
rect 8109 -28980 8115 -28928
rect 7165 -28981 8115 -28980
rect 6067 -28985 8115 -28981
rect 8182 -28976 8914 -28923
rect 9929 -28929 10000 -28927
rect 6067 -28990 6073 -28985
rect 5992 -28996 6073 -28990
rect 7321 -29018 7393 -29013
rect 8182 -29018 8248 -28976
rect 6429 -29056 6516 -29047
rect 6429 -29125 6438 -29056
rect 6507 -29125 6516 -29056
rect 7321 -29084 7327 -29018
rect 7393 -29084 8248 -29018
rect 8424 -29011 8493 -29005
rect 8861 -29024 8914 -28976
rect 8989 -28987 8998 -28931
rect 9054 -28987 9063 -28931
rect 9923 -28985 9935 -28929
rect 9991 -28985 10000 -28929
rect 10256 -28980 10336 -28974
rect 9929 -28991 9993 -28985
rect 8541 -29056 8600 -29052
rect 8493 -29061 8605 -29056
rect 8493 -29063 8541 -29061
rect 7321 -29090 7393 -29084
rect 8424 -29120 8541 -29063
rect 8600 -29120 8605 -29061
rect 8861 -29077 8989 -29024
rect 9042 -29077 9048 -29024
rect 10256 -29049 10262 -28980
rect 10331 -29049 10336 -28980
rect 10256 -29056 10336 -29049
rect 10405 -28990 10860 -28924
rect 10926 -28990 10932 -28924
rect 8424 -29125 8605 -29120
rect 6429 -29134 6516 -29125
rect 8541 -29129 8600 -29125
rect 10405 -29134 10471 -28990
rect 5448 -29243 5454 -29177
rect 5520 -29243 8986 -29177
rect 9052 -29243 9058 -29177
rect 9792 -29200 9798 -29134
rect 9864 -29200 10471 -29134
rect 10536 -29084 10858 -29018
rect 10924 -29084 10930 -29018
rect 12187 -29038 12189 -28835
rect 12187 -29049 12198 -29038
rect 12420 -29049 12441 -28827
rect 12187 -29060 12431 -29049
rect 4860 -29273 4919 -29272
rect 4860 -29278 9917 -29273
rect 4919 -29337 9917 -29278
rect 4860 -29339 9917 -29337
rect 9983 -29339 9989 -29273
rect 4860 -29343 4919 -29339
rect 5732 -29390 7106 -29379
rect 4414 -29438 7106 -29390
rect 5732 -29445 7106 -29438
rect 7172 -29445 7178 -29379
rect 10536 -29382 10602 -29084
rect 8812 -29448 8818 -29382
rect 8884 -29448 10602 -29382
rect 10659 -29178 10850 -29112
rect 10915 -29178 10921 -29112
rect 5732 -29500 8050 -29483
rect 4306 -29548 8050 -29500
rect 5732 -29549 8050 -29548
rect 8116 -29549 8122 -29483
rect 10659 -29636 10725 -29178
rect 7866 -29702 7872 -29636
rect 7938 -29702 10725 -29636
rect 7156 -29981 11207 -29909
rect 7156 -30159 7227 -29981
rect 7405 -30159 8162 -29981
rect 8340 -30159 9098 -29981
rect 9276 -30158 10029 -29981
rect 10206 -30158 10956 -29981
rect 9276 -30159 10956 -30158
rect 11134 -30159 11207 -29981
rect 7156 -30230 11207 -30159
rect 12414 -30400 12821 -30288
rect 12128 -30404 12821 -30400
rect 7847 -30495 7853 -30429
rect 7919 -30495 10121 -30429
rect 4122 -30585 5856 -30562
rect 4122 -30651 8989 -30585
rect 9055 -30651 9061 -30585
rect 4122 -30666 5856 -30651
rect 10055 -30707 10121 -30495
rect 12128 -30430 13042 -30404
rect 12128 -30492 13186 -30430
rect 12128 -30611 12233 -30492
rect 12352 -30533 13186 -30492
rect 12352 -30611 12960 -30533
rect 12128 -30652 12960 -30611
rect 13079 -30652 13186 -30533
rect 5732 -30722 9917 -30707
rect 3956 -30770 9917 -30722
rect 5732 -30773 9917 -30770
rect 9983 -30773 9989 -30707
rect 10055 -30773 10704 -30707
rect 12128 -30717 13186 -30652
rect 3818 -30871 7102 -30805
rect 7168 -30871 7174 -30805
rect 3818 -30874 3902 -30871
rect 8831 -30905 8837 -30839
rect 8903 -30905 10588 -30839
rect 3656 -30992 8050 -30926
rect 8116 -30992 8122 -30926
rect 3656 -30994 3740 -30992
rect 9801 -30997 9807 -30933
rect 9873 -30997 10453 -30933
rect 8396 -31028 8470 -31022
rect 6780 -31047 6849 -31041
rect 6849 -31100 8206 -31061
rect 8396 -31063 8405 -31028
rect 8461 -31063 8470 -31028
rect 8396 -31092 8401 -31063
rect 6780 -31122 6849 -31116
rect 6066 -31150 6132 -31144
rect 6132 -31159 8139 -31150
rect 6132 -31211 8079 -31159
rect 8131 -31211 8139 -31159
rect 8167 -31169 8206 -31100
rect 8465 -31092 8470 -31063
rect 8615 -31122 8993 -31056
rect 9059 -31122 9065 -31056
rect 10264 -31063 10324 -31057
rect 10257 -31121 10264 -31065
rect 10324 -31121 10331 -31065
rect 8401 -31133 8465 -31127
rect 8616 -31169 8655 -31122
rect 10264 -31129 10324 -31123
rect 8167 -31208 8655 -31169
rect 6132 -31216 8139 -31211
rect 8992 -31216 9001 -31150
rect 9067 -31216 9076 -31150
rect 9931 -31215 9937 -31149
rect 10003 -31215 10012 -31149
rect 10387 -31150 10453 -30997
rect 10522 -31056 10588 -30905
rect 10638 -30962 10704 -30773
rect 12467 -30876 13186 -30717
rect 12796 -30909 13186 -30876
rect 10638 -31028 10850 -30962
rect 10916 -31028 10922 -30962
rect 10522 -31122 10888 -31056
rect 10954 -31122 10963 -31056
rect 10387 -31216 10859 -31150
rect 10925 -31216 10931 -31150
rect 6066 -31222 6132 -31216
rect 6934 -31310 6941 -31244
rect 7007 -31253 10062 -31244
rect 7007 -31305 8063 -31253
rect 8128 -31305 8992 -31253
rect 9057 -31305 9951 -31253
rect 10016 -31305 10062 -31253
rect 7007 -31310 10062 -31305
rect 6941 -31316 7007 -31310
rect 11883 -31529 12147 -31518
rect 11883 -31771 11894 -31529
rect 12136 -31771 12147 -31529
rect 11883 -31782 12147 -31771
rect 5558 -32149 5627 -32096
rect 5554 -32208 5563 -32149
rect 5622 -32208 5631 -32149
rect 5998 -32164 6067 -32096
rect 6438 -32131 6507 -32096
rect 5558 -32345 5627 -32208
rect 5994 -32223 6003 -32164
rect 6062 -32223 6071 -32164
rect 5998 -32345 6067 -32223
rect 6438 -32345 6507 -32201
rect 5552 -32414 5558 -32345
rect 5627 -32414 5633 -32345
rect 5992 -32414 5998 -32345
rect 6067 -32414 6073 -32345
rect 6432 -32414 6438 -32345
rect 6507 -32414 6513 -32345
rect 5901 -32799 7113 -32730
rect 5901 -32910 5970 -32799
rect 5703 -32994 5823 -32966
rect 5901 -32985 5970 -32979
rect 6158 -32975 6236 -32965
rect 5703 -33050 5732 -32994
rect 5788 -33050 5823 -32994
rect 6158 -33031 6170 -32975
rect 6226 -33031 6236 -32975
rect 6335 -32981 6341 -32912
rect 6410 -32981 6416 -32912
rect 6580 -32966 6700 -32950
rect 6158 -33046 6236 -33031
rect 5703 -33079 5823 -33050
rect 6341 -33191 6410 -32981
rect 6580 -33022 6610 -32966
rect 6666 -33022 6700 -32966
rect 6580 -33063 6700 -33022
rect 6299 -33250 6410 -33191
rect 6299 -33349 6367 -33250
rect 6295 -33407 6304 -33349
rect 6362 -33407 6371 -33349
rect 7044 -33354 7113 -32799
rect 7044 -33363 10140 -33354
rect 6299 -33412 6367 -33407
rect 7044 -33415 7106 -33363
rect 7158 -33364 9002 -33363
rect 7158 -33415 8069 -33364
rect 7044 -33416 8069 -33415
rect 8122 -33415 9002 -33364
rect 9055 -33415 9933 -33363
rect 9986 -33415 10140 -33363
rect 8122 -33416 10140 -33415
rect 7044 -33423 10140 -33416
rect 12187 -33355 12431 -33344
rect 12187 -33363 12198 -33355
rect 5992 -33449 6073 -33443
rect 5992 -33518 5998 -33449
rect 6067 -33454 6073 -33449
rect 6067 -33456 8115 -33454
rect 6067 -33457 8057 -33456
rect 6067 -33509 7113 -33457
rect 7165 -33508 8057 -33457
rect 8109 -33508 8115 -33456
rect 7165 -33509 8115 -33508
rect 6067 -33513 8115 -33509
rect 8182 -33504 8914 -33451
rect 9929 -33457 10000 -33455
rect 6067 -33518 6073 -33513
rect 5992 -33524 6073 -33518
rect 7321 -33546 7393 -33541
rect 8182 -33546 8248 -33504
rect 6429 -33584 6516 -33575
rect 6429 -33653 6438 -33584
rect 6507 -33653 6516 -33584
rect 7321 -33612 7327 -33546
rect 7393 -33612 8248 -33546
rect 8424 -33539 8493 -33533
rect 8861 -33552 8914 -33504
rect 8989 -33515 8998 -33459
rect 9054 -33515 9063 -33459
rect 9923 -33513 9935 -33457
rect 9991 -33513 10000 -33457
rect 10256 -33508 10336 -33502
rect 9929 -33519 9993 -33513
rect 8541 -33584 8600 -33580
rect 8493 -33589 8605 -33584
rect 8493 -33591 8541 -33589
rect 7321 -33618 7393 -33612
rect 8424 -33648 8541 -33591
rect 8600 -33648 8605 -33589
rect 8861 -33605 8989 -33552
rect 9042 -33605 9048 -33552
rect 10256 -33577 10262 -33508
rect 10331 -33577 10336 -33508
rect 10256 -33584 10336 -33577
rect 10405 -33518 10860 -33452
rect 10926 -33518 10932 -33452
rect 8424 -33653 8605 -33648
rect 6429 -33662 6516 -33653
rect 8541 -33657 8600 -33653
rect 10405 -33662 10471 -33518
rect 5419 -33771 5425 -33705
rect 5491 -33771 8986 -33705
rect 9052 -33771 9058 -33705
rect 9792 -33728 9798 -33662
rect 9864 -33728 10471 -33662
rect 10536 -33612 10858 -33546
rect 10924 -33612 10930 -33546
rect 12187 -33566 12189 -33363
rect 12187 -33577 12198 -33566
rect 12420 -33577 12441 -33355
rect 12187 -33588 12431 -33577
rect 3657 -33867 3663 -33801
rect 3729 -33867 9917 -33801
rect 9983 -33867 9989 -33801
rect 3510 -33958 7106 -33907
rect 3511 -33973 7106 -33958
rect 7172 -33973 7178 -33907
rect 10536 -33910 10602 -33612
rect 8812 -33976 8818 -33910
rect 8884 -33976 10602 -33910
rect 10659 -33706 10850 -33640
rect 10915 -33706 10921 -33640
rect 3424 -34077 8050 -34011
rect 8116 -34077 8122 -34011
rect 3424 -34082 3756 -34077
rect 10659 -34164 10725 -33706
rect 7866 -34230 7872 -34164
rect 7938 -34230 10725 -34164
rect 7156 -34509 11207 -34437
rect 7156 -34687 7227 -34509
rect 7405 -34687 8162 -34509
rect 8340 -34687 9098 -34509
rect 9276 -34686 10029 -34509
rect 10206 -34686 10956 -34509
rect 9276 -34687 10956 -34686
rect 11134 -34687 11207 -34509
rect 7156 -34758 11207 -34687
rect 12414 -34928 12821 -34816
rect 12128 -34932 12821 -34928
rect 7847 -35023 7853 -34957
rect 7919 -35023 10121 -34957
rect 3025 -35179 8989 -35113
rect 9055 -35179 9061 -35113
rect 10055 -35235 10121 -35023
rect 12128 -34958 13042 -34932
rect 12128 -35020 13186 -34958
rect 12128 -35139 12233 -35020
rect 12352 -35061 13186 -35020
rect 12352 -35139 12960 -35061
rect 12128 -35180 12960 -35139
rect 13079 -35180 13186 -35061
rect 2789 -35301 9917 -35235
rect 9983 -35301 9989 -35235
rect 10055 -35301 10704 -35235
rect 12128 -35245 13186 -35180
rect 2612 -35399 7102 -35333
rect 7168 -35399 7174 -35333
rect 2612 -35400 2696 -35399
rect 8831 -35433 8837 -35367
rect 8903 -35433 10588 -35367
rect 2328 -35520 8050 -35454
rect 8116 -35520 8122 -35454
rect 9801 -35525 9807 -35461
rect 9873 -35525 10453 -35461
rect 8396 -35556 8470 -35550
rect 6780 -35575 6849 -35569
rect 6849 -35628 8206 -35589
rect 8396 -35591 8405 -35556
rect 8461 -35591 8470 -35556
rect 8396 -35620 8401 -35591
rect 6780 -35650 6849 -35644
rect 6066 -35678 6132 -35672
rect 6132 -35687 8139 -35678
rect 6132 -35739 8079 -35687
rect 8131 -35739 8139 -35687
rect 8167 -35697 8206 -35628
rect 8465 -35620 8470 -35591
rect 8615 -35650 8993 -35584
rect 9059 -35650 9065 -35584
rect 10264 -35591 10324 -35585
rect 10257 -35649 10264 -35593
rect 10324 -35649 10331 -35593
rect 8401 -35661 8465 -35655
rect 8616 -35697 8655 -35650
rect 10264 -35657 10324 -35651
rect 8167 -35736 8655 -35697
rect 6132 -35744 8139 -35739
rect 8992 -35744 9001 -35678
rect 9067 -35744 9076 -35678
rect 9931 -35743 9937 -35677
rect 10003 -35743 10012 -35677
rect 10387 -35678 10453 -35525
rect 10522 -35584 10588 -35433
rect 10638 -35490 10704 -35301
rect 12467 -35404 13186 -35245
rect 12796 -35437 13186 -35404
rect 10638 -35556 10850 -35490
rect 10916 -35556 10922 -35490
rect 10522 -35650 10888 -35584
rect 10954 -35650 10963 -35584
rect 10387 -35744 10859 -35678
rect 10925 -35744 10931 -35678
rect 6066 -35750 6132 -35744
rect 6934 -35838 6941 -35772
rect 7007 -35781 10062 -35772
rect 7007 -35833 8063 -35781
rect 8128 -35833 8992 -35781
rect 9057 -35833 9951 -35781
rect 10016 -35833 10062 -35781
rect 7007 -35838 10062 -35833
rect 6941 -35844 7007 -35838
rect 12549 -35955 12646 -35946
rect 11883 -36057 12147 -36046
rect 11883 -36299 11894 -36057
rect 12136 -36299 12147 -36057
rect 12549 -36061 12646 -36052
rect 13558 -35959 13662 -35950
rect 13558 -36072 13662 -36063
rect 11883 -36310 12147 -36299
<< via2 >>
rect -22627 7013 -22565 7075
rect -27520 4457 -27441 4536
rect -24000 4445 -22878 4517
rect -21811 6730 -21732 6809
rect -19307 6588 -19245 6650
rect -18524 6417 -18445 6496
rect -16014 6242 -15952 6304
rect 1841 6169 2963 6241
rect -15226 6071 -15147 6150
rect 3447 6169 4569 6241
rect 5151 6167 6273 6239
rect -12737 5911 -12675 5973
rect -11936 5705 -11857 5784
rect -9434 5546 -9372 5608
rect -8636 5402 -8557 5481
rect -6161 5274 -6101 5334
rect -5353 5123 -5268 5202
rect -2870 4961 -2808 5023
rect -2054 4797 -1975 4876
rect -20709 4445 -19587 4517
rect -17418 4445 -16296 4517
rect -14127 4445 -13005 4517
rect -10836 4445 -9714 4517
rect -7546 4445 -6424 4517
rect -4255 4445 -3133 4517
rect 2301 4789 2361 4849
rect 430 4684 492 4721
rect 430 4659 492 4684
rect -964 4445 158 4517
rect -23398 3065 -23338 3125
rect -24670 2661 -23548 2733
rect -23111 2661 -21989 2733
rect -24210 1281 -24150 1341
rect -24412 929 -24156 1001
rect -24046 518 -23963 666
rect -24336 255 -24001 259
rect -24336 203 -24001 255
rect -20107 3065 -20047 3125
rect -21379 2661 -20257 2733
rect -19820 2661 -18698 2733
rect -22651 1281 -22591 1341
rect -23123 929 -22867 1001
rect -22406 929 -22150 1001
rect -22628 375 -22483 450
rect -23100 188 -23038 250
rect -22235 223 -22179 225
rect -22235 171 -22233 223
rect -22233 171 -22181 223
rect -22181 171 -22179 223
rect -22235 169 -22179 171
rect -20919 1281 -20859 1341
rect -21121 929 -20865 1001
rect -20755 518 -20672 666
rect -21045 255 -20710 259
rect -21045 203 -20710 255
rect -16816 3065 -16756 3125
rect -18088 2661 -16966 2733
rect -16529 2661 -15407 2733
rect -19360 1281 -19300 1341
rect -19832 929 -19576 1001
rect -19115 929 -18859 1001
rect -19337 375 -19192 450
rect -19809 188 -19747 250
rect -18944 223 -18888 225
rect -18944 171 -18942 223
rect -18942 171 -18890 223
rect -18890 171 -18888 223
rect -18944 169 -18888 171
rect -17628 1281 -17568 1341
rect -17830 929 -17574 1001
rect -17464 518 -17381 666
rect -17754 255 -17419 259
rect -17754 203 -17419 255
rect -13525 3065 -13465 3125
rect -14797 2661 -13675 2733
rect -13238 2661 -12116 2733
rect -16069 1281 -16009 1341
rect -16541 929 -16285 1001
rect -15824 929 -15568 1001
rect -16046 375 -15901 450
rect -16518 188 -16456 250
rect -15653 223 -15597 225
rect -15653 171 -15651 223
rect -15651 171 -15599 223
rect -15599 171 -15597 223
rect -15653 169 -15597 171
rect -14337 1281 -14277 1341
rect -14539 929 -14283 1001
rect -14173 518 -14090 666
rect -14463 255 -14128 259
rect -14463 203 -14128 255
rect -10234 3065 -10174 3125
rect -11506 2661 -10384 2733
rect -9947 2661 -8825 2733
rect -12778 1281 -12718 1341
rect -13250 929 -12994 1001
rect -12533 929 -12277 1001
rect -12755 375 -12610 450
rect -13227 188 -13165 250
rect -12362 223 -12306 225
rect -12362 171 -12360 223
rect -12360 171 -12308 223
rect -12308 171 -12306 223
rect -12362 169 -12306 171
rect -11046 1281 -10986 1341
rect -11248 929 -10992 1001
rect -10882 518 -10799 666
rect -11172 255 -10837 259
rect -11172 203 -10837 255
rect -6944 3065 -6884 3125
rect -8216 2661 -7094 2733
rect -6657 2661 -5535 2733
rect -9487 1281 -9427 1341
rect -9959 929 -9703 1001
rect -9242 929 -8986 1001
rect -9464 375 -9319 450
rect -9936 188 -9874 250
rect -9071 223 -9015 225
rect -9071 171 -9069 223
rect -9069 171 -9017 223
rect -9017 171 -9015 223
rect -9071 169 -9015 171
rect -7756 1281 -7696 1341
rect -7958 929 -7702 1001
rect -7592 518 -7509 666
rect -7882 255 -7547 259
rect -7882 203 -7547 255
rect -3653 3065 -3593 3125
rect -4925 2661 -3803 2733
rect -3366 2661 -2244 2733
rect -6197 1281 -6137 1341
rect -6669 929 -6413 1001
rect -5952 929 -5696 1001
rect -6174 375 -6029 450
rect -6646 188 -6584 250
rect -5781 223 -5725 225
rect -5781 171 -5779 223
rect -5779 171 -5727 223
rect -5727 171 -5725 223
rect -5781 169 -5725 171
rect -4465 1281 -4405 1341
rect -4667 929 -4411 1001
rect -4301 518 -4218 666
rect -4591 255 -4256 259
rect -4591 203 -4256 255
rect -362 3065 -302 3125
rect -1634 2661 -512 2733
rect -75 2661 1047 2733
rect -2906 1281 -2846 1341
rect -3378 929 -3122 1001
rect -2661 929 -2405 1001
rect -2883 375 -2738 450
rect -3355 188 -3293 250
rect -2490 223 -2434 225
rect -2490 171 -2488 223
rect -2488 171 -2436 223
rect -2436 171 -2434 223
rect -2490 169 -2434 171
rect -1174 1281 -1114 1341
rect -1376 929 -1120 1001
rect -1010 518 -927 666
rect -1300 255 -965 259
rect -1300 203 -965 255
rect 385 1281 445 1341
rect -87 929 169 1001
rect 630 929 886 1001
rect 408 375 553 450
rect -64 188 -2 250
rect 801 223 857 225
rect 801 171 803 223
rect 803 171 855 223
rect 855 171 857 223
rect 801 169 857 171
rect 3907 4789 3967 4849
rect 5611 4787 5671 4847
rect 5558 4029 5627 4099
rect 5998 4029 6067 4099
rect 6445 4022 6504 4081
rect 5732 3228 5788 3230
rect 5732 3176 5734 3228
rect 5734 3176 5786 3228
rect 5786 3176 5788 3228
rect 5732 3174 5788 3176
rect 6170 3247 6226 3249
rect 6170 3195 6172 3247
rect 6172 3195 6224 3247
rect 6224 3195 6226 3247
rect 6170 3193 6226 3195
rect 6610 3256 6666 3258
rect 6610 3204 6612 3256
rect 6612 3204 6664 3256
rect 6664 3204 6666 3256
rect 6610 3202 6666 3204
rect 6304 2817 6362 2875
rect 12198 2861 12420 2869
rect 6438 2571 6507 2640
rect 8998 2763 9054 2765
rect 8998 2711 9000 2763
rect 9000 2711 9052 2763
rect 9052 2711 9054 2763
rect 8998 2709 9054 2711
rect 9935 2763 9991 2767
rect 9935 2711 9987 2763
rect 9987 2711 9991 2763
rect 8541 2576 8600 2635
rect 10267 2652 10326 2711
rect 12198 2658 12410 2861
rect 12410 2658 12420 2861
rect 12198 2647 12420 2658
rect 7227 1537 7405 1715
rect 8162 1537 8340 1715
rect 9098 1537 9276 1715
rect 10029 1538 10206 1715
rect 10956 1537 11134 1715
rect 12233 1085 12352 1204
rect 12960 1044 13079 1163
rect 8405 633 8461 668
rect 8405 612 8461 633
rect 10266 575 10322 631
rect 9001 480 9067 542
rect 9947 481 10003 542
rect 11894 -75 12136 167
rect 5563 -509 5622 -450
rect 6003 -483 6062 -424
rect 6443 -514 6502 -455
rect 5732 -1300 5788 -1298
rect 5732 -1352 5734 -1300
rect 5734 -1352 5786 -1300
rect 5786 -1352 5788 -1300
rect 5732 -1354 5788 -1352
rect 6170 -1281 6226 -1279
rect 6170 -1333 6172 -1281
rect 6172 -1333 6224 -1281
rect 6224 -1333 6226 -1281
rect 6170 -1335 6226 -1333
rect 6610 -1272 6666 -1270
rect 6610 -1324 6612 -1272
rect 6612 -1324 6664 -1272
rect 6664 -1324 6666 -1272
rect 6610 -1326 6666 -1324
rect 6304 -1711 6362 -1653
rect 12198 -1667 12420 -1659
rect 6438 -1957 6507 -1888
rect 8998 -1765 9054 -1763
rect 8998 -1817 9000 -1765
rect 9000 -1817 9052 -1765
rect 9052 -1817 9054 -1765
rect 8998 -1819 9054 -1817
rect 9935 -1765 9991 -1761
rect 9935 -1817 9987 -1765
rect 9987 -1817 9991 -1765
rect 8541 -1952 8600 -1893
rect 10267 -1876 10326 -1817
rect 12198 -1870 12410 -1667
rect 12410 -1870 12420 -1667
rect 12198 -1881 12420 -1870
rect -23605 -2304 -23436 -2225
rect -24410 -2467 -23856 -2327
rect -25216 -2591 -25155 -2529
rect -21585 -2304 -21416 -2225
rect -22373 -2467 -21819 -2327
rect -19844 -2304 -19675 -2225
rect -20643 -2467 -20089 -2327
rect -24550 -3165 -24428 -2987
rect -24184 -3057 -23844 -2983
rect -23601 -2974 -23452 -2878
rect -22594 -3080 -22431 -2852
rect -22147 -3057 -21807 -2983
rect -21581 -2974 -21432 -2878
rect -18065 -2304 -17896 -2225
rect -18883 -2467 -18329 -2327
rect -20917 -3165 -20741 -3042
rect -20417 -3057 -20077 -2983
rect -19840 -2974 -19691 -2878
rect -19241 -3087 -19043 -2934
rect -18657 -3057 -18317 -2983
rect -18061 -2974 -17912 -2878
rect -22600 -3848 -22476 -3742
rect -24807 -4337 -24618 -4064
rect -23561 -4116 -23392 -4037
rect -24359 -4279 -23805 -4139
rect -21823 -4116 -21654 -4037
rect -22623 -4279 -22069 -4139
rect -23195 -4594 -23064 -4480
rect -24133 -4869 -23793 -4795
rect -23557 -4786 -23408 -4690
rect -22397 -4869 -22057 -4795
rect -21819 -4786 -21670 -4690
rect -20603 -3899 -19481 -3827
rect -19044 -3899 -17922 -3827
rect -25504 -5097 -25442 -5035
rect -23563 -5408 -23394 -5329
rect -24359 -5571 -23805 -5431
rect -21829 -5408 -21660 -5329
rect -22623 -5571 -22069 -5431
rect -24612 -6247 -24466 -6049
rect -24133 -6161 -23793 -6087
rect -23559 -6078 -23410 -5982
rect -22862 -6046 -22773 -5995
rect -22862 -6441 -22773 -6046
rect -22397 -6161 -22057 -6087
rect -21825 -6078 -21676 -5982
rect -20143 -5279 -20083 -5219
rect -20345 -5631 -20089 -5559
rect -19979 -6042 -19896 -5894
rect -20269 -6305 -19934 -6301
rect -20269 -6357 -19934 -6305
rect -17312 -3899 -16190 -3827
rect -15753 -3899 -14631 -3827
rect -18584 -5279 -18524 -5219
rect -19056 -5631 -18800 -5559
rect -18339 -5631 -18083 -5559
rect -18561 -6185 -18416 -6110
rect -19033 -6372 -18971 -6310
rect -18168 -6337 -18112 -6335
rect -18168 -6389 -18166 -6337
rect -18166 -6389 -18114 -6337
rect -18114 -6389 -18112 -6337
rect -18168 -6391 -18112 -6389
rect -16852 -5279 -16792 -5219
rect -17054 -5631 -16798 -5559
rect -16688 -6042 -16605 -5894
rect -16978 -6305 -16643 -6301
rect -16978 -6357 -16643 -6305
rect -14021 -3899 -12899 -3827
rect -12462 -3899 -11340 -3827
rect -15293 -5279 -15233 -5219
rect -15765 -5631 -15509 -5559
rect -15048 -5631 -14792 -5559
rect -15270 -6185 -15125 -6110
rect -15742 -6372 -15680 -6310
rect -14877 -6337 -14821 -6335
rect -14877 -6389 -14875 -6337
rect -14875 -6389 -14823 -6337
rect -14823 -6389 -14821 -6337
rect -14877 -6391 -14821 -6389
rect -13561 -5279 -13501 -5219
rect -13763 -5631 -13507 -5559
rect -13397 -6042 -13314 -5894
rect -13687 -6305 -13352 -6301
rect -13687 -6357 -13352 -6305
rect -25655 -6832 -25576 -6751
rect -24619 -6824 -24490 -6684
rect -21515 -6818 -21386 -6678
rect -23562 -7381 -23393 -7302
rect -24359 -7544 -23805 -7404
rect -21827 -7381 -21658 -7302
rect -22622 -7544 -22068 -7404
rect -23198 -7745 -23067 -7743
rect -23198 -7857 -23064 -7745
rect -23195 -7859 -23064 -7857
rect -24133 -8134 -23793 -8060
rect -23558 -8051 -23409 -7955
rect -22396 -8134 -22056 -8060
rect -21823 -8051 -21674 -7955
rect -20603 -7164 -19481 -7092
rect -19044 -7164 -17922 -7092
rect -10730 -3899 -9608 -3827
rect -9171 -3899 -8049 -3827
rect -12002 -5279 -11942 -5219
rect -12474 -5631 -12218 -5559
rect -11757 -5631 -11501 -5559
rect -11979 -6185 -11834 -6110
rect -12451 -6372 -12389 -6310
rect -11586 -6337 -11530 -6335
rect -11586 -6389 -11584 -6337
rect -11584 -6389 -11532 -6337
rect -11532 -6389 -11530 -6337
rect -11586 -6391 -11530 -6389
rect -10270 -5279 -10210 -5219
rect -10472 -5631 -10216 -5559
rect -10106 -6042 -10023 -5894
rect -10396 -6305 -10061 -6301
rect -10396 -6357 -10061 -6305
rect -8711 -5279 -8651 -5219
rect -9183 -5631 -8927 -5559
rect -8466 -5631 -8210 -5559
rect -8688 -6185 -8543 -6110
rect -9160 -6372 -9098 -6310
rect -8295 -6337 -8239 -6335
rect -8295 -6389 -8293 -6337
rect -8293 -6389 -8241 -6337
rect -8241 -6389 -8239 -6337
rect -8295 -6391 -8239 -6389
rect -25809 -8362 -25749 -8302
rect -23560 -8673 -23391 -8594
rect -24359 -8836 -23805 -8696
rect -21823 -8673 -21654 -8594
rect -22623 -8836 -22069 -8696
rect -24612 -9512 -24466 -9314
rect -24133 -9426 -23793 -9352
rect -23556 -9343 -23407 -9247
rect -22866 -9260 -22777 -9239
rect -22866 -9303 -22773 -9260
rect -22866 -9685 -22773 -9303
rect -22397 -9426 -22057 -9352
rect -21819 -9343 -21670 -9247
rect -22862 -9706 -22773 -9685
rect -20143 -8544 -20083 -8484
rect -20345 -8896 -20089 -8824
rect -19979 -9307 -19896 -9159
rect -20269 -9570 -19934 -9566
rect -20269 -9622 -19934 -9570
rect -17312 -7164 -16190 -7092
rect -15753 -7164 -14631 -7092
rect -18584 -8544 -18524 -8484
rect -19056 -8896 -18800 -8824
rect -18339 -8896 -18083 -8824
rect -18561 -9450 -18416 -9375
rect -19033 -9637 -18971 -9575
rect -18168 -9602 -18112 -9600
rect -18168 -9654 -18166 -9602
rect -18166 -9654 -18114 -9602
rect -18114 -9654 -18112 -9602
rect -18168 -9656 -18112 -9654
rect -16852 -8544 -16792 -8484
rect -17054 -8896 -16798 -8824
rect -16688 -9307 -16605 -9159
rect -16978 -9570 -16643 -9566
rect -16978 -9622 -16643 -9570
rect -14021 -7164 -12899 -7092
rect -12462 -7164 -11340 -7092
rect -15293 -8544 -15233 -8484
rect -15765 -8896 -15509 -8824
rect -15048 -8896 -14792 -8824
rect -15270 -9450 -15125 -9375
rect -15742 -9637 -15680 -9575
rect -14877 -9602 -14821 -9600
rect -14877 -9654 -14875 -9602
rect -14875 -9654 -14823 -9602
rect -14823 -9654 -14821 -9602
rect -14877 -9656 -14821 -9654
rect -13561 -8544 -13501 -8484
rect -13763 -8896 -13507 -8824
rect -13397 -9307 -13314 -9159
rect -25978 -10241 -25899 -10160
rect -23560 -10645 -23391 -10566
rect -24359 -10808 -23805 -10668
rect -25365 -11055 -25286 -10976
rect -21827 -10645 -21658 -10566
rect -22622 -10808 -22068 -10668
rect -23198 -11121 -23061 -11007
rect -23195 -11123 -23064 -11121
rect -24133 -11398 -23793 -11324
rect -23556 -11315 -23407 -11219
rect -22396 -11398 -22056 -11324
rect -21823 -11315 -21674 -11219
rect -20603 -10428 -19481 -10356
rect -19044 -10428 -17922 -10356
rect -26164 -11653 -26102 -11591
rect -23560 -11937 -23391 -11858
rect -24359 -12100 -23805 -11960
rect -21831 -11937 -21662 -11858
rect -22622 -12100 -22068 -11960
rect -24612 -12776 -24466 -12578
rect -24133 -12690 -23793 -12616
rect -23556 -12607 -23407 -12511
rect -22866 -12518 -22777 -12503
rect -22869 -12524 -22777 -12518
rect -22869 -12964 -22773 -12524
rect -22396 -12690 -22056 -12616
rect -21827 -12607 -21678 -12511
rect -22862 -12970 -22773 -12964
rect -20143 -11808 -20083 -11748
rect -20345 -12160 -20089 -12088
rect -19979 -12571 -19896 -12423
rect -20269 -12834 -19934 -12830
rect -20269 -12886 -19934 -12834
rect -13687 -9570 -13352 -9566
rect -13687 -9622 -13352 -9570
rect -10730 -7164 -9608 -7092
rect -9171 -7164 -8049 -7092
rect -12002 -8544 -11942 -8484
rect -12474 -8896 -12218 -8824
rect -11757 -8896 -11501 -8824
rect -11979 -9450 -11834 -9375
rect -12451 -9637 -12389 -9575
rect -11586 -9602 -11530 -9600
rect -11586 -9654 -11584 -9602
rect -11584 -9654 -11532 -9602
rect -11532 -9654 -11530 -9602
rect -11586 -9656 -11530 -9654
rect -10270 -8544 -10210 -8484
rect -10472 -8896 -10216 -8824
rect -10106 -9307 -10023 -9159
rect -10396 -9570 -10061 -9566
rect -10396 -9622 -10061 -9570
rect -17312 -10428 -16190 -10356
rect -15753 -10428 -14631 -10356
rect -8711 -8544 -8651 -8484
rect -9183 -8896 -8927 -8824
rect -8466 -8896 -8210 -8824
rect -8688 -9450 -8543 -9375
rect -9160 -9637 -9098 -9575
rect -8295 -9602 -8239 -9600
rect -8295 -9654 -8293 -9602
rect -8293 -9654 -8241 -9602
rect -8241 -9654 -8239 -9602
rect -8295 -9656 -8239 -9654
rect -18584 -11808 -18524 -11748
rect -19056 -12160 -18800 -12088
rect -18339 -12160 -18083 -12088
rect -18561 -12714 -18416 -12639
rect -19033 -12901 -18971 -12839
rect -18168 -12866 -18112 -12864
rect -18168 -12918 -18166 -12866
rect -18166 -12918 -18114 -12866
rect -18114 -12918 -18112 -12866
rect -18168 -12920 -18112 -12918
rect -16852 -11808 -16792 -11748
rect -17054 -12160 -16798 -12088
rect -16688 -12571 -16605 -12423
rect -16978 -12834 -16643 -12830
rect -16978 -12886 -16643 -12834
rect -26327 -13144 -26248 -13063
rect -14021 -10428 -12899 -10356
rect -12462 -10428 -11340 -10356
rect -15293 -11808 -15233 -11748
rect -15765 -12160 -15509 -12088
rect -15048 -12160 -14792 -12088
rect -15270 -12714 -15125 -12639
rect -15742 -12901 -15680 -12839
rect -14877 -12866 -14821 -12864
rect -14877 -12918 -14875 -12866
rect -14875 -12918 -14823 -12866
rect -14823 -12918 -14821 -12866
rect -14877 -12920 -14821 -12918
rect -13561 -11808 -13501 -11748
rect -13763 -12160 -13507 -12088
rect -13397 -12571 -13314 -12423
rect -13687 -12834 -13352 -12830
rect -13687 -12886 -13352 -12834
rect -10730 -10428 -9608 -10356
rect -9171 -10428 -8049 -10356
rect -12002 -11808 -11942 -11748
rect -12474 -12160 -12218 -12088
rect -11757 -12160 -11501 -12088
rect -11979 -12714 -11834 -12639
rect -12451 -12901 -12389 -12839
rect -11586 -12866 -11530 -12864
rect -11586 -12918 -11584 -12866
rect -11584 -12918 -11532 -12866
rect -11532 -12918 -11530 -12866
rect -11586 -12920 -11530 -12918
rect -10270 -11808 -10210 -11748
rect -10472 -12160 -10216 -12088
rect -10106 -12571 -10023 -12423
rect -10396 -12834 -10061 -12830
rect -10396 -12886 -10061 -12834
rect -8711 -11808 -8651 -11748
rect -9183 -12160 -8927 -12088
rect -8466 -12160 -8210 -12088
rect -8688 -12714 -8543 -12639
rect -9160 -12901 -9098 -12839
rect -8295 -12866 -8239 -12864
rect -8295 -12918 -8293 -12866
rect -8293 -12918 -8241 -12866
rect -8241 -12918 -8239 -12866
rect -8295 -12920 -8239 -12918
rect -23421 -15176 -23320 -15075
rect -24839 -15290 -24743 -15194
rect -24916 -15658 -24844 -15586
rect -24903 -15828 -24812 -15739
rect -24835 -16464 -24739 -16368
rect -23378 -16372 -23277 -16271
rect -24908 -16842 -24836 -16770
rect -24915 -17012 -24836 -16923
rect -23369 -17584 -23268 -17483
rect -24829 -17696 -24733 -17600
rect -24921 -18054 -24851 -17984
rect 7227 -2991 7405 -2813
rect 8162 -2991 8340 -2813
rect 9098 -2991 9276 -2813
rect 10029 -2990 10206 -2813
rect 10956 -2991 11134 -2813
rect -24917 -18217 -24824 -18128
rect -21933 -18117 -21873 -18113
rect -21933 -18169 -21929 -18117
rect -21929 -18169 -21877 -18117
rect -21877 -18169 -21873 -18117
rect -21933 -18173 -21873 -18169
rect -20643 -18174 -20554 -18085
rect 12233 -3443 12352 -3324
rect 12960 -3484 13079 -3365
rect -24815 -18810 -24719 -18714
rect -23361 -18725 -23260 -18624
rect -21939 -18626 -21879 -18622
rect -21939 -18678 -21935 -18626
rect -21935 -18678 -21883 -18626
rect -21883 -18678 -21879 -18626
rect -21939 -18682 -21879 -18678
rect -20650 -18667 -20561 -18578
rect -18072 -15355 -17998 -15281
rect -16909 -15330 -16849 -15326
rect -16909 -15382 -16905 -15330
rect -16905 -15382 -16853 -15330
rect -16853 -15382 -16849 -15330
rect -16909 -15386 -16849 -15382
rect -12473 -15345 -12401 -14223
rect 8405 -3895 8461 -3860
rect 8405 -3916 8461 -3895
rect 10266 -3953 10322 -3897
rect 9001 -4048 9067 -3986
rect 9947 -4047 10003 -3986
rect 11894 -4603 12136 -4361
rect 5563 -4919 5622 -4860
rect 6003 -4939 6062 -4880
rect 6442 -4948 6501 -4889
rect 5732 -5728 5788 -5726
rect 5732 -5780 5734 -5728
rect 5734 -5780 5786 -5728
rect 5786 -5780 5788 -5728
rect 5732 -5782 5788 -5780
rect 6170 -5709 6226 -5707
rect 6170 -5761 6172 -5709
rect 6172 -5761 6224 -5709
rect 6224 -5761 6226 -5709
rect 6170 -5763 6226 -5761
rect 6610 -5700 6666 -5698
rect 6610 -5752 6612 -5700
rect 6612 -5752 6664 -5700
rect 6664 -5752 6666 -5700
rect 6610 -5754 6666 -5752
rect 6304 -6139 6362 -6081
rect 12198 -6095 12420 -6087
rect 6438 -6385 6507 -6316
rect 8998 -6193 9054 -6191
rect 8998 -6245 9000 -6193
rect 9000 -6245 9052 -6193
rect 9052 -6245 9054 -6193
rect 8998 -6247 9054 -6245
rect 9935 -6193 9991 -6189
rect 9935 -6245 9987 -6193
rect 9987 -6245 9991 -6193
rect 8541 -6380 8600 -6321
rect 10267 -6304 10326 -6245
rect 12198 -6298 12410 -6095
rect 12410 -6298 12420 -6095
rect 12198 -6309 12420 -6298
rect 7227 -7419 7405 -7241
rect 8162 -7419 8340 -7241
rect 9098 -7419 9276 -7241
rect 10029 -7418 10206 -7241
rect 10956 -7419 11134 -7241
rect 12233 -7871 12352 -7752
rect 12960 -7912 13079 -7793
rect 8405 -8323 8461 -8288
rect 8405 -8344 8461 -8323
rect 10266 -8381 10322 -8325
rect 9001 -8476 9067 -8414
rect 9947 -8475 10003 -8414
rect 11894 -9031 12136 -8789
rect 5563 -9582 5622 -9523
rect 6003 -9587 6062 -9528
rect 6445 -9573 6504 -9514
rect 5732 -10356 5788 -10354
rect 5732 -10408 5734 -10356
rect 5734 -10408 5786 -10356
rect 5786 -10408 5788 -10356
rect 5732 -10410 5788 -10408
rect 6170 -10337 6226 -10335
rect 6170 -10389 6172 -10337
rect 6172 -10389 6224 -10337
rect 6224 -10389 6226 -10337
rect 6170 -10391 6226 -10389
rect 6610 -10328 6666 -10326
rect 6610 -10380 6612 -10328
rect 6612 -10380 6664 -10328
rect 6664 -10380 6666 -10328
rect 6610 -10382 6666 -10380
rect 6304 -10767 6362 -10709
rect 12198 -10723 12420 -10715
rect 6438 -11013 6507 -10944
rect 8998 -10821 9054 -10819
rect 8998 -10873 9000 -10821
rect 9000 -10873 9052 -10821
rect 9052 -10873 9054 -10821
rect 8998 -10875 9054 -10873
rect 9935 -10821 9991 -10817
rect 9935 -10873 9987 -10821
rect 9987 -10873 9991 -10821
rect 8541 -11008 8600 -10949
rect 10267 -10932 10326 -10873
rect 12198 -10926 12410 -10723
rect 12410 -10926 12420 -10723
rect 12198 -10937 12420 -10926
rect 7227 -12047 7405 -11869
rect 8162 -12047 8340 -11869
rect 9098 -12047 9276 -11869
rect 10029 -12046 10206 -11869
rect 10956 -12047 11134 -11869
rect 12233 -12499 12352 -12380
rect 12960 -12540 13079 -12421
rect -11081 -14885 -11021 -14825
rect -17961 -15653 -17899 -15591
rect -12719 -15653 -12657 -15591
rect -18118 -15822 -18039 -15743
rect -12555 -15837 -12456 -15738
rect -5021 -14365 -4915 -14259
rect -5003 -14561 -4941 -14499
rect 8405 -12951 8461 -12916
rect 8405 -12972 8461 -12951
rect 10266 -13009 10322 -12953
rect 9001 -13104 9067 -13042
rect 9947 -13103 10003 -13042
rect -2304 -14167 -2200 -14063
rect -1288 -14171 -1191 -14074
rect -4004 -14347 -3907 -14250
rect -2283 -14561 -2221 -14499
rect -5020 -14991 -4916 -14887
rect -4004 -14980 -3907 -14883
rect -2304 -14986 -2200 -14882
rect -1288 -14990 -1191 -14893
rect -8494 -15429 -8434 -15425
rect -8494 -15481 -8490 -15429
rect -8490 -15481 -8438 -15429
rect -8438 -15481 -8434 -15429
rect -8494 -15485 -8434 -15481
rect -7204 -15486 -7115 -15397
rect -8671 -15563 -8609 -15501
rect -4961 -15373 -4899 -15311
rect -2259 -15373 -2197 -15311
rect -24870 -19175 -24798 -19103
rect -21939 -19109 -21879 -19105
rect -21939 -19161 -21935 -19109
rect -21935 -19161 -21883 -19109
rect -21883 -19161 -21879 -19109
rect -21939 -19165 -21879 -19161
rect -20651 -19153 -20562 -19064
rect -24875 -19345 -24796 -19256
rect -8500 -15938 -8440 -15934
rect -8500 -15990 -8496 -15938
rect -8496 -15990 -8444 -15938
rect -8444 -15990 -8440 -15938
rect -8500 -15994 -8440 -15990
rect -7211 -15979 -7122 -15890
rect -5020 -15810 -4916 -15706
rect -4004 -15799 -3907 -15702
rect -2304 -15805 -2200 -15701
rect -1288 -15809 -1191 -15712
rect 11894 -13659 12136 -13417
rect 5563 -14109 5622 -14050
rect 6003 -14093 6062 -14034
rect 6442 -14076 6501 -14017
rect 5732 -14884 5788 -14882
rect 5732 -14936 5734 -14884
rect 5734 -14936 5786 -14884
rect 5786 -14936 5788 -14884
rect 5732 -14938 5788 -14936
rect 6170 -14865 6226 -14863
rect 6170 -14917 6172 -14865
rect 6172 -14917 6224 -14865
rect 6224 -14917 6226 -14865
rect 6170 -14919 6226 -14917
rect 6610 -14856 6666 -14854
rect 6610 -14908 6612 -14856
rect 6612 -14908 6664 -14856
rect 6664 -14908 6666 -14856
rect 6610 -14910 6666 -14908
rect 6304 -15295 6362 -15237
rect 12198 -15251 12420 -15243
rect 6438 -15541 6507 -15472
rect 8998 -15349 9054 -15347
rect 8998 -15401 9000 -15349
rect 9000 -15401 9052 -15349
rect 9052 -15401 9054 -15349
rect 8998 -15403 9054 -15401
rect 9935 -15349 9991 -15345
rect 9935 -15401 9987 -15349
rect 9987 -15401 9991 -15349
rect 8541 -15536 8600 -15477
rect 10267 -15460 10326 -15401
rect 12198 -15454 12410 -15251
rect 12410 -15454 12420 -15251
rect 12198 -15465 12420 -15454
rect -8549 -16219 -8487 -16157
rect -4990 -16190 -4930 -16130
rect -2280 -16190 -2220 -16130
rect -8500 -16421 -8440 -16417
rect -8500 -16473 -8496 -16421
rect -8496 -16473 -8444 -16421
rect -8444 -16473 -8440 -16421
rect -8500 -16477 -8440 -16473
rect -7212 -16465 -7123 -16376
rect -5020 -16629 -4916 -16525
rect -4004 -16618 -3907 -16521
rect -2304 -16624 -2200 -16520
rect -1288 -16628 -1191 -16531
rect 7227 -16575 7405 -16397
rect 8162 -16575 8340 -16397
rect 9098 -16575 9276 -16397
rect 10029 -16574 10206 -16397
rect 10956 -16575 11134 -16397
rect -18084 -16757 -18010 -16683
rect -16909 -16735 -16849 -16732
rect -16909 -16789 -16906 -16735
rect -16906 -16789 -16852 -16735
rect -16852 -16789 -16849 -16735
rect -16909 -16792 -16849 -16789
rect -8551 -16754 -8482 -16685
rect -18077 -17047 -18015 -16985
rect -8500 -16943 -8440 -16939
rect -8500 -16995 -8496 -16943
rect -8496 -16995 -8444 -16943
rect -8444 -16995 -8440 -16943
rect -8500 -16999 -8440 -16995
rect -7216 -16972 -7127 -16883
rect -4997 -17018 -4941 -16962
rect -2288 -17018 -2232 -16962
rect -18085 -17197 -18005 -17118
rect -16342 -17988 -16282 -17984
rect -16342 -18040 -16338 -17988
rect -16338 -18040 -16286 -17988
rect -16286 -18040 -16282 -17988
rect -16342 -18044 -16282 -18040
rect -15052 -18045 -14963 -17956
rect -18088 -18143 -18014 -18069
rect -17040 -18167 -16980 -18163
rect -17040 -18219 -17036 -18167
rect -17036 -18219 -16984 -18167
rect -16984 -18219 -16980 -18167
rect -17040 -18223 -16980 -18219
rect -12471 -18161 -12399 -17039
rect 12233 -17027 12352 -16908
rect 12960 -17068 13079 -16949
rect 16285 -16995 16543 -16737
rect -8549 -17274 -8480 -17205
rect -8497 -17412 -8437 -17408
rect -8497 -17464 -8493 -17412
rect -8493 -17464 -8441 -17412
rect -8441 -17464 -8437 -17412
rect -8497 -17468 -8437 -17464
rect -7215 -17447 -7126 -17358
rect -5020 -17448 -4916 -17344
rect -4004 -17437 -3907 -17340
rect -2304 -17443 -2200 -17339
rect -1288 -17447 -1191 -17350
rect -11079 -17701 -11019 -17641
rect -8554 -17684 -8485 -17615
rect -8495 -17869 -8435 -17865
rect -8495 -17921 -8491 -17869
rect -8491 -17921 -8439 -17869
rect -8439 -17921 -8435 -17869
rect -8495 -17925 -8435 -17921
rect -7210 -17899 -7121 -17810
rect -4977 -17839 -4921 -17783
rect -2267 -17839 -2211 -17783
rect 8405 -17479 8461 -17444
rect 8405 -17500 8461 -17479
rect -8554 -18166 -8485 -18097
rect -18060 -18450 -18000 -18390
rect -8493 -18334 -8433 -18330
rect -8493 -18386 -8489 -18334
rect -8489 -18386 -8437 -18334
rect -8437 -18386 -8433 -18334
rect -8493 -18390 -8433 -18386
rect -7210 -18341 -7121 -18252
rect -5020 -18267 -4916 -18163
rect -4004 -18256 -3907 -18159
rect -2304 -18262 -2200 -18158
rect -1288 -18266 -1191 -18169
rect -18094 -18599 -18015 -18520
rect -16348 -18497 -16288 -18493
rect -16348 -18549 -16344 -18497
rect -16344 -18549 -16292 -18497
rect -16292 -18549 -16288 -18497
rect -16348 -18553 -16288 -18549
rect -15059 -18538 -14970 -18449
rect -12661 -18463 -12599 -18401
rect -12628 -18657 -12549 -18578
rect -8554 -18636 -8485 -18567
rect -5001 -18649 -4939 -18587
rect -2289 -18649 -2227 -18587
rect -16348 -18980 -16288 -18976
rect -16348 -19032 -16344 -18980
rect -16344 -19032 -16292 -18980
rect -16292 -19032 -16288 -18980
rect -16348 -19036 -16288 -19032
rect -15060 -19024 -14971 -18935
rect -18086 -19549 -18012 -19475
rect -16348 -19502 -16288 -19498
rect -16348 -19554 -16344 -19502
rect -16344 -19554 -16292 -19502
rect -16292 -19554 -16288 -19502
rect -16348 -19558 -16288 -19554
rect -15064 -19531 -14975 -19442
rect -21939 -19631 -21879 -19627
rect -21939 -19683 -21935 -19631
rect -21935 -19683 -21883 -19631
rect -21883 -19683 -21879 -19631
rect -21939 -19687 -21879 -19683
rect -20655 -19660 -20566 -19571
rect -18013 -19682 -17957 -19626
rect -16925 -19622 -16865 -19618
rect -16925 -19674 -16921 -19622
rect -16921 -19674 -16869 -19622
rect -16869 -19674 -16865 -19622
rect -16925 -19678 -16865 -19674
rect -8489 -18815 -8429 -18811
rect -8489 -18867 -8485 -18815
rect -8485 -18867 -8433 -18815
rect -8433 -18867 -8429 -18815
rect -8489 -18871 -8429 -18867
rect -7216 -18822 -7127 -18733
rect -5020 -19086 -4916 -18982
rect -4004 -19075 -3907 -18978
rect -2304 -19081 -2200 -18977
rect -1288 -19085 -1191 -18988
rect -8579 -19165 -8517 -19103
rect -5009 -19497 -4947 -19435
rect -2295 -19497 -2233 -19435
rect -23338 -19897 -23237 -19796
rect -24815 -20004 -24719 -19908
rect -17981 -19973 -17920 -19912
rect -16345 -19971 -16285 -19967
rect -16345 -20023 -16341 -19971
rect -16341 -20023 -16289 -19971
rect -16289 -20023 -16285 -19971
rect -16345 -20027 -16285 -20023
rect -15063 -20006 -14974 -19917
rect -21936 -20100 -21876 -20096
rect -21936 -20152 -21932 -20100
rect -21932 -20152 -21880 -20100
rect -21880 -20152 -21876 -20100
rect -21936 -20156 -21876 -20152
rect -20654 -20135 -20565 -20046
rect -24936 -20363 -24864 -20291
rect -24902 -20533 -24811 -20444
rect -21934 -20557 -21874 -20553
rect -21934 -20609 -21930 -20557
rect -21930 -20609 -21878 -20557
rect -21878 -20609 -21874 -20557
rect -21934 -20613 -21874 -20609
rect -20649 -20587 -20560 -20498
rect -24815 -21200 -24719 -21104
rect -23329 -21095 -23228 -20994
rect -21932 -21022 -21872 -21018
rect -21932 -21074 -21928 -21022
rect -21928 -21074 -21876 -21022
rect -21876 -21074 -21872 -21022
rect -21932 -21078 -21872 -21074
rect -20649 -21029 -20560 -20940
rect -24914 -21569 -24852 -21497
rect -21928 -21503 -21868 -21499
rect -21928 -21555 -21924 -21503
rect -21924 -21555 -21872 -21503
rect -21872 -21555 -21868 -21503
rect -21928 -21559 -21868 -21555
rect -20655 -21510 -20566 -21421
rect -24913 -21739 -24823 -21650
rect -16343 -20428 -16283 -20424
rect -16343 -20480 -16339 -20428
rect -16339 -20480 -16287 -20428
rect -16287 -20480 -16283 -20428
rect -16343 -20484 -16283 -20480
rect -15058 -20458 -14969 -20369
rect -18090 -20943 -18016 -20869
rect -16341 -20893 -16281 -20889
rect -16341 -20945 -16337 -20893
rect -16337 -20945 -16285 -20893
rect -16285 -20945 -16281 -20893
rect -16341 -20949 -16281 -20945
rect -15058 -20900 -14969 -20811
rect -16916 -21075 -16854 -21013
rect -12471 -21118 -12399 -19996
rect -5020 -19905 -4916 -19801
rect -4004 -19894 -3907 -19797
rect -2304 -19900 -2200 -19796
rect -1288 -19904 -1191 -19807
rect -5161 -20123 -5099 -20061
rect -2415 -20123 -2353 -20061
rect 10266 -17537 10322 -17481
rect 9001 -17632 9067 -17570
rect 9947 -17631 10003 -17570
rect 11894 -18187 12136 -17945
rect 17526 -18154 17659 -18021
rect 5563 -18615 5622 -18556
rect 6003 -18633 6062 -18574
rect 6440 -18626 6499 -18567
rect 15551 -18658 15695 -18514
rect 17977 -18940 18048 -18869
rect 5732 -19412 5788 -19410
rect 5732 -19464 5734 -19412
rect 5734 -19464 5786 -19412
rect 5786 -19464 5788 -19412
rect 5732 -19466 5788 -19464
rect 6170 -19393 6226 -19391
rect 6170 -19445 6172 -19393
rect 6172 -19445 6224 -19393
rect 6224 -19445 6226 -19393
rect 6170 -19447 6226 -19445
rect 6610 -19384 6666 -19382
rect 6610 -19436 6612 -19384
rect 6612 -19436 6664 -19384
rect 6664 -19436 6666 -19384
rect 6610 -19438 6666 -19436
rect 6304 -19823 6362 -19765
rect 12198 -19779 12420 -19771
rect 6438 -20069 6507 -20000
rect 8998 -19877 9054 -19875
rect 8998 -19929 9000 -19877
rect 9000 -19929 9052 -19877
rect 9052 -19929 9054 -19877
rect 8998 -19931 9054 -19929
rect 9935 -19877 9991 -19873
rect 9935 -19929 9987 -19877
rect 9987 -19929 9991 -19877
rect 8541 -20064 8600 -20005
rect 10267 -19988 10326 -19929
rect 12198 -19982 12410 -19779
rect 12410 -19982 12420 -19779
rect 12198 -19993 12420 -19982
rect -11079 -20658 -11019 -20598
rect -18051 -21235 -17995 -21179
rect -17964 -21400 -17908 -21344
rect -16337 -21374 -16277 -21370
rect -16337 -21426 -16333 -21374
rect -16333 -21426 -16281 -21374
rect -16281 -21426 -16277 -21374
rect -16337 -21430 -16277 -21426
rect -15064 -21381 -14975 -21292
rect -12604 -21432 -12544 -21372
rect -12623 -21611 -12544 -21532
rect -16726 -22047 -16662 -21983
rect -2305 -20528 -2199 -20422
rect -1288 -20537 -1191 -20440
rect 16231 -20436 16480 -20177
rect -5020 -20724 -4916 -20620
rect -4004 -20713 -3907 -20616
rect 7227 -21103 7405 -20925
rect 8162 -21103 8340 -20925
rect 9098 -21103 9276 -20925
rect 10029 -21102 10206 -20925
rect 10956 -21103 11134 -20925
rect 12233 -21555 12352 -21436
rect 12960 -21596 13079 -21477
rect -23332 -22389 -23231 -22288
rect -18088 -22347 -18014 -22273
rect -24805 -22508 -24709 -22412
rect -18061 -22666 -17995 -22600
rect -24890 -22870 -24818 -22798
rect -18067 -22829 -17987 -22750
rect -24913 -23040 -24819 -22951
rect -16688 -23445 -16610 -23367
rect -23372 -23705 -23271 -23604
rect -24825 -23814 -24729 -23718
rect -18090 -23749 -18016 -23675
rect -12471 -23697 -12399 -22575
rect -11079 -23237 -11019 -23177
rect -18037 -24053 -17975 -23991
rect -12673 -24011 -12617 -23955
rect -24926 -24180 -24864 -24108
rect -18058 -24215 -17979 -24136
rect -12681 -24158 -12619 -24097
rect -24907 -24350 -24813 -24261
rect -16688 -24849 -16614 -24775
rect -18084 -25129 -18010 -25055
rect -17951 -25417 -17889 -25355
rect -17971 -25637 -17892 -25558
rect -12471 -26465 -12399 -25343
rect -11079 -26005 -11019 -25945
rect -12741 -26803 -12685 -26747
rect -12744 -26994 -12688 -26938
rect -12471 -29098 -12399 -27976
rect -11079 -28638 -11019 -28578
rect -12719 -29441 -12657 -29379
rect -12723 -29621 -12643 -29542
rect -12471 -31707 -12399 -30585
rect -11079 -31247 -11019 -31187
rect -12753 -31985 -12691 -31923
rect -12787 -32171 -12707 -32092
rect -12473 -34327 -12401 -33205
rect -11081 -33867 -11021 -33807
rect -12577 -34571 -12515 -34509
rect -12721 -34755 -12642 -34676
rect 8405 -22007 8461 -21972
rect 8405 -22028 8461 -22007
rect 10266 -22065 10322 -22009
rect 9001 -22160 9067 -22098
rect 9947 -22159 10003 -22098
rect 11894 -22715 12136 -22473
rect 5563 -23159 5622 -23100
rect 6003 -23149 6062 -23090
rect 6448 -23124 6507 -23065
rect 5732 -23940 5788 -23938
rect 5732 -23992 5734 -23940
rect 5734 -23992 5786 -23940
rect 5786 -23992 5788 -23940
rect 5732 -23994 5788 -23992
rect 6170 -23921 6226 -23919
rect 6170 -23973 6172 -23921
rect 6172 -23973 6224 -23921
rect 6224 -23973 6226 -23921
rect 6170 -23975 6226 -23973
rect 6610 -23912 6666 -23910
rect 6610 -23964 6612 -23912
rect 6612 -23964 6664 -23912
rect 6664 -23964 6666 -23912
rect 6610 -23966 6666 -23964
rect 6304 -24351 6362 -24293
rect 12198 -24307 12420 -24299
rect 6438 -24597 6507 -24528
rect 8998 -24405 9054 -24403
rect 8998 -24457 9000 -24405
rect 9000 -24457 9052 -24405
rect 9052 -24457 9054 -24405
rect 8998 -24459 9054 -24457
rect 9935 -24405 9991 -24401
rect 9935 -24457 9987 -24405
rect 9987 -24457 9991 -24405
rect 8541 -24592 8600 -24533
rect 10267 -24516 10326 -24457
rect 12198 -24510 12410 -24307
rect 12410 -24510 12420 -24307
rect 12198 -24521 12420 -24510
rect 7227 -25631 7405 -25453
rect 8162 -25631 8340 -25453
rect 9098 -25631 9276 -25453
rect 10029 -25630 10206 -25453
rect 10956 -25631 11134 -25453
rect 12233 -26083 12352 -25964
rect 12960 -26124 13079 -26005
rect 8405 -26535 8461 -26500
rect 8405 -26556 8461 -26535
rect 10266 -26593 10322 -26537
rect 9001 -26688 9067 -26626
rect 9947 -26687 10003 -26626
rect 11894 -27243 12136 -27001
rect 5563 -27699 5622 -27640
rect 6003 -27694 6062 -27635
rect 6438 -27640 6497 -27581
rect 5732 -28468 5788 -28466
rect 5732 -28520 5734 -28468
rect 5734 -28520 5786 -28468
rect 5786 -28520 5788 -28468
rect 5732 -28522 5788 -28520
rect 6170 -28449 6226 -28447
rect 6170 -28501 6172 -28449
rect 6172 -28501 6224 -28449
rect 6224 -28501 6226 -28449
rect 6170 -28503 6226 -28501
rect 6610 -28440 6666 -28438
rect 6610 -28492 6612 -28440
rect 6612 -28492 6664 -28440
rect 6664 -28492 6666 -28440
rect 6610 -28494 6666 -28492
rect 6304 -28879 6362 -28821
rect 12198 -28835 12420 -28827
rect 6438 -29125 6507 -29056
rect 8998 -28933 9054 -28931
rect 8998 -28985 9000 -28933
rect 9000 -28985 9052 -28933
rect 9052 -28985 9054 -28933
rect 8998 -28987 9054 -28985
rect 9935 -28933 9991 -28929
rect 9935 -28985 9987 -28933
rect 9987 -28985 9991 -28933
rect 8541 -29120 8600 -29061
rect 10267 -29044 10326 -28985
rect 12198 -29038 12410 -28835
rect 12410 -29038 12420 -28835
rect 12198 -29049 12420 -29038
rect 7227 -30159 7405 -29981
rect 8162 -30159 8340 -29981
rect 9098 -30159 9276 -29981
rect 10029 -30158 10206 -29981
rect 10956 -30159 11134 -29981
rect 12233 -30611 12352 -30492
rect 12960 -30652 13079 -30533
rect 8405 -31063 8461 -31028
rect 8405 -31084 8461 -31063
rect 10266 -31121 10322 -31065
rect 9001 -31216 9067 -31154
rect 9947 -31215 10003 -31154
rect 11894 -31771 12136 -31529
rect 5563 -32208 5622 -32149
rect 6003 -32223 6062 -32164
rect 6438 -32201 6507 -32131
rect 5732 -32996 5788 -32994
rect 5732 -33048 5734 -32996
rect 5734 -33048 5786 -32996
rect 5786 -33048 5788 -32996
rect 5732 -33050 5788 -33048
rect 6170 -32977 6226 -32975
rect 6170 -33029 6172 -32977
rect 6172 -33029 6224 -32977
rect 6224 -33029 6226 -32977
rect 6170 -33031 6226 -33029
rect 6610 -32968 6666 -32966
rect 6610 -33020 6612 -32968
rect 6612 -33020 6664 -32968
rect 6664 -33020 6666 -32968
rect 6610 -33022 6666 -33020
rect 6304 -33407 6362 -33349
rect 12198 -33363 12420 -33355
rect 6438 -33653 6507 -33584
rect 8998 -33461 9054 -33459
rect 8998 -33513 9000 -33461
rect 9000 -33513 9052 -33461
rect 9052 -33513 9054 -33461
rect 8998 -33515 9054 -33513
rect 9935 -33461 9991 -33457
rect 9935 -33513 9987 -33461
rect 9987 -33513 9991 -33461
rect 8541 -33648 8600 -33589
rect 10267 -33572 10326 -33513
rect 12198 -33566 12410 -33363
rect 12410 -33566 12420 -33363
rect 12198 -33577 12420 -33566
rect 7227 -34687 7405 -34509
rect 8162 -34687 8340 -34509
rect 9098 -34687 9276 -34509
rect 10029 -34686 10206 -34509
rect 10956 -34687 11134 -34509
rect 12233 -35139 12352 -35020
rect 12960 -35180 13079 -35061
rect 8405 -35591 8461 -35556
rect 8405 -35612 8461 -35591
rect 10266 -35649 10322 -35593
rect 9001 -35744 9067 -35682
rect 9947 -35743 10003 -35682
rect 11894 -36299 12136 -36057
rect 12549 -36052 12646 -35955
rect 13558 -36063 13662 -35959
<< metal3 >>
rect -27376 7075 -22560 7080
rect -27376 7013 -22627 7075
rect -22565 7013 -22560 7075
rect -27376 7008 -22560 7013
rect -27525 4536 -27436 4541
rect -27525 4457 -27520 4536
rect -27441 4457 -27436 4536
rect -27525 -24260 -27436 4457
rect -27376 -24108 -27304 7008
rect -27210 6809 -21727 6814
rect -27210 6730 -21811 6809
rect -21732 6730 -21727 6809
rect -27210 6725 -21727 6730
rect -27210 6717 -27121 6725
rect -27210 -22950 -27131 6717
rect -27070 6650 -19240 6655
rect -27070 6588 -19307 6650
rect -19245 6588 -19240 6650
rect -27070 6583 -19240 6588
rect -27070 -22798 -26998 6583
rect -26921 6496 -18440 6501
rect -26921 6417 -18524 6496
rect -18445 6417 -18440 6496
rect -26921 6412 -18440 6417
rect -26921 6411 -26832 6412
rect -26921 -21642 -26842 6411
rect -26782 6304 -15947 6309
rect -26782 6242 -16014 6304
rect -15952 6242 -15947 6304
rect -26782 6237 -15947 6242
rect 1795 6241 3005 6269
rect -26782 -21497 -26710 6237
rect 1795 6169 1841 6241
rect 2963 6169 3005 6241
rect -26650 6150 -15142 6155
rect -26650 6071 -15226 6150
rect -15147 6071 -15142 6150
rect 1795 6143 3005 6169
rect 3401 6241 4611 6269
rect 3401 6169 3447 6241
rect 4569 6169 4611 6241
rect 3401 6143 4611 6169
rect 5105 6239 6315 6267
rect 5105 6167 5151 6239
rect 6273 6167 6315 6239
rect 5105 6141 6315 6167
rect -26650 6066 -15142 6071
rect -26650 -20443 -26564 6066
rect -26500 5973 -12670 5978
rect -26500 5911 -12737 5973
rect -12675 5911 -12670 5973
rect -26500 5906 -12670 5911
rect -26500 -20291 -26428 5906
rect -26332 5784 -11852 5789
rect -26332 5705 -11936 5784
rect -11857 5705 -11852 5784
rect -26332 5700 -11852 5705
rect -26332 -13063 -26243 5700
rect -26332 -13144 -26327 -13063
rect -26248 -13144 -26243 -13063
rect -26332 -19255 -26243 -13144
rect -26169 5608 -9367 5613
rect -26169 5546 -9434 5608
rect -9372 5546 -9367 5608
rect -26169 5541 -9367 5546
rect -26169 -11591 -26097 5541
rect -9298 5481 -8552 5486
rect -9298 5479 -8636 5481
rect -26169 -11653 -26164 -11591
rect -26102 -11653 -26097 -11591
rect -26169 -19103 -26097 -11653
rect -25983 5402 -8636 5479
rect -8557 5402 -8552 5481
rect -25983 5397 -8552 5402
rect -25983 -10160 -25894 5397
rect -8489 5336 -6096 5339
rect -25983 -10241 -25978 -10160
rect -25899 -10241 -25894 -10160
rect -25983 -18127 -25894 -10241
rect -25814 5334 -6096 5336
rect -25814 5274 -6161 5334
rect -6101 5274 -6096 5334
rect -25814 5269 -6096 5274
rect -25814 -8302 -25744 5269
rect -25814 -8362 -25809 -8302
rect -25749 -8362 -25744 -8302
rect -25814 -17984 -25744 -8362
rect -25660 5202 -5263 5207
rect -25660 5123 -5353 5202
rect -5268 5123 -5263 5202
rect -25660 5118 -5263 5123
rect -25660 -6751 -25571 5118
rect -25660 -6832 -25655 -6751
rect -25576 -6832 -25571 -6751
rect -25660 -16922 -25571 -6832
rect -25509 5023 -2803 5028
rect -25509 4961 -2870 5023
rect -2808 4961 -2803 5023
rect -25509 4956 -2803 4961
rect -25509 -5035 -25437 4956
rect -25509 -5097 -25504 -5035
rect -25442 -5097 -25437 -5035
rect -25509 -16770 -25437 -5097
rect -25370 4876 -1970 4881
rect -25370 4797 -2054 4876
rect -1975 4797 -1970 4876
rect -25370 4792 -1970 4797
rect 2276 4854 2402 4860
rect -25370 -10976 -25281 4792
rect 2276 4784 2296 4854
rect 2366 4784 2402 4854
rect 2276 4769 2402 4784
rect 3882 4854 4008 4860
rect 3882 4784 3902 4854
rect 3972 4784 4008 4854
rect 3882 4769 4008 4784
rect 5586 4852 5712 4858
rect 5586 4782 5606 4852
rect 5676 4782 5712 4852
rect 5586 4767 5712 4782
rect -25370 -11055 -25365 -10976
rect -25286 -11055 -25281 -10976
rect -25370 -15738 -25281 -11055
rect -25221 4721 497 4726
rect -25221 4659 430 4721
rect 492 4659 497 4721
rect -25221 4654 497 4659
rect -25221 -2529 -25150 4654
rect -24042 4517 -22832 4545
rect -24042 4445 -24000 4517
rect -22878 4445 -22832 4517
rect -24042 4419 -22832 4445
rect -20751 4517 -19541 4545
rect -20751 4445 -20709 4517
rect -19587 4445 -19541 4517
rect -20751 4419 -19541 4445
rect -17460 4517 -16250 4545
rect -17460 4445 -17418 4517
rect -16296 4445 -16250 4517
rect -17460 4419 -16250 4445
rect -14169 4517 -12959 4545
rect -14169 4445 -14127 4517
rect -13005 4445 -12959 4517
rect -14169 4419 -12959 4445
rect -10878 4517 -9668 4545
rect -10878 4445 -10836 4517
rect -9714 4445 -9668 4517
rect -10878 4419 -9668 4445
rect -7588 4517 -6378 4545
rect -7588 4445 -7546 4517
rect -6424 4445 -6378 4517
rect -7588 4419 -6378 4445
rect -4297 4517 -3087 4545
rect -4297 4445 -4255 4517
rect -3133 4445 -3087 4517
rect -4297 4419 -3087 4445
rect -1006 4517 204 4545
rect -1006 4445 -964 4517
rect 158 4445 204 4517
rect -1006 4419 204 4445
rect 5553 4099 5632 4104
rect 5553 4029 5558 4099
rect 5627 4029 5632 4099
rect 5553 4024 5632 4029
rect 5993 4099 6072 4104
rect 5993 4029 5998 4099
rect 6067 4029 6072 4099
rect 5993 4024 6072 4029
rect 6440 4081 6509 4086
rect -23439 3130 -23313 3136
rect -23439 3060 -23403 3130
rect -23333 3060 -23313 3130
rect -23439 3045 -23313 3060
rect -20148 3130 -20022 3136
rect -20148 3060 -20112 3130
rect -20042 3060 -20022 3130
rect -20148 3045 -20022 3060
rect -16857 3130 -16731 3136
rect -16857 3060 -16821 3130
rect -16751 3060 -16731 3130
rect -16857 3045 -16731 3060
rect -13566 3130 -13440 3136
rect -13566 3060 -13530 3130
rect -13460 3060 -13440 3130
rect -13566 3045 -13440 3060
rect -10275 3130 -10149 3136
rect -10275 3060 -10239 3130
rect -10169 3060 -10149 3130
rect -10275 3045 -10149 3060
rect -6985 3130 -6859 3136
rect -6985 3060 -6949 3130
rect -6879 3060 -6859 3130
rect -6985 3045 -6859 3060
rect -3694 3130 -3568 3136
rect -3694 3060 -3658 3130
rect -3588 3060 -3568 3130
rect -3694 3045 -3568 3060
rect -403 3130 -277 3136
rect -403 3060 -367 3130
rect -297 3060 -277 3130
rect -403 3045 -277 3060
rect -24716 2733 -23506 2761
rect -24716 2661 -24670 2733
rect -23548 2661 -23506 2733
rect -24716 2635 -23506 2661
rect -23157 2733 -21947 2761
rect -23157 2661 -23111 2733
rect -21989 2661 -21947 2733
rect -23157 2635 -21947 2661
rect -21425 2733 -20215 2761
rect -21425 2661 -21379 2733
rect -20257 2661 -20215 2733
rect -21425 2635 -20215 2661
rect -19866 2733 -18656 2761
rect -19866 2661 -19820 2733
rect -18698 2661 -18656 2733
rect -19866 2635 -18656 2661
rect -18134 2733 -16924 2761
rect -18134 2661 -18088 2733
rect -16966 2661 -16924 2733
rect -18134 2635 -16924 2661
rect -16575 2733 -15365 2761
rect -16575 2661 -16529 2733
rect -15407 2661 -15365 2733
rect -16575 2635 -15365 2661
rect -14843 2733 -13633 2761
rect -14843 2661 -14797 2733
rect -13675 2661 -13633 2733
rect -14843 2635 -13633 2661
rect -13284 2733 -12074 2761
rect -13284 2661 -13238 2733
rect -12116 2661 -12074 2733
rect -13284 2635 -12074 2661
rect -11552 2733 -10342 2761
rect -11552 2661 -11506 2733
rect -10384 2661 -10342 2733
rect -11552 2635 -10342 2661
rect -9993 2733 -8783 2761
rect -9993 2661 -9947 2733
rect -8825 2661 -8783 2733
rect -9993 2635 -8783 2661
rect -8262 2733 -7052 2761
rect -8262 2661 -8216 2733
rect -7094 2661 -7052 2733
rect -8262 2635 -7052 2661
rect -6703 2733 -5493 2761
rect -6703 2661 -6657 2733
rect -5535 2661 -5493 2733
rect -6703 2635 -5493 2661
rect -4971 2733 -3761 2761
rect -4971 2661 -4925 2733
rect -3803 2661 -3761 2733
rect -4971 2635 -3761 2661
rect -3412 2733 -2202 2761
rect -3412 2661 -3366 2733
rect -2244 2661 -2202 2733
rect -3412 2635 -2202 2661
rect -1680 2733 -470 2761
rect -1680 2661 -1634 2733
rect -512 2661 -470 2733
rect -1680 2635 -470 2661
rect -121 2733 1089 2761
rect -121 2661 -75 2733
rect 1047 2661 1089 2733
rect -121 2635 1089 2661
rect -24235 1346 -24109 1352
rect -24235 1276 -24215 1346
rect -24145 1276 -24109 1346
rect -24235 1261 -24109 1276
rect -22676 1346 -22550 1352
rect -22676 1276 -22656 1346
rect -22586 1276 -22550 1346
rect -22676 1261 -22550 1276
rect -20944 1346 -20818 1352
rect -20944 1276 -20924 1346
rect -20854 1276 -20818 1346
rect -20944 1261 -20818 1276
rect -19385 1346 -19259 1352
rect -19385 1276 -19365 1346
rect -19295 1276 -19259 1346
rect -19385 1261 -19259 1276
rect -17653 1346 -17527 1352
rect -17653 1276 -17633 1346
rect -17563 1276 -17527 1346
rect -17653 1261 -17527 1276
rect -16094 1346 -15968 1352
rect -16094 1276 -16074 1346
rect -16004 1276 -15968 1346
rect -16094 1261 -15968 1276
rect -14362 1346 -14236 1352
rect -14362 1276 -14342 1346
rect -14272 1276 -14236 1346
rect -14362 1261 -14236 1276
rect -12803 1346 -12677 1352
rect -12803 1276 -12783 1346
rect -12713 1276 -12677 1346
rect -12803 1261 -12677 1276
rect -11071 1346 -10945 1352
rect -11071 1276 -11051 1346
rect -10981 1276 -10945 1346
rect -11071 1261 -10945 1276
rect -9512 1346 -9386 1352
rect -9512 1276 -9492 1346
rect -9422 1276 -9386 1346
rect -9512 1261 -9386 1276
rect -7781 1346 -7655 1352
rect -7781 1276 -7761 1346
rect -7691 1276 -7655 1346
rect -7781 1261 -7655 1276
rect -6222 1346 -6096 1352
rect -6222 1276 -6202 1346
rect -6132 1276 -6096 1346
rect -6222 1261 -6096 1276
rect -4490 1346 -4364 1352
rect -4490 1276 -4470 1346
rect -4400 1276 -4364 1346
rect -4490 1261 -4364 1276
rect -2931 1346 -2805 1352
rect -2931 1276 -2911 1346
rect -2841 1276 -2805 1346
rect -2931 1261 -2805 1276
rect -1199 1346 -1073 1352
rect -1199 1276 -1179 1346
rect -1109 1276 -1073 1346
rect -1199 1261 -1073 1276
rect 360 1346 486 1352
rect 360 1276 380 1346
rect 450 1276 486 1346
rect 360 1261 486 1276
rect -24421 1001 -24147 1010
rect -24421 929 -24412 1001
rect -24156 929 -24147 1001
rect -24421 920 -24147 929
rect -23132 1001 -22858 1010
rect -23132 929 -23123 1001
rect -22867 929 -22858 1001
rect -23132 920 -22858 929
rect -22415 1001 -22141 1010
rect -22415 929 -22406 1001
rect -22150 929 -22141 1001
rect -22415 920 -22141 929
rect -21130 1001 -20856 1010
rect -21130 929 -21121 1001
rect -20865 929 -20856 1001
rect -21130 920 -20856 929
rect -19841 1001 -19567 1010
rect -19841 929 -19832 1001
rect -19576 929 -19567 1001
rect -19841 920 -19567 929
rect -19124 1001 -18850 1010
rect -19124 929 -19115 1001
rect -18859 929 -18850 1001
rect -19124 920 -18850 929
rect -17839 1001 -17565 1010
rect -17839 929 -17830 1001
rect -17574 929 -17565 1001
rect -17839 920 -17565 929
rect -16550 1001 -16276 1010
rect -16550 929 -16541 1001
rect -16285 929 -16276 1001
rect -16550 920 -16276 929
rect -15833 1001 -15559 1010
rect -15833 929 -15824 1001
rect -15568 929 -15559 1001
rect -15833 920 -15559 929
rect -14548 1001 -14274 1010
rect -14548 929 -14539 1001
rect -14283 929 -14274 1001
rect -14548 920 -14274 929
rect -13259 1001 -12985 1010
rect -13259 929 -13250 1001
rect -12994 929 -12985 1001
rect -13259 920 -12985 929
rect -12542 1001 -12268 1010
rect -12542 929 -12533 1001
rect -12277 929 -12268 1001
rect -12542 920 -12268 929
rect -11257 1001 -10983 1010
rect -11257 929 -11248 1001
rect -10992 929 -10983 1001
rect -11257 920 -10983 929
rect -9968 1001 -9694 1010
rect -9968 929 -9959 1001
rect -9703 929 -9694 1001
rect -9968 920 -9694 929
rect -9251 1001 -8977 1010
rect -9251 929 -9242 1001
rect -8986 929 -8977 1001
rect -9251 920 -8977 929
rect -7967 1001 -7693 1010
rect -7967 929 -7958 1001
rect -7702 929 -7693 1001
rect -7967 920 -7693 929
rect -6678 1001 -6404 1010
rect -6678 929 -6669 1001
rect -6413 929 -6404 1001
rect -6678 920 -6404 929
rect -5961 1001 -5687 1010
rect -5961 929 -5952 1001
rect -5696 929 -5687 1001
rect -5961 920 -5687 929
rect -4676 1001 -4402 1010
rect -4676 929 -4667 1001
rect -4411 929 -4402 1001
rect -4676 920 -4402 929
rect -3387 1001 -3113 1010
rect -3387 929 -3378 1001
rect -3122 929 -3113 1001
rect -3387 920 -3113 929
rect -2670 1001 -2396 1010
rect -2670 929 -2661 1001
rect -2405 929 -2396 1001
rect -2670 920 -2396 929
rect -1385 1001 -1111 1010
rect -1385 929 -1376 1001
rect -1120 929 -1111 1001
rect -1385 920 -1111 929
rect -96 1001 178 1010
rect -96 929 -87 1001
rect 169 929 178 1001
rect -96 920 178 929
rect 621 1001 895 1010
rect 621 929 630 1001
rect 886 929 895 1001
rect 621 920 895 929
rect -24063 666 -23941 699
rect -24063 518 -24046 666
rect -23963 518 -23941 666
rect -24063 465 -23941 518
rect -20772 666 -20650 699
rect -20772 518 -20755 666
rect -20672 518 -20650 666
rect -20772 465 -20650 518
rect -17481 666 -17359 699
rect -17481 518 -17464 666
rect -17381 518 -17359 666
rect -17481 465 -17359 518
rect -14190 666 -14068 699
rect -14190 518 -14173 666
rect -14090 518 -14068 666
rect -14190 465 -14068 518
rect -10899 666 -10777 699
rect -10899 518 -10882 666
rect -10799 518 -10777 666
rect -10899 465 -10777 518
rect -7609 666 -7487 699
rect -7609 518 -7592 666
rect -7509 518 -7487 666
rect -7609 465 -7487 518
rect -4318 666 -4196 699
rect -4318 518 -4301 666
rect -4218 518 -4196 666
rect -4318 465 -4196 518
rect -1027 666 -905 699
rect -1027 518 -1010 666
rect -927 518 -905 666
rect -1027 465 -905 518
rect -24063 450 -22462 465
rect -24063 375 -22628 450
rect -22483 375 -22462 450
rect -24063 363 -22462 375
rect -20772 450 -19171 465
rect -20772 375 -19337 450
rect -19192 375 -19171 450
rect -20772 363 -19171 375
rect -17481 450 -15880 465
rect -17481 375 -16046 450
rect -15901 375 -15880 450
rect -17481 363 -15880 375
rect -14190 450 -12589 465
rect -14190 375 -12755 450
rect -12610 375 -12589 450
rect -14190 363 -12589 375
rect -10899 450 -9298 465
rect -10899 375 -9464 450
rect -9319 375 -9298 450
rect -10899 363 -9298 375
rect -7609 450 -6008 465
rect -7609 375 -6174 450
rect -6029 375 -6008 450
rect -7609 363 -6008 375
rect -4318 450 -2717 465
rect -4318 375 -2883 450
rect -2738 375 -2717 450
rect -4318 363 -2717 375
rect -1027 450 574 465
rect -1027 375 408 450
rect 553 375 574 450
rect -1027 363 574 375
rect -24345 267 -23992 268
rect -24345 203 -24336 267
rect -24001 203 -23992 267
rect -24345 194 -23992 203
rect -23125 255 -23013 269
rect -23125 183 -23105 255
rect -23033 183 -23013 255
rect -21054 267 -20701 268
rect -23125 172 -23013 183
rect -22258 230 -22155 244
rect -22258 164 -22240 230
rect -22174 164 -22155 230
rect -21054 203 -21045 267
rect -20710 203 -20701 267
rect -21054 194 -20701 203
rect -19834 255 -19722 269
rect -19834 183 -19814 255
rect -19742 183 -19722 255
rect -17763 267 -17410 268
rect -19834 172 -19722 183
rect -18967 230 -18864 244
rect -22258 146 -22155 164
rect -18967 164 -18949 230
rect -18883 164 -18864 230
rect -17763 203 -17754 267
rect -17419 203 -17410 267
rect -17763 194 -17410 203
rect -16543 255 -16431 269
rect -16543 183 -16523 255
rect -16451 183 -16431 255
rect -14472 267 -14119 268
rect -16543 172 -16431 183
rect -15676 230 -15573 244
rect -18967 146 -18864 164
rect -15676 164 -15658 230
rect -15592 164 -15573 230
rect -14472 203 -14463 267
rect -14128 203 -14119 267
rect -14472 194 -14119 203
rect -13252 255 -13140 269
rect -13252 183 -13232 255
rect -13160 183 -13140 255
rect -11181 267 -10828 268
rect -13252 172 -13140 183
rect -12385 230 -12282 244
rect -15676 146 -15573 164
rect -12385 164 -12367 230
rect -12301 164 -12282 230
rect -11181 203 -11172 267
rect -10837 203 -10828 267
rect -11181 194 -10828 203
rect -9961 255 -9849 269
rect -9961 183 -9941 255
rect -9869 183 -9849 255
rect -7891 267 -7538 268
rect -9961 172 -9849 183
rect -9094 230 -8991 244
rect -12385 146 -12282 164
rect -9094 164 -9076 230
rect -9010 164 -8991 230
rect -7891 203 -7882 267
rect -7547 203 -7538 267
rect -7891 194 -7538 203
rect -6671 255 -6559 269
rect -6671 183 -6651 255
rect -6579 183 -6559 255
rect -4600 267 -4247 268
rect -6671 172 -6559 183
rect -5804 230 -5701 244
rect -9094 146 -8991 164
rect -5804 164 -5786 230
rect -5720 164 -5701 230
rect -4600 203 -4591 267
rect -4256 203 -4247 267
rect -4600 194 -4247 203
rect -3380 255 -3268 269
rect -3380 183 -3360 255
rect -3288 183 -3268 255
rect -1309 267 -956 268
rect -3380 172 -3268 183
rect -2513 230 -2410 244
rect -5804 146 -5701 164
rect -2513 164 -2495 230
rect -2429 164 -2410 230
rect -1309 203 -1300 267
rect -965 203 -956 267
rect -1309 194 -956 203
rect -89 255 23 269
rect -89 183 -69 255
rect 3 183 23 255
rect -89 172 23 183
rect 778 230 881 244
rect -2513 146 -2410 164
rect 778 164 796 230
rect 862 164 881 230
rect 778 146 881 164
rect 5558 -450 5627 4024
rect 5707 3235 5827 3259
rect 5707 3169 5727 3235
rect 5793 3169 5827 3235
rect 5707 3146 5827 3169
rect 5558 -509 5563 -450
rect 5622 -509 5627 -450
rect -25221 -2591 -25216 -2529
rect -25155 -2591 -25150 -2529
rect -25221 -15586 -25150 -2591
rect -24861 -1976 -24679 -1972
rect -24861 -2141 -19075 -1976
rect -24861 -3997 -24679 -2141
rect -23628 -2225 -23414 -2203
rect -24448 -2327 -23814 -2293
rect -23628 -2304 -23605 -2225
rect -23436 -2304 -23414 -2225
rect -21608 -2225 -21394 -2203
rect -23628 -2323 -23414 -2304
rect -24448 -2467 -24410 -2327
rect -23856 -2467 -23814 -2327
rect -24448 -2506 -23814 -2467
rect -22411 -2327 -21777 -2293
rect -21608 -2304 -21585 -2225
rect -21416 -2304 -21394 -2225
rect -19867 -2225 -19653 -2203
rect -21608 -2323 -21394 -2304
rect -22411 -2467 -22373 -2327
rect -21819 -2467 -21777 -2327
rect -22411 -2506 -21777 -2467
rect -20681 -2327 -20047 -2293
rect -19867 -2304 -19844 -2225
rect -19675 -2304 -19653 -2225
rect -19867 -2323 -19653 -2304
rect -20681 -2467 -20643 -2327
rect -20089 -2467 -20047 -2327
rect -20681 -2506 -20047 -2467
rect -24588 -2940 -24398 -2859
rect -23628 -2878 -23428 -2850
rect -24603 -2987 -24394 -2940
rect -24603 -3165 -24550 -2987
rect -24428 -3165 -24394 -2987
rect -24213 -2983 -23813 -2955
rect -24213 -3057 -24184 -2983
rect -23844 -3057 -23813 -2983
rect -23628 -2974 -23601 -2878
rect -23452 -2974 -23428 -2878
rect -23628 -3000 -23428 -2974
rect -22627 -2852 -22400 -2819
rect -24213 -3078 -23813 -3057
rect -24603 -3194 -24394 -3165
rect -22627 -3080 -22594 -2852
rect -22431 -3080 -22400 -2852
rect -21608 -2878 -21408 -2850
rect -22176 -2983 -21776 -2955
rect -22176 -3057 -22147 -2983
rect -21807 -3057 -21776 -2983
rect -21608 -2974 -21581 -2878
rect -21432 -2974 -21408 -2878
rect -19867 -2878 -19667 -2850
rect -21608 -3000 -21408 -2974
rect -20446 -2983 -20046 -2955
rect -22176 -3078 -21776 -3057
rect -20944 -3042 -20726 -3021
rect -22627 -3113 -22400 -3080
rect -24586 -3395 -24402 -3194
rect -24586 -3399 -22754 -3395
rect -24586 -3595 -22752 -3399
rect -24861 -4064 -24578 -3997
rect -24861 -4337 -24807 -4064
rect -24618 -4337 -24578 -4064
rect -23584 -4037 -23370 -4015
rect -24397 -4139 -23763 -4105
rect -23584 -4116 -23561 -4037
rect -23392 -4116 -23370 -4037
rect -23584 -4135 -23370 -4116
rect -24397 -4279 -24359 -4139
rect -23805 -4279 -23763 -4139
rect -24397 -4318 -23763 -4279
rect -24861 -4379 -24578 -4337
rect -23210 -4480 -23051 -4435
rect -23210 -4594 -23195 -4480
rect -23064 -4594 -23051 -4480
rect -23584 -4690 -23384 -4662
rect -24162 -4795 -23762 -4767
rect -24162 -4869 -24133 -4795
rect -23793 -4869 -23762 -4795
rect -23584 -4786 -23557 -4690
rect -23408 -4786 -23384 -4690
rect -23584 -4812 -23384 -4786
rect -24162 -4890 -23762 -4869
rect -23586 -5329 -23372 -5307
rect -24397 -5431 -23763 -5397
rect -23586 -5408 -23563 -5329
rect -23394 -5408 -23372 -5329
rect -23586 -5427 -23372 -5408
rect -24397 -5571 -24359 -5431
rect -23805 -5571 -23763 -5431
rect -24397 -5610 -23763 -5571
rect -24651 -6020 -24460 -5899
rect -23586 -5982 -23386 -5954
rect -24651 -6049 -24439 -6020
rect -24651 -6247 -24612 -6049
rect -24466 -6247 -24439 -6049
rect -24162 -6087 -23762 -6059
rect -24162 -6161 -24133 -6087
rect -23793 -6161 -23762 -6087
rect -23586 -6078 -23559 -5982
rect -23410 -6078 -23386 -5982
rect -23586 -6104 -23386 -6078
rect -24162 -6182 -23762 -6161
rect -24651 -6262 -24439 -6247
rect -24651 -6684 -24460 -6262
rect -24651 -6824 -24619 -6684
rect -24490 -6824 -24460 -6684
rect -24651 -9285 -24460 -6824
rect -23585 -7302 -23371 -7280
rect -24397 -7404 -23763 -7370
rect -23585 -7381 -23562 -7302
rect -23393 -7381 -23371 -7302
rect -23585 -7400 -23371 -7381
rect -24397 -7544 -24359 -7404
rect -23805 -7544 -23763 -7404
rect -24397 -7583 -23763 -7544
rect -23210 -7743 -23051 -4594
rect -23210 -7857 -23198 -7743
rect -23067 -7745 -23051 -7743
rect -23210 -7859 -23195 -7857
rect -23064 -7859 -23051 -7745
rect -23585 -7955 -23385 -7927
rect -24162 -8060 -23762 -8032
rect -24162 -8134 -24133 -8060
rect -23793 -8134 -23762 -8060
rect -23585 -8051 -23558 -7955
rect -23409 -8051 -23385 -7955
rect -23585 -8077 -23385 -8051
rect -24162 -8155 -23762 -8134
rect -23583 -8594 -23369 -8572
rect -24397 -8696 -23763 -8662
rect -23583 -8673 -23560 -8594
rect -23391 -8673 -23369 -8594
rect -23583 -8692 -23369 -8673
rect -24397 -8836 -24359 -8696
rect -23805 -8836 -23763 -8696
rect -24397 -8875 -23763 -8836
rect -23583 -9247 -23383 -9219
rect -24651 -9314 -24439 -9285
rect -24651 -9512 -24612 -9314
rect -24466 -9512 -24439 -9314
rect -24162 -9352 -23762 -9324
rect -24162 -9426 -24133 -9352
rect -23793 -9426 -23762 -9352
rect -23583 -9343 -23556 -9247
rect -23407 -9343 -23383 -9247
rect -23583 -9369 -23383 -9343
rect -24162 -9447 -23762 -9426
rect -24651 -9527 -24439 -9512
rect -24651 -12549 -24460 -9527
rect -23583 -10566 -23369 -10544
rect -24397 -10668 -23763 -10634
rect -23583 -10645 -23560 -10566
rect -23391 -10645 -23369 -10566
rect -23583 -10664 -23369 -10645
rect -24397 -10808 -24359 -10668
rect -23805 -10808 -23763 -10668
rect -24397 -10847 -23763 -10808
rect -23210 -11007 -23051 -7859
rect -23210 -11121 -23198 -11007
rect -23061 -11121 -23051 -11007
rect -23210 -11123 -23195 -11121
rect -23064 -11123 -23051 -11121
rect -23210 -11132 -23051 -11123
rect -22937 -5995 -22752 -3595
rect -22627 -3742 -22459 -3113
rect -20944 -3165 -20917 -3042
rect -20741 -3165 -20726 -3042
rect -20446 -3057 -20417 -2983
rect -20077 -3057 -20046 -2983
rect -19867 -2974 -19840 -2878
rect -19691 -2974 -19667 -2878
rect -19867 -3000 -19667 -2974
rect -19292 -2908 -19075 -2141
rect -18088 -2225 -17874 -2203
rect -18921 -2327 -18287 -2293
rect -18088 -2304 -18065 -2225
rect -17896 -2304 -17874 -2225
rect -18088 -2323 -17874 -2304
rect -18921 -2467 -18883 -2327
rect -18329 -2467 -18287 -2327
rect -18921 -2506 -18287 -2467
rect -18088 -2878 -17888 -2850
rect -19292 -2934 -19012 -2908
rect -20446 -3078 -20046 -3057
rect -19292 -3087 -19241 -2934
rect -19043 -3087 -19012 -2934
rect -18686 -2983 -18286 -2955
rect -18686 -3057 -18657 -2983
rect -18317 -3057 -18286 -2983
rect -18088 -2974 -18061 -2878
rect -17912 -2974 -17888 -2878
rect -18088 -3000 -17888 -2974
rect -18686 -3078 -18286 -3057
rect -19292 -3115 -19012 -3087
rect -20944 -3179 -20726 -3165
rect -21524 -3186 -20726 -3179
rect -21524 -3198 -20773 -3186
rect -22627 -3848 -22600 -3742
rect -22476 -3848 -22459 -3742
rect -22627 -3869 -22459 -3848
rect -21525 -3363 -20773 -3198
rect -21525 -3373 -20779 -3363
rect -21846 -4037 -21632 -4015
rect -22661 -4139 -22027 -4105
rect -21846 -4116 -21823 -4037
rect -21654 -4116 -21632 -4037
rect -21846 -4135 -21632 -4116
rect -22661 -4279 -22623 -4139
rect -22069 -4279 -22027 -4139
rect -22661 -4318 -22027 -4279
rect -21846 -4690 -21646 -4662
rect -22426 -4795 -22026 -4767
rect -22426 -4869 -22397 -4795
rect -22057 -4869 -22026 -4795
rect -21846 -4786 -21819 -4690
rect -21670 -4786 -21646 -4690
rect -21846 -4812 -21646 -4786
rect -22426 -4890 -22026 -4869
rect -21852 -5329 -21638 -5307
rect -22661 -5431 -22027 -5397
rect -21852 -5408 -21829 -5329
rect -21660 -5408 -21638 -5329
rect -21852 -5427 -21638 -5408
rect -22661 -5571 -22623 -5431
rect -22069 -5571 -22027 -5431
rect -22661 -5610 -22027 -5571
rect -22937 -6441 -22862 -5995
rect -22773 -6441 -22752 -5995
rect -21852 -5982 -21652 -5954
rect -22426 -6087 -22026 -6059
rect -22426 -6161 -22397 -6087
rect -22057 -6161 -22026 -6087
rect -21852 -6078 -21825 -5982
rect -21676 -6078 -21652 -5982
rect -21852 -6104 -21652 -6078
rect -22426 -6182 -22026 -6161
rect -22937 -9239 -22752 -6441
rect -21525 -6678 -21345 -3373
rect -20649 -3827 -19439 -3799
rect -20649 -3899 -20603 -3827
rect -19481 -3899 -19439 -3827
rect -20649 -3925 -19439 -3899
rect -19090 -3827 -17880 -3799
rect -19090 -3899 -19044 -3827
rect -17922 -3899 -17880 -3827
rect -19090 -3925 -17880 -3899
rect -17358 -3827 -16148 -3799
rect -17358 -3899 -17312 -3827
rect -16190 -3899 -16148 -3827
rect -17358 -3925 -16148 -3899
rect -15799 -3827 -14589 -3799
rect -15799 -3899 -15753 -3827
rect -14631 -3899 -14589 -3827
rect -15799 -3925 -14589 -3899
rect -14067 -3827 -12857 -3799
rect -14067 -3899 -14021 -3827
rect -12899 -3899 -12857 -3827
rect -14067 -3925 -12857 -3899
rect -12508 -3827 -11298 -3799
rect -12508 -3899 -12462 -3827
rect -11340 -3899 -11298 -3827
rect -12508 -3925 -11298 -3899
rect -10776 -3827 -9566 -3799
rect -10776 -3899 -10730 -3827
rect -9608 -3899 -9566 -3827
rect -10776 -3925 -9566 -3899
rect -9217 -3827 -8007 -3799
rect -9217 -3899 -9171 -3827
rect -8049 -3899 -8007 -3827
rect -9217 -3925 -8007 -3899
rect 5558 -4860 5627 -509
rect 5998 -424 6067 4024
rect 6440 4022 6445 4081
rect 6504 4022 6509 4081
rect 6144 3254 6264 3280
rect 6144 3188 6165 3254
rect 6231 3188 6264 3254
rect 6144 3167 6264 3188
rect 6440 3020 6509 4022
rect 6579 3263 6699 3281
rect 6579 3197 6605 3263
rect 6671 3197 6699 3263
rect 6579 3168 6699 3197
rect 6144 2951 6509 3020
rect 6144 302 6213 2951
rect 6299 2875 6367 2880
rect 6299 2817 6304 2875
rect 6362 2817 6367 2875
rect 6299 2774 6367 2817
rect 12187 2874 12431 2880
rect 6299 2767 10002 2774
rect 6299 2765 9935 2767
rect 6299 2709 8998 2765
rect 9054 2711 9935 2765
rect 9991 2711 10002 2767
rect 9054 2709 10002 2711
rect 6299 2706 10002 2709
rect 6299 547 6365 2706
rect 6573 2704 10002 2706
rect 10262 2711 10331 2716
rect 10262 2652 10267 2711
rect 10326 2652 10331 2711
rect 6433 2640 6512 2645
rect 10262 2640 10331 2652
rect 6433 2571 6438 2640
rect 6507 2635 10331 2640
rect 12187 2642 12193 2874
rect 12425 2642 12431 2874
rect 12187 2636 12431 2642
rect 6507 2576 8541 2635
rect 8600 2576 10331 2635
rect 6507 2571 10331 2576
rect 6433 2566 6512 2571
rect 6433 2493 6507 2566
rect 6440 667 6500 2493
rect 7156 1720 11207 1787
rect 7156 1532 7222 1720
rect 7410 1532 8157 1720
rect 8345 1532 9093 1720
rect 9281 1533 10024 1720
rect 10211 1533 10951 1720
rect 9281 1532 10951 1533
rect 11139 1532 11207 1720
rect 7156 1466 11207 1532
rect 12414 1296 12821 1408
rect 12128 1292 12821 1296
rect 12128 1266 13042 1292
rect 12128 1209 13186 1266
rect 12128 1080 12228 1209
rect 12357 1168 13186 1209
rect 12357 1080 12955 1168
rect 12128 1039 12955 1080
rect 13084 1039 13186 1168
rect 12128 979 13186 1039
rect 12467 820 13186 979
rect 12796 787 13186 820
rect 8398 668 8471 673
rect 8398 667 8405 668
rect 6440 612 8405 667
rect 8461 667 8471 668
rect 8461 636 10324 667
rect 8461 631 10327 636
rect 8461 612 10266 631
rect 6440 607 10266 612
rect 10261 575 10266 607
rect 10322 575 10327 631
rect 10261 570 10327 575
rect 6299 542 10021 547
rect 6299 481 9001 542
rect 8996 480 9001 481
rect 9067 481 9947 542
rect 10003 481 10021 542
rect 9067 480 9072 481
rect 8996 475 9072 480
rect 9942 476 10021 481
rect 6144 233 6507 302
rect 5998 -483 6003 -424
rect 6062 -483 6067 -424
rect 5707 -1293 5827 -1269
rect 5707 -1359 5727 -1293
rect 5793 -1359 5827 -1293
rect 5707 -1382 5827 -1359
rect 5558 -4919 5563 -4860
rect 5622 -4919 5627 -4860
rect -20168 -5214 -20042 -5208
rect -20168 -5284 -20148 -5214
rect -20078 -5284 -20042 -5214
rect -20168 -5299 -20042 -5284
rect -18609 -5214 -18483 -5208
rect -18609 -5284 -18589 -5214
rect -18519 -5284 -18483 -5214
rect -18609 -5299 -18483 -5284
rect -16877 -5214 -16751 -5208
rect -16877 -5284 -16857 -5214
rect -16787 -5284 -16751 -5214
rect -16877 -5299 -16751 -5284
rect -15318 -5214 -15192 -5208
rect -15318 -5284 -15298 -5214
rect -15228 -5284 -15192 -5214
rect -15318 -5299 -15192 -5284
rect -13586 -5214 -13460 -5208
rect -13586 -5284 -13566 -5214
rect -13496 -5284 -13460 -5214
rect -13586 -5299 -13460 -5284
rect -12027 -5214 -11901 -5208
rect -12027 -5284 -12007 -5214
rect -11937 -5284 -11901 -5214
rect -12027 -5299 -11901 -5284
rect -10295 -5214 -10169 -5208
rect -10295 -5284 -10275 -5214
rect -10205 -5284 -10169 -5214
rect -10295 -5299 -10169 -5284
rect -8736 -5214 -8610 -5208
rect -8736 -5284 -8716 -5214
rect -8646 -5284 -8610 -5214
rect -8736 -5299 -8610 -5284
rect -20354 -5559 -20080 -5550
rect -20354 -5631 -20345 -5559
rect -20089 -5631 -20080 -5559
rect -20354 -5640 -20080 -5631
rect -19065 -5559 -18791 -5550
rect -19065 -5631 -19056 -5559
rect -18800 -5631 -18791 -5559
rect -19065 -5640 -18791 -5631
rect -18348 -5559 -18074 -5550
rect -18348 -5631 -18339 -5559
rect -18083 -5631 -18074 -5559
rect -18348 -5640 -18074 -5631
rect -17063 -5559 -16789 -5550
rect -17063 -5631 -17054 -5559
rect -16798 -5631 -16789 -5559
rect -17063 -5640 -16789 -5631
rect -15774 -5559 -15500 -5550
rect -15774 -5631 -15765 -5559
rect -15509 -5631 -15500 -5559
rect -15774 -5640 -15500 -5631
rect -15057 -5559 -14783 -5550
rect -15057 -5631 -15048 -5559
rect -14792 -5631 -14783 -5559
rect -15057 -5640 -14783 -5631
rect -13772 -5559 -13498 -5550
rect -13772 -5631 -13763 -5559
rect -13507 -5631 -13498 -5559
rect -13772 -5640 -13498 -5631
rect -12483 -5559 -12209 -5550
rect -12483 -5631 -12474 -5559
rect -12218 -5631 -12209 -5559
rect -12483 -5640 -12209 -5631
rect -11766 -5559 -11492 -5550
rect -11766 -5631 -11757 -5559
rect -11501 -5631 -11492 -5559
rect -11766 -5640 -11492 -5631
rect -10481 -5559 -10207 -5550
rect -10481 -5631 -10472 -5559
rect -10216 -5631 -10207 -5559
rect -10481 -5640 -10207 -5631
rect -9192 -5559 -8918 -5550
rect -9192 -5631 -9183 -5559
rect -8927 -5631 -8918 -5559
rect -9192 -5640 -8918 -5631
rect -8475 -5559 -8201 -5550
rect -8475 -5631 -8466 -5559
rect -8210 -5631 -8201 -5559
rect -8475 -5640 -8201 -5631
rect -19996 -5894 -19874 -5861
rect -19996 -6042 -19979 -5894
rect -19896 -6042 -19874 -5894
rect -19996 -6095 -19874 -6042
rect -16705 -5894 -16583 -5861
rect -16705 -6042 -16688 -5894
rect -16605 -6042 -16583 -5894
rect -16705 -6095 -16583 -6042
rect -13414 -5894 -13292 -5861
rect -13414 -6042 -13397 -5894
rect -13314 -6042 -13292 -5894
rect -13414 -6095 -13292 -6042
rect -10123 -5894 -10001 -5861
rect -10123 -6042 -10106 -5894
rect -10023 -6042 -10001 -5894
rect -10123 -6095 -10001 -6042
rect -19996 -6110 -18395 -6095
rect -19996 -6185 -18561 -6110
rect -18416 -6185 -18395 -6110
rect -19996 -6197 -18395 -6185
rect -16705 -6110 -15104 -6095
rect -16705 -6185 -15270 -6110
rect -15125 -6185 -15104 -6110
rect -16705 -6197 -15104 -6185
rect -13414 -6110 -11813 -6095
rect -13414 -6185 -11979 -6110
rect -11834 -6185 -11813 -6110
rect -13414 -6197 -11813 -6185
rect -10123 -6110 -8522 -6095
rect -10123 -6185 -8688 -6110
rect -8543 -6185 -8522 -6110
rect -10123 -6197 -8522 -6185
rect -20278 -6293 -19925 -6292
rect -20278 -6357 -20269 -6293
rect -19934 -6357 -19925 -6293
rect -20278 -6366 -19925 -6357
rect -19058 -6305 -18946 -6291
rect -19058 -6377 -19038 -6305
rect -18966 -6377 -18946 -6305
rect -16987 -6293 -16634 -6292
rect -19058 -6388 -18946 -6377
rect -18191 -6330 -18088 -6316
rect -18191 -6396 -18173 -6330
rect -18107 -6396 -18088 -6330
rect -16987 -6357 -16978 -6293
rect -16643 -6357 -16634 -6293
rect -16987 -6366 -16634 -6357
rect -15767 -6305 -15655 -6291
rect -15767 -6377 -15747 -6305
rect -15675 -6377 -15655 -6305
rect -13696 -6293 -13343 -6292
rect -15767 -6388 -15655 -6377
rect -14900 -6330 -14797 -6316
rect -18191 -6414 -18088 -6396
rect -14900 -6396 -14882 -6330
rect -14816 -6396 -14797 -6330
rect -13696 -6357 -13687 -6293
rect -13352 -6357 -13343 -6293
rect -13696 -6366 -13343 -6357
rect -12476 -6305 -12364 -6291
rect -12476 -6377 -12456 -6305
rect -12384 -6377 -12364 -6305
rect -10405 -6293 -10052 -6292
rect -12476 -6388 -12364 -6377
rect -11609 -6330 -11506 -6316
rect -14900 -6414 -14797 -6396
rect -11609 -6396 -11591 -6330
rect -11525 -6396 -11506 -6330
rect -10405 -6357 -10396 -6293
rect -10061 -6357 -10052 -6293
rect -10405 -6366 -10052 -6357
rect -9185 -6305 -9073 -6291
rect -9185 -6377 -9165 -6305
rect -9093 -6377 -9073 -6305
rect -9185 -6388 -9073 -6377
rect -8318 -6330 -8215 -6316
rect -11609 -6414 -11506 -6396
rect -8318 -6396 -8300 -6330
rect -8234 -6396 -8215 -6330
rect -8318 -6414 -8215 -6396
rect -21525 -6818 -21515 -6678
rect -21386 -6818 -21345 -6678
rect -21525 -6854 -21345 -6818
rect -20649 -7092 -19439 -7064
rect -20649 -7164 -20603 -7092
rect -19481 -7164 -19439 -7092
rect -20649 -7190 -19439 -7164
rect -19090 -7092 -17880 -7064
rect -19090 -7164 -19044 -7092
rect -17922 -7164 -17880 -7092
rect -19090 -7190 -17880 -7164
rect -17358 -7092 -16148 -7064
rect -17358 -7164 -17312 -7092
rect -16190 -7164 -16148 -7092
rect -17358 -7190 -16148 -7164
rect -15799 -7092 -14589 -7064
rect -15799 -7164 -15753 -7092
rect -14631 -7164 -14589 -7092
rect -15799 -7190 -14589 -7164
rect -14067 -7092 -12857 -7064
rect -14067 -7164 -14021 -7092
rect -12899 -7164 -12857 -7092
rect -14067 -7190 -12857 -7164
rect -12508 -7092 -11298 -7064
rect -12508 -7164 -12462 -7092
rect -11340 -7164 -11298 -7092
rect -12508 -7190 -11298 -7164
rect -10776 -7092 -9566 -7064
rect -10776 -7164 -10730 -7092
rect -9608 -7164 -9566 -7092
rect -10776 -7190 -9566 -7164
rect -9217 -7092 -8007 -7064
rect -9217 -7164 -9171 -7092
rect -8049 -7164 -8007 -7092
rect -9217 -7190 -8007 -7164
rect -21850 -7302 -21636 -7280
rect -22660 -7404 -22026 -7370
rect -21850 -7381 -21827 -7302
rect -21658 -7381 -21636 -7302
rect -21850 -7400 -21636 -7381
rect -22660 -7544 -22622 -7404
rect -22068 -7544 -22026 -7404
rect -22660 -7583 -22026 -7544
rect -21850 -7955 -21650 -7927
rect -22425 -8060 -22025 -8032
rect -22425 -8134 -22396 -8060
rect -22056 -8134 -22025 -8060
rect -21850 -8051 -21823 -7955
rect -21674 -8051 -21650 -7955
rect -21850 -8077 -21650 -8051
rect -22425 -8155 -22025 -8134
rect -20168 -8479 -20042 -8473
rect -20168 -8549 -20148 -8479
rect -20078 -8549 -20042 -8479
rect -20168 -8564 -20042 -8549
rect -18609 -8479 -18483 -8473
rect -18609 -8549 -18589 -8479
rect -18519 -8549 -18483 -8479
rect -18609 -8564 -18483 -8549
rect -16877 -8479 -16751 -8473
rect -16877 -8549 -16857 -8479
rect -16787 -8549 -16751 -8479
rect -16877 -8564 -16751 -8549
rect -15318 -8479 -15192 -8473
rect -15318 -8549 -15298 -8479
rect -15228 -8549 -15192 -8479
rect -15318 -8564 -15192 -8549
rect -13586 -8479 -13460 -8473
rect -13586 -8549 -13566 -8479
rect -13496 -8549 -13460 -8479
rect -13586 -8564 -13460 -8549
rect -12027 -8479 -11901 -8473
rect -12027 -8549 -12007 -8479
rect -11937 -8549 -11901 -8479
rect -12027 -8564 -11901 -8549
rect -10295 -8479 -10169 -8473
rect -10295 -8549 -10275 -8479
rect -10205 -8549 -10169 -8479
rect -10295 -8564 -10169 -8549
rect -8736 -8479 -8610 -8473
rect -8736 -8549 -8716 -8479
rect -8646 -8549 -8610 -8479
rect -8736 -8564 -8610 -8549
rect -21846 -8594 -21632 -8572
rect -22661 -8696 -22027 -8662
rect -21846 -8673 -21823 -8594
rect -21654 -8673 -21632 -8594
rect -21846 -8692 -21632 -8673
rect -22661 -8836 -22623 -8696
rect -22069 -8836 -22027 -8696
rect -22661 -8875 -22027 -8836
rect -20354 -8824 -20080 -8815
rect -20354 -8896 -20345 -8824
rect -20089 -8896 -20080 -8824
rect -20354 -8905 -20080 -8896
rect -19065 -8824 -18791 -8815
rect -19065 -8896 -19056 -8824
rect -18800 -8896 -18791 -8824
rect -19065 -8905 -18791 -8896
rect -18348 -8824 -18074 -8815
rect -18348 -8896 -18339 -8824
rect -18083 -8896 -18074 -8824
rect -18348 -8905 -18074 -8896
rect -17063 -8824 -16789 -8815
rect -17063 -8896 -17054 -8824
rect -16798 -8896 -16789 -8824
rect -17063 -8905 -16789 -8896
rect -15774 -8824 -15500 -8815
rect -15774 -8896 -15765 -8824
rect -15509 -8896 -15500 -8824
rect -15774 -8905 -15500 -8896
rect -15057 -8824 -14783 -8815
rect -15057 -8896 -15048 -8824
rect -14792 -8896 -14783 -8824
rect -15057 -8905 -14783 -8896
rect -13772 -8824 -13498 -8815
rect -13772 -8896 -13763 -8824
rect -13507 -8896 -13498 -8824
rect -13772 -8905 -13498 -8896
rect -12483 -8824 -12209 -8815
rect -12483 -8896 -12474 -8824
rect -12218 -8896 -12209 -8824
rect -12483 -8905 -12209 -8896
rect -11766 -8824 -11492 -8815
rect -11766 -8896 -11757 -8824
rect -11501 -8896 -11492 -8824
rect -11766 -8905 -11492 -8896
rect -10481 -8824 -10207 -8815
rect -10481 -8896 -10472 -8824
rect -10216 -8896 -10207 -8824
rect -10481 -8905 -10207 -8896
rect -9192 -8824 -8918 -8815
rect -9192 -8896 -9183 -8824
rect -8927 -8896 -8918 -8824
rect -9192 -8905 -8918 -8896
rect -8475 -8824 -8201 -8815
rect -8475 -8896 -8466 -8824
rect -8210 -8896 -8201 -8824
rect -8475 -8905 -8201 -8896
rect -19996 -9159 -19874 -9126
rect -22937 -9685 -22866 -9239
rect -22777 -9260 -22752 -9239
rect -22937 -9706 -22862 -9685
rect -22773 -9706 -22752 -9260
rect -21846 -9247 -21646 -9219
rect -22426 -9352 -22026 -9324
rect -22426 -9426 -22397 -9352
rect -22057 -9426 -22026 -9352
rect -21846 -9343 -21819 -9247
rect -21670 -9343 -21646 -9247
rect -21846 -9369 -21646 -9343
rect -19996 -9307 -19979 -9159
rect -19896 -9307 -19874 -9159
rect -19996 -9360 -19874 -9307
rect -16705 -9159 -16583 -9126
rect -16705 -9307 -16688 -9159
rect -16605 -9307 -16583 -9159
rect -16705 -9360 -16583 -9307
rect -13414 -9159 -13292 -9126
rect -13414 -9307 -13397 -9159
rect -13314 -9307 -13292 -9159
rect -13414 -9360 -13292 -9307
rect -10123 -9159 -10001 -9126
rect -10123 -9307 -10106 -9159
rect -10023 -9307 -10001 -9159
rect -10123 -9360 -10001 -9307
rect -22426 -9447 -22026 -9426
rect -19996 -9375 -18395 -9360
rect -19996 -9450 -18561 -9375
rect -18416 -9450 -18395 -9375
rect -19996 -9462 -18395 -9450
rect -16705 -9375 -15104 -9360
rect -16705 -9450 -15270 -9375
rect -15125 -9450 -15104 -9375
rect -16705 -9462 -15104 -9450
rect -13414 -9375 -11813 -9360
rect -13414 -9450 -11979 -9375
rect -11834 -9450 -11813 -9375
rect -13414 -9462 -11813 -9450
rect -10123 -9375 -8522 -9360
rect -10123 -9450 -8688 -9375
rect -8543 -9450 -8522 -9375
rect -10123 -9462 -8522 -9450
rect 5558 -9523 5627 -4919
rect 5998 -4880 6067 -483
rect 6438 -455 6507 233
rect 11883 172 12147 178
rect 11883 -80 11889 172
rect 12141 -80 12147 172
rect 11883 -86 12147 -80
rect 6438 -514 6443 -455
rect 6502 -514 6507 -455
rect 6144 -1274 6264 -1248
rect 6144 -1340 6165 -1274
rect 6231 -1340 6264 -1274
rect 6144 -1361 6264 -1340
rect 6438 -1465 6507 -514
rect 6579 -1265 6699 -1247
rect 6579 -1331 6605 -1265
rect 6671 -1331 6699 -1265
rect 6579 -1360 6699 -1331
rect 6168 -1534 6507 -1465
rect 6168 -4240 6237 -1534
rect 6299 -1653 6367 -1648
rect 6299 -1711 6304 -1653
rect 6362 -1711 6367 -1653
rect 6299 -1754 6367 -1711
rect 12187 -1654 12431 -1648
rect 6299 -1761 10002 -1754
rect 6299 -1763 9935 -1761
rect 6299 -1819 8998 -1763
rect 9054 -1817 9935 -1763
rect 9991 -1817 10002 -1761
rect 9054 -1819 10002 -1817
rect 6299 -1822 10002 -1819
rect 6299 -3981 6365 -1822
rect 6573 -1824 10002 -1822
rect 10262 -1817 10331 -1812
rect 10262 -1876 10267 -1817
rect 10326 -1876 10331 -1817
rect 6433 -1888 6512 -1883
rect 10262 -1888 10331 -1876
rect 6433 -1957 6438 -1888
rect 6507 -1893 10331 -1888
rect 12187 -1886 12193 -1654
rect 12425 -1886 12431 -1654
rect 12187 -1892 12431 -1886
rect 6507 -1952 8541 -1893
rect 8600 -1952 10331 -1893
rect 6507 -1957 10331 -1952
rect 6433 -1962 6512 -1957
rect 6433 -2035 6507 -1962
rect 6440 -3861 6500 -2035
rect 7156 -2808 11207 -2741
rect 7156 -2996 7222 -2808
rect 7410 -2996 8157 -2808
rect 8345 -2996 9093 -2808
rect 9281 -2995 10024 -2808
rect 10211 -2995 10951 -2808
rect 9281 -2996 10951 -2995
rect 11139 -2996 11207 -2808
rect 7156 -3062 11207 -2996
rect 12414 -3232 12821 -3120
rect 12128 -3236 12821 -3232
rect 12128 -3262 13042 -3236
rect 12128 -3319 13186 -3262
rect 12128 -3448 12228 -3319
rect 12357 -3360 13186 -3319
rect 12357 -3448 12955 -3360
rect 12128 -3489 12955 -3448
rect 13084 -3489 13186 -3360
rect 12128 -3549 13186 -3489
rect 12467 -3708 13186 -3549
rect 12796 -3741 13186 -3708
rect 8398 -3860 8471 -3855
rect 8398 -3861 8405 -3860
rect 6440 -3916 8405 -3861
rect 8461 -3861 8471 -3860
rect 8461 -3892 10324 -3861
rect 8461 -3897 10327 -3892
rect 8461 -3916 10266 -3897
rect 6440 -3921 10266 -3916
rect 10261 -3953 10266 -3921
rect 10322 -3953 10327 -3897
rect 10261 -3958 10327 -3953
rect 6299 -3986 10021 -3981
rect 6299 -4047 9001 -3986
rect 8996 -4048 9001 -4047
rect 9067 -4047 9947 -3986
rect 10003 -4047 10021 -3986
rect 9067 -4048 9072 -4047
rect 8996 -4053 9072 -4048
rect 9942 -4052 10021 -4047
rect 6168 -4309 6506 -4240
rect 5998 -4939 6003 -4880
rect 6062 -4939 6067 -4880
rect 5707 -5721 5827 -5697
rect 5707 -5787 5727 -5721
rect 5793 -5787 5827 -5721
rect 5707 -5810 5827 -5787
rect -20278 -9558 -19925 -9557
rect -20278 -9622 -20269 -9558
rect -19934 -9622 -19925 -9558
rect -20278 -9631 -19925 -9622
rect -19058 -9570 -18946 -9556
rect -19058 -9642 -19038 -9570
rect -18966 -9642 -18946 -9570
rect -16987 -9558 -16634 -9557
rect -19058 -9653 -18946 -9642
rect -18191 -9595 -18088 -9581
rect -18191 -9661 -18173 -9595
rect -18107 -9661 -18088 -9595
rect -16987 -9622 -16978 -9558
rect -16643 -9622 -16634 -9558
rect -16987 -9631 -16634 -9622
rect -15767 -9570 -15655 -9556
rect -15767 -9642 -15747 -9570
rect -15675 -9642 -15655 -9570
rect -13696 -9558 -13343 -9557
rect -15767 -9653 -15655 -9642
rect -14900 -9595 -14797 -9581
rect -18191 -9679 -18088 -9661
rect -14900 -9661 -14882 -9595
rect -14816 -9661 -14797 -9595
rect -13696 -9622 -13687 -9558
rect -13352 -9622 -13343 -9558
rect -13696 -9631 -13343 -9622
rect -12476 -9570 -12364 -9556
rect -12476 -9642 -12456 -9570
rect -12384 -9642 -12364 -9570
rect -10405 -9558 -10052 -9557
rect -12476 -9653 -12364 -9642
rect -11609 -9595 -11506 -9581
rect -14900 -9679 -14797 -9661
rect -11609 -9661 -11591 -9595
rect -11525 -9661 -11506 -9595
rect -10405 -9622 -10396 -9558
rect -10061 -9622 -10052 -9558
rect -10405 -9631 -10052 -9622
rect -9185 -9570 -9073 -9556
rect -9185 -9642 -9165 -9570
rect -9093 -9642 -9073 -9570
rect -9185 -9653 -9073 -9642
rect -8318 -9595 -8215 -9581
rect -11609 -9679 -11506 -9661
rect -8318 -9661 -8300 -9595
rect -8234 -9661 -8215 -9595
rect -8318 -9679 -8215 -9661
rect 5558 -9582 5563 -9523
rect 5622 -9582 5627 -9523
rect -22937 -11019 -22752 -9706
rect -20649 -10356 -19439 -10328
rect -20649 -10428 -20603 -10356
rect -19481 -10428 -19439 -10356
rect -20649 -10454 -19439 -10428
rect -19090 -10356 -17880 -10328
rect -19090 -10428 -19044 -10356
rect -17922 -10428 -17880 -10356
rect -19090 -10454 -17880 -10428
rect -17358 -10356 -16148 -10328
rect -17358 -10428 -17312 -10356
rect -16190 -10428 -16148 -10356
rect -17358 -10454 -16148 -10428
rect -15799 -10356 -14589 -10328
rect -15799 -10428 -15753 -10356
rect -14631 -10428 -14589 -10356
rect -15799 -10454 -14589 -10428
rect -14067 -10356 -12857 -10328
rect -14067 -10428 -14021 -10356
rect -12899 -10428 -12857 -10356
rect -14067 -10454 -12857 -10428
rect -12508 -10356 -11298 -10328
rect -12508 -10428 -12462 -10356
rect -11340 -10428 -11298 -10356
rect -12508 -10454 -11298 -10428
rect -10776 -10356 -9566 -10328
rect -10776 -10428 -10730 -10356
rect -9608 -10428 -9566 -10356
rect -10776 -10454 -9566 -10428
rect -9217 -10356 -8007 -10328
rect -9217 -10428 -9171 -10356
rect -8049 -10428 -8007 -10356
rect -9217 -10454 -8007 -10428
rect -21850 -10566 -21636 -10544
rect -22660 -10668 -22026 -10634
rect -21850 -10645 -21827 -10566
rect -21658 -10645 -21636 -10566
rect -21850 -10664 -21636 -10645
rect -22660 -10808 -22622 -10668
rect -22068 -10808 -22026 -10668
rect -22660 -10847 -22026 -10808
rect -22937 -11113 -22650 -11019
rect -22937 -11179 -22752 -11113
rect -23583 -11219 -23383 -11191
rect -24162 -11324 -23762 -11296
rect -24162 -11398 -24133 -11324
rect -23793 -11398 -23762 -11324
rect -23583 -11315 -23556 -11219
rect -23407 -11315 -23383 -11219
rect -23583 -11341 -23383 -11315
rect -22937 -11275 -22644 -11179
rect -21850 -11219 -21650 -11191
rect -24162 -11419 -23762 -11398
rect -23583 -11858 -23369 -11836
rect -24397 -11960 -23763 -11926
rect -23583 -11937 -23560 -11858
rect -23391 -11937 -23369 -11858
rect -23583 -11956 -23369 -11937
rect -24397 -12100 -24359 -11960
rect -23805 -12100 -23763 -11960
rect -24397 -12139 -23763 -12100
rect -23583 -12511 -23383 -12483
rect -24651 -12578 -24439 -12549
rect -24651 -12776 -24612 -12578
rect -24466 -12776 -24439 -12578
rect -24162 -12616 -23762 -12588
rect -24162 -12690 -24133 -12616
rect -23793 -12690 -23762 -12616
rect -23583 -12607 -23556 -12511
rect -23407 -12607 -23383 -12511
rect -23583 -12633 -23383 -12607
rect -22937 -12503 -22752 -11275
rect -22425 -11324 -22025 -11296
rect -22425 -11398 -22396 -11324
rect -22056 -11398 -22025 -11324
rect -21850 -11315 -21823 -11219
rect -21674 -11315 -21650 -11219
rect -21850 -11341 -21650 -11315
rect -22425 -11419 -22025 -11398
rect -20168 -11743 -20042 -11737
rect -20168 -11813 -20148 -11743
rect -20078 -11813 -20042 -11743
rect -20168 -11828 -20042 -11813
rect -18609 -11743 -18483 -11737
rect -18609 -11813 -18589 -11743
rect -18519 -11813 -18483 -11743
rect -18609 -11828 -18483 -11813
rect -16877 -11743 -16751 -11737
rect -16877 -11813 -16857 -11743
rect -16787 -11813 -16751 -11743
rect -16877 -11828 -16751 -11813
rect -15318 -11743 -15192 -11737
rect -15318 -11813 -15298 -11743
rect -15228 -11813 -15192 -11743
rect -15318 -11828 -15192 -11813
rect -13586 -11743 -13460 -11737
rect -13586 -11813 -13566 -11743
rect -13496 -11813 -13460 -11743
rect -13586 -11828 -13460 -11813
rect -12027 -11743 -11901 -11737
rect -12027 -11813 -12007 -11743
rect -11937 -11813 -11901 -11743
rect -12027 -11828 -11901 -11813
rect -10295 -11743 -10169 -11737
rect -10295 -11813 -10275 -11743
rect -10205 -11813 -10169 -11743
rect -10295 -11828 -10169 -11813
rect -8736 -11743 -8610 -11737
rect -8736 -11813 -8716 -11743
rect -8646 -11813 -8610 -11743
rect -8736 -11828 -8610 -11813
rect -21854 -11858 -21640 -11836
rect -22660 -11960 -22026 -11926
rect -21854 -11937 -21831 -11858
rect -21662 -11937 -21640 -11858
rect -21854 -11956 -21640 -11937
rect -22660 -12100 -22622 -11960
rect -22068 -12100 -22026 -11960
rect -22660 -12139 -22026 -12100
rect -20354 -12088 -20080 -12079
rect -20354 -12160 -20345 -12088
rect -20089 -12160 -20080 -12088
rect -20354 -12169 -20080 -12160
rect -19065 -12088 -18791 -12079
rect -19065 -12160 -19056 -12088
rect -18800 -12160 -18791 -12088
rect -19065 -12169 -18791 -12160
rect -18348 -12088 -18074 -12079
rect -18348 -12160 -18339 -12088
rect -18083 -12160 -18074 -12088
rect -18348 -12169 -18074 -12160
rect -17063 -12088 -16789 -12079
rect -17063 -12160 -17054 -12088
rect -16798 -12160 -16789 -12088
rect -17063 -12169 -16789 -12160
rect -15774 -12088 -15500 -12079
rect -15774 -12160 -15765 -12088
rect -15509 -12160 -15500 -12088
rect -15774 -12169 -15500 -12160
rect -15057 -12088 -14783 -12079
rect -15057 -12160 -15048 -12088
rect -14792 -12160 -14783 -12088
rect -15057 -12169 -14783 -12160
rect -13772 -12088 -13498 -12079
rect -13772 -12160 -13763 -12088
rect -13507 -12160 -13498 -12088
rect -13772 -12169 -13498 -12160
rect -12483 -12088 -12209 -12079
rect -12483 -12160 -12474 -12088
rect -12218 -12160 -12209 -12088
rect -12483 -12169 -12209 -12160
rect -11766 -12088 -11492 -12079
rect -11766 -12160 -11757 -12088
rect -11501 -12160 -11492 -12088
rect -11766 -12169 -11492 -12160
rect -10481 -12088 -10207 -12079
rect -10481 -12160 -10472 -12088
rect -10216 -12160 -10207 -12088
rect -10481 -12169 -10207 -12160
rect -9192 -12088 -8918 -12079
rect -9192 -12160 -9183 -12088
rect -8927 -12160 -8918 -12088
rect -9192 -12169 -8918 -12160
rect -8475 -12088 -8201 -12079
rect -8475 -12160 -8466 -12088
rect -8210 -12160 -8201 -12088
rect -8475 -12169 -8201 -12160
rect -19996 -12423 -19874 -12390
rect -22937 -12518 -22866 -12503
rect -24162 -12711 -23762 -12690
rect -24651 -12791 -24439 -12776
rect -24651 -13003 -24460 -12791
rect -22937 -12964 -22869 -12518
rect -22777 -12524 -22752 -12503
rect -22937 -12970 -22862 -12964
rect -22773 -12970 -22752 -12524
rect -21854 -12511 -21654 -12483
rect -22425 -12616 -22025 -12588
rect -22425 -12690 -22396 -12616
rect -22056 -12690 -22025 -12616
rect -21854 -12607 -21827 -12511
rect -21678 -12607 -21654 -12511
rect -21854 -12633 -21654 -12607
rect -19996 -12571 -19979 -12423
rect -19896 -12571 -19874 -12423
rect -19996 -12624 -19874 -12571
rect -16705 -12423 -16583 -12390
rect -16705 -12571 -16688 -12423
rect -16605 -12571 -16583 -12423
rect -16705 -12624 -16583 -12571
rect -13414 -12423 -13292 -12390
rect -13414 -12571 -13397 -12423
rect -13314 -12571 -13292 -12423
rect -13414 -12624 -13292 -12571
rect -10123 -12423 -10001 -12390
rect -10123 -12571 -10106 -12423
rect -10023 -12571 -10001 -12423
rect -10123 -12624 -10001 -12571
rect -22425 -12711 -22025 -12690
rect -19996 -12639 -18395 -12624
rect -19996 -12714 -18561 -12639
rect -18416 -12714 -18395 -12639
rect -19996 -12726 -18395 -12714
rect -16705 -12639 -15104 -12624
rect -16705 -12714 -15270 -12639
rect -15125 -12714 -15104 -12639
rect -16705 -12726 -15104 -12714
rect -13414 -12639 -11813 -12624
rect -13414 -12714 -11979 -12639
rect -11834 -12714 -11813 -12639
rect -13414 -12726 -11813 -12714
rect -10123 -12639 -8522 -12624
rect -10123 -12714 -8688 -12639
rect -8543 -12714 -8522 -12639
rect -10123 -12726 -8522 -12714
rect -20278 -12822 -19925 -12821
rect -20278 -12886 -20269 -12822
rect -19934 -12886 -19925 -12822
rect -20278 -12895 -19925 -12886
rect -19058 -12834 -18946 -12820
rect -19058 -12906 -19038 -12834
rect -18966 -12906 -18946 -12834
rect -16987 -12822 -16634 -12821
rect -19058 -12917 -18946 -12906
rect -18191 -12859 -18088 -12845
rect -18191 -12925 -18173 -12859
rect -18107 -12925 -18088 -12859
rect -16987 -12886 -16978 -12822
rect -16643 -12886 -16634 -12822
rect -16987 -12895 -16634 -12886
rect -15767 -12834 -15655 -12820
rect -15767 -12906 -15747 -12834
rect -15675 -12906 -15655 -12834
rect -13696 -12822 -13343 -12821
rect -15767 -12917 -15655 -12906
rect -14900 -12859 -14797 -12845
rect -18191 -12943 -18088 -12925
rect -14900 -12925 -14882 -12859
rect -14816 -12925 -14797 -12859
rect -13696 -12886 -13687 -12822
rect -13352 -12886 -13343 -12822
rect -13696 -12895 -13343 -12886
rect -12476 -12834 -12364 -12820
rect -12476 -12906 -12456 -12834
rect -12384 -12906 -12364 -12834
rect -10405 -12822 -10052 -12821
rect -12476 -12917 -12364 -12906
rect -11609 -12859 -11506 -12845
rect -14900 -12943 -14797 -12925
rect -11609 -12925 -11591 -12859
rect -11525 -12925 -11506 -12859
rect -10405 -12886 -10396 -12822
rect -10061 -12886 -10052 -12822
rect -10405 -12895 -10052 -12886
rect -9185 -12834 -9073 -12820
rect -9185 -12906 -9165 -12834
rect -9093 -12906 -9073 -12834
rect -9185 -12917 -9073 -12906
rect -8318 -12859 -8215 -12845
rect -11609 -12943 -11506 -12925
rect -8318 -12925 -8300 -12859
rect -8234 -12925 -8215 -12859
rect -8318 -12943 -8215 -12925
rect -22937 -13013 -22752 -12970
rect 5558 -14050 5627 -9582
rect 5998 -9528 6067 -4939
rect 6437 -4889 6506 -4309
rect 11883 -4356 12147 -4350
rect 11883 -4608 11889 -4356
rect 12141 -4608 12147 -4356
rect 11883 -4614 12147 -4608
rect 6437 -4948 6442 -4889
rect 6501 -4948 6506 -4889
rect 6144 -5702 6264 -5676
rect 6144 -5768 6165 -5702
rect 6231 -5768 6264 -5702
rect 6144 -5789 6264 -5768
rect 6437 -5912 6506 -4948
rect 6579 -5693 6699 -5675
rect 6579 -5759 6605 -5693
rect 6671 -5759 6699 -5693
rect 6579 -5788 6699 -5759
rect 6165 -5981 6506 -5912
rect 6165 -9037 6234 -5981
rect 6299 -6081 6367 -6076
rect 6299 -6139 6304 -6081
rect 6362 -6139 6367 -6081
rect 6299 -6182 6367 -6139
rect 12187 -6082 12431 -6076
rect 6299 -6189 10002 -6182
rect 6299 -6191 9935 -6189
rect 6299 -6247 8998 -6191
rect 9054 -6245 9935 -6191
rect 9991 -6245 10002 -6189
rect 9054 -6247 10002 -6245
rect 6299 -6250 10002 -6247
rect 6299 -8409 6365 -6250
rect 6573 -6252 10002 -6250
rect 10262 -6245 10331 -6240
rect 10262 -6304 10267 -6245
rect 10326 -6304 10331 -6245
rect 6433 -6316 6512 -6311
rect 10262 -6316 10331 -6304
rect 6433 -6385 6438 -6316
rect 6507 -6321 10331 -6316
rect 12187 -6314 12193 -6082
rect 12425 -6314 12431 -6082
rect 12187 -6320 12431 -6314
rect 6507 -6380 8541 -6321
rect 8600 -6380 10331 -6321
rect 6507 -6385 10331 -6380
rect 6433 -6390 6512 -6385
rect 6433 -6463 6507 -6390
rect 6440 -8289 6500 -6463
rect 7156 -7236 11207 -7169
rect 7156 -7424 7222 -7236
rect 7410 -7424 8157 -7236
rect 8345 -7424 9093 -7236
rect 9281 -7423 10024 -7236
rect 10211 -7423 10951 -7236
rect 9281 -7424 10951 -7423
rect 11139 -7424 11207 -7236
rect 7156 -7490 11207 -7424
rect 12414 -7660 12821 -7548
rect 12128 -7664 12821 -7660
rect 12128 -7690 13042 -7664
rect 12128 -7747 13186 -7690
rect 12128 -7876 12228 -7747
rect 12357 -7788 13186 -7747
rect 12357 -7876 12955 -7788
rect 12128 -7917 12955 -7876
rect 13084 -7917 13186 -7788
rect 12128 -7977 13186 -7917
rect 12467 -8136 13186 -7977
rect 12796 -8169 13186 -8136
rect 8398 -8288 8471 -8283
rect 8398 -8289 8405 -8288
rect 6440 -8344 8405 -8289
rect 8461 -8289 8471 -8288
rect 8461 -8320 10324 -8289
rect 8461 -8325 10327 -8320
rect 8461 -8344 10266 -8325
rect 6440 -8349 10266 -8344
rect 10261 -8381 10266 -8349
rect 10322 -8381 10327 -8325
rect 10261 -8386 10327 -8381
rect 6299 -8414 10021 -8409
rect 6299 -8475 9001 -8414
rect 8996 -8476 9001 -8475
rect 9067 -8475 9947 -8414
rect 10003 -8475 10021 -8414
rect 9067 -8476 9072 -8475
rect 8996 -8481 9072 -8476
rect 9942 -8480 10021 -8475
rect 11883 -8784 12147 -8778
rect 11883 -9036 11889 -8784
rect 12141 -9036 12147 -8784
rect 6165 -9106 6509 -9037
rect 11883 -9042 12147 -9036
rect 5998 -9587 6003 -9528
rect 6062 -9587 6067 -9528
rect 5707 -10349 5827 -10325
rect 5707 -10415 5727 -10349
rect 5793 -10415 5827 -10349
rect 5707 -10438 5827 -10415
rect -2315 -14172 -2309 -14058
rect -2195 -14172 -2189 -14058
rect -1299 -14176 -1293 -14069
rect -1186 -14176 -1180 -14069
rect 5558 -14109 5563 -14050
rect 5622 -14109 5627 -14050
rect -12501 -14223 -12375 -14181
rect -23450 -15070 -23287 -15051
rect -23450 -15181 -23426 -15070
rect -23315 -15181 -23287 -15070
rect -24851 -15189 -24731 -15182
rect -24851 -15295 -24844 -15189
rect -24738 -15295 -24731 -15189
rect -23450 -15207 -23287 -15181
rect -24851 -15302 -24731 -15295
rect -18084 -15276 -17986 -15269
rect -18084 -15360 -18077 -15276
rect -17993 -15360 -17986 -15276
rect -18084 -15367 -17986 -15360
rect -16938 -15321 -16822 -15295
rect -16938 -15391 -16914 -15321
rect -16844 -15391 -16822 -15321
rect -12501 -15345 -12473 -14223
rect -12401 -15345 -12375 -14223
rect -5026 -14255 -4910 -14254
rect -5031 -14369 -5025 -14255
rect -4911 -14369 -4905 -14255
rect -4015 -14352 -4009 -14245
rect -3902 -14352 -3896 -14245
rect -5026 -14370 -4910 -14369
rect -6212 -14496 -2216 -14494
rect -6780 -14499 -2216 -14496
rect -6780 -14561 -5003 -14499
rect -4941 -14561 -2283 -14499
rect -2221 -14561 -2216 -14499
rect -6780 -14566 -2216 -14561
rect -6780 -14568 -6124 -14566
rect -11092 -14820 -11001 -14784
rect -11092 -14890 -11086 -14820
rect -11016 -14890 -11001 -14820
rect -11092 -14910 -11001 -14890
rect -12501 -15391 -12375 -15345
rect -16938 -15417 -16822 -15391
rect -8533 -15420 -8408 -15374
rect -8533 -15490 -8499 -15420
rect -8429 -15490 -8408 -15420
rect -8676 -15501 -8604 -15496
rect -8676 -15563 -8671 -15501
rect -8609 -15563 -8604 -15501
rect -8533 -15540 -8408 -15490
rect -7209 -15392 -7110 -15386
rect -7209 -15497 -7110 -15491
rect -24921 -15586 -24839 -15581
rect -12730 -15586 -12656 -15570
rect -25221 -15658 -24916 -15586
rect -24844 -15591 -9810 -15586
rect -24844 -15653 -17961 -15591
rect -17899 -15653 -12719 -15591
rect -12657 -15632 -9810 -15591
rect -8676 -15632 -8604 -15563
rect -6780 -15632 -6708 -14568
rect -5031 -14996 -5025 -14882
rect -4911 -14996 -4905 -14882
rect -4015 -14985 -4009 -14878
rect -3902 -14985 -3896 -14878
rect -2315 -14991 -2309 -14877
rect -2195 -14991 -2189 -14877
rect -1299 -14995 -1293 -14888
rect -1186 -14995 -1180 -14888
rect -6596 -15311 -2184 -15306
rect -6596 -15373 -4961 -15311
rect -4899 -15373 -2259 -15311
rect -2197 -15373 -2184 -15311
rect -6596 -15378 -2184 -15373
rect -12657 -15653 -6688 -15632
rect -24844 -15658 -6688 -15653
rect -24921 -15663 -24839 -15658
rect -12730 -15666 -12656 -15658
rect -9882 -15704 -6688 -15658
rect -9882 -15708 -9810 -15704
rect -24908 -15738 -24807 -15734
rect -12560 -15738 -12451 -15733
rect -25370 -15739 -12555 -15738
rect -25370 -15827 -24903 -15739
rect -24908 -15828 -24903 -15827
rect -24812 -15743 -12555 -15739
rect -24812 -15822 -18118 -15743
rect -18039 -15822 -12555 -15743
rect -24812 -15827 -12555 -15822
rect -24812 -15828 -24807 -15827
rect -24908 -15833 -24807 -15828
rect -12560 -15837 -12555 -15827
rect -12456 -15827 -10774 -15738
rect -12456 -15837 -12451 -15827
rect -12560 -15842 -12451 -15837
rect -8535 -15929 -8408 -15882
rect -8535 -15999 -8505 -15929
rect -8435 -15999 -8408 -15929
rect -7216 -15885 -7117 -15879
rect -7216 -15990 -7117 -15984
rect -8535 -16037 -8408 -15999
rect -6596 -16152 -6524 -15378
rect -5031 -15815 -5025 -15701
rect -4911 -15815 -4905 -15701
rect -4015 -15804 -4009 -15697
rect -3902 -15804 -3896 -15697
rect -2315 -15810 -2309 -15696
rect -2195 -15810 -2189 -15696
rect -1299 -15814 -1293 -15707
rect -1186 -15814 -1180 -15707
rect -6209 -16130 -2203 -16125
rect -10052 -16157 -6510 -16152
rect -10052 -16219 -8549 -16157
rect -8487 -16219 -6510 -16157
rect -10052 -16224 -6510 -16219
rect -6209 -16190 -4990 -16130
rect -4930 -16190 -2280 -16130
rect -2220 -16190 -2203 -16130
rect -6209 -16195 -2203 -16190
rect -23407 -16266 -23244 -16247
rect -24847 -16363 -24727 -16356
rect -24847 -16469 -24840 -16363
rect -24734 -16469 -24727 -16363
rect -23407 -16377 -23383 -16266
rect -23272 -16377 -23244 -16266
rect -23407 -16403 -23244 -16377
rect -24847 -16476 -24727 -16469
rect -18096 -16678 -17998 -16671
rect -18096 -16762 -18089 -16678
rect -18005 -16762 -17998 -16678
rect -24913 -16770 -24831 -16765
rect -18096 -16769 -17998 -16762
rect -16938 -16727 -16822 -16699
rect -25509 -16842 -24908 -16770
rect -24836 -16842 -18526 -16770
rect -16938 -16797 -16914 -16727
rect -16844 -16797 -16822 -16727
rect -16938 -16821 -16822 -16797
rect -24913 -16847 -24831 -16842
rect -24920 -16922 -24831 -16918
rect -25660 -16923 -18736 -16922
rect -25660 -17011 -24915 -16923
rect -24920 -17012 -24915 -17011
rect -24836 -17011 -18736 -16923
rect -24836 -17012 -24831 -17011
rect -24920 -17017 -24831 -17012
rect -18825 -17113 -18736 -17011
rect -18598 -16980 -18526 -16842
rect -18598 -16985 -13076 -16980
rect -18598 -17047 -18077 -16985
rect -18015 -17047 -13076 -16985
rect -18598 -17052 -13076 -17047
rect -18825 -17118 -17178 -17113
rect -18825 -17197 -18085 -17118
rect -18005 -17155 -17178 -17118
rect -18005 -17197 -13292 -17155
rect -18825 -17202 -13292 -17197
rect -17304 -17244 -13292 -17202
rect -23398 -17478 -23235 -17459
rect -24841 -17595 -24721 -17588
rect -24841 -17701 -24834 -17595
rect -24728 -17701 -24721 -17595
rect -23398 -17589 -23374 -17478
rect -23263 -17589 -23235 -17478
rect -23398 -17615 -23235 -17589
rect -24841 -17708 -24721 -17701
rect -22395 -17977 -18413 -17907
rect -24926 -17984 -24846 -17979
rect -22395 -17984 -22325 -17977
rect -25814 -18054 -24921 -17984
rect -24851 -18054 -22325 -17984
rect -24926 -18059 -24846 -18054
rect -21972 -18108 -21847 -18062
rect -24922 -18127 -24819 -18123
rect -25983 -18128 -22118 -18127
rect -25983 -18216 -24917 -18128
rect -24922 -18217 -24917 -18216
rect -24824 -18216 -22118 -18128
rect -24824 -18217 -24819 -18216
rect -24922 -18222 -24819 -18217
rect -22207 -18315 -22118 -18216
rect -21972 -18178 -21938 -18108
rect -21868 -18178 -21847 -18108
rect -21972 -18228 -21847 -18178
rect -20648 -18080 -20549 -18074
rect -20648 -18185 -20549 -18179
rect -22207 -18404 -18592 -18315
rect -18681 -18515 -18592 -18404
rect -18483 -18385 -18413 -17977
rect -16381 -17979 -16256 -17933
rect -16381 -18049 -16347 -17979
rect -16277 -18049 -16256 -17979
rect -18100 -18064 -18002 -18057
rect -18100 -18148 -18093 -18064
rect -18009 -18148 -18002 -18064
rect -16381 -18099 -16256 -18049
rect -15057 -17951 -14958 -17945
rect -15057 -18056 -14958 -18050
rect -18100 -18155 -18002 -18148
rect -17074 -18158 -16948 -18133
rect -17074 -18228 -17045 -18158
rect -16975 -18228 -16948 -18158
rect -17074 -18255 -16948 -18228
rect -16571 -18301 -13459 -18231
rect -16571 -18385 -16501 -18301
rect -18483 -18390 -16501 -18385
rect -18483 -18450 -18060 -18390
rect -18000 -18450 -16501 -18390
rect -18483 -18455 -16501 -18450
rect -16383 -18488 -16256 -18441
rect -18681 -18520 -16570 -18515
rect -23390 -18619 -23227 -18600
rect -24827 -18709 -24707 -18702
rect -24827 -18815 -24820 -18709
rect -24714 -18815 -24707 -18709
rect -23390 -18730 -23366 -18619
rect -23255 -18730 -23227 -18619
rect -21974 -18617 -21847 -18570
rect -21974 -18687 -21944 -18617
rect -21874 -18687 -21847 -18617
rect -20655 -18573 -20556 -18567
rect -18681 -18599 -18094 -18520
rect -18015 -18599 -16570 -18520
rect -16383 -18558 -16353 -18488
rect -16283 -18558 -16256 -18488
rect -15064 -18444 -14965 -18438
rect -15064 -18549 -14965 -18543
rect -16383 -18596 -16256 -18558
rect -18681 -18604 -16570 -18599
rect -20655 -18678 -20556 -18672
rect -21974 -18725 -21847 -18687
rect -16659 -18695 -16570 -18604
rect -23390 -18756 -23227 -18730
rect -16659 -18784 -13618 -18695
rect -24827 -18822 -24707 -18815
rect -13707 -18903 -13618 -18784
rect -13529 -18769 -13459 -18301
rect -13381 -18573 -13292 -17244
rect -13148 -18396 -13076 -17052
rect -12499 -17039 -12373 -16997
rect -12499 -18161 -12471 -17039
rect -12399 -18161 -12373 -17039
rect -11090 -17636 -10999 -17600
rect -11090 -17706 -11084 -17636
rect -11014 -17706 -10999 -17636
rect -11090 -17726 -10999 -17706
rect -12499 -18207 -12373 -18161
rect -10052 -18396 -9980 -16224
rect -8535 -16412 -8408 -16356
rect -8535 -16482 -8505 -16412
rect -8435 -16482 -8408 -16412
rect -7217 -16371 -7118 -16365
rect -7217 -16476 -7118 -16470
rect -8535 -16525 -8408 -16482
rect -8556 -16685 -8477 -16680
rect -8556 -16687 -8551 -16685
rect -13148 -18401 -9980 -18396
rect -13148 -18463 -12661 -18401
rect -12599 -18463 -9980 -18401
rect -13148 -18468 -9980 -18463
rect -9825 -16754 -8551 -16687
rect -8482 -16687 -8477 -16685
rect -6209 -16687 -6139 -16195
rect -5031 -16634 -5025 -16520
rect -4911 -16634 -4905 -16520
rect -4015 -16623 -4009 -16516
rect -3902 -16623 -3896 -16516
rect -2315 -16629 -2309 -16515
rect -2195 -16629 -2189 -16515
rect -1299 -16633 -1293 -16526
rect -1186 -16633 -1180 -16526
rect -8482 -16754 -6139 -16687
rect -9825 -16757 -6139 -16754
rect -13381 -18578 -12544 -18573
rect -13381 -18657 -12628 -18578
rect -12549 -18657 -12544 -18578
rect -13381 -18662 -12544 -18657
rect -13529 -18839 -12679 -18769
rect -22106 -18980 -18438 -18908
rect -16383 -18971 -16256 -18915
rect -24875 -19103 -24793 -19098
rect -22106 -19103 -22034 -18980
rect -26169 -19175 -24870 -19103
rect -24798 -19175 -22034 -19103
rect -21974 -19100 -21847 -19044
rect -21974 -19170 -21944 -19100
rect -21874 -19170 -21847 -19100
rect -20656 -19059 -20557 -19053
rect -20656 -19164 -20557 -19158
rect -24875 -19180 -24793 -19175
rect -21974 -19213 -21847 -19170
rect -24880 -19255 -24791 -19251
rect -26332 -19256 -22060 -19255
rect -26332 -19344 -24875 -19256
rect -24880 -19345 -24875 -19344
rect -24796 -19344 -22060 -19256
rect -24796 -19345 -24791 -19344
rect -24880 -19350 -24791 -19345
rect -22149 -19385 -22060 -19344
rect -22149 -19474 -18636 -19385
rect -20660 -19566 -20561 -19560
rect -21974 -19622 -21847 -19578
rect -21974 -19692 -21944 -19622
rect -21874 -19692 -21847 -19622
rect -20660 -19671 -20561 -19665
rect -21974 -19729 -21847 -19692
rect -23367 -19791 -23204 -19772
rect -24827 -19903 -24707 -19896
rect -24827 -20009 -24820 -19903
rect -24714 -20009 -24707 -19903
rect -23367 -19902 -23343 -19791
rect -23232 -19902 -23204 -19791
rect -23367 -19928 -23204 -19902
rect -18725 -19907 -18636 -19474
rect -18506 -19780 -18442 -18980
rect -16383 -19041 -16353 -18971
rect -16283 -19041 -16256 -18971
rect -15065 -18930 -14966 -18924
rect -13707 -18992 -12844 -18903
rect -15065 -19035 -14966 -19029
rect -16383 -19084 -16256 -19041
rect -15069 -19437 -14970 -19431
rect -18098 -19470 -18000 -19463
rect -18098 -19554 -18091 -19470
rect -18007 -19554 -18000 -19470
rect -18098 -19561 -18000 -19554
rect -16383 -19493 -16256 -19449
rect -16383 -19563 -16353 -19493
rect -16283 -19563 -16256 -19493
rect -15069 -19542 -14970 -19536
rect -16952 -19613 -16838 -19589
rect -16383 -19600 -16256 -19563
rect -18018 -19626 -17952 -19621
rect -18018 -19682 -18013 -19626
rect -17957 -19682 -17952 -19626
rect -18018 -19687 -17952 -19682
rect -16952 -19683 -16930 -19613
rect -16860 -19683 -16838 -19613
rect -18017 -19780 -17954 -19687
rect -16952 -19703 -16838 -19683
rect -18506 -19843 -13041 -19780
rect -18506 -19844 -18442 -19843
rect -18725 -19912 -16507 -19907
rect -18725 -19973 -17981 -19912
rect -17920 -19973 -16507 -19912
rect -15068 -19912 -14969 -19906
rect -18725 -19978 -16507 -19973
rect -24827 -20016 -24707 -20009
rect -20659 -20041 -20560 -20035
rect -21964 -20091 -21847 -20044
rect -21964 -20161 -21941 -20091
rect -21871 -20161 -21847 -20091
rect -20659 -20146 -20560 -20140
rect -16578 -20132 -16507 -19978
rect -16373 -19962 -16256 -19915
rect -16373 -20032 -16350 -19962
rect -16280 -20032 -16256 -19962
rect -15068 -20017 -14969 -20011
rect -16373 -20070 -16256 -20032
rect -21964 -20199 -21847 -20161
rect -16578 -20203 -13191 -20132
rect -24941 -20291 -24859 -20286
rect -26500 -20363 -24936 -20291
rect -24864 -20363 -18314 -20291
rect -24941 -20368 -24859 -20363
rect -24907 -20443 -24806 -20439
rect -26650 -20444 -22144 -20443
rect -26650 -20532 -24902 -20444
rect -24907 -20533 -24902 -20532
rect -24811 -20532 -22144 -20444
rect -20654 -20493 -20555 -20487
rect -24811 -20533 -24806 -20532
rect -24907 -20538 -24806 -20533
rect -22233 -20717 -22144 -20532
rect -21959 -20548 -21848 -20526
rect -21959 -20618 -21939 -20548
rect -21869 -20618 -21848 -20548
rect -20654 -20598 -20555 -20592
rect -21959 -20641 -21848 -20618
rect -22233 -20806 -18498 -20717
rect -20654 -20935 -20555 -20929
rect -23358 -20989 -23195 -20970
rect -24827 -21099 -24707 -21092
rect -24827 -21205 -24820 -21099
rect -24714 -21205 -24707 -21099
rect -23358 -21100 -23334 -20989
rect -23223 -21100 -23195 -20989
rect -23358 -21126 -23195 -21100
rect -21952 -21013 -21852 -20994
rect -21952 -21083 -21937 -21013
rect -21867 -21083 -21852 -21013
rect -20654 -21040 -20555 -21034
rect -21952 -21105 -21852 -21083
rect -24827 -21212 -24707 -21205
rect -18587 -21340 -18498 -20806
rect -18380 -21177 -18319 -20363
rect -15063 -20364 -14964 -20358
rect -16368 -20419 -16257 -20397
rect -16368 -20489 -16348 -20419
rect -16278 -20489 -16257 -20419
rect -15063 -20469 -14964 -20463
rect -16368 -20512 -16257 -20489
rect -15063 -20806 -14964 -20800
rect -18102 -20864 -18004 -20857
rect -18102 -20948 -18095 -20864
rect -18011 -20948 -18004 -20864
rect -18102 -20955 -18004 -20948
rect -16361 -20884 -16261 -20865
rect -16361 -20954 -16346 -20884
rect -16276 -20954 -16261 -20884
rect -15063 -20911 -14964 -20905
rect -16361 -20976 -16261 -20954
rect -16938 -21008 -16830 -20989
rect -16938 -21080 -16921 -21008
rect -16849 -21080 -16830 -21008
rect -16938 -21099 -16830 -21080
rect -18056 -21177 -17990 -21174
rect -16037 -21177 -13362 -21120
rect -18380 -21179 -13362 -21177
rect -18380 -21235 -18051 -21179
rect -17995 -21181 -13362 -21179
rect -17995 -21235 -15976 -21181
rect -18380 -21238 -15976 -21235
rect -18056 -21240 -17990 -21238
rect -15091 -21287 -14944 -21261
rect -17969 -21340 -17903 -21339
rect -18587 -21344 -16574 -21340
rect -18587 -21350 -17964 -21344
rect -20682 -21416 -20535 -21390
rect -18574 -21400 -17964 -21350
rect -17908 -21400 -16574 -21344
rect -18574 -21404 -16574 -21400
rect -17969 -21405 -17903 -21404
rect -24919 -21497 -24847 -21492
rect -21969 -21494 -21830 -21441
rect -26782 -21569 -24914 -21497
rect -24852 -21569 -22110 -21497
rect -24919 -21574 -24847 -21569
rect -26921 -21649 -26832 -21642
rect -24918 -21649 -24818 -21645
rect -26921 -21650 -22298 -21649
rect -26921 -21738 -24913 -21650
rect -24918 -21739 -24913 -21738
rect -24823 -21738 -22298 -21650
rect -24823 -21739 -24818 -21738
rect -24918 -21744 -24818 -21739
rect -23361 -22283 -23198 -22264
rect -23361 -22394 -23337 -22283
rect -23226 -22394 -23198 -22283
rect -24817 -22407 -24697 -22400
rect -24817 -22513 -24810 -22407
rect -24704 -22513 -24697 -22407
rect -23361 -22420 -23198 -22394
rect -24817 -22520 -24697 -22513
rect -22387 -22745 -22298 -21738
rect -22182 -22586 -22110 -21569
rect -21969 -21564 -21933 -21494
rect -21863 -21564 -21830 -21494
rect -20682 -21515 -20660 -21416
rect -20561 -21515 -20535 -21416
rect -20682 -21540 -20535 -21515
rect -21969 -21605 -21830 -21564
rect -16638 -21578 -16574 -21404
rect -16378 -21365 -16239 -21312
rect -16378 -21435 -16342 -21365
rect -16272 -21435 -16239 -21365
rect -15091 -21386 -15069 -21287
rect -14970 -21386 -14944 -21287
rect -15091 -21411 -14944 -21386
rect -16378 -21476 -16239 -21435
rect -16638 -21642 -13506 -21578
rect -16744 -21978 -16644 -21967
rect -16744 -22052 -16731 -21978
rect -16657 -22052 -16644 -21978
rect -16744 -22065 -16644 -22052
rect -18100 -22268 -18002 -22261
rect -18100 -22352 -18093 -22268
rect -18009 -22352 -18002 -22268
rect -18100 -22359 -18002 -22352
rect -22182 -22600 -13654 -22586
rect -22182 -22658 -18061 -22600
rect -18066 -22666 -18061 -22658
rect -17995 -22658 -13654 -22600
rect -17995 -22666 -17990 -22658
rect -18066 -22671 -17990 -22666
rect -22387 -22750 -13824 -22745
rect -24895 -22798 -24813 -22793
rect -27070 -22870 -24890 -22798
rect -24818 -22870 -22488 -22798
rect -22387 -22829 -18067 -22750
rect -17987 -22829 -13824 -22750
rect -22387 -22834 -13824 -22829
rect -24895 -22875 -24813 -22870
rect -24918 -22950 -24814 -22946
rect -27210 -22951 -22674 -22950
rect -27210 -23039 -24913 -22951
rect -24918 -23040 -24913 -23039
rect -24819 -23039 -22674 -22951
rect -24819 -23040 -24814 -23039
rect -24918 -23045 -24814 -23040
rect -23401 -23599 -23238 -23580
rect -24837 -23713 -24717 -23706
rect -24837 -23819 -24830 -23713
rect -24724 -23819 -24717 -23713
rect -23401 -23710 -23377 -23599
rect -23266 -23710 -23238 -23599
rect -23401 -23736 -23238 -23710
rect -24837 -23826 -24717 -23819
rect -24931 -24108 -24859 -24103
rect -27376 -24180 -24926 -24108
rect -24864 -24180 -22986 -24108
rect -24931 -24185 -24859 -24180
rect -24934 -24260 -24778 -24252
rect -27525 -24261 -23124 -24260
rect -27525 -24349 -24907 -24261
rect -24934 -24350 -24907 -24349
rect -24813 -24349 -23124 -24261
rect -24813 -24350 -24778 -24349
rect -24934 -24360 -24778 -24350
rect -23213 -25553 -23124 -24349
rect -23058 -25350 -22986 -24180
rect -22763 -24131 -22674 -23039
rect -22560 -23986 -22488 -22870
rect -16706 -23362 -16596 -23349
rect -16706 -23450 -16693 -23362
rect -16605 -23450 -16596 -23362
rect -16706 -23459 -16596 -23450
rect -18102 -23670 -18004 -23663
rect -18102 -23754 -18095 -23670
rect -18011 -23754 -18004 -23670
rect -18102 -23761 -18004 -23754
rect -22560 -23991 -14032 -23986
rect -22560 -24053 -18037 -23991
rect -17975 -24053 -14032 -23991
rect -22560 -24058 -14032 -24053
rect -22763 -24136 -14178 -24131
rect -22763 -24215 -18058 -24136
rect -17979 -24215 -14178 -24136
rect -22763 -24220 -14178 -24215
rect -16704 -24770 -16598 -24759
rect -16704 -24854 -16693 -24770
rect -16609 -24854 -16598 -24770
rect -16704 -24865 -16598 -24854
rect -18096 -25050 -17998 -25043
rect -18096 -25134 -18089 -25050
rect -18005 -25134 -17998 -25050
rect -18096 -25141 -17998 -25134
rect -23058 -25355 -14392 -25350
rect -23058 -25417 -17951 -25355
rect -17889 -25417 -14392 -25355
rect -23058 -25422 -14392 -25417
rect -23213 -25558 -14534 -25553
rect -23213 -25637 -17971 -25558
rect -17892 -25637 -14534 -25558
rect -23213 -25642 -14534 -25637
rect -14623 -34671 -14534 -25642
rect -14464 -34504 -14392 -25422
rect -14267 -32087 -14178 -24220
rect -14104 -31918 -14032 -24058
rect -13913 -29537 -13824 -22834
rect -13726 -29374 -13654 -22658
rect -13570 -26934 -13506 -21642
rect -13423 -26745 -13362 -21181
rect -13262 -24092 -13191 -20203
rect -13104 -23952 -13041 -19843
rect -12933 -21527 -12844 -18992
rect -12749 -21367 -12679 -18839
rect -12499 -19996 -12373 -19954
rect -12499 -21118 -12471 -19996
rect -12399 -21118 -12373 -19996
rect -11090 -20593 -10999 -20557
rect -11090 -20663 -11084 -20593
rect -11014 -20663 -10999 -20593
rect -11090 -20683 -10999 -20663
rect -12499 -21164 -12373 -21118
rect -12749 -21372 -9935 -21367
rect -12749 -21432 -12604 -21372
rect -12544 -21385 -9935 -21372
rect -9825 -21385 -9755 -16757
rect -8556 -16759 -8477 -16757
rect -7221 -16878 -7122 -16872
rect -8535 -16934 -8408 -16890
rect -8535 -17004 -8505 -16934
rect -8435 -17004 -8408 -16934
rect -5002 -16959 -4936 -16957
rect -2293 -16959 -2227 -16957
rect -7221 -16983 -7122 -16977
rect -5941 -16962 -2195 -16959
rect -8535 -17041 -8408 -17004
rect -5941 -17018 -4997 -16962
rect -4941 -17018 -2288 -16962
rect -2232 -17018 -2195 -16962
rect -5941 -17022 -2195 -17018
rect -8554 -17205 -8475 -17200
rect -8554 -17209 -8549 -17205
rect -12544 -21432 -9755 -21385
rect -12749 -21437 -9755 -21432
rect -10035 -21455 -9755 -21437
rect -9648 -17272 -8549 -17209
rect -12933 -21532 -12486 -21527
rect -12933 -21611 -12623 -21532
rect -12544 -21611 -12486 -21532
rect -12933 -21616 -12486 -21611
rect -12499 -22575 -12373 -22533
rect -12499 -23697 -12471 -22575
rect -12399 -23697 -12373 -22575
rect -11090 -23172 -10999 -23136
rect -11090 -23242 -11084 -23172
rect -11014 -23242 -10999 -23172
rect -11090 -23262 -10999 -23242
rect -12499 -23743 -12373 -23697
rect -12688 -23952 -12602 -23946
rect -9648 -23952 -9585 -17272
rect -8554 -17274 -8549 -17272
rect -8480 -17209 -8475 -17205
rect -5941 -17209 -5878 -17022
rect -5002 -17023 -4936 -17022
rect -2293 -17023 -2227 -17022
rect -8480 -17272 -5875 -17209
rect -8480 -17274 -8475 -17272
rect -8554 -17279 -8475 -17274
rect -7220 -17353 -7121 -17347
rect -8525 -17403 -8408 -17356
rect -8525 -17473 -8502 -17403
rect -8432 -17473 -8408 -17403
rect -7220 -17458 -7121 -17452
rect -5031 -17453 -5025 -17339
rect -4911 -17453 -4905 -17339
rect -4015 -17442 -4009 -17335
rect -3902 -17442 -3896 -17335
rect -2315 -17448 -2309 -17334
rect -2195 -17448 -2189 -17334
rect -1299 -17452 -1293 -17345
rect -1186 -17452 -1180 -17345
rect -8525 -17511 -8408 -17473
rect -8559 -17615 -8480 -17610
rect -8559 -17616 -8554 -17615
rect -13104 -23955 -9585 -23952
rect -13104 -24011 -12673 -23955
rect -12617 -24011 -9585 -23955
rect -13104 -24015 -9585 -24011
rect -9457 -17677 -8554 -17616
rect -12678 -24016 -12612 -24015
rect -12738 -24092 -12574 -24076
rect -13262 -24097 -12523 -24092
rect -13262 -24158 -12681 -24097
rect -12619 -24158 -12523 -24097
rect -13262 -24163 -12523 -24158
rect -12738 -24164 -12574 -24163
rect -12499 -25343 -12373 -25301
rect -12499 -26465 -12471 -25343
rect -12399 -26465 -12373 -25343
rect -11090 -25940 -10999 -25904
rect -11090 -26010 -11084 -25940
rect -11014 -26010 -10999 -25940
rect -11090 -26030 -10999 -26010
rect -12499 -26511 -12373 -26465
rect -12770 -26745 -12612 -26742
rect -9457 -26745 -9396 -17677
rect -8559 -17684 -8554 -17677
rect -8485 -17616 -8480 -17615
rect -8485 -17677 -5420 -17616
rect -8485 -17684 -8480 -17677
rect -8559 -17689 -8480 -17684
rect -5481 -17781 -5420 -17677
rect -4982 -17781 -4916 -17778
rect -2272 -17781 -2206 -17778
rect -5481 -17783 -2196 -17781
rect -7215 -17805 -7116 -17799
rect -8520 -17860 -8409 -17838
rect -8520 -17930 -8500 -17860
rect -8430 -17930 -8409 -17860
rect -5481 -17839 -4977 -17783
rect -4921 -17839 -2267 -17783
rect -2211 -17839 -2196 -17783
rect -5481 -17842 -2196 -17839
rect -4982 -17844 -4916 -17842
rect -2272 -17844 -2206 -17842
rect -7215 -17910 -7116 -17904
rect -8520 -17953 -8409 -17930
rect -8559 -18094 -8480 -18092
rect -13423 -26747 -9396 -26745
rect -13423 -26803 -12741 -26747
rect -12685 -26803 -9396 -26747
rect -13423 -26806 -9396 -26803
rect -9308 -18097 -5472 -18094
rect -9308 -18166 -8554 -18097
rect -8485 -18166 -5472 -18097
rect -12746 -26808 -12680 -26806
rect -12749 -26934 -12683 -26933
rect -13570 -26938 -12532 -26934
rect -13570 -26994 -12744 -26938
rect -12688 -26994 -12532 -26938
rect -13570 -26998 -12532 -26994
rect -12749 -26999 -12683 -26998
rect -12499 -27976 -12373 -27934
rect -12499 -29098 -12471 -27976
rect -12399 -29098 -12373 -27976
rect -11090 -28573 -10999 -28537
rect -11090 -28643 -11084 -28573
rect -11014 -28643 -10999 -28573
rect -11090 -28663 -10999 -28643
rect -12499 -29144 -12373 -29098
rect -9308 -29374 -9236 -18166
rect -8559 -18171 -8480 -18166
rect -7215 -18247 -7116 -18241
rect -8513 -18325 -8413 -18306
rect -8513 -18395 -8498 -18325
rect -8428 -18395 -8413 -18325
rect -7215 -18352 -7116 -18346
rect -8513 -18417 -8413 -18395
rect -13726 -29379 -9236 -29374
rect -13726 -29441 -12719 -29379
rect -12657 -29441 -9236 -29379
rect -13726 -29446 -9236 -29441
rect -9076 -18567 -5782 -18562
rect -9076 -18634 -8554 -18567
rect -13913 -29542 -12094 -29537
rect -13913 -29621 -12723 -29542
rect -12643 -29621 -12094 -29542
rect -13913 -29626 -12094 -29621
rect -12499 -30585 -12373 -30543
rect -12499 -31707 -12471 -30585
rect -12399 -31707 -12373 -30585
rect -11090 -31182 -10999 -31146
rect -11090 -31252 -11084 -31182
rect -11014 -31252 -10999 -31182
rect -11090 -31272 -10999 -31252
rect -12499 -31753 -12373 -31707
rect -12834 -31918 -12670 -31900
rect -9076 -31918 -9004 -18634
rect -8559 -18636 -8554 -18634
rect -8485 -18634 -5782 -18567
rect -8485 -18636 -8480 -18634
rect -8559 -18641 -8480 -18636
rect -7243 -18728 -7096 -18702
rect -8530 -18806 -8391 -18753
rect -8530 -18876 -8494 -18806
rect -8424 -18876 -8391 -18806
rect -7243 -18827 -7221 -18728
rect -7122 -18827 -7096 -18728
rect -7243 -18852 -7096 -18827
rect -8530 -18917 -8391 -18876
rect -14104 -31923 -9004 -31918
rect -14104 -31985 -12753 -31923
rect -12691 -31985 -9004 -31923
rect -14104 -31990 -9004 -31985
rect -8828 -19103 -5924 -19098
rect -8828 -19165 -8579 -19103
rect -8517 -19165 -5924 -19103
rect -8828 -19170 -5924 -19165
rect -14267 -32092 -12460 -32087
rect -14267 -32171 -12787 -32092
rect -12707 -32171 -12460 -32092
rect -14267 -32176 -12460 -32171
rect -12501 -33205 -12375 -33163
rect -12501 -34327 -12473 -33205
rect -12401 -34327 -12375 -33205
rect -11092 -33802 -11001 -33766
rect -11092 -33872 -11086 -33802
rect -11016 -33872 -11001 -33802
rect -11092 -33892 -11001 -33872
rect -12501 -34373 -12375 -34327
rect -8828 -34504 -8756 -19170
rect -5996 -20056 -5924 -19170
rect -5854 -19430 -5782 -18634
rect -5544 -18582 -5472 -18166
rect -5031 -18272 -5025 -18158
rect -4911 -18272 -4905 -18158
rect -4015 -18261 -4009 -18154
rect -3902 -18261 -3896 -18154
rect -2315 -18267 -2309 -18153
rect -2195 -18267 -2189 -18153
rect -1299 -18271 -1293 -18164
rect -1186 -18271 -1180 -18164
rect 5558 -18556 5627 -14109
rect 5998 -14034 6067 -9587
rect 6440 -9514 6509 -9106
rect 6440 -9573 6445 -9514
rect 6504 -9573 6509 -9514
rect 6144 -10330 6264 -10304
rect 6144 -10396 6165 -10330
rect 6231 -10396 6264 -10330
rect 6144 -10417 6264 -10396
rect 6440 -10527 6509 -9573
rect 6579 -10321 6699 -10303
rect 6579 -10387 6605 -10321
rect 6671 -10387 6699 -10321
rect 6579 -10416 6699 -10387
rect 6166 -10596 6509 -10527
rect 6166 -13281 6235 -10596
rect 6299 -10709 6367 -10704
rect 6299 -10767 6304 -10709
rect 6362 -10767 6367 -10709
rect 6299 -10810 6367 -10767
rect 12187 -10710 12431 -10704
rect 6299 -10817 10002 -10810
rect 6299 -10819 9935 -10817
rect 6299 -10875 8998 -10819
rect 9054 -10873 9935 -10819
rect 9991 -10873 10002 -10817
rect 9054 -10875 10002 -10873
rect 6299 -10878 10002 -10875
rect 6299 -13037 6365 -10878
rect 6573 -10880 10002 -10878
rect 10262 -10873 10331 -10868
rect 10262 -10932 10267 -10873
rect 10326 -10932 10331 -10873
rect 6433 -10944 6512 -10939
rect 10262 -10944 10331 -10932
rect 6433 -11013 6438 -10944
rect 6507 -10949 10331 -10944
rect 12187 -10942 12193 -10710
rect 12425 -10942 12431 -10710
rect 12187 -10948 12431 -10942
rect 6507 -11008 8541 -10949
rect 8600 -11008 10331 -10949
rect 6507 -11013 10331 -11008
rect 6433 -11018 6512 -11013
rect 6433 -11091 6507 -11018
rect 6440 -12917 6500 -11091
rect 7156 -11864 11207 -11797
rect 7156 -12052 7222 -11864
rect 7410 -12052 8157 -11864
rect 8345 -12052 9093 -11864
rect 9281 -12051 10024 -11864
rect 10211 -12051 10951 -11864
rect 9281 -12052 10951 -12051
rect 11139 -12052 11207 -11864
rect 7156 -12118 11207 -12052
rect 12414 -12288 12821 -12176
rect 12128 -12292 12821 -12288
rect 12128 -12318 13042 -12292
rect 12128 -12375 13186 -12318
rect 12128 -12504 12228 -12375
rect 12357 -12416 13186 -12375
rect 12357 -12504 12955 -12416
rect 12128 -12545 12955 -12504
rect 13084 -12545 13186 -12416
rect 12128 -12605 13186 -12545
rect 12467 -12764 13186 -12605
rect 12796 -12797 13186 -12764
rect 8398 -12916 8471 -12911
rect 8398 -12917 8405 -12916
rect 6440 -12972 8405 -12917
rect 8461 -12917 8471 -12916
rect 8461 -12948 10324 -12917
rect 8461 -12953 10327 -12948
rect 8461 -12972 10266 -12953
rect 6440 -12977 10266 -12972
rect 10261 -13009 10266 -12977
rect 10322 -13009 10327 -12953
rect 10261 -13014 10327 -13009
rect 6299 -13042 10021 -13037
rect 6299 -13103 9001 -13042
rect 8996 -13104 9001 -13103
rect 9067 -13103 9947 -13042
rect 10003 -13103 10021 -13042
rect 9067 -13104 9072 -13103
rect 8996 -13109 9072 -13104
rect 9942 -13108 10021 -13103
rect 6166 -13350 6506 -13281
rect 5998 -14093 6003 -14034
rect 6062 -14093 6067 -14034
rect 5707 -14877 5827 -14853
rect 5707 -14943 5727 -14877
rect 5793 -14943 5827 -14877
rect 5707 -14966 5827 -14943
rect -5544 -18587 -2222 -18582
rect -5544 -18649 -5001 -18587
rect -4939 -18649 -2289 -18587
rect -2227 -18649 -2222 -18587
rect -5544 -18654 -2222 -18649
rect 5558 -18615 5563 -18556
rect 5622 -18615 5627 -18556
rect -5031 -19091 -5025 -18977
rect -4911 -19091 -4905 -18977
rect -4015 -19080 -4009 -18973
rect -3902 -19080 -3896 -18973
rect -2315 -19086 -2309 -18972
rect -2195 -19086 -2189 -18972
rect -1299 -19090 -1293 -18983
rect -1186 -19090 -1180 -18983
rect -5854 -19435 -2216 -19430
rect -5854 -19497 -5009 -19435
rect -4947 -19497 -2295 -19435
rect -2233 -19497 -2216 -19435
rect -5854 -19502 -2216 -19497
rect -5031 -19910 -5025 -19796
rect -4911 -19910 -4905 -19796
rect -4015 -19899 -4009 -19792
rect -3902 -19899 -3896 -19792
rect -2315 -19905 -2309 -19791
rect -2195 -19905 -2189 -19791
rect -1299 -19909 -1293 -19802
rect -1186 -19909 -1180 -19802
rect -5996 -20061 -2348 -20056
rect -5996 -20123 -5161 -20061
rect -5099 -20123 -2415 -20061
rect -2353 -20123 -2348 -20061
rect -5996 -20128 -2348 -20123
rect -2310 -20418 -2194 -20417
rect -2315 -20532 -2309 -20418
rect -2195 -20532 -2189 -20418
rect -2310 -20533 -2194 -20532
rect -1299 -20542 -1293 -20435
rect -1186 -20542 -1180 -20435
rect -5031 -20729 -5025 -20615
rect -4911 -20729 -4905 -20615
rect -4015 -20718 -4009 -20611
rect -3902 -20718 -3896 -20611
rect 5558 -23100 5627 -18615
rect 5998 -18574 6067 -14093
rect 6437 -14017 6506 -13350
rect 11883 -13412 12147 -13406
rect 11883 -13664 11889 -13412
rect 12141 -13664 12147 -13412
rect 11883 -13670 12147 -13664
rect 6437 -14076 6442 -14017
rect 6501 -14076 6506 -14017
rect 6144 -14858 6264 -14832
rect 6144 -14924 6165 -14858
rect 6231 -14924 6264 -14858
rect 6144 -14945 6264 -14924
rect 6437 -15089 6506 -14076
rect 6579 -14849 6699 -14831
rect 6579 -14915 6605 -14849
rect 6671 -14915 6699 -14849
rect 6579 -14944 6699 -14915
rect 6155 -15158 6506 -15089
rect 6155 -17862 6224 -15158
rect 6299 -15237 6367 -15232
rect 6299 -15295 6304 -15237
rect 6362 -15295 6367 -15237
rect 6299 -15338 6367 -15295
rect 12187 -15238 12431 -15232
rect 6299 -15345 10002 -15338
rect 6299 -15347 9935 -15345
rect 6299 -15403 8998 -15347
rect 9054 -15401 9935 -15347
rect 9991 -15401 10002 -15345
rect 9054 -15403 10002 -15401
rect 6299 -15406 10002 -15403
rect 6299 -17565 6365 -15406
rect 6573 -15408 10002 -15406
rect 10262 -15401 10331 -15396
rect 10262 -15460 10267 -15401
rect 10326 -15460 10331 -15401
rect 6433 -15472 6512 -15467
rect 10262 -15472 10331 -15460
rect 6433 -15541 6438 -15472
rect 6507 -15477 10331 -15472
rect 12187 -15470 12193 -15238
rect 12425 -15470 12431 -15238
rect 12187 -15476 12431 -15470
rect 6507 -15536 8541 -15477
rect 8600 -15536 10331 -15477
rect 6507 -15541 10331 -15536
rect 6433 -15546 6512 -15541
rect 6433 -15619 6507 -15546
rect 6440 -17445 6500 -15619
rect 7156 -16392 11207 -16325
rect 7156 -16580 7222 -16392
rect 7410 -16580 8157 -16392
rect 8345 -16580 9093 -16392
rect 9281 -16579 10024 -16392
rect 10211 -16579 10951 -16392
rect 9281 -16580 10951 -16579
rect 11139 -16580 11207 -16392
rect 7156 -16646 11207 -16580
rect 12414 -16816 12821 -16704
rect 12128 -16820 12821 -16816
rect 16250 -16732 16588 -16694
rect 12128 -16846 13042 -16820
rect 12128 -16903 13186 -16846
rect 12128 -17032 12228 -16903
rect 12357 -16944 13186 -16903
rect 12357 -17032 12955 -16944
rect 12128 -17073 12955 -17032
rect 13084 -17073 13186 -16944
rect 16250 -17000 16280 -16732
rect 16548 -17000 16588 -16732
rect 16250 -17028 16588 -17000
rect 12128 -17133 13186 -17073
rect 12467 -17292 13186 -17133
rect 12796 -17325 13186 -17292
rect 8398 -17444 8471 -17439
rect 8398 -17445 8405 -17444
rect 6440 -17500 8405 -17445
rect 8461 -17445 8471 -17444
rect 8461 -17476 10324 -17445
rect 8461 -17481 10327 -17476
rect 8461 -17500 10266 -17481
rect 6440 -17505 10266 -17500
rect 10261 -17537 10266 -17505
rect 10322 -17537 10327 -17481
rect 10261 -17542 10327 -17537
rect 6299 -17570 10021 -17565
rect 6299 -17631 9001 -17570
rect 8996 -17632 9001 -17631
rect 9067 -17631 9947 -17570
rect 10003 -17631 10021 -17570
rect 9067 -17632 9072 -17631
rect 8996 -17637 9072 -17632
rect 9942 -17636 10021 -17631
rect 6155 -17931 6504 -17862
rect 5998 -18633 6003 -18574
rect 6062 -18633 6067 -18574
rect 5707 -19405 5827 -19381
rect 5707 -19471 5727 -19405
rect 5793 -19471 5827 -19405
rect 5707 -19494 5827 -19471
rect 5558 -23159 5563 -23100
rect 5622 -23159 5627 -23100
rect 5558 -27640 5627 -23159
rect 5998 -23090 6067 -18633
rect 6435 -18567 6504 -17931
rect 11883 -17940 12147 -17934
rect 11883 -18192 11889 -17940
rect 12141 -18192 12147 -17940
rect 17515 -18016 17672 -18008
rect 17515 -18159 17521 -18016
rect 17664 -18159 17672 -18016
rect 17515 -18165 17672 -18159
rect 11883 -18198 12147 -18192
rect 6435 -18626 6440 -18567
rect 6499 -18626 6504 -18567
rect 6144 -19386 6264 -19360
rect 6144 -19452 6165 -19386
rect 6231 -19452 6264 -19386
rect 6144 -19473 6264 -19452
rect 6435 -19597 6504 -18626
rect 15538 -18509 15708 -18501
rect 15538 -18663 15546 -18509
rect 15700 -18663 15708 -18509
rect 15538 -18671 15708 -18663
rect 17951 -18864 18077 -18845
rect 17951 -18945 17972 -18864
rect 18053 -18945 18077 -18864
rect 17951 -18965 18077 -18945
rect 6579 -19377 6699 -19359
rect 6579 -19443 6605 -19377
rect 6671 -19443 6699 -19377
rect 6579 -19472 6699 -19443
rect 6166 -19666 6504 -19597
rect 6166 -22390 6235 -19666
rect 6299 -19765 6367 -19760
rect 6299 -19823 6304 -19765
rect 6362 -19823 6367 -19765
rect 6299 -19866 6367 -19823
rect 12187 -19766 12431 -19760
rect 6299 -19873 10002 -19866
rect 6299 -19875 9935 -19873
rect 6299 -19931 8998 -19875
rect 9054 -19929 9935 -19875
rect 9991 -19929 10002 -19873
rect 9054 -19931 10002 -19929
rect 6299 -19934 10002 -19931
rect 6299 -22093 6365 -19934
rect 6573 -19936 10002 -19934
rect 10262 -19929 10331 -19924
rect 10262 -19988 10267 -19929
rect 10326 -19988 10331 -19929
rect 6433 -20000 6512 -19995
rect 10262 -20000 10331 -19988
rect 6433 -20069 6438 -20000
rect 6507 -20005 10331 -20000
rect 12187 -19998 12193 -19766
rect 12425 -19998 12431 -19766
rect 12187 -20004 12431 -19998
rect 6507 -20064 8541 -20005
rect 8600 -20064 10331 -20005
rect 6507 -20069 10331 -20064
rect 6433 -20074 6512 -20069
rect 6433 -20147 6507 -20074
rect 6440 -21973 6500 -20147
rect 16196 -20172 16516 -20147
rect 16196 -20441 16226 -20172
rect 16485 -20441 16516 -20172
rect 16196 -20467 16516 -20441
rect 7156 -20920 11207 -20853
rect 7156 -21108 7222 -20920
rect 7410 -21108 8157 -20920
rect 8345 -21108 9093 -20920
rect 9281 -21107 10024 -20920
rect 10211 -21107 10951 -20920
rect 9281 -21108 10951 -21107
rect 11139 -21108 11207 -20920
rect 7156 -21174 11207 -21108
rect 12414 -21344 12821 -21232
rect 12128 -21348 12821 -21344
rect 12128 -21374 13042 -21348
rect 12128 -21431 13186 -21374
rect 12128 -21560 12228 -21431
rect 12357 -21472 13186 -21431
rect 12357 -21560 12955 -21472
rect 12128 -21601 12955 -21560
rect 13084 -21601 13186 -21472
rect 12128 -21661 13186 -21601
rect 12467 -21820 13186 -21661
rect 12796 -21853 13186 -21820
rect 8398 -21972 8471 -21967
rect 8398 -21973 8405 -21972
rect 6440 -22028 8405 -21973
rect 8461 -21973 8471 -21972
rect 8461 -22004 10324 -21973
rect 8461 -22009 10327 -22004
rect 8461 -22028 10266 -22009
rect 6440 -22033 10266 -22028
rect 10261 -22065 10266 -22033
rect 10322 -22065 10327 -22009
rect 10261 -22070 10327 -22065
rect 6299 -22098 10021 -22093
rect 6299 -22159 9001 -22098
rect 8996 -22160 9001 -22159
rect 9067 -22159 9947 -22098
rect 10003 -22159 10021 -22098
rect 9067 -22160 9072 -22159
rect 8996 -22165 9072 -22160
rect 9942 -22164 10021 -22159
rect 6166 -22459 6512 -22390
rect 5998 -23149 6003 -23090
rect 6062 -23149 6067 -23090
rect 5707 -23933 5827 -23909
rect 5707 -23999 5727 -23933
rect 5793 -23999 5827 -23933
rect 5707 -24022 5827 -23999
rect 5558 -27699 5563 -27640
rect 5622 -27699 5627 -27640
rect 5558 -32149 5627 -27699
rect 5998 -27635 6067 -23149
rect 6443 -23065 6512 -22459
rect 11883 -22468 12147 -22462
rect 11883 -22720 11889 -22468
rect 12141 -22720 12147 -22468
rect 11883 -22726 12147 -22720
rect 6443 -23124 6448 -23065
rect 6507 -23124 6512 -23065
rect 6144 -23914 6264 -23888
rect 6144 -23980 6165 -23914
rect 6231 -23980 6264 -23914
rect 6144 -24001 6264 -23980
rect 6443 -24122 6512 -23124
rect 6579 -23905 6699 -23887
rect 6579 -23971 6605 -23905
rect 6671 -23971 6699 -23905
rect 6579 -24000 6699 -23971
rect 6155 -24191 6512 -24122
rect 6155 -26902 6224 -24191
rect 6299 -24293 6367 -24288
rect 6299 -24351 6304 -24293
rect 6362 -24351 6367 -24293
rect 6299 -24394 6367 -24351
rect 12187 -24294 12431 -24288
rect 6299 -24401 10002 -24394
rect 6299 -24403 9935 -24401
rect 6299 -24459 8998 -24403
rect 9054 -24457 9935 -24403
rect 9991 -24457 10002 -24401
rect 9054 -24459 10002 -24457
rect 6299 -24462 10002 -24459
rect 6299 -26621 6365 -24462
rect 6573 -24464 10002 -24462
rect 10262 -24457 10331 -24452
rect 10262 -24516 10267 -24457
rect 10326 -24516 10331 -24457
rect 6433 -24528 6512 -24523
rect 10262 -24528 10331 -24516
rect 6433 -24597 6438 -24528
rect 6507 -24533 10331 -24528
rect 12187 -24526 12193 -24294
rect 12425 -24526 12431 -24294
rect 12187 -24532 12431 -24526
rect 6507 -24592 8541 -24533
rect 8600 -24592 10331 -24533
rect 6507 -24597 10331 -24592
rect 6433 -24602 6512 -24597
rect 6433 -24675 6507 -24602
rect 6440 -26501 6500 -24675
rect 7156 -25448 11207 -25381
rect 7156 -25636 7222 -25448
rect 7410 -25636 8157 -25448
rect 8345 -25636 9093 -25448
rect 9281 -25635 10024 -25448
rect 10211 -25635 10951 -25448
rect 9281 -25636 10951 -25635
rect 11139 -25636 11207 -25448
rect 7156 -25702 11207 -25636
rect 12414 -25872 12821 -25760
rect 12128 -25876 12821 -25872
rect 12128 -25902 13042 -25876
rect 12128 -25959 13186 -25902
rect 12128 -26088 12228 -25959
rect 12357 -26000 13186 -25959
rect 12357 -26088 12955 -26000
rect 12128 -26129 12955 -26088
rect 13084 -26129 13186 -26000
rect 12128 -26189 13186 -26129
rect 12467 -26348 13186 -26189
rect 12796 -26381 13186 -26348
rect 8398 -26500 8471 -26495
rect 8398 -26501 8405 -26500
rect 6440 -26556 8405 -26501
rect 8461 -26501 8471 -26500
rect 8461 -26532 10324 -26501
rect 8461 -26537 10327 -26532
rect 8461 -26556 10266 -26537
rect 6440 -26561 10266 -26556
rect 10261 -26593 10266 -26561
rect 10322 -26593 10327 -26537
rect 10261 -26598 10327 -26593
rect 6299 -26626 10021 -26621
rect 6299 -26687 9001 -26626
rect 8996 -26688 9001 -26687
rect 9067 -26687 9947 -26626
rect 10003 -26687 10021 -26626
rect 9067 -26688 9072 -26687
rect 8996 -26693 9072 -26688
rect 9942 -26692 10021 -26687
rect 6155 -26971 6502 -26902
rect 5998 -27694 6003 -27635
rect 6062 -27694 6067 -27635
rect 5707 -28461 5827 -28437
rect 5707 -28527 5727 -28461
rect 5793 -28527 5827 -28461
rect 5707 -28550 5827 -28527
rect 5558 -32208 5563 -32149
rect 5622 -32208 5627 -32149
rect 5558 -32279 5627 -32208
rect 5998 -32164 6067 -27694
rect 6433 -27581 6502 -26971
rect 11883 -26996 12147 -26990
rect 11883 -27248 11889 -26996
rect 12141 -27248 12147 -26996
rect 11883 -27254 12147 -27248
rect 6433 -27640 6438 -27581
rect 6497 -27640 6502 -27581
rect 6144 -28442 6264 -28416
rect 6144 -28508 6165 -28442
rect 6231 -28508 6264 -28442
rect 6144 -28529 6264 -28508
rect 6433 -28684 6502 -27640
rect 6579 -28433 6699 -28415
rect 6579 -28499 6605 -28433
rect 6671 -28499 6699 -28433
rect 6579 -28528 6699 -28499
rect 6145 -28753 6502 -28684
rect 6145 -31454 6214 -28753
rect 6299 -28821 6367 -28816
rect 6299 -28879 6304 -28821
rect 6362 -28879 6367 -28821
rect 6299 -28922 6367 -28879
rect 12187 -28822 12431 -28816
rect 6299 -28929 10002 -28922
rect 6299 -28931 9935 -28929
rect 6299 -28987 8998 -28931
rect 9054 -28985 9935 -28931
rect 9991 -28985 10002 -28929
rect 9054 -28987 10002 -28985
rect 6299 -28990 10002 -28987
rect 6299 -31149 6365 -28990
rect 6573 -28992 10002 -28990
rect 10262 -28985 10331 -28980
rect 10262 -29044 10267 -28985
rect 10326 -29044 10331 -28985
rect 6433 -29056 6512 -29051
rect 10262 -29056 10331 -29044
rect 6433 -29125 6438 -29056
rect 6507 -29061 10331 -29056
rect 12187 -29054 12193 -28822
rect 12425 -29054 12431 -28822
rect 12187 -29060 12431 -29054
rect 6507 -29120 8541 -29061
rect 8600 -29120 10331 -29061
rect 6507 -29125 10331 -29120
rect 6433 -29130 6512 -29125
rect 6433 -29203 6507 -29130
rect 6440 -31029 6500 -29203
rect 7156 -29976 11207 -29909
rect 7156 -30164 7222 -29976
rect 7410 -30164 8157 -29976
rect 8345 -30164 9093 -29976
rect 9281 -30163 10024 -29976
rect 10211 -30163 10951 -29976
rect 9281 -30164 10951 -30163
rect 11139 -30164 11207 -29976
rect 7156 -30230 11207 -30164
rect 12414 -30400 12821 -30288
rect 12128 -30404 12821 -30400
rect 12128 -30430 13042 -30404
rect 12128 -30487 13186 -30430
rect 12128 -30616 12228 -30487
rect 12357 -30528 13186 -30487
rect 12357 -30616 12955 -30528
rect 12128 -30657 12955 -30616
rect 13084 -30657 13186 -30528
rect 12128 -30717 13186 -30657
rect 12467 -30876 13186 -30717
rect 12796 -30909 13186 -30876
rect 8398 -31028 8471 -31023
rect 8398 -31029 8405 -31028
rect 6440 -31084 8405 -31029
rect 8461 -31029 8471 -31028
rect 8461 -31060 10324 -31029
rect 8461 -31065 10327 -31060
rect 8461 -31084 10266 -31065
rect 6440 -31089 10266 -31084
rect 10261 -31121 10266 -31089
rect 10322 -31121 10327 -31065
rect 10261 -31126 10327 -31121
rect 6299 -31154 10021 -31149
rect 6299 -31215 9001 -31154
rect 8996 -31216 9001 -31215
rect 9067 -31215 9947 -31154
rect 10003 -31215 10021 -31154
rect 9067 -31216 9072 -31215
rect 8996 -31221 9072 -31216
rect 9942 -31220 10021 -31215
rect 6145 -31523 6507 -31454
rect 6438 -32126 6507 -31523
rect 11883 -31524 12147 -31518
rect 11883 -31776 11889 -31524
rect 12141 -31776 12147 -31524
rect 11883 -31782 12147 -31776
rect 5998 -32223 6003 -32164
rect 6062 -32223 6067 -32164
rect 6433 -32131 6512 -32126
rect 6433 -32201 6438 -32131
rect 6507 -32201 6512 -32131
rect 6433 -32206 6512 -32201
rect 5998 -32228 6067 -32223
rect 5707 -32989 5827 -32965
rect 5707 -33055 5727 -32989
rect 5793 -33055 5827 -32989
rect 5707 -33078 5827 -33055
rect 6144 -32970 6264 -32944
rect 6144 -33036 6165 -32970
rect 6231 -33036 6264 -32970
rect 6144 -33057 6264 -33036
rect 6579 -32961 6699 -32943
rect 6579 -33027 6605 -32961
rect 6671 -33027 6699 -32961
rect 6579 -33056 6699 -33027
rect -14464 -34509 -8756 -34504
rect -14464 -34571 -12577 -34509
rect -12515 -34571 -8756 -34509
rect -14464 -34576 -8756 -34571
rect 6299 -33349 6367 -33344
rect 6299 -33407 6304 -33349
rect 6362 -33407 6367 -33349
rect 6299 -33450 6367 -33407
rect 12187 -33350 12431 -33344
rect 6299 -33457 10002 -33450
rect 6299 -33459 9935 -33457
rect 6299 -33515 8998 -33459
rect 9054 -33513 9935 -33459
rect 9991 -33513 10002 -33457
rect 9054 -33515 10002 -33513
rect 6299 -33518 10002 -33515
rect -14623 -34676 -12520 -34671
rect -14623 -34755 -12721 -34676
rect -12642 -34755 -12520 -34676
rect -14623 -34760 -12520 -34755
rect 6299 -35677 6365 -33518
rect 6573 -33520 10002 -33518
rect 10262 -33513 10331 -33508
rect 10262 -33572 10267 -33513
rect 10326 -33572 10331 -33513
rect 6433 -33584 6512 -33579
rect 10262 -33584 10331 -33572
rect 6433 -33653 6438 -33584
rect 6507 -33589 10331 -33584
rect 12187 -33582 12193 -33350
rect 12425 -33582 12431 -33350
rect 12187 -33588 12431 -33582
rect 6507 -33648 8541 -33589
rect 8600 -33648 10331 -33589
rect 6507 -33653 10331 -33648
rect 6433 -33658 6512 -33653
rect 6433 -33731 6507 -33658
rect 6440 -35557 6500 -33731
rect 7156 -34504 11207 -34437
rect 7156 -34692 7222 -34504
rect 7410 -34692 8157 -34504
rect 8345 -34692 9093 -34504
rect 9281 -34691 10024 -34504
rect 10211 -34691 10951 -34504
rect 9281 -34692 10951 -34691
rect 11139 -34692 11207 -34504
rect 7156 -34758 11207 -34692
rect 12414 -34928 12821 -34816
rect 12128 -34932 12821 -34928
rect 12128 -34958 13042 -34932
rect 12128 -35015 13186 -34958
rect 12128 -35144 12228 -35015
rect 12357 -35056 13186 -35015
rect 12357 -35144 12955 -35056
rect 12128 -35185 12955 -35144
rect 13084 -35185 13186 -35056
rect 12128 -35245 13186 -35185
rect 12467 -35404 13186 -35245
rect 12796 -35437 13186 -35404
rect 8398 -35556 8471 -35551
rect 8398 -35557 8405 -35556
rect 6440 -35612 8405 -35557
rect 8461 -35557 8471 -35556
rect 8461 -35588 10324 -35557
rect 8461 -35593 10327 -35588
rect 8461 -35612 10266 -35593
rect 6440 -35617 10266 -35612
rect 10261 -35649 10266 -35617
rect 10322 -35649 10327 -35593
rect 10261 -35654 10327 -35649
rect 6299 -35682 10021 -35677
rect 6299 -35743 9001 -35682
rect 8996 -35744 9001 -35743
rect 9067 -35743 9947 -35682
rect 10003 -35743 10021 -35682
rect 9067 -35744 9072 -35743
rect 8996 -35749 9072 -35744
rect 9942 -35748 10021 -35743
rect 11883 -36052 12147 -36046
rect 11883 -36304 11889 -36052
rect 12141 -36304 12147 -36052
rect 12538 -36057 12544 -35950
rect 12651 -36057 12657 -35950
rect 13547 -36068 13553 -35954
rect 13667 -36068 13673 -35954
rect 11883 -36310 12147 -36304
<< via3 >>
rect 1841 6169 2963 6241
rect 3447 6169 4569 6241
rect 5151 6167 6273 6239
rect 2296 4849 2366 4854
rect 2296 4789 2301 4849
rect 2301 4789 2361 4849
rect 2361 4789 2366 4849
rect 2296 4784 2366 4789
rect 3902 4849 3972 4854
rect 3902 4789 3907 4849
rect 3907 4789 3967 4849
rect 3967 4789 3972 4849
rect 3902 4784 3972 4789
rect 5606 4847 5676 4852
rect 5606 4787 5611 4847
rect 5611 4787 5671 4847
rect 5671 4787 5676 4847
rect 5606 4782 5676 4787
rect -24000 4445 -22878 4517
rect -20709 4445 -19587 4517
rect -17418 4445 -16296 4517
rect -14127 4445 -13005 4517
rect -10836 4445 -9714 4517
rect -7546 4445 -6424 4517
rect -4255 4445 -3133 4517
rect -964 4445 158 4517
rect -23403 3125 -23333 3130
rect -23403 3065 -23398 3125
rect -23398 3065 -23338 3125
rect -23338 3065 -23333 3125
rect -23403 3060 -23333 3065
rect -20112 3125 -20042 3130
rect -20112 3065 -20107 3125
rect -20107 3065 -20047 3125
rect -20047 3065 -20042 3125
rect -20112 3060 -20042 3065
rect -16821 3125 -16751 3130
rect -16821 3065 -16816 3125
rect -16816 3065 -16756 3125
rect -16756 3065 -16751 3125
rect -16821 3060 -16751 3065
rect -13530 3125 -13460 3130
rect -13530 3065 -13525 3125
rect -13525 3065 -13465 3125
rect -13465 3065 -13460 3125
rect -13530 3060 -13460 3065
rect -10239 3125 -10169 3130
rect -10239 3065 -10234 3125
rect -10234 3065 -10174 3125
rect -10174 3065 -10169 3125
rect -10239 3060 -10169 3065
rect -6949 3125 -6879 3130
rect -6949 3065 -6944 3125
rect -6944 3065 -6884 3125
rect -6884 3065 -6879 3125
rect -6949 3060 -6879 3065
rect -3658 3125 -3588 3130
rect -3658 3065 -3653 3125
rect -3653 3065 -3593 3125
rect -3593 3065 -3588 3125
rect -3658 3060 -3588 3065
rect -367 3125 -297 3130
rect -367 3065 -362 3125
rect -362 3065 -302 3125
rect -302 3065 -297 3125
rect -367 3060 -297 3065
rect -24670 2661 -23548 2733
rect -23111 2661 -21989 2733
rect -21379 2661 -20257 2733
rect -19820 2661 -18698 2733
rect -18088 2661 -16966 2733
rect -16529 2661 -15407 2733
rect -14797 2661 -13675 2733
rect -13238 2661 -12116 2733
rect -11506 2661 -10384 2733
rect -9947 2661 -8825 2733
rect -8216 2661 -7094 2733
rect -6657 2661 -5535 2733
rect -4925 2661 -3803 2733
rect -3366 2661 -2244 2733
rect -1634 2661 -512 2733
rect -75 2661 1047 2733
rect -24215 1341 -24145 1346
rect -24215 1281 -24210 1341
rect -24210 1281 -24150 1341
rect -24150 1281 -24145 1341
rect -24215 1276 -24145 1281
rect -22656 1341 -22586 1346
rect -22656 1281 -22651 1341
rect -22651 1281 -22591 1341
rect -22591 1281 -22586 1341
rect -22656 1276 -22586 1281
rect -20924 1341 -20854 1346
rect -20924 1281 -20919 1341
rect -20919 1281 -20859 1341
rect -20859 1281 -20854 1341
rect -20924 1276 -20854 1281
rect -19365 1341 -19295 1346
rect -19365 1281 -19360 1341
rect -19360 1281 -19300 1341
rect -19300 1281 -19295 1341
rect -19365 1276 -19295 1281
rect -17633 1341 -17563 1346
rect -17633 1281 -17628 1341
rect -17628 1281 -17568 1341
rect -17568 1281 -17563 1341
rect -17633 1276 -17563 1281
rect -16074 1341 -16004 1346
rect -16074 1281 -16069 1341
rect -16069 1281 -16009 1341
rect -16009 1281 -16004 1341
rect -16074 1276 -16004 1281
rect -14342 1341 -14272 1346
rect -14342 1281 -14337 1341
rect -14337 1281 -14277 1341
rect -14277 1281 -14272 1341
rect -14342 1276 -14272 1281
rect -12783 1341 -12713 1346
rect -12783 1281 -12778 1341
rect -12778 1281 -12718 1341
rect -12718 1281 -12713 1341
rect -12783 1276 -12713 1281
rect -11051 1341 -10981 1346
rect -11051 1281 -11046 1341
rect -11046 1281 -10986 1341
rect -10986 1281 -10981 1341
rect -11051 1276 -10981 1281
rect -9492 1341 -9422 1346
rect -9492 1281 -9487 1341
rect -9487 1281 -9427 1341
rect -9427 1281 -9422 1341
rect -9492 1276 -9422 1281
rect -7761 1341 -7691 1346
rect -7761 1281 -7756 1341
rect -7756 1281 -7696 1341
rect -7696 1281 -7691 1341
rect -7761 1276 -7691 1281
rect -6202 1341 -6132 1346
rect -6202 1281 -6197 1341
rect -6197 1281 -6137 1341
rect -6137 1281 -6132 1341
rect -6202 1276 -6132 1281
rect -4470 1341 -4400 1346
rect -4470 1281 -4465 1341
rect -4465 1281 -4405 1341
rect -4405 1281 -4400 1341
rect -4470 1276 -4400 1281
rect -2911 1341 -2841 1346
rect -2911 1281 -2906 1341
rect -2906 1281 -2846 1341
rect -2846 1281 -2841 1341
rect -2911 1276 -2841 1281
rect -1179 1341 -1109 1346
rect -1179 1281 -1174 1341
rect -1174 1281 -1114 1341
rect -1114 1281 -1109 1341
rect -1179 1276 -1109 1281
rect 380 1341 450 1346
rect 380 1281 385 1341
rect 385 1281 445 1341
rect 445 1281 450 1341
rect 380 1276 450 1281
rect -24412 929 -24156 1001
rect -23123 929 -22867 1001
rect -22406 929 -22150 1001
rect -21121 929 -20865 1001
rect -19832 929 -19576 1001
rect -19115 929 -18859 1001
rect -17830 929 -17574 1001
rect -16541 929 -16285 1001
rect -15824 929 -15568 1001
rect -14539 929 -14283 1001
rect -13250 929 -12994 1001
rect -12533 929 -12277 1001
rect -11248 929 -10992 1001
rect -9959 929 -9703 1001
rect -9242 929 -8986 1001
rect -7958 929 -7702 1001
rect -6669 929 -6413 1001
rect -5952 929 -5696 1001
rect -4667 929 -4411 1001
rect -3378 929 -3122 1001
rect -2661 929 -2405 1001
rect -1376 929 -1120 1001
rect -87 929 169 1001
rect 630 929 886 1001
rect -24336 259 -24001 267
rect -24336 203 -24001 259
rect -23105 250 -23033 255
rect -23105 188 -23100 250
rect -23100 188 -23038 250
rect -23038 188 -23033 250
rect -23105 183 -23033 188
rect -22240 225 -22174 230
rect -22240 169 -22235 225
rect -22235 169 -22179 225
rect -22179 169 -22174 225
rect -22240 164 -22174 169
rect -21045 259 -20710 267
rect -21045 203 -20710 259
rect -19814 250 -19742 255
rect -19814 188 -19809 250
rect -19809 188 -19747 250
rect -19747 188 -19742 250
rect -19814 183 -19742 188
rect -18949 225 -18883 230
rect -18949 169 -18944 225
rect -18944 169 -18888 225
rect -18888 169 -18883 225
rect -18949 164 -18883 169
rect -17754 259 -17419 267
rect -17754 203 -17419 259
rect -16523 250 -16451 255
rect -16523 188 -16518 250
rect -16518 188 -16456 250
rect -16456 188 -16451 250
rect -16523 183 -16451 188
rect -15658 225 -15592 230
rect -15658 169 -15653 225
rect -15653 169 -15597 225
rect -15597 169 -15592 225
rect -15658 164 -15592 169
rect -14463 259 -14128 267
rect -14463 203 -14128 259
rect -13232 250 -13160 255
rect -13232 188 -13227 250
rect -13227 188 -13165 250
rect -13165 188 -13160 250
rect -13232 183 -13160 188
rect -12367 225 -12301 230
rect -12367 169 -12362 225
rect -12362 169 -12306 225
rect -12306 169 -12301 225
rect -12367 164 -12301 169
rect -11172 259 -10837 267
rect -11172 203 -10837 259
rect -9941 250 -9869 255
rect -9941 188 -9936 250
rect -9936 188 -9874 250
rect -9874 188 -9869 250
rect -9941 183 -9869 188
rect -9076 225 -9010 230
rect -9076 169 -9071 225
rect -9071 169 -9015 225
rect -9015 169 -9010 225
rect -9076 164 -9010 169
rect -7882 259 -7547 267
rect -7882 203 -7547 259
rect -6651 250 -6579 255
rect -6651 188 -6646 250
rect -6646 188 -6584 250
rect -6584 188 -6579 250
rect -6651 183 -6579 188
rect -5786 225 -5720 230
rect -5786 169 -5781 225
rect -5781 169 -5725 225
rect -5725 169 -5720 225
rect -5786 164 -5720 169
rect -4591 259 -4256 267
rect -4591 203 -4256 259
rect -3360 250 -3288 255
rect -3360 188 -3355 250
rect -3355 188 -3293 250
rect -3293 188 -3288 250
rect -3360 183 -3288 188
rect -2495 225 -2429 230
rect -2495 169 -2490 225
rect -2490 169 -2434 225
rect -2434 169 -2429 225
rect -2495 164 -2429 169
rect -1300 259 -965 267
rect -1300 203 -965 259
rect -69 250 3 255
rect -69 188 -64 250
rect -64 188 -2 250
rect -2 188 3 250
rect -69 183 3 188
rect 796 225 862 230
rect 796 169 801 225
rect 801 169 857 225
rect 857 169 862 225
rect 796 164 862 169
rect 5727 3230 5793 3235
rect 5727 3174 5732 3230
rect 5732 3174 5788 3230
rect 5788 3174 5793 3230
rect 5727 3169 5793 3174
rect -23605 -2304 -23436 -2225
rect -24410 -2467 -23856 -2327
rect -21585 -2304 -21416 -2225
rect -22373 -2467 -21819 -2327
rect -19844 -2304 -19675 -2225
rect -20643 -2467 -20089 -2327
rect -24184 -3057 -23844 -2983
rect -23601 -2974 -23452 -2878
rect -22147 -3057 -21807 -2983
rect -21581 -2974 -21432 -2878
rect -23561 -4116 -23392 -4037
rect -24359 -4279 -23805 -4139
rect -24133 -4869 -23793 -4795
rect -23557 -4786 -23408 -4690
rect -23563 -5408 -23394 -5329
rect -24359 -5571 -23805 -5431
rect -24133 -6161 -23793 -6087
rect -23559 -6078 -23410 -5982
rect -23562 -7381 -23393 -7302
rect -24359 -7544 -23805 -7404
rect -24133 -8134 -23793 -8060
rect -23558 -8051 -23409 -7955
rect -23560 -8673 -23391 -8594
rect -24359 -8836 -23805 -8696
rect -24133 -9426 -23793 -9352
rect -23556 -9343 -23407 -9247
rect -23560 -10645 -23391 -10566
rect -24359 -10808 -23805 -10668
rect -20417 -3057 -20077 -2983
rect -19840 -2974 -19691 -2878
rect -18065 -2304 -17896 -2225
rect -18883 -2467 -18329 -2327
rect -18657 -3057 -18317 -2983
rect -18061 -2974 -17912 -2878
rect -21823 -4116 -21654 -4037
rect -22623 -4279 -22069 -4139
rect -22397 -4869 -22057 -4795
rect -21819 -4786 -21670 -4690
rect -21829 -5408 -21660 -5329
rect -22623 -5571 -22069 -5431
rect -22397 -6161 -22057 -6087
rect -21825 -6078 -21676 -5982
rect -20603 -3899 -19481 -3827
rect -19044 -3899 -17922 -3827
rect -17312 -3899 -16190 -3827
rect -15753 -3899 -14631 -3827
rect -14021 -3899 -12899 -3827
rect -12462 -3899 -11340 -3827
rect -10730 -3899 -9608 -3827
rect -9171 -3899 -8049 -3827
rect 6165 3249 6231 3254
rect 6165 3193 6170 3249
rect 6170 3193 6226 3249
rect 6226 3193 6231 3249
rect 6165 3188 6231 3193
rect 6605 3258 6671 3263
rect 6605 3202 6610 3258
rect 6610 3202 6666 3258
rect 6666 3202 6671 3258
rect 6605 3197 6671 3202
rect 12193 2869 12425 2874
rect 12193 2647 12198 2869
rect 12198 2647 12420 2869
rect 12420 2647 12425 2869
rect 12193 2642 12425 2647
rect 7222 1715 7410 1720
rect 7222 1537 7227 1715
rect 7227 1537 7405 1715
rect 7405 1537 7410 1715
rect 7222 1532 7410 1537
rect 8157 1715 8345 1720
rect 8157 1537 8162 1715
rect 8162 1537 8340 1715
rect 8340 1537 8345 1715
rect 8157 1532 8345 1537
rect 9093 1715 9281 1720
rect 9093 1537 9098 1715
rect 9098 1537 9276 1715
rect 9276 1537 9281 1715
rect 9093 1532 9281 1537
rect 10024 1715 10211 1720
rect 10024 1538 10029 1715
rect 10029 1538 10206 1715
rect 10206 1538 10211 1715
rect 10024 1533 10211 1538
rect 10951 1715 11139 1720
rect 10951 1537 10956 1715
rect 10956 1537 11134 1715
rect 11134 1537 11139 1715
rect 10951 1532 11139 1537
rect 12228 1204 12357 1209
rect 12228 1085 12233 1204
rect 12233 1085 12352 1204
rect 12352 1085 12357 1204
rect 12228 1080 12357 1085
rect 12955 1163 13084 1168
rect 12955 1044 12960 1163
rect 12960 1044 13079 1163
rect 13079 1044 13084 1163
rect 12955 1039 13084 1044
rect 5727 -1298 5793 -1293
rect 5727 -1354 5732 -1298
rect 5732 -1354 5788 -1298
rect 5788 -1354 5793 -1298
rect 5727 -1359 5793 -1354
rect -20148 -5219 -20078 -5214
rect -20148 -5279 -20143 -5219
rect -20143 -5279 -20083 -5219
rect -20083 -5279 -20078 -5219
rect -20148 -5284 -20078 -5279
rect -18589 -5219 -18519 -5214
rect -18589 -5279 -18584 -5219
rect -18584 -5279 -18524 -5219
rect -18524 -5279 -18519 -5219
rect -18589 -5284 -18519 -5279
rect -16857 -5219 -16787 -5214
rect -16857 -5279 -16852 -5219
rect -16852 -5279 -16792 -5219
rect -16792 -5279 -16787 -5219
rect -16857 -5284 -16787 -5279
rect -15298 -5219 -15228 -5214
rect -15298 -5279 -15293 -5219
rect -15293 -5279 -15233 -5219
rect -15233 -5279 -15228 -5219
rect -15298 -5284 -15228 -5279
rect -13566 -5219 -13496 -5214
rect -13566 -5279 -13561 -5219
rect -13561 -5279 -13501 -5219
rect -13501 -5279 -13496 -5219
rect -13566 -5284 -13496 -5279
rect -12007 -5219 -11937 -5214
rect -12007 -5279 -12002 -5219
rect -12002 -5279 -11942 -5219
rect -11942 -5279 -11937 -5219
rect -12007 -5284 -11937 -5279
rect -10275 -5219 -10205 -5214
rect -10275 -5279 -10270 -5219
rect -10270 -5279 -10210 -5219
rect -10210 -5279 -10205 -5219
rect -10275 -5284 -10205 -5279
rect -8716 -5219 -8646 -5214
rect -8716 -5279 -8711 -5219
rect -8711 -5279 -8651 -5219
rect -8651 -5279 -8646 -5219
rect -8716 -5284 -8646 -5279
rect -20345 -5631 -20089 -5559
rect -19056 -5631 -18800 -5559
rect -18339 -5631 -18083 -5559
rect -17054 -5631 -16798 -5559
rect -15765 -5631 -15509 -5559
rect -15048 -5631 -14792 -5559
rect -13763 -5631 -13507 -5559
rect -12474 -5631 -12218 -5559
rect -11757 -5631 -11501 -5559
rect -10472 -5631 -10216 -5559
rect -9183 -5631 -8927 -5559
rect -8466 -5631 -8210 -5559
rect -20269 -6301 -19934 -6293
rect -20269 -6357 -19934 -6301
rect -19038 -6310 -18966 -6305
rect -19038 -6372 -19033 -6310
rect -19033 -6372 -18971 -6310
rect -18971 -6372 -18966 -6310
rect -19038 -6377 -18966 -6372
rect -18173 -6335 -18107 -6330
rect -18173 -6391 -18168 -6335
rect -18168 -6391 -18112 -6335
rect -18112 -6391 -18107 -6335
rect -18173 -6396 -18107 -6391
rect -16978 -6301 -16643 -6293
rect -16978 -6357 -16643 -6301
rect -15747 -6310 -15675 -6305
rect -15747 -6372 -15742 -6310
rect -15742 -6372 -15680 -6310
rect -15680 -6372 -15675 -6310
rect -15747 -6377 -15675 -6372
rect -14882 -6335 -14816 -6330
rect -14882 -6391 -14877 -6335
rect -14877 -6391 -14821 -6335
rect -14821 -6391 -14816 -6335
rect -14882 -6396 -14816 -6391
rect -13687 -6301 -13352 -6293
rect -13687 -6357 -13352 -6301
rect -12456 -6310 -12384 -6305
rect -12456 -6372 -12451 -6310
rect -12451 -6372 -12389 -6310
rect -12389 -6372 -12384 -6310
rect -12456 -6377 -12384 -6372
rect -11591 -6335 -11525 -6330
rect -11591 -6391 -11586 -6335
rect -11586 -6391 -11530 -6335
rect -11530 -6391 -11525 -6335
rect -11591 -6396 -11525 -6391
rect -10396 -6301 -10061 -6293
rect -10396 -6357 -10061 -6301
rect -9165 -6310 -9093 -6305
rect -9165 -6372 -9160 -6310
rect -9160 -6372 -9098 -6310
rect -9098 -6372 -9093 -6310
rect -9165 -6377 -9093 -6372
rect -8300 -6335 -8234 -6330
rect -8300 -6391 -8295 -6335
rect -8295 -6391 -8239 -6335
rect -8239 -6391 -8234 -6335
rect -8300 -6396 -8234 -6391
rect -20603 -7164 -19481 -7092
rect -19044 -7164 -17922 -7092
rect -17312 -7164 -16190 -7092
rect -15753 -7164 -14631 -7092
rect -14021 -7164 -12899 -7092
rect -12462 -7164 -11340 -7092
rect -10730 -7164 -9608 -7092
rect -9171 -7164 -8049 -7092
rect -21827 -7381 -21658 -7302
rect -22622 -7544 -22068 -7404
rect -22396 -8134 -22056 -8060
rect -21823 -8051 -21674 -7955
rect -20148 -8484 -20078 -8479
rect -20148 -8544 -20143 -8484
rect -20143 -8544 -20083 -8484
rect -20083 -8544 -20078 -8484
rect -20148 -8549 -20078 -8544
rect -18589 -8484 -18519 -8479
rect -18589 -8544 -18584 -8484
rect -18584 -8544 -18524 -8484
rect -18524 -8544 -18519 -8484
rect -18589 -8549 -18519 -8544
rect -16857 -8484 -16787 -8479
rect -16857 -8544 -16852 -8484
rect -16852 -8544 -16792 -8484
rect -16792 -8544 -16787 -8484
rect -16857 -8549 -16787 -8544
rect -15298 -8484 -15228 -8479
rect -15298 -8544 -15293 -8484
rect -15293 -8544 -15233 -8484
rect -15233 -8544 -15228 -8484
rect -15298 -8549 -15228 -8544
rect -13566 -8484 -13496 -8479
rect -13566 -8544 -13561 -8484
rect -13561 -8544 -13501 -8484
rect -13501 -8544 -13496 -8484
rect -13566 -8549 -13496 -8544
rect -12007 -8484 -11937 -8479
rect -12007 -8544 -12002 -8484
rect -12002 -8544 -11942 -8484
rect -11942 -8544 -11937 -8484
rect -12007 -8549 -11937 -8544
rect -10275 -8484 -10205 -8479
rect -10275 -8544 -10270 -8484
rect -10270 -8544 -10210 -8484
rect -10210 -8544 -10205 -8484
rect -10275 -8549 -10205 -8544
rect -8716 -8484 -8646 -8479
rect -8716 -8544 -8711 -8484
rect -8711 -8544 -8651 -8484
rect -8651 -8544 -8646 -8484
rect -8716 -8549 -8646 -8544
rect -21823 -8673 -21654 -8594
rect -22623 -8836 -22069 -8696
rect -20345 -8896 -20089 -8824
rect -19056 -8896 -18800 -8824
rect -18339 -8896 -18083 -8824
rect -17054 -8896 -16798 -8824
rect -15765 -8896 -15509 -8824
rect -15048 -8896 -14792 -8824
rect -13763 -8896 -13507 -8824
rect -12474 -8896 -12218 -8824
rect -11757 -8896 -11501 -8824
rect -10472 -8896 -10216 -8824
rect -9183 -8896 -8927 -8824
rect -8466 -8896 -8210 -8824
rect -22397 -9426 -22057 -9352
rect -21819 -9343 -21670 -9247
rect 11889 167 12141 172
rect 11889 -75 11894 167
rect 11894 -75 12136 167
rect 12136 -75 12141 167
rect 11889 -80 12141 -75
rect 6165 -1279 6231 -1274
rect 6165 -1335 6170 -1279
rect 6170 -1335 6226 -1279
rect 6226 -1335 6231 -1279
rect 6165 -1340 6231 -1335
rect 6605 -1270 6671 -1265
rect 6605 -1326 6610 -1270
rect 6610 -1326 6666 -1270
rect 6666 -1326 6671 -1270
rect 6605 -1331 6671 -1326
rect 12193 -1659 12425 -1654
rect 12193 -1881 12198 -1659
rect 12198 -1881 12420 -1659
rect 12420 -1881 12425 -1659
rect 12193 -1886 12425 -1881
rect 7222 -2813 7410 -2808
rect 7222 -2991 7227 -2813
rect 7227 -2991 7405 -2813
rect 7405 -2991 7410 -2813
rect 7222 -2996 7410 -2991
rect 8157 -2813 8345 -2808
rect 8157 -2991 8162 -2813
rect 8162 -2991 8340 -2813
rect 8340 -2991 8345 -2813
rect 8157 -2996 8345 -2991
rect 9093 -2813 9281 -2808
rect 9093 -2991 9098 -2813
rect 9098 -2991 9276 -2813
rect 9276 -2991 9281 -2813
rect 9093 -2996 9281 -2991
rect 10024 -2813 10211 -2808
rect 10024 -2990 10029 -2813
rect 10029 -2990 10206 -2813
rect 10206 -2990 10211 -2813
rect 10024 -2995 10211 -2990
rect 10951 -2813 11139 -2808
rect 10951 -2991 10956 -2813
rect 10956 -2991 11134 -2813
rect 11134 -2991 11139 -2813
rect 10951 -2996 11139 -2991
rect 12228 -3324 12357 -3319
rect 12228 -3443 12233 -3324
rect 12233 -3443 12352 -3324
rect 12352 -3443 12357 -3324
rect 12228 -3448 12357 -3443
rect 12955 -3365 13084 -3360
rect 12955 -3484 12960 -3365
rect 12960 -3484 13079 -3365
rect 13079 -3484 13084 -3365
rect 12955 -3489 13084 -3484
rect 5727 -5726 5793 -5721
rect 5727 -5782 5732 -5726
rect 5732 -5782 5788 -5726
rect 5788 -5782 5793 -5726
rect 5727 -5787 5793 -5782
rect -20269 -9566 -19934 -9558
rect -20269 -9622 -19934 -9566
rect -19038 -9575 -18966 -9570
rect -19038 -9637 -19033 -9575
rect -19033 -9637 -18971 -9575
rect -18971 -9637 -18966 -9575
rect -19038 -9642 -18966 -9637
rect -18173 -9600 -18107 -9595
rect -18173 -9656 -18168 -9600
rect -18168 -9656 -18112 -9600
rect -18112 -9656 -18107 -9600
rect -18173 -9661 -18107 -9656
rect -16978 -9566 -16643 -9558
rect -16978 -9622 -16643 -9566
rect -15747 -9575 -15675 -9570
rect -15747 -9637 -15742 -9575
rect -15742 -9637 -15680 -9575
rect -15680 -9637 -15675 -9575
rect -15747 -9642 -15675 -9637
rect -14882 -9600 -14816 -9595
rect -14882 -9656 -14877 -9600
rect -14877 -9656 -14821 -9600
rect -14821 -9656 -14816 -9600
rect -14882 -9661 -14816 -9656
rect -13687 -9566 -13352 -9558
rect -13687 -9622 -13352 -9566
rect -12456 -9575 -12384 -9570
rect -12456 -9637 -12451 -9575
rect -12451 -9637 -12389 -9575
rect -12389 -9637 -12384 -9575
rect -12456 -9642 -12384 -9637
rect -11591 -9600 -11525 -9595
rect -11591 -9656 -11586 -9600
rect -11586 -9656 -11530 -9600
rect -11530 -9656 -11525 -9600
rect -11591 -9661 -11525 -9656
rect -10396 -9566 -10061 -9558
rect -10396 -9622 -10061 -9566
rect -9165 -9575 -9093 -9570
rect -9165 -9637 -9160 -9575
rect -9160 -9637 -9098 -9575
rect -9098 -9637 -9093 -9575
rect -9165 -9642 -9093 -9637
rect -8300 -9600 -8234 -9595
rect -8300 -9656 -8295 -9600
rect -8295 -9656 -8239 -9600
rect -8239 -9656 -8234 -9600
rect -8300 -9661 -8234 -9656
rect -20603 -10428 -19481 -10356
rect -19044 -10428 -17922 -10356
rect -17312 -10428 -16190 -10356
rect -15753 -10428 -14631 -10356
rect -14021 -10428 -12899 -10356
rect -12462 -10428 -11340 -10356
rect -10730 -10428 -9608 -10356
rect -9171 -10428 -8049 -10356
rect -21827 -10645 -21658 -10566
rect -22622 -10808 -22068 -10668
rect -24133 -11398 -23793 -11324
rect -23556 -11315 -23407 -11219
rect -23560 -11937 -23391 -11858
rect -24359 -12100 -23805 -11960
rect -24133 -12690 -23793 -12616
rect -23556 -12607 -23407 -12511
rect -22396 -11398 -22056 -11324
rect -21823 -11315 -21674 -11219
rect -20148 -11748 -20078 -11743
rect -20148 -11808 -20143 -11748
rect -20143 -11808 -20083 -11748
rect -20083 -11808 -20078 -11748
rect -20148 -11813 -20078 -11808
rect -18589 -11748 -18519 -11743
rect -18589 -11808 -18584 -11748
rect -18584 -11808 -18524 -11748
rect -18524 -11808 -18519 -11748
rect -18589 -11813 -18519 -11808
rect -16857 -11748 -16787 -11743
rect -16857 -11808 -16852 -11748
rect -16852 -11808 -16792 -11748
rect -16792 -11808 -16787 -11748
rect -16857 -11813 -16787 -11808
rect -15298 -11748 -15228 -11743
rect -15298 -11808 -15293 -11748
rect -15293 -11808 -15233 -11748
rect -15233 -11808 -15228 -11748
rect -15298 -11813 -15228 -11808
rect -13566 -11748 -13496 -11743
rect -13566 -11808 -13561 -11748
rect -13561 -11808 -13501 -11748
rect -13501 -11808 -13496 -11748
rect -13566 -11813 -13496 -11808
rect -12007 -11748 -11937 -11743
rect -12007 -11808 -12002 -11748
rect -12002 -11808 -11942 -11748
rect -11942 -11808 -11937 -11748
rect -12007 -11813 -11937 -11808
rect -10275 -11748 -10205 -11743
rect -10275 -11808 -10270 -11748
rect -10270 -11808 -10210 -11748
rect -10210 -11808 -10205 -11748
rect -10275 -11813 -10205 -11808
rect -8716 -11748 -8646 -11743
rect -8716 -11808 -8711 -11748
rect -8711 -11808 -8651 -11748
rect -8651 -11808 -8646 -11748
rect -8716 -11813 -8646 -11808
rect -21831 -11937 -21662 -11858
rect -22622 -12100 -22068 -11960
rect -20345 -12160 -20089 -12088
rect -19056 -12160 -18800 -12088
rect -18339 -12160 -18083 -12088
rect -17054 -12160 -16798 -12088
rect -15765 -12160 -15509 -12088
rect -15048 -12160 -14792 -12088
rect -13763 -12160 -13507 -12088
rect -12474 -12160 -12218 -12088
rect -11757 -12160 -11501 -12088
rect -10472 -12160 -10216 -12088
rect -9183 -12160 -8927 -12088
rect -8466 -12160 -8210 -12088
rect -22396 -12690 -22056 -12616
rect -21827 -12607 -21678 -12511
rect -20269 -12830 -19934 -12822
rect -20269 -12886 -19934 -12830
rect -19038 -12839 -18966 -12834
rect -19038 -12901 -19033 -12839
rect -19033 -12901 -18971 -12839
rect -18971 -12901 -18966 -12839
rect -19038 -12906 -18966 -12901
rect -18173 -12864 -18107 -12859
rect -18173 -12920 -18168 -12864
rect -18168 -12920 -18112 -12864
rect -18112 -12920 -18107 -12864
rect -18173 -12925 -18107 -12920
rect -16978 -12830 -16643 -12822
rect -16978 -12886 -16643 -12830
rect -15747 -12839 -15675 -12834
rect -15747 -12901 -15742 -12839
rect -15742 -12901 -15680 -12839
rect -15680 -12901 -15675 -12839
rect -15747 -12906 -15675 -12901
rect -14882 -12864 -14816 -12859
rect -14882 -12920 -14877 -12864
rect -14877 -12920 -14821 -12864
rect -14821 -12920 -14816 -12864
rect -14882 -12925 -14816 -12920
rect -13687 -12830 -13352 -12822
rect -13687 -12886 -13352 -12830
rect -12456 -12839 -12384 -12834
rect -12456 -12901 -12451 -12839
rect -12451 -12901 -12389 -12839
rect -12389 -12901 -12384 -12839
rect -12456 -12906 -12384 -12901
rect -11591 -12864 -11525 -12859
rect -11591 -12920 -11586 -12864
rect -11586 -12920 -11530 -12864
rect -11530 -12920 -11525 -12864
rect -11591 -12925 -11525 -12920
rect -10396 -12830 -10061 -12822
rect -10396 -12886 -10061 -12830
rect -9165 -12839 -9093 -12834
rect -9165 -12901 -9160 -12839
rect -9160 -12901 -9098 -12839
rect -9098 -12901 -9093 -12839
rect -9165 -12906 -9093 -12901
rect -8300 -12864 -8234 -12859
rect -8300 -12920 -8295 -12864
rect -8295 -12920 -8239 -12864
rect -8239 -12920 -8234 -12864
rect -8300 -12925 -8234 -12920
rect 11889 -4361 12141 -4356
rect 11889 -4603 11894 -4361
rect 11894 -4603 12136 -4361
rect 12136 -4603 12141 -4361
rect 11889 -4608 12141 -4603
rect 6165 -5707 6231 -5702
rect 6165 -5763 6170 -5707
rect 6170 -5763 6226 -5707
rect 6226 -5763 6231 -5707
rect 6165 -5768 6231 -5763
rect 6605 -5698 6671 -5693
rect 6605 -5754 6610 -5698
rect 6610 -5754 6666 -5698
rect 6666 -5754 6671 -5698
rect 6605 -5759 6671 -5754
rect 12193 -6087 12425 -6082
rect 12193 -6309 12198 -6087
rect 12198 -6309 12420 -6087
rect 12420 -6309 12425 -6087
rect 12193 -6314 12425 -6309
rect 7222 -7241 7410 -7236
rect 7222 -7419 7227 -7241
rect 7227 -7419 7405 -7241
rect 7405 -7419 7410 -7241
rect 7222 -7424 7410 -7419
rect 8157 -7241 8345 -7236
rect 8157 -7419 8162 -7241
rect 8162 -7419 8340 -7241
rect 8340 -7419 8345 -7241
rect 8157 -7424 8345 -7419
rect 9093 -7241 9281 -7236
rect 9093 -7419 9098 -7241
rect 9098 -7419 9276 -7241
rect 9276 -7419 9281 -7241
rect 9093 -7424 9281 -7419
rect 10024 -7241 10211 -7236
rect 10024 -7418 10029 -7241
rect 10029 -7418 10206 -7241
rect 10206 -7418 10211 -7241
rect 10024 -7423 10211 -7418
rect 10951 -7241 11139 -7236
rect 10951 -7419 10956 -7241
rect 10956 -7419 11134 -7241
rect 11134 -7419 11139 -7241
rect 10951 -7424 11139 -7419
rect 12228 -7752 12357 -7747
rect 12228 -7871 12233 -7752
rect 12233 -7871 12352 -7752
rect 12352 -7871 12357 -7752
rect 12228 -7876 12357 -7871
rect 12955 -7793 13084 -7788
rect 12955 -7912 12960 -7793
rect 12960 -7912 13079 -7793
rect 13079 -7912 13084 -7793
rect 12955 -7917 13084 -7912
rect 11889 -8789 12141 -8784
rect 11889 -9031 11894 -8789
rect 11894 -9031 12136 -8789
rect 12136 -9031 12141 -8789
rect 11889 -9036 12141 -9031
rect 5727 -10354 5793 -10349
rect 5727 -10410 5732 -10354
rect 5732 -10410 5788 -10354
rect 5788 -10410 5793 -10354
rect 5727 -10415 5793 -10410
rect -2309 -14063 -2195 -14058
rect -2309 -14167 -2304 -14063
rect -2304 -14167 -2200 -14063
rect -2200 -14167 -2195 -14063
rect -2309 -14172 -2195 -14167
rect -1293 -14074 -1186 -14069
rect -1293 -14171 -1288 -14074
rect -1288 -14171 -1191 -14074
rect -1191 -14171 -1186 -14074
rect -1293 -14176 -1186 -14171
rect -23426 -15075 -23315 -15070
rect -23426 -15176 -23421 -15075
rect -23421 -15176 -23320 -15075
rect -23320 -15176 -23315 -15075
rect -23426 -15181 -23315 -15176
rect -24844 -15194 -24738 -15189
rect -24844 -15290 -24839 -15194
rect -24839 -15290 -24743 -15194
rect -24743 -15290 -24738 -15194
rect -24844 -15295 -24738 -15290
rect -18077 -15281 -17993 -15276
rect -18077 -15355 -18072 -15281
rect -18072 -15355 -17998 -15281
rect -17998 -15355 -17993 -15281
rect -18077 -15360 -17993 -15355
rect -16914 -15326 -16844 -15321
rect -16914 -15386 -16909 -15326
rect -16909 -15386 -16849 -15326
rect -16849 -15386 -16844 -15326
rect -16914 -15391 -16844 -15386
rect -12473 -15345 -12401 -14223
rect -5025 -14259 -4911 -14255
rect -5025 -14365 -5021 -14259
rect -5021 -14365 -4915 -14259
rect -4915 -14365 -4911 -14259
rect -5025 -14369 -4911 -14365
rect -4009 -14250 -3902 -14245
rect -4009 -14347 -4004 -14250
rect -4004 -14347 -3907 -14250
rect -3907 -14347 -3902 -14250
rect -4009 -14352 -3902 -14347
rect -11086 -14825 -11016 -14820
rect -11086 -14885 -11081 -14825
rect -11081 -14885 -11021 -14825
rect -11021 -14885 -11016 -14825
rect -11086 -14890 -11016 -14885
rect -8499 -15425 -8429 -15420
rect -8499 -15485 -8494 -15425
rect -8494 -15485 -8434 -15425
rect -8434 -15485 -8429 -15425
rect -8499 -15490 -8429 -15485
rect -7209 -15397 -7110 -15392
rect -7209 -15486 -7204 -15397
rect -7204 -15486 -7115 -15397
rect -7115 -15486 -7110 -15397
rect -7209 -15491 -7110 -15486
rect -5025 -14887 -4911 -14882
rect -5025 -14991 -5020 -14887
rect -5020 -14991 -4916 -14887
rect -4916 -14991 -4911 -14887
rect -5025 -14996 -4911 -14991
rect -4009 -14883 -3902 -14878
rect -4009 -14980 -4004 -14883
rect -4004 -14980 -3907 -14883
rect -3907 -14980 -3902 -14883
rect -4009 -14985 -3902 -14980
rect -2309 -14882 -2195 -14877
rect -2309 -14986 -2304 -14882
rect -2304 -14986 -2200 -14882
rect -2200 -14986 -2195 -14882
rect -2309 -14991 -2195 -14986
rect -1293 -14893 -1186 -14888
rect -1293 -14990 -1288 -14893
rect -1288 -14990 -1191 -14893
rect -1191 -14990 -1186 -14893
rect -1293 -14995 -1186 -14990
rect -8505 -15934 -8435 -15929
rect -8505 -15994 -8500 -15934
rect -8500 -15994 -8440 -15934
rect -8440 -15994 -8435 -15934
rect -8505 -15999 -8435 -15994
rect -7216 -15890 -7117 -15885
rect -7216 -15979 -7211 -15890
rect -7211 -15979 -7122 -15890
rect -7122 -15979 -7117 -15890
rect -7216 -15984 -7117 -15979
rect -5025 -15706 -4911 -15701
rect -5025 -15810 -5020 -15706
rect -5020 -15810 -4916 -15706
rect -4916 -15810 -4911 -15706
rect -5025 -15815 -4911 -15810
rect -4009 -15702 -3902 -15697
rect -4009 -15799 -4004 -15702
rect -4004 -15799 -3907 -15702
rect -3907 -15799 -3902 -15702
rect -4009 -15804 -3902 -15799
rect -2309 -15701 -2195 -15696
rect -2309 -15805 -2304 -15701
rect -2304 -15805 -2200 -15701
rect -2200 -15805 -2195 -15701
rect -2309 -15810 -2195 -15805
rect -1293 -15712 -1186 -15707
rect -1293 -15809 -1288 -15712
rect -1288 -15809 -1191 -15712
rect -1191 -15809 -1186 -15712
rect -1293 -15814 -1186 -15809
rect -24840 -16368 -24734 -16363
rect -24840 -16464 -24835 -16368
rect -24835 -16464 -24739 -16368
rect -24739 -16464 -24734 -16368
rect -24840 -16469 -24734 -16464
rect -23383 -16271 -23272 -16266
rect -23383 -16372 -23378 -16271
rect -23378 -16372 -23277 -16271
rect -23277 -16372 -23272 -16271
rect -23383 -16377 -23272 -16372
rect -18089 -16683 -18005 -16678
rect -18089 -16757 -18084 -16683
rect -18084 -16757 -18010 -16683
rect -18010 -16757 -18005 -16683
rect -18089 -16762 -18005 -16757
rect -16914 -16732 -16844 -16727
rect -16914 -16792 -16909 -16732
rect -16909 -16792 -16849 -16732
rect -16849 -16792 -16844 -16732
rect -16914 -16797 -16844 -16792
rect -24834 -17600 -24728 -17595
rect -24834 -17696 -24829 -17600
rect -24829 -17696 -24733 -17600
rect -24733 -17696 -24728 -17600
rect -24834 -17701 -24728 -17696
rect -23374 -17483 -23263 -17478
rect -23374 -17584 -23369 -17483
rect -23369 -17584 -23268 -17483
rect -23268 -17584 -23263 -17483
rect -23374 -17589 -23263 -17584
rect -21938 -18113 -21868 -18108
rect -21938 -18173 -21933 -18113
rect -21933 -18173 -21873 -18113
rect -21873 -18173 -21868 -18113
rect -21938 -18178 -21868 -18173
rect -20648 -18085 -20549 -18080
rect -20648 -18174 -20643 -18085
rect -20643 -18174 -20554 -18085
rect -20554 -18174 -20549 -18085
rect -20648 -18179 -20549 -18174
rect -16347 -17984 -16277 -17979
rect -16347 -18044 -16342 -17984
rect -16342 -18044 -16282 -17984
rect -16282 -18044 -16277 -17984
rect -16347 -18049 -16277 -18044
rect -18093 -18069 -18009 -18064
rect -18093 -18143 -18088 -18069
rect -18088 -18143 -18014 -18069
rect -18014 -18143 -18009 -18069
rect -18093 -18148 -18009 -18143
rect -15057 -17956 -14958 -17951
rect -15057 -18045 -15052 -17956
rect -15052 -18045 -14963 -17956
rect -14963 -18045 -14958 -17956
rect -15057 -18050 -14958 -18045
rect -17045 -18163 -16975 -18158
rect -17045 -18223 -17040 -18163
rect -17040 -18223 -16980 -18163
rect -16980 -18223 -16975 -18163
rect -17045 -18228 -16975 -18223
rect -24820 -18714 -24714 -18709
rect -24820 -18810 -24815 -18714
rect -24815 -18810 -24719 -18714
rect -24719 -18810 -24714 -18714
rect -24820 -18815 -24714 -18810
rect -23366 -18624 -23255 -18619
rect -23366 -18725 -23361 -18624
rect -23361 -18725 -23260 -18624
rect -23260 -18725 -23255 -18624
rect -23366 -18730 -23255 -18725
rect -21944 -18622 -21874 -18617
rect -21944 -18682 -21939 -18622
rect -21939 -18682 -21879 -18622
rect -21879 -18682 -21874 -18622
rect -21944 -18687 -21874 -18682
rect -20655 -18578 -20556 -18573
rect -20655 -18667 -20650 -18578
rect -20650 -18667 -20561 -18578
rect -20561 -18667 -20556 -18578
rect -16353 -18493 -16283 -18488
rect -16353 -18553 -16348 -18493
rect -16348 -18553 -16288 -18493
rect -16288 -18553 -16283 -18493
rect -16353 -18558 -16283 -18553
rect -15064 -18449 -14965 -18444
rect -15064 -18538 -15059 -18449
rect -15059 -18538 -14970 -18449
rect -14970 -18538 -14965 -18449
rect -15064 -18543 -14965 -18538
rect -20655 -18672 -20556 -18667
rect -12471 -18161 -12399 -17039
rect -11084 -17641 -11014 -17636
rect -11084 -17701 -11079 -17641
rect -11079 -17701 -11019 -17641
rect -11019 -17701 -11014 -17641
rect -11084 -17706 -11014 -17701
rect -8505 -16417 -8435 -16412
rect -8505 -16477 -8500 -16417
rect -8500 -16477 -8440 -16417
rect -8440 -16477 -8435 -16417
rect -8505 -16482 -8435 -16477
rect -7217 -16376 -7118 -16371
rect -7217 -16465 -7212 -16376
rect -7212 -16465 -7123 -16376
rect -7123 -16465 -7118 -16376
rect -7217 -16470 -7118 -16465
rect -5025 -16525 -4911 -16520
rect -5025 -16629 -5020 -16525
rect -5020 -16629 -4916 -16525
rect -4916 -16629 -4911 -16525
rect -5025 -16634 -4911 -16629
rect -4009 -16521 -3902 -16516
rect -4009 -16618 -4004 -16521
rect -4004 -16618 -3907 -16521
rect -3907 -16618 -3902 -16521
rect -4009 -16623 -3902 -16618
rect -2309 -16520 -2195 -16515
rect -2309 -16624 -2304 -16520
rect -2304 -16624 -2200 -16520
rect -2200 -16624 -2195 -16520
rect -2309 -16629 -2195 -16624
rect -1293 -16531 -1186 -16526
rect -1293 -16628 -1288 -16531
rect -1288 -16628 -1191 -16531
rect -1191 -16628 -1186 -16531
rect -1293 -16633 -1186 -16628
rect -21944 -19105 -21874 -19100
rect -21944 -19165 -21939 -19105
rect -21939 -19165 -21879 -19105
rect -21879 -19165 -21874 -19105
rect -21944 -19170 -21874 -19165
rect -20656 -19064 -20557 -19059
rect -20656 -19153 -20651 -19064
rect -20651 -19153 -20562 -19064
rect -20562 -19153 -20557 -19064
rect -20656 -19158 -20557 -19153
rect -20660 -19571 -20561 -19566
rect -21944 -19627 -21874 -19622
rect -21944 -19687 -21939 -19627
rect -21939 -19687 -21879 -19627
rect -21879 -19687 -21874 -19627
rect -21944 -19692 -21874 -19687
rect -20660 -19660 -20655 -19571
rect -20655 -19660 -20566 -19571
rect -20566 -19660 -20561 -19571
rect -20660 -19665 -20561 -19660
rect -24820 -19908 -24714 -19903
rect -24820 -20004 -24815 -19908
rect -24815 -20004 -24719 -19908
rect -24719 -20004 -24714 -19908
rect -24820 -20009 -24714 -20004
rect -23343 -19796 -23232 -19791
rect -23343 -19897 -23338 -19796
rect -23338 -19897 -23237 -19796
rect -23237 -19897 -23232 -19796
rect -23343 -19902 -23232 -19897
rect -16353 -18976 -16283 -18971
rect -16353 -19036 -16348 -18976
rect -16348 -19036 -16288 -18976
rect -16288 -19036 -16283 -18976
rect -16353 -19041 -16283 -19036
rect -15065 -18935 -14966 -18930
rect -15065 -19024 -15060 -18935
rect -15060 -19024 -14971 -18935
rect -14971 -19024 -14966 -18935
rect -15065 -19029 -14966 -19024
rect -15069 -19442 -14970 -19437
rect -18091 -19475 -18007 -19470
rect -18091 -19549 -18086 -19475
rect -18086 -19549 -18012 -19475
rect -18012 -19549 -18007 -19475
rect -18091 -19554 -18007 -19549
rect -16353 -19498 -16283 -19493
rect -16353 -19558 -16348 -19498
rect -16348 -19558 -16288 -19498
rect -16288 -19558 -16283 -19498
rect -16353 -19563 -16283 -19558
rect -15069 -19531 -15064 -19442
rect -15064 -19531 -14975 -19442
rect -14975 -19531 -14970 -19442
rect -15069 -19536 -14970 -19531
rect -16930 -19618 -16860 -19613
rect -16930 -19678 -16925 -19618
rect -16925 -19678 -16865 -19618
rect -16865 -19678 -16860 -19618
rect -16930 -19683 -16860 -19678
rect -21941 -20096 -21871 -20091
rect -21941 -20156 -21936 -20096
rect -21936 -20156 -21876 -20096
rect -21876 -20156 -21871 -20096
rect -21941 -20161 -21871 -20156
rect -20659 -20046 -20560 -20041
rect -20659 -20135 -20654 -20046
rect -20654 -20135 -20565 -20046
rect -20565 -20135 -20560 -20046
rect -20659 -20140 -20560 -20135
rect -16350 -19967 -16280 -19962
rect -16350 -20027 -16345 -19967
rect -16345 -20027 -16285 -19967
rect -16285 -20027 -16280 -19967
rect -16350 -20032 -16280 -20027
rect -15068 -19917 -14969 -19912
rect -15068 -20006 -15063 -19917
rect -15063 -20006 -14974 -19917
rect -14974 -20006 -14969 -19917
rect -15068 -20011 -14969 -20006
rect -20654 -20498 -20555 -20493
rect -21939 -20553 -21869 -20548
rect -21939 -20613 -21934 -20553
rect -21934 -20613 -21874 -20553
rect -21874 -20613 -21869 -20553
rect -21939 -20618 -21869 -20613
rect -20654 -20587 -20649 -20498
rect -20649 -20587 -20560 -20498
rect -20560 -20587 -20555 -20498
rect -20654 -20592 -20555 -20587
rect -20654 -20940 -20555 -20935
rect -24820 -21104 -24714 -21099
rect -24820 -21200 -24815 -21104
rect -24815 -21200 -24719 -21104
rect -24719 -21200 -24714 -21104
rect -24820 -21205 -24714 -21200
rect -23334 -20994 -23223 -20989
rect -23334 -21095 -23329 -20994
rect -23329 -21095 -23228 -20994
rect -23228 -21095 -23223 -20994
rect -23334 -21100 -23223 -21095
rect -21937 -21018 -21867 -21013
rect -21937 -21078 -21932 -21018
rect -21932 -21078 -21872 -21018
rect -21872 -21078 -21867 -21018
rect -21937 -21083 -21867 -21078
rect -20654 -21029 -20649 -20940
rect -20649 -21029 -20560 -20940
rect -20560 -21029 -20555 -20940
rect -20654 -21034 -20555 -21029
rect -15063 -20369 -14964 -20364
rect -16348 -20424 -16278 -20419
rect -16348 -20484 -16343 -20424
rect -16343 -20484 -16283 -20424
rect -16283 -20484 -16278 -20424
rect -16348 -20489 -16278 -20484
rect -15063 -20458 -15058 -20369
rect -15058 -20458 -14969 -20369
rect -14969 -20458 -14964 -20369
rect -15063 -20463 -14964 -20458
rect -15063 -20811 -14964 -20806
rect -18095 -20869 -18011 -20864
rect -18095 -20943 -18090 -20869
rect -18090 -20943 -18016 -20869
rect -18016 -20943 -18011 -20869
rect -18095 -20948 -18011 -20943
rect -16346 -20889 -16276 -20884
rect -16346 -20949 -16341 -20889
rect -16341 -20949 -16281 -20889
rect -16281 -20949 -16276 -20889
rect -16346 -20954 -16276 -20949
rect -15063 -20900 -15058 -20811
rect -15058 -20900 -14969 -20811
rect -14969 -20900 -14964 -20811
rect -15063 -20905 -14964 -20900
rect -16921 -21013 -16849 -21008
rect -16921 -21075 -16916 -21013
rect -16916 -21075 -16854 -21013
rect -16854 -21075 -16849 -21013
rect -16921 -21080 -16849 -21075
rect -23337 -22288 -23226 -22283
rect -23337 -22389 -23332 -22288
rect -23332 -22389 -23231 -22288
rect -23231 -22389 -23226 -22288
rect -23337 -22394 -23226 -22389
rect -24810 -22412 -24704 -22407
rect -24810 -22508 -24805 -22412
rect -24805 -22508 -24709 -22412
rect -24709 -22508 -24704 -22412
rect -24810 -22513 -24704 -22508
rect -21933 -21499 -21863 -21494
rect -21933 -21559 -21928 -21499
rect -21928 -21559 -21868 -21499
rect -21868 -21559 -21863 -21499
rect -21933 -21564 -21863 -21559
rect -20660 -21421 -20561 -21416
rect -20660 -21510 -20655 -21421
rect -20655 -21510 -20566 -21421
rect -20566 -21510 -20561 -21421
rect -20660 -21515 -20561 -21510
rect -16342 -21370 -16272 -21365
rect -16342 -21430 -16337 -21370
rect -16337 -21430 -16277 -21370
rect -16277 -21430 -16272 -21370
rect -16342 -21435 -16272 -21430
rect -15069 -21292 -14970 -21287
rect -15069 -21381 -15064 -21292
rect -15064 -21381 -14975 -21292
rect -14975 -21381 -14970 -21292
rect -15069 -21386 -14970 -21381
rect -16731 -21983 -16657 -21978
rect -16731 -22047 -16726 -21983
rect -16726 -22047 -16662 -21983
rect -16662 -22047 -16657 -21983
rect -16731 -22052 -16657 -22047
rect -18093 -22273 -18009 -22268
rect -18093 -22347 -18088 -22273
rect -18088 -22347 -18014 -22273
rect -18014 -22347 -18009 -22273
rect -18093 -22352 -18009 -22347
rect -24830 -23718 -24724 -23713
rect -24830 -23814 -24825 -23718
rect -24825 -23814 -24729 -23718
rect -24729 -23814 -24724 -23718
rect -24830 -23819 -24724 -23814
rect -23377 -23604 -23266 -23599
rect -23377 -23705 -23372 -23604
rect -23372 -23705 -23271 -23604
rect -23271 -23705 -23266 -23604
rect -23377 -23710 -23266 -23705
rect -16693 -23367 -16605 -23362
rect -16693 -23445 -16688 -23367
rect -16688 -23445 -16610 -23367
rect -16610 -23445 -16605 -23367
rect -16693 -23450 -16605 -23445
rect -18095 -23675 -18011 -23670
rect -18095 -23749 -18090 -23675
rect -18090 -23749 -18016 -23675
rect -18016 -23749 -18011 -23675
rect -18095 -23754 -18011 -23749
rect -16693 -24775 -16609 -24770
rect -16693 -24849 -16688 -24775
rect -16688 -24849 -16614 -24775
rect -16614 -24849 -16609 -24775
rect -16693 -24854 -16609 -24849
rect -18089 -25055 -18005 -25050
rect -18089 -25129 -18084 -25055
rect -18084 -25129 -18010 -25055
rect -18010 -25129 -18005 -25055
rect -18089 -25134 -18005 -25129
rect -12471 -21118 -12399 -19996
rect -11084 -20598 -11014 -20593
rect -11084 -20658 -11079 -20598
rect -11079 -20658 -11019 -20598
rect -11019 -20658 -11014 -20598
rect -11084 -20663 -11014 -20658
rect -7221 -16883 -7122 -16878
rect -8505 -16939 -8435 -16934
rect -8505 -16999 -8500 -16939
rect -8500 -16999 -8440 -16939
rect -8440 -16999 -8435 -16939
rect -8505 -17004 -8435 -16999
rect -7221 -16972 -7216 -16883
rect -7216 -16972 -7127 -16883
rect -7127 -16972 -7122 -16883
rect -7221 -16977 -7122 -16972
rect -12471 -23697 -12399 -22575
rect -11084 -23177 -11014 -23172
rect -11084 -23237 -11079 -23177
rect -11079 -23237 -11019 -23177
rect -11019 -23237 -11014 -23177
rect -11084 -23242 -11014 -23237
rect -8502 -17408 -8432 -17403
rect -8502 -17468 -8497 -17408
rect -8497 -17468 -8437 -17408
rect -8437 -17468 -8432 -17408
rect -8502 -17473 -8432 -17468
rect -7220 -17358 -7121 -17353
rect -7220 -17447 -7215 -17358
rect -7215 -17447 -7126 -17358
rect -7126 -17447 -7121 -17358
rect -7220 -17452 -7121 -17447
rect -5025 -17344 -4911 -17339
rect -5025 -17448 -5020 -17344
rect -5020 -17448 -4916 -17344
rect -4916 -17448 -4911 -17344
rect -5025 -17453 -4911 -17448
rect -4009 -17340 -3902 -17335
rect -4009 -17437 -4004 -17340
rect -4004 -17437 -3907 -17340
rect -3907 -17437 -3902 -17340
rect -4009 -17442 -3902 -17437
rect -2309 -17339 -2195 -17334
rect -2309 -17443 -2304 -17339
rect -2304 -17443 -2200 -17339
rect -2200 -17443 -2195 -17339
rect -2309 -17448 -2195 -17443
rect -1293 -17350 -1186 -17345
rect -1293 -17447 -1288 -17350
rect -1288 -17447 -1191 -17350
rect -1191 -17447 -1186 -17350
rect -1293 -17452 -1186 -17447
rect -12471 -26465 -12399 -25343
rect -11084 -25945 -11014 -25940
rect -11084 -26005 -11079 -25945
rect -11079 -26005 -11019 -25945
rect -11019 -26005 -11014 -25945
rect -11084 -26010 -11014 -26005
rect -7215 -17810 -7116 -17805
rect -8500 -17865 -8430 -17860
rect -8500 -17925 -8495 -17865
rect -8495 -17925 -8435 -17865
rect -8435 -17925 -8430 -17865
rect -8500 -17930 -8430 -17925
rect -7215 -17899 -7210 -17810
rect -7210 -17899 -7121 -17810
rect -7121 -17899 -7116 -17810
rect -7215 -17904 -7116 -17899
rect -12471 -29098 -12399 -27976
rect -11084 -28578 -11014 -28573
rect -11084 -28638 -11079 -28578
rect -11079 -28638 -11019 -28578
rect -11019 -28638 -11014 -28578
rect -11084 -28643 -11014 -28638
rect -7215 -18252 -7116 -18247
rect -8498 -18330 -8428 -18325
rect -8498 -18390 -8493 -18330
rect -8493 -18390 -8433 -18330
rect -8433 -18390 -8428 -18330
rect -8498 -18395 -8428 -18390
rect -7215 -18341 -7210 -18252
rect -7210 -18341 -7121 -18252
rect -7121 -18341 -7116 -18252
rect -7215 -18346 -7116 -18341
rect -12471 -31707 -12399 -30585
rect -11084 -31187 -11014 -31182
rect -11084 -31247 -11079 -31187
rect -11079 -31247 -11019 -31187
rect -11019 -31247 -11014 -31187
rect -11084 -31252 -11014 -31247
rect -8494 -18811 -8424 -18806
rect -8494 -18871 -8489 -18811
rect -8489 -18871 -8429 -18811
rect -8429 -18871 -8424 -18811
rect -8494 -18876 -8424 -18871
rect -7221 -18733 -7122 -18728
rect -7221 -18822 -7216 -18733
rect -7216 -18822 -7127 -18733
rect -7127 -18822 -7122 -18733
rect -7221 -18827 -7122 -18822
rect -12473 -34327 -12401 -33205
rect -11086 -33807 -11016 -33802
rect -11086 -33867 -11081 -33807
rect -11081 -33867 -11021 -33807
rect -11021 -33867 -11016 -33807
rect -11086 -33872 -11016 -33867
rect -5025 -18163 -4911 -18158
rect -5025 -18267 -5020 -18163
rect -5020 -18267 -4916 -18163
rect -4916 -18267 -4911 -18163
rect -5025 -18272 -4911 -18267
rect -4009 -18159 -3902 -18154
rect -4009 -18256 -4004 -18159
rect -4004 -18256 -3907 -18159
rect -3907 -18256 -3902 -18159
rect -4009 -18261 -3902 -18256
rect -2309 -18158 -2195 -18153
rect -2309 -18262 -2304 -18158
rect -2304 -18262 -2200 -18158
rect -2200 -18262 -2195 -18158
rect -2309 -18267 -2195 -18262
rect -1293 -18169 -1186 -18164
rect -1293 -18266 -1288 -18169
rect -1288 -18266 -1191 -18169
rect -1191 -18266 -1186 -18169
rect -1293 -18271 -1186 -18266
rect 6165 -10335 6231 -10330
rect 6165 -10391 6170 -10335
rect 6170 -10391 6226 -10335
rect 6226 -10391 6231 -10335
rect 6165 -10396 6231 -10391
rect 6605 -10326 6671 -10321
rect 6605 -10382 6610 -10326
rect 6610 -10382 6666 -10326
rect 6666 -10382 6671 -10326
rect 6605 -10387 6671 -10382
rect 12193 -10715 12425 -10710
rect 12193 -10937 12198 -10715
rect 12198 -10937 12420 -10715
rect 12420 -10937 12425 -10715
rect 12193 -10942 12425 -10937
rect 7222 -11869 7410 -11864
rect 7222 -12047 7227 -11869
rect 7227 -12047 7405 -11869
rect 7405 -12047 7410 -11869
rect 7222 -12052 7410 -12047
rect 8157 -11869 8345 -11864
rect 8157 -12047 8162 -11869
rect 8162 -12047 8340 -11869
rect 8340 -12047 8345 -11869
rect 8157 -12052 8345 -12047
rect 9093 -11869 9281 -11864
rect 9093 -12047 9098 -11869
rect 9098 -12047 9276 -11869
rect 9276 -12047 9281 -11869
rect 9093 -12052 9281 -12047
rect 10024 -11869 10211 -11864
rect 10024 -12046 10029 -11869
rect 10029 -12046 10206 -11869
rect 10206 -12046 10211 -11869
rect 10024 -12051 10211 -12046
rect 10951 -11869 11139 -11864
rect 10951 -12047 10956 -11869
rect 10956 -12047 11134 -11869
rect 11134 -12047 11139 -11869
rect 10951 -12052 11139 -12047
rect 12228 -12380 12357 -12375
rect 12228 -12499 12233 -12380
rect 12233 -12499 12352 -12380
rect 12352 -12499 12357 -12380
rect 12228 -12504 12357 -12499
rect 12955 -12421 13084 -12416
rect 12955 -12540 12960 -12421
rect 12960 -12540 13079 -12421
rect 13079 -12540 13084 -12421
rect 12955 -12545 13084 -12540
rect 5727 -14882 5793 -14877
rect 5727 -14938 5732 -14882
rect 5732 -14938 5788 -14882
rect 5788 -14938 5793 -14882
rect 5727 -14943 5793 -14938
rect -5025 -18982 -4911 -18977
rect -5025 -19086 -5020 -18982
rect -5020 -19086 -4916 -18982
rect -4916 -19086 -4911 -18982
rect -5025 -19091 -4911 -19086
rect -4009 -18978 -3902 -18973
rect -4009 -19075 -4004 -18978
rect -4004 -19075 -3907 -18978
rect -3907 -19075 -3902 -18978
rect -4009 -19080 -3902 -19075
rect -2309 -18977 -2195 -18972
rect -2309 -19081 -2304 -18977
rect -2304 -19081 -2200 -18977
rect -2200 -19081 -2195 -18977
rect -2309 -19086 -2195 -19081
rect -1293 -18988 -1186 -18983
rect -1293 -19085 -1288 -18988
rect -1288 -19085 -1191 -18988
rect -1191 -19085 -1186 -18988
rect -1293 -19090 -1186 -19085
rect -5025 -19801 -4911 -19796
rect -5025 -19905 -5020 -19801
rect -5020 -19905 -4916 -19801
rect -4916 -19905 -4911 -19801
rect -5025 -19910 -4911 -19905
rect -4009 -19797 -3902 -19792
rect -4009 -19894 -4004 -19797
rect -4004 -19894 -3907 -19797
rect -3907 -19894 -3902 -19797
rect -4009 -19899 -3902 -19894
rect -2309 -19796 -2195 -19791
rect -2309 -19900 -2304 -19796
rect -2304 -19900 -2200 -19796
rect -2200 -19900 -2195 -19796
rect -2309 -19905 -2195 -19900
rect -1293 -19807 -1186 -19802
rect -1293 -19904 -1288 -19807
rect -1288 -19904 -1191 -19807
rect -1191 -19904 -1186 -19807
rect -1293 -19909 -1186 -19904
rect -2309 -20422 -2195 -20418
rect -2309 -20528 -2305 -20422
rect -2305 -20528 -2199 -20422
rect -2199 -20528 -2195 -20422
rect -2309 -20532 -2195 -20528
rect -1293 -20440 -1186 -20435
rect -1293 -20537 -1288 -20440
rect -1288 -20537 -1191 -20440
rect -1191 -20537 -1186 -20440
rect -1293 -20542 -1186 -20537
rect -5025 -20620 -4911 -20615
rect -5025 -20724 -5020 -20620
rect -5020 -20724 -4916 -20620
rect -4916 -20724 -4911 -20620
rect -5025 -20729 -4911 -20724
rect -4009 -20616 -3902 -20611
rect -4009 -20713 -4004 -20616
rect -4004 -20713 -3907 -20616
rect -3907 -20713 -3902 -20616
rect -4009 -20718 -3902 -20713
rect 11889 -13417 12141 -13412
rect 11889 -13659 11894 -13417
rect 11894 -13659 12136 -13417
rect 12136 -13659 12141 -13417
rect 11889 -13664 12141 -13659
rect 6165 -14863 6231 -14858
rect 6165 -14919 6170 -14863
rect 6170 -14919 6226 -14863
rect 6226 -14919 6231 -14863
rect 6165 -14924 6231 -14919
rect 6605 -14854 6671 -14849
rect 6605 -14910 6610 -14854
rect 6610 -14910 6666 -14854
rect 6666 -14910 6671 -14854
rect 6605 -14915 6671 -14910
rect 12193 -15243 12425 -15238
rect 12193 -15465 12198 -15243
rect 12198 -15465 12420 -15243
rect 12420 -15465 12425 -15243
rect 12193 -15470 12425 -15465
rect 7222 -16397 7410 -16392
rect 7222 -16575 7227 -16397
rect 7227 -16575 7405 -16397
rect 7405 -16575 7410 -16397
rect 7222 -16580 7410 -16575
rect 8157 -16397 8345 -16392
rect 8157 -16575 8162 -16397
rect 8162 -16575 8340 -16397
rect 8340 -16575 8345 -16397
rect 8157 -16580 8345 -16575
rect 9093 -16397 9281 -16392
rect 9093 -16575 9098 -16397
rect 9098 -16575 9276 -16397
rect 9276 -16575 9281 -16397
rect 9093 -16580 9281 -16575
rect 10024 -16397 10211 -16392
rect 10024 -16574 10029 -16397
rect 10029 -16574 10206 -16397
rect 10206 -16574 10211 -16397
rect 10024 -16579 10211 -16574
rect 10951 -16397 11139 -16392
rect 10951 -16575 10956 -16397
rect 10956 -16575 11134 -16397
rect 11134 -16575 11139 -16397
rect 10951 -16580 11139 -16575
rect 12228 -16908 12357 -16903
rect 12228 -17027 12233 -16908
rect 12233 -17027 12352 -16908
rect 12352 -17027 12357 -16908
rect 12228 -17032 12357 -17027
rect 12955 -16949 13084 -16944
rect 12955 -17068 12960 -16949
rect 12960 -17068 13079 -16949
rect 13079 -17068 13084 -16949
rect 12955 -17073 13084 -17068
rect 16280 -16737 16548 -16732
rect 16280 -16995 16285 -16737
rect 16285 -16995 16543 -16737
rect 16543 -16995 16548 -16737
rect 16280 -17000 16548 -16995
rect 5727 -19410 5793 -19405
rect 5727 -19466 5732 -19410
rect 5732 -19466 5788 -19410
rect 5788 -19466 5793 -19410
rect 5727 -19471 5793 -19466
rect 11889 -17945 12141 -17940
rect 11889 -18187 11894 -17945
rect 11894 -18187 12136 -17945
rect 12136 -18187 12141 -17945
rect 11889 -18192 12141 -18187
rect 17521 -18021 17664 -18016
rect 17521 -18154 17526 -18021
rect 17526 -18154 17659 -18021
rect 17659 -18154 17664 -18021
rect 17521 -18159 17664 -18154
rect 6165 -19391 6231 -19386
rect 6165 -19447 6170 -19391
rect 6170 -19447 6226 -19391
rect 6226 -19447 6231 -19391
rect 6165 -19452 6231 -19447
rect 15546 -18514 15700 -18509
rect 15546 -18658 15551 -18514
rect 15551 -18658 15695 -18514
rect 15695 -18658 15700 -18514
rect 15546 -18663 15700 -18658
rect 17972 -18869 18053 -18864
rect 17972 -18940 17977 -18869
rect 17977 -18940 18048 -18869
rect 18048 -18940 18053 -18869
rect 17972 -18945 18053 -18940
rect 6605 -19382 6671 -19377
rect 6605 -19438 6610 -19382
rect 6610 -19438 6666 -19382
rect 6666 -19438 6671 -19382
rect 6605 -19443 6671 -19438
rect 12193 -19771 12425 -19766
rect 12193 -19993 12198 -19771
rect 12198 -19993 12420 -19771
rect 12420 -19993 12425 -19771
rect 12193 -19998 12425 -19993
rect 16226 -20177 16485 -20172
rect 16226 -20436 16231 -20177
rect 16231 -20436 16480 -20177
rect 16480 -20436 16485 -20177
rect 16226 -20441 16485 -20436
rect 7222 -20925 7410 -20920
rect 7222 -21103 7227 -20925
rect 7227 -21103 7405 -20925
rect 7405 -21103 7410 -20925
rect 7222 -21108 7410 -21103
rect 8157 -20925 8345 -20920
rect 8157 -21103 8162 -20925
rect 8162 -21103 8340 -20925
rect 8340 -21103 8345 -20925
rect 8157 -21108 8345 -21103
rect 9093 -20925 9281 -20920
rect 9093 -21103 9098 -20925
rect 9098 -21103 9276 -20925
rect 9276 -21103 9281 -20925
rect 9093 -21108 9281 -21103
rect 10024 -20925 10211 -20920
rect 10024 -21102 10029 -20925
rect 10029 -21102 10206 -20925
rect 10206 -21102 10211 -20925
rect 10024 -21107 10211 -21102
rect 10951 -20925 11139 -20920
rect 10951 -21103 10956 -20925
rect 10956 -21103 11134 -20925
rect 11134 -21103 11139 -20925
rect 10951 -21108 11139 -21103
rect 12228 -21436 12357 -21431
rect 12228 -21555 12233 -21436
rect 12233 -21555 12352 -21436
rect 12352 -21555 12357 -21436
rect 12228 -21560 12357 -21555
rect 12955 -21477 13084 -21472
rect 12955 -21596 12960 -21477
rect 12960 -21596 13079 -21477
rect 13079 -21596 13084 -21477
rect 12955 -21601 13084 -21596
rect 5727 -23938 5793 -23933
rect 5727 -23994 5732 -23938
rect 5732 -23994 5788 -23938
rect 5788 -23994 5793 -23938
rect 5727 -23999 5793 -23994
rect 11889 -22473 12141 -22468
rect 11889 -22715 11894 -22473
rect 11894 -22715 12136 -22473
rect 12136 -22715 12141 -22473
rect 11889 -22720 12141 -22715
rect 6165 -23919 6231 -23914
rect 6165 -23975 6170 -23919
rect 6170 -23975 6226 -23919
rect 6226 -23975 6231 -23919
rect 6165 -23980 6231 -23975
rect 6605 -23910 6671 -23905
rect 6605 -23966 6610 -23910
rect 6610 -23966 6666 -23910
rect 6666 -23966 6671 -23910
rect 6605 -23971 6671 -23966
rect 12193 -24299 12425 -24294
rect 12193 -24521 12198 -24299
rect 12198 -24521 12420 -24299
rect 12420 -24521 12425 -24299
rect 12193 -24526 12425 -24521
rect 7222 -25453 7410 -25448
rect 7222 -25631 7227 -25453
rect 7227 -25631 7405 -25453
rect 7405 -25631 7410 -25453
rect 7222 -25636 7410 -25631
rect 8157 -25453 8345 -25448
rect 8157 -25631 8162 -25453
rect 8162 -25631 8340 -25453
rect 8340 -25631 8345 -25453
rect 8157 -25636 8345 -25631
rect 9093 -25453 9281 -25448
rect 9093 -25631 9098 -25453
rect 9098 -25631 9276 -25453
rect 9276 -25631 9281 -25453
rect 9093 -25636 9281 -25631
rect 10024 -25453 10211 -25448
rect 10024 -25630 10029 -25453
rect 10029 -25630 10206 -25453
rect 10206 -25630 10211 -25453
rect 10024 -25635 10211 -25630
rect 10951 -25453 11139 -25448
rect 10951 -25631 10956 -25453
rect 10956 -25631 11134 -25453
rect 11134 -25631 11139 -25453
rect 10951 -25636 11139 -25631
rect 12228 -25964 12357 -25959
rect 12228 -26083 12233 -25964
rect 12233 -26083 12352 -25964
rect 12352 -26083 12357 -25964
rect 12228 -26088 12357 -26083
rect 12955 -26005 13084 -26000
rect 12955 -26124 12960 -26005
rect 12960 -26124 13079 -26005
rect 13079 -26124 13084 -26005
rect 12955 -26129 13084 -26124
rect 5727 -28466 5793 -28461
rect 5727 -28522 5732 -28466
rect 5732 -28522 5788 -28466
rect 5788 -28522 5793 -28466
rect 5727 -28527 5793 -28522
rect 11889 -27001 12141 -26996
rect 11889 -27243 11894 -27001
rect 11894 -27243 12136 -27001
rect 12136 -27243 12141 -27001
rect 11889 -27248 12141 -27243
rect 6165 -28447 6231 -28442
rect 6165 -28503 6170 -28447
rect 6170 -28503 6226 -28447
rect 6226 -28503 6231 -28447
rect 6165 -28508 6231 -28503
rect 6605 -28438 6671 -28433
rect 6605 -28494 6610 -28438
rect 6610 -28494 6666 -28438
rect 6666 -28494 6671 -28438
rect 6605 -28499 6671 -28494
rect 12193 -28827 12425 -28822
rect 12193 -29049 12198 -28827
rect 12198 -29049 12420 -28827
rect 12420 -29049 12425 -28827
rect 12193 -29054 12425 -29049
rect 7222 -29981 7410 -29976
rect 7222 -30159 7227 -29981
rect 7227 -30159 7405 -29981
rect 7405 -30159 7410 -29981
rect 7222 -30164 7410 -30159
rect 8157 -29981 8345 -29976
rect 8157 -30159 8162 -29981
rect 8162 -30159 8340 -29981
rect 8340 -30159 8345 -29981
rect 8157 -30164 8345 -30159
rect 9093 -29981 9281 -29976
rect 9093 -30159 9098 -29981
rect 9098 -30159 9276 -29981
rect 9276 -30159 9281 -29981
rect 9093 -30164 9281 -30159
rect 10024 -29981 10211 -29976
rect 10024 -30158 10029 -29981
rect 10029 -30158 10206 -29981
rect 10206 -30158 10211 -29981
rect 10024 -30163 10211 -30158
rect 10951 -29981 11139 -29976
rect 10951 -30159 10956 -29981
rect 10956 -30159 11134 -29981
rect 11134 -30159 11139 -29981
rect 10951 -30164 11139 -30159
rect 12228 -30492 12357 -30487
rect 12228 -30611 12233 -30492
rect 12233 -30611 12352 -30492
rect 12352 -30611 12357 -30492
rect 12228 -30616 12357 -30611
rect 12955 -30533 13084 -30528
rect 12955 -30652 12960 -30533
rect 12960 -30652 13079 -30533
rect 13079 -30652 13084 -30533
rect 12955 -30657 13084 -30652
rect 11889 -31529 12141 -31524
rect 11889 -31771 11894 -31529
rect 11894 -31771 12136 -31529
rect 12136 -31771 12141 -31529
rect 11889 -31776 12141 -31771
rect 5727 -32994 5793 -32989
rect 5727 -33050 5732 -32994
rect 5732 -33050 5788 -32994
rect 5788 -33050 5793 -32994
rect 5727 -33055 5793 -33050
rect 6165 -32975 6231 -32970
rect 6165 -33031 6170 -32975
rect 6170 -33031 6226 -32975
rect 6226 -33031 6231 -32975
rect 6165 -33036 6231 -33031
rect 6605 -32966 6671 -32961
rect 6605 -33022 6610 -32966
rect 6610 -33022 6666 -32966
rect 6666 -33022 6671 -32966
rect 6605 -33027 6671 -33022
rect 12193 -33355 12425 -33350
rect 12193 -33577 12198 -33355
rect 12198 -33577 12420 -33355
rect 12420 -33577 12425 -33355
rect 12193 -33582 12425 -33577
rect 7222 -34509 7410 -34504
rect 7222 -34687 7227 -34509
rect 7227 -34687 7405 -34509
rect 7405 -34687 7410 -34509
rect 7222 -34692 7410 -34687
rect 8157 -34509 8345 -34504
rect 8157 -34687 8162 -34509
rect 8162 -34687 8340 -34509
rect 8340 -34687 8345 -34509
rect 8157 -34692 8345 -34687
rect 9093 -34509 9281 -34504
rect 9093 -34687 9098 -34509
rect 9098 -34687 9276 -34509
rect 9276 -34687 9281 -34509
rect 9093 -34692 9281 -34687
rect 10024 -34509 10211 -34504
rect 10024 -34686 10029 -34509
rect 10029 -34686 10206 -34509
rect 10206 -34686 10211 -34509
rect 10024 -34691 10211 -34686
rect 10951 -34509 11139 -34504
rect 10951 -34687 10956 -34509
rect 10956 -34687 11134 -34509
rect 11134 -34687 11139 -34509
rect 10951 -34692 11139 -34687
rect 12228 -35020 12357 -35015
rect 12228 -35139 12233 -35020
rect 12233 -35139 12352 -35020
rect 12352 -35139 12357 -35020
rect 12228 -35144 12357 -35139
rect 12955 -35061 13084 -35056
rect 12955 -35180 12960 -35061
rect 12960 -35180 13079 -35061
rect 13079 -35180 13084 -35061
rect 12955 -35185 13084 -35180
rect 11889 -36057 12141 -36052
rect 11889 -36299 11894 -36057
rect 11894 -36299 12136 -36057
rect 12136 -36299 12141 -36057
rect 11889 -36304 12141 -36299
rect 12544 -35955 12651 -35950
rect 12544 -36052 12549 -35955
rect 12549 -36052 12646 -35955
rect 12646 -36052 12651 -35955
rect 12544 -36057 12651 -36052
rect 13553 -35959 13667 -35954
rect 13553 -36063 13558 -35959
rect 13558 -36063 13662 -35959
rect 13662 -36063 13667 -35959
rect 13553 -36068 13667 -36063
<< metal4 >>
rect -208 6241 6474 6352
rect -208 6169 1841 6241
rect 2963 6169 3447 6241
rect 4569 6239 6474 6241
rect 4569 6169 5151 6239
rect -208 6167 5151 6169
rect 6273 6167 6474 6239
rect -208 6040 6474 6167
rect -208 4679 104 6040
rect -24310 4517 375 4679
rect -24310 4445 -24000 4517
rect -22878 4445 -20709 4517
rect -19587 4445 -17418 4517
rect -16296 4445 -14127 4517
rect -13005 4445 -10836 4517
rect -9714 4445 -7546 4517
rect -6424 4445 -4255 4517
rect -3133 4445 -964 4517
rect 158 4445 375 4517
rect 6162 4462 6474 6040
rect -24310 4367 375 4445
rect -24225 2775 -24099 4367
rect -20934 2775 -20808 4367
rect -17643 2775 -17517 4367
rect -14352 2775 -14226 4367
rect -11061 2775 -10935 4367
rect -7771 2775 -7645 4367
rect -4480 2775 -4354 4367
rect -1189 2775 -1063 4367
rect 5006 4200 6474 4462
rect 5006 3668 6834 4200
rect -24225 2761 -22550 2775
rect -20934 2761 -19259 2775
rect -17643 2761 -15968 2775
rect -14352 2761 -12677 2775
rect -11061 2761 -9386 2775
rect -7771 2761 -6096 2775
rect -4480 2761 -2805 2775
rect -1189 2761 486 2775
rect -24716 2733 -21947 2761
rect -24716 2661 -24670 2733
rect -23548 2661 -23111 2733
rect -21989 2661 -21947 2733
rect -24716 2649 -21947 2661
rect -24716 2635 -23506 2649
rect -23404 1010 -23226 2649
rect -23157 2635 -21947 2649
rect -21425 2733 -18656 2761
rect -21425 2661 -21379 2733
rect -20257 2661 -19820 2733
rect -18698 2661 -18656 2733
rect -21425 2649 -18656 2661
rect -21425 2635 -20215 2649
rect -20113 1010 -19935 2649
rect -19866 2635 -18656 2649
rect -18134 2733 -15365 2761
rect -18134 2661 -18088 2733
rect -16966 2661 -16529 2733
rect -15407 2661 -15365 2733
rect -18134 2649 -15365 2661
rect -18134 2635 -16924 2649
rect -16822 1010 -16644 2649
rect -16575 2635 -15365 2649
rect -14843 2733 -12074 2761
rect -14843 2661 -14797 2733
rect -13675 2661 -13238 2733
rect -12116 2661 -12074 2733
rect -14843 2649 -12074 2661
rect -14843 2635 -13633 2649
rect -13531 1010 -13353 2649
rect -13284 2635 -12074 2649
rect -11552 2733 -8783 2761
rect -11552 2661 -11506 2733
rect -10384 2661 -9947 2733
rect -8825 2661 -8783 2733
rect -11552 2649 -8783 2661
rect -11552 2635 -10342 2649
rect -10240 1010 -10062 2649
rect -9993 2635 -8783 2649
rect -8262 2733 -5493 2761
rect -8262 2661 -8216 2733
rect -7094 2661 -6657 2733
rect -5535 2661 -5493 2733
rect -8262 2649 -5493 2661
rect -8262 2635 -7052 2649
rect -6950 1010 -6772 2649
rect -6703 2635 -5493 2649
rect -4971 2733 -2202 2761
rect -4971 2661 -4925 2733
rect -3803 2661 -3366 2733
rect -2244 2661 -2202 2733
rect -4971 2649 -2202 2661
rect -4971 2635 -3761 2649
rect -3659 1010 -3481 2649
rect -3412 2635 -2202 2649
rect -1680 2733 1089 2761
rect -1680 2661 -1634 2733
rect -512 2661 -75 2733
rect 1047 2661 1089 2733
rect -1680 2649 1089 2661
rect -1680 2635 -470 2649
rect -368 1010 -190 2649
rect -121 2635 1089 2649
rect -24421 1001 -22141 1010
rect -24421 929 -24412 1001
rect -24156 929 -23123 1001
rect -22867 929 -22406 1001
rect -22150 929 -22141 1001
rect -24421 920 -22141 929
rect -21130 1001 -18850 1010
rect -21130 929 -21121 1001
rect -20865 929 -19832 1001
rect -19576 929 -19115 1001
rect -18859 929 -18850 1001
rect -21130 920 -18850 929
rect -17839 1001 -15559 1010
rect -17839 929 -17830 1001
rect -17574 929 -16541 1001
rect -16285 929 -15824 1001
rect -15568 929 -15559 1001
rect -17839 920 -15559 929
rect -14548 1001 -12268 1010
rect -14548 929 -14539 1001
rect -14283 929 -13250 1001
rect -12994 929 -12533 1001
rect -12277 929 -12268 1001
rect -14548 920 -12268 929
rect -11257 1001 -8977 1010
rect -11257 929 -11248 1001
rect -10992 929 -9959 1001
rect -9703 929 -9242 1001
rect -8986 929 -8977 1001
rect -11257 920 -8977 929
rect -7967 1001 -5687 1010
rect -7967 929 -7958 1001
rect -7702 929 -6669 1001
rect -6413 929 -5952 1001
rect -5696 929 -5687 1001
rect -7967 920 -5687 929
rect -4676 1001 -2396 1010
rect -4676 929 -4667 1001
rect -4411 929 -3378 1001
rect -3122 929 -2661 1001
rect -2405 929 -2396 1001
rect -4676 920 -2396 929
rect -1385 1001 895 1010
rect -1385 929 -1376 1001
rect -1120 929 -87 1001
rect 169 929 630 1001
rect 886 929 895 1001
rect -1385 920 895 929
rect -24345 203 -24336 268
rect -24001 203 -23992 268
rect -24345 194 -23992 203
rect -21054 203 -21045 268
rect -20710 203 -20701 268
rect -21054 194 -20701 203
rect -20361 -2089 -20271 920
rect -17763 203 -17754 268
rect -17419 203 -17410 268
rect -17763 194 -17410 203
rect -14472 203 -14463 268
rect -14128 203 -14119 268
rect -14472 194 -14119 203
rect -11181 203 -11172 268
rect -10837 203 -10828 268
rect -11181 194 -10828 203
rect -7891 203 -7882 268
rect -7547 203 -7538 268
rect -7891 194 -7538 203
rect -4600 203 -4591 268
rect -4256 203 -4247 268
rect -4600 194 -4247 203
rect -1309 203 -1300 268
rect -965 203 -956 268
rect -1309 194 -956 203
rect 5006 -428 5318 3668
rect 5581 3366 6823 3399
rect 5581 3357 6502 3366
rect 5581 3338 6062 3357
rect 5581 3066 5624 3338
rect 5896 3085 6062 3338
rect 6334 3094 6502 3357
rect 6774 3094 6823 3366
rect 6334 3085 6823 3094
rect 5896 3066 6823 3085
rect 5581 3032 6823 3066
rect 12121 2970 12450 3036
rect 12121 2874 13912 2970
rect 12121 2856 12193 2874
rect 11317 2642 12193 2856
rect 12425 2642 13912 2874
rect 11317 2634 13912 2642
rect 11317 2527 12450 2634
rect 7156 1763 11207 1787
rect 7156 1762 9982 1763
rect 7156 1490 7180 1762
rect 7452 1490 8115 1762
rect 8387 1490 9051 1762
rect 9323 1491 9982 1762
rect 10254 1762 11207 1763
rect 10254 1491 10909 1762
rect 9323 1490 10909 1491
rect 11181 1490 11207 1762
rect 7156 1466 11207 1490
rect 11317 834 11646 2527
rect 12414 1296 12821 1408
rect 12128 1292 12821 1296
rect 12128 1281 13042 1292
rect 12128 1009 12157 1281
rect 12429 1266 13042 1281
rect 12429 1240 13186 1266
rect 12429 1009 12884 1240
rect 12128 979 12884 1009
rect 12467 968 12884 979
rect 13156 968 13186 1240
rect 11317 505 11889 834
rect 12467 820 13186 968
rect 12796 787 13186 820
rect 11560 241 11889 505
rect 11560 208 12159 241
rect 13576 208 13912 2634
rect 11560 172 13912 208
rect 11560 -80 11889 172
rect 12141 -80 13912 172
rect 11560 -128 13912 -80
rect 5006 -740 6890 -428
rect 5006 -1450 5318 -740
rect 5581 -1162 6823 -1129
rect 5581 -1171 6502 -1162
rect 5581 -1190 6062 -1171
rect 5006 -1560 5518 -1450
rect 5581 -1462 5624 -1190
rect 5896 -1443 6062 -1190
rect 6334 -1434 6502 -1171
rect 6774 -1434 6823 -1162
rect 6334 -1443 6823 -1434
rect 5896 -1462 6823 -1443
rect 12098 -1450 12410 -128
rect 5581 -1496 6823 -1462
rect 6892 -1492 12410 -1450
rect 6892 -1538 12450 -1492
rect 6892 -1560 12502 -1538
rect 5006 -1654 12502 -1560
rect 5006 -1762 12193 -1654
rect -24449 -2090 -17781 -2089
rect -24449 -2225 -17354 -2090
rect -24449 -2304 -23605 -2225
rect -23436 -2304 -21585 -2225
rect -21416 -2304 -19844 -2225
rect -19675 -2304 -18065 -2225
rect -17896 -2304 -17354 -2225
rect -24449 -2327 -17354 -2304
rect -24449 -2467 -24410 -2327
rect -23856 -2467 -22373 -2327
rect -21819 -2467 -20643 -2327
rect -20089 -2467 -18883 -2327
rect -18329 -2467 -17354 -2327
rect -24449 -2506 -17354 -2467
rect -24248 -2878 -21372 -2785
rect -24248 -2883 -23601 -2878
rect -23452 -2883 -21581 -2878
rect -24248 -2983 -23987 -2883
rect -21717 -2974 -21581 -2883
rect -21432 -2974 -21372 -2878
rect -24248 -3057 -24184 -2983
rect -24248 -3191 -23987 -3057
rect -21717 -3191 -21372 -2974
rect -24248 -3249 -21372 -3191
rect -21095 -3707 -20762 -2506
rect -17801 -2507 -17354 -2506
rect -20485 -2878 -17851 -2819
rect -20485 -2914 -19840 -2878
rect -19691 -2914 -18061 -2878
rect -20485 -2983 -20247 -2914
rect -17912 -2974 -17851 -2878
rect -20485 -3057 -20417 -2983
rect -20485 -3222 -20247 -3057
rect -17977 -3222 -17851 -2974
rect -20485 -3297 -17851 -3222
rect -17690 -3707 -17357 -2507
rect -21628 -3732 -7975 -3707
rect -24399 -3827 -7975 -3732
rect -24399 -3899 -20603 -3827
rect -19481 -3899 -19044 -3827
rect -17922 -3899 -17312 -3827
rect -16190 -3899 -15753 -3827
rect -14631 -3899 -14021 -3827
rect -12899 -3899 -12462 -3827
rect -11340 -3899 -10730 -3827
rect -9608 -3899 -9171 -3827
rect -8049 -3899 -7975 -3827
rect -24399 -3926 -7975 -3899
rect -24399 -4037 -21594 -3926
rect -24399 -4116 -23561 -4037
rect -23392 -4116 -21823 -4037
rect -21654 -4116 -21594 -4037
rect -24399 -4139 -21594 -4116
rect -24399 -4279 -24359 -4139
rect -23805 -4279 -22623 -4139
rect -22069 -4279 -21594 -4139
rect -24399 -4319 -21594 -4279
rect -24210 -4612 -21613 -4527
rect -24210 -4795 -24007 -4612
rect -21737 -4690 -21613 -4612
rect -21670 -4786 -21613 -4690
rect -24210 -4869 -24133 -4795
rect -24210 -4920 -24007 -4869
rect -21737 -4920 -21613 -4786
rect -24210 -4984 -21613 -4920
rect -24403 -5329 -21636 -5306
rect -24403 -5408 -23563 -5329
rect -23394 -5408 -21829 -5329
rect -21660 -5408 -21636 -5329
rect -24403 -5431 -21636 -5408
rect -24403 -5547 -24359 -5431
rect -24406 -5571 -24359 -5547
rect -23805 -5571 -22623 -5431
rect -22069 -5547 -21636 -5431
rect -21095 -5547 -20762 -3926
rect -19337 -5547 -19159 -3926
rect -17690 -5547 -17357 -3926
rect -16046 -5547 -15868 -3926
rect -14421 -5547 -14088 -3926
rect -12755 -5547 -12577 -3926
rect -11116 -5547 -10783 -3926
rect -9464 -5547 -9286 -3926
rect 5006 -4832 5318 -1762
rect 11317 -1886 12193 -1762
rect 12425 -1730 12502 -1654
rect 13576 -1730 13912 -128
rect 12425 -1886 13912 -1730
rect 11317 -2001 13912 -1886
rect 7156 -2765 11207 -2741
rect 7156 -2766 9982 -2765
rect 7156 -3038 7180 -2766
rect 7452 -3038 8115 -2766
rect 8387 -3038 9051 -2766
rect 9323 -3037 9982 -2766
rect 10254 -2766 11207 -2765
rect 10254 -3037 10909 -2766
rect 9323 -3038 10909 -3037
rect 11181 -3038 11207 -2766
rect 7156 -3062 11207 -3038
rect 11317 -3694 11646 -2001
rect 12098 -2030 13912 -2001
rect 12166 -2066 13912 -2030
rect 12414 -3232 12821 -3120
rect 12128 -3236 12821 -3232
rect 12128 -3247 13042 -3236
rect 12128 -3519 12157 -3247
rect 12429 -3262 13042 -3247
rect 12429 -3288 13186 -3262
rect 12429 -3519 12884 -3288
rect 12128 -3549 12884 -3519
rect 12467 -3560 12884 -3549
rect 13156 -3560 13186 -3288
rect 11317 -4023 11889 -3694
rect 12467 -3708 13186 -3560
rect 12796 -3741 13186 -3708
rect 11560 -4287 11889 -4023
rect 11560 -4328 12159 -4287
rect 13576 -4328 13912 -2066
rect 11560 -4356 13912 -4328
rect 11560 -4608 11889 -4356
rect 12141 -4608 13912 -4356
rect 11560 -4656 13912 -4608
rect 11866 -4664 13912 -4656
rect 5006 -5144 6820 -4832
rect -22069 -5559 -8201 -5547
rect -22069 -5571 -20345 -5559
rect -24406 -5631 -20345 -5571
rect -20089 -5631 -19056 -5559
rect -18800 -5631 -18339 -5559
rect -18083 -5631 -17054 -5559
rect -16798 -5631 -15765 -5559
rect -15509 -5631 -15048 -5559
rect -14792 -5631 -13763 -5559
rect -13507 -5631 -12474 -5559
rect -12218 -5631 -11757 -5559
rect -11501 -5631 -10472 -5559
rect -10216 -5631 -9183 -5559
rect -8927 -5631 -8466 -5559
rect -8210 -5631 -8201 -5559
rect -24406 -5696 -8201 -5631
rect -24207 -5976 -21610 -5892
rect -24207 -6087 -24008 -5976
rect -21738 -5982 -21610 -5976
rect -21676 -6078 -21610 -5982
rect -24207 -6161 -24133 -6087
rect -24207 -6284 -24008 -6161
rect -21738 -6284 -21610 -6078
rect -24207 -6349 -21610 -6284
rect -21095 -7005 -20762 -5696
rect -20278 -6357 -20269 -6292
rect -19934 -6357 -19925 -6292
rect -20278 -6366 -19925 -6357
rect -17690 -7005 -17357 -5696
rect -16987 -6357 -16978 -6292
rect -16643 -6357 -16634 -6292
rect -16987 -6366 -16634 -6357
rect -14421 -7005 -14088 -5696
rect -13696 -6357 -13687 -6292
rect -13352 -6357 -13343 -6292
rect -13696 -6366 -13343 -6357
rect -11116 -7005 -10783 -5696
rect -10405 -6357 -10396 -6292
rect -10061 -6357 -10052 -6292
rect -10405 -6366 -10052 -6357
rect -24403 -7092 -7993 -7005
rect -24403 -7164 -20603 -7092
rect -19481 -7164 -19044 -7092
rect -17922 -7164 -17312 -7092
rect -16190 -7164 -15753 -7092
rect -14631 -7164 -14021 -7092
rect -12899 -7164 -12462 -7092
rect -11340 -7164 -10730 -7092
rect -9608 -7164 -9171 -7092
rect -8049 -7164 -7993 -7092
rect -24403 -7262 -7993 -7164
rect -24403 -7302 -21632 -7262
rect -24403 -7381 -23562 -7302
rect -23393 -7381 -21827 -7302
rect -21658 -7381 -21632 -7302
rect -24403 -7404 -21632 -7381
rect -24403 -7544 -24359 -7404
rect -23805 -7544 -22622 -7404
rect -22068 -7544 -21632 -7404
rect -24403 -7583 -21632 -7544
rect -24207 -7870 -21610 -7803
rect -24207 -8060 -24046 -7870
rect -21776 -7955 -21610 -7870
rect -21674 -8051 -21610 -7955
rect -24207 -8134 -24133 -8060
rect -24207 -8178 -24046 -8134
rect -21776 -8178 -21610 -8051
rect -24207 -8260 -21610 -8178
rect -24398 -8594 -21631 -8572
rect -24398 -8673 -23560 -8594
rect -23391 -8673 -21823 -8594
rect -21654 -8673 -21631 -8594
rect -24398 -8696 -21631 -8673
rect -24398 -8836 -24359 -8696
rect -23805 -8836 -22623 -8696
rect -22069 -8815 -21631 -8696
rect -21095 -8815 -20762 -7262
rect -19337 -8815 -19159 -7262
rect -17690 -8815 -17357 -7262
rect -16046 -8815 -15868 -7262
rect -14421 -8815 -14088 -7262
rect -12755 -8815 -12577 -7262
rect -11116 -8815 -10783 -7262
rect -9464 -8815 -9286 -7262
rect -22069 -8824 -8193 -8815
rect -22069 -8836 -20345 -8824
rect -24398 -8896 -20345 -8836
rect -20089 -8896 -19056 -8824
rect -18800 -8896 -18339 -8824
rect -18083 -8896 -17054 -8824
rect -16798 -8896 -15765 -8824
rect -15509 -8896 -15048 -8824
rect -14792 -8896 -13763 -8824
rect -13507 -8896 -12474 -8824
rect -12218 -8896 -11757 -8824
rect -11501 -8896 -10472 -8824
rect -10216 -8896 -9183 -8824
rect -8927 -8896 -8466 -8824
rect -8210 -8896 -8193 -8824
rect -24398 -8964 -8193 -8896
rect -24200 -9247 -21603 -9178
rect -24200 -9248 -23556 -9247
rect -23407 -9248 -21819 -9247
rect -24200 -9352 -24060 -9248
rect -21670 -9343 -21603 -9247
rect -24200 -9426 -24133 -9352
rect -24200 -9556 -24060 -9426
rect -21790 -9556 -21603 -9343
rect -24200 -9635 -21603 -9556
rect -24400 -10274 -21629 -10271
rect -21095 -10274 -20762 -8964
rect -20278 -9622 -20269 -9557
rect -19934 -9622 -19925 -9557
rect -20278 -9631 -19925 -9622
rect -17690 -10274 -17357 -8964
rect -16987 -9622 -16978 -9557
rect -16643 -9622 -16634 -9557
rect -16987 -9631 -16634 -9622
rect -14421 -10274 -14088 -8964
rect -13696 -9622 -13687 -9557
rect -13352 -9622 -13343 -9557
rect -13696 -9631 -13343 -9622
rect -11116 -10274 -10783 -8964
rect -10405 -9622 -10396 -9557
rect 5006 -9450 5318 -5144
rect 5581 -5590 6823 -5557
rect 5581 -5599 6502 -5590
rect 5581 -5618 6062 -5599
rect 5581 -5890 5624 -5618
rect 5896 -5871 6062 -5618
rect 6334 -5862 6502 -5599
rect 6774 -5862 6823 -5590
rect 6334 -5871 6823 -5862
rect 5896 -5890 6823 -5871
rect 5581 -5924 6823 -5890
rect 12121 -6000 12450 -5920
rect 13576 -6000 13912 -4664
rect 12028 -6082 13912 -6000
rect 12028 -6100 12193 -6082
rect 11317 -6314 12193 -6100
rect 12425 -6314 13912 -6082
rect 11317 -6336 13912 -6314
rect 11317 -6429 12450 -6336
rect 7156 -7193 11207 -7169
rect 7156 -7194 9982 -7193
rect 7156 -7466 7180 -7194
rect 7452 -7466 8115 -7194
rect 8387 -7466 9051 -7194
rect 9323 -7465 9982 -7194
rect 10254 -7194 11207 -7193
rect 10254 -7465 10909 -7194
rect 9323 -7466 10909 -7465
rect 11181 -7466 11207 -7194
rect 7156 -7490 11207 -7466
rect 11317 -8122 11646 -6429
rect 12414 -7660 12821 -7548
rect 12128 -7664 12821 -7660
rect 12128 -7675 13042 -7664
rect 12128 -7947 12157 -7675
rect 12429 -7690 13042 -7675
rect 12429 -7716 13186 -7690
rect 12429 -7947 12884 -7716
rect 12128 -7977 12884 -7947
rect 12467 -7988 12884 -7977
rect 13156 -7988 13186 -7716
rect 11317 -8451 11889 -8122
rect 12467 -8136 13186 -7988
rect 12796 -8169 13186 -8136
rect 11560 -8715 11889 -8451
rect 11560 -8750 12159 -8715
rect 13576 -8750 13912 -6336
rect 11560 -8784 13912 -8750
rect 11560 -9036 11889 -8784
rect 12141 -9036 13912 -8784
rect 11560 -9084 13912 -9036
rect 11866 -9086 13912 -9084
rect -10061 -9622 -10052 -9557
rect -10405 -9631 -10052 -9622
rect 5006 -9762 7020 -9450
rect -24400 -10356 -8005 -10274
rect -24400 -10428 -20603 -10356
rect -19481 -10428 -19044 -10356
rect -17922 -10428 -17312 -10356
rect -16190 -10428 -15753 -10356
rect -14631 -10428 -14021 -10356
rect -12899 -10428 -12462 -10356
rect -11340 -10428 -10730 -10356
rect -9608 -10428 -9171 -10356
rect -8049 -10428 -8005 -10356
rect -24400 -10531 -8005 -10428
rect -24400 -10566 -21629 -10531
rect -24400 -10645 -23560 -10566
rect -23391 -10645 -21827 -10566
rect -21658 -10645 -21629 -10566
rect -24400 -10668 -21629 -10645
rect -24400 -10808 -24359 -10668
rect -23805 -10808 -22622 -10668
rect -22068 -10808 -21629 -10668
rect -24400 -10849 -21629 -10808
rect -24207 -11202 -21610 -11138
rect -24207 -11324 -24018 -11202
rect -21748 -11219 -21610 -11202
rect -21674 -11315 -21610 -11219
rect -24207 -11398 -24133 -11324
rect -24207 -11510 -24018 -11398
rect -21748 -11510 -21610 -11315
rect -24207 -11595 -21610 -11510
rect -24397 -11858 -21630 -11834
rect -24397 -11937 -23560 -11858
rect -23391 -11937 -21831 -11858
rect -21662 -11937 -21630 -11858
rect -24397 -11960 -21630 -11937
rect -24397 -12076 -24359 -11960
rect -24399 -12100 -24359 -12076
rect -23805 -12100 -22622 -11960
rect -22068 -12076 -21630 -11960
rect -21095 -12076 -20762 -10531
rect -19337 -12076 -19159 -10531
rect -17690 -12076 -17357 -10531
rect -16046 -12076 -15868 -10531
rect -14421 -12076 -14088 -10531
rect -12755 -12076 -12577 -10531
rect -11116 -12076 -10783 -10531
rect -9464 -12076 -9286 -10531
rect -22068 -12088 -8194 -12076
rect -22068 -12100 -20345 -12088
rect -24399 -12160 -20345 -12100
rect -20089 -12160 -19056 -12088
rect -18800 -12160 -18339 -12088
rect -18083 -12160 -17054 -12088
rect -16798 -12160 -15765 -12088
rect -15509 -12160 -15048 -12088
rect -14792 -12160 -13763 -12088
rect -13507 -12160 -12474 -12088
rect -12218 -12160 -11757 -12088
rect -11501 -12160 -10472 -12088
rect -10216 -12160 -9183 -12088
rect -8927 -12160 -8466 -12088
rect -8210 -12160 -8194 -12088
rect -24399 -12225 -8194 -12160
rect -24174 -12511 -21636 -12445
rect -24174 -12535 -23556 -12511
rect -23407 -12535 -21827 -12511
rect -24174 -12616 -24029 -12535
rect -21678 -12607 -21636 -12511
rect -24174 -12690 -24133 -12616
rect -24174 -12843 -24029 -12690
rect -21759 -12843 -21636 -12607
rect -24174 -12912 -21636 -12843
rect -24936 -15189 -24666 -14968
rect -24936 -15295 -24844 -15189
rect -24738 -15295 -24666 -15189
rect -24936 -15679 -24666 -15295
rect -21095 -15679 -20762 -12225
rect -20278 -12886 -20269 -12821
rect -19934 -12886 -19925 -12821
rect -20278 -12895 -19925 -12886
rect -16987 -12886 -16978 -12821
rect -16643 -12886 -16634 -12821
rect -16987 -12895 -16634 -12886
rect -13696 -12886 -13687 -12821
rect -13352 -12886 -13343 -12821
rect -13696 -12895 -13343 -12886
rect -10405 -12886 -10396 -12821
rect -10061 -12886 -10052 -12821
rect -10405 -12895 -10052 -12886
rect -5026 -13504 -2152 -13388
rect -12501 -14223 -12375 -14181
rect -18248 -15276 -17860 -15053
rect -18248 -15360 -18077 -15276
rect -17993 -15360 -17860 -15276
rect -18248 -15679 -17860 -15360
rect -12501 -15345 -12473 -14223
rect -12401 -15345 -12375 -14223
rect -5026 -14255 -4910 -13504
rect -2268 -14057 -2152 -13504
rect 5006 -13946 5318 -9762
rect 5581 -10218 6823 -10185
rect 5581 -10227 6502 -10218
rect 5581 -10246 6062 -10227
rect 5581 -10518 5624 -10246
rect 5896 -10499 6062 -10246
rect 6334 -10490 6502 -10227
rect 6774 -10490 6823 -10218
rect 6334 -10499 6823 -10490
rect 5896 -10518 6823 -10499
rect 5581 -10552 6823 -10518
rect 12121 -10584 12450 -10548
rect 13576 -10584 13912 -9086
rect 12014 -10710 13912 -10584
rect 12014 -10728 12193 -10710
rect 11317 -10942 12193 -10728
rect 12425 -10920 13912 -10710
rect 12425 -10942 12450 -10920
rect 11317 -11057 12450 -10942
rect 7156 -11821 11207 -11797
rect 7156 -11822 9982 -11821
rect 7156 -12094 7180 -11822
rect 7452 -12094 8115 -11822
rect 8387 -12094 9051 -11822
rect 9323 -12093 9982 -11822
rect 10254 -11822 11207 -11821
rect 10254 -12093 10909 -11822
rect 9323 -12094 10909 -12093
rect 11181 -12094 11207 -11822
rect 7156 -12118 11207 -12094
rect 11317 -12750 11646 -11057
rect 12414 -12288 12821 -12176
rect 12128 -12292 12821 -12288
rect 12128 -12303 13042 -12292
rect 12128 -12575 12157 -12303
rect 12429 -12318 13042 -12303
rect 12429 -12344 13186 -12318
rect 12429 -12575 12884 -12344
rect 12128 -12605 12884 -12575
rect 12467 -12616 12884 -12605
rect 13156 -12616 13186 -12344
rect 11317 -13079 11889 -12750
rect 12467 -12764 13186 -12616
rect 12796 -12797 13186 -12764
rect 11560 -13326 11889 -13079
rect 13576 -13326 13912 -10920
rect 11560 -13412 13912 -13326
rect 11560 -13664 11889 -13412
rect 12141 -13662 13912 -13412
rect 12141 -13664 12159 -13662
rect 11560 -13712 12159 -13664
rect -2310 -14058 -2152 -14057
rect -5026 -14369 -5025 -14255
rect -4911 -14369 -4910 -14255
rect -5026 -14707 -4910 -14369
rect -2310 -14172 -2309 -14058
rect -2195 -14172 -2152 -14058
rect -8554 -14870 -4910 -14707
rect -2310 -14530 -2152 -14172
rect 5006 -14258 6904 -13946
rect -24936 -15865 -17860 -15679
rect -12501 -15865 -12375 -15345
rect -8554 -15420 -8391 -14870
rect -5026 -14882 -4910 -14870
rect -5026 -14996 -5025 -14882
rect -4911 -14996 -4910 -14882
rect -8554 -15490 -8499 -15420
rect -8429 -15490 -8391 -15420
rect -8554 -15865 -8391 -15490
rect -5026 -15701 -4910 -14996
rect -2310 -14877 -2194 -14530
rect -2310 -14991 -2309 -14877
rect -2195 -14991 -2194 -14877
rect -24936 -15929 -8391 -15865
rect -24936 -15949 -8505 -15929
rect -24936 -16363 -24666 -15949
rect -24936 -16469 -24840 -16363
rect -24734 -16469 -24666 -16363
rect -24936 -17595 -24666 -16469
rect -24936 -17701 -24834 -17595
rect -24728 -17701 -24666 -17595
rect -24936 -18709 -24666 -17701
rect -21891 -18062 -21621 -15949
rect -18248 -15999 -8505 -15949
rect -8435 -15999 -8391 -15929
rect -18248 -16135 -8391 -15999
rect -5026 -15815 -5025 -15701
rect -4911 -15815 -4910 -15701
rect -18248 -16678 -17860 -16135
rect -18248 -16762 -18089 -16678
rect -18005 -16762 -17860 -16678
rect -21993 -18108 -21621 -18062
rect -21993 -18178 -21938 -18108
rect -21868 -18178 -21621 -18108
rect -24936 -18815 -24820 -18709
rect -24714 -18815 -24666 -18709
rect -24936 -19903 -24666 -18815
rect -21993 -18617 -21621 -18178
rect -18248 -18064 -17860 -16762
rect -12501 -16997 -12375 -16135
rect -8554 -16412 -8391 -16135
rect -8554 -16482 -8505 -16412
rect -8435 -16482 -8391 -16412
rect -8554 -16934 -8391 -16482
rect -5026 -16520 -4910 -15815
rect -2310 -15696 -2194 -14991
rect -2310 -15810 -2309 -15696
rect -2195 -15810 -2194 -15696
rect -5026 -16634 -5025 -16520
rect -4911 -16634 -4910 -16520
rect -12501 -17039 -12373 -16997
rect -16402 -17935 -16256 -17933
rect -16402 -17979 -16239 -17935
rect -18248 -18148 -18093 -18064
rect -18009 -18148 -17860 -18064
rect -21993 -18687 -21944 -18617
rect -21874 -18687 -21621 -18617
rect -21993 -19100 -21621 -18687
rect -21993 -19170 -21944 -19100
rect -21874 -19170 -21621 -19100
rect -21993 -19622 -21621 -19170
rect -24936 -20009 -24820 -19903
rect -24714 -20009 -24666 -19903
rect -21993 -19692 -21944 -19622
rect -21874 -19692 -21621 -19622
rect -24936 -21099 -24666 -20009
rect -21993 -20091 -21621 -19692
rect -18248 -19470 -17860 -18148
rect -16402 -18049 -16347 -17979
rect -16277 -18049 -16239 -17979
rect -18248 -19554 -18091 -19470
rect -18007 -19554 -17860 -19470
rect -16402 -18488 -16239 -18049
rect -12501 -18161 -12471 -17039
rect -12399 -18161 -12373 -17039
rect -8554 -17004 -8505 -16934
rect -8435 -17004 -8391 -16934
rect -8554 -17403 -8391 -17004
rect -8554 -17473 -8502 -17403
rect -8432 -17473 -8391 -17403
rect -12501 -18207 -12373 -18161
rect -8554 -17860 -8391 -17473
rect -5026 -17339 -4910 -16634
rect -2310 -16515 -2194 -15810
rect -2310 -16629 -2309 -16515
rect -2195 -16629 -2194 -16515
rect -5026 -17453 -5025 -17339
rect -4911 -17453 -4910 -17339
rect -8554 -17930 -8500 -17860
rect -8430 -17930 -8391 -17860
rect -16402 -18558 -16353 -18488
rect -16283 -18558 -16239 -18488
rect -16402 -18971 -16239 -18558
rect -16402 -19041 -16353 -18971
rect -16283 -19041 -16239 -18971
rect -21993 -20161 -21941 -20091
rect -21871 -20161 -21621 -20091
rect -21993 -20548 -21621 -20161
rect -18248 -20155 -17860 -19554
rect -16402 -19493 -16239 -19041
rect -16402 -19563 -16353 -19493
rect -16283 -19563 -16239 -19493
rect -16402 -19962 -16239 -19563
rect -16402 -20032 -16350 -19962
rect -16280 -20032 -16239 -19962
rect -16402 -20155 -16239 -20032
rect -12501 -19954 -12375 -18207
rect -8554 -18325 -8391 -17930
rect -8554 -18395 -8498 -18325
rect -8428 -18395 -8391 -18325
rect -8554 -18806 -8391 -18395
rect -5026 -18158 -4910 -17453
rect -2310 -17334 -2194 -16629
rect -2310 -17448 -2309 -17334
rect -2195 -17448 -2194 -17334
rect -5026 -18272 -5025 -18158
rect -4911 -18272 -4910 -18158
rect -8554 -18876 -8494 -18806
rect -8424 -18876 -8391 -18806
rect -8554 -18917 -8391 -18876
rect -5026 -18977 -4910 -18272
rect -2310 -18153 -2194 -17448
rect -2310 -18267 -2309 -18153
rect -2195 -18267 -2194 -18153
rect -5026 -19091 -5025 -18977
rect -4911 -19091 -4910 -18977
rect -5026 -19796 -4910 -19091
rect -2310 -18972 -2194 -18267
rect 5006 -18520 5318 -14258
rect 5581 -14746 6823 -14713
rect 5581 -14755 6502 -14746
rect 5581 -14774 6062 -14755
rect 5581 -15046 5624 -14774
rect 5896 -15027 6062 -14774
rect 6334 -15018 6502 -14755
rect 6774 -15018 6823 -14746
rect 6334 -15027 6823 -15018
rect 5896 -15046 6823 -15027
rect 5581 -15080 6823 -15046
rect 12121 -15146 12450 -15076
rect 13576 -15146 13912 -13662
rect 12121 -15238 13912 -15146
rect 12121 -15256 12193 -15238
rect 11317 -15470 12193 -15256
rect 12425 -15470 13912 -15238
rect 11317 -15482 13912 -15470
rect 11317 -15585 12450 -15482
rect 7156 -16349 11207 -16325
rect 7156 -16350 9982 -16349
rect 7156 -16622 7180 -16350
rect 7452 -16622 8115 -16350
rect 8387 -16622 9051 -16350
rect 9323 -16621 9982 -16350
rect 10254 -16350 11207 -16349
rect 10254 -16621 10909 -16350
rect 9323 -16622 10909 -16621
rect 11181 -16622 11207 -16350
rect 7156 -16646 11207 -16622
rect 11317 -17278 11646 -15585
rect 12414 -16816 12821 -16704
rect 12128 -16820 12821 -16816
rect 12128 -16831 13042 -16820
rect 12128 -17103 12157 -16831
rect 12429 -16846 13042 -16831
rect 12429 -16872 13186 -16846
rect 12429 -17103 12884 -16872
rect 12128 -17133 12884 -17103
rect 12467 -17144 12884 -17133
rect 13156 -17144 13186 -16872
rect 11317 -17607 11889 -17278
rect 12467 -17292 13186 -17144
rect 12796 -17325 13186 -17292
rect 11560 -17871 11889 -17607
rect 11560 -17878 12159 -17871
rect 11560 -17940 12264 -17878
rect 11560 -18192 11889 -17940
rect 12141 -18112 12264 -17940
rect 13576 -18112 13912 -15482
rect 17292 -17998 17830 -17876
rect 12141 -18192 13912 -18112
rect 15682 -18016 17830 -17998
rect 15682 -18159 17521 -18016
rect 17664 -18159 17830 -18016
rect 15682 -18170 17830 -18159
rect 11560 -18240 13912 -18192
rect 11928 -18448 13912 -18240
rect 13576 -18480 13912 -18448
rect 17292 -18212 17830 -18170
rect 17292 -18480 17628 -18212
rect 13576 -18509 17628 -18480
rect 5006 -18832 6920 -18520
rect 13576 -18663 15546 -18509
rect 15700 -18663 17628 -18509
rect 13576 -18816 17628 -18663
rect -2310 -19086 -2309 -18972
rect -2195 -19086 -2194 -18972
rect -5026 -19910 -5025 -19796
rect -4911 -19910 -4910 -19796
rect -12501 -19996 -12373 -19954
rect -21993 -20618 -21939 -20548
rect -21869 -20618 -21621 -20548
rect -24936 -21205 -24820 -21099
rect -24714 -21205 -24666 -21099
rect -21993 -21013 -21621 -20618
rect -18248 -20419 -16239 -20155
rect -18248 -20435 -16348 -20419
rect -21993 -21083 -21937 -21013
rect -21867 -21083 -21621 -21013
rect -24936 -22407 -24666 -21205
rect -21993 -21494 -21621 -21083
rect -18248 -20864 -17860 -20435
rect -18248 -20948 -18095 -20864
rect -18011 -20948 -17860 -20864
rect -16402 -20489 -16348 -20435
rect -16278 -20489 -16239 -20419
rect -16402 -20884 -16239 -20489
rect -21993 -21564 -21933 -21494
rect -21863 -21564 -21621 -21494
rect -21993 -21605 -21621 -21564
rect -21891 -21721 -21621 -21605
rect -24936 -22513 -24810 -22407
rect -24704 -22513 -24666 -22407
rect -18248 -22268 -17860 -20948
rect -16402 -20954 -16346 -20884
rect -16276 -20954 -16239 -20884
rect -16402 -21365 -16239 -20954
rect -12501 -21118 -12471 -19996
rect -12399 -21118 -12373 -19996
rect -5026 -20615 -4910 -19910
rect -2310 -19791 -2194 -19086
rect -2310 -19905 -2309 -19791
rect -2195 -19905 -2194 -19791
rect -2310 -20418 -2194 -19905
rect -5026 -20729 -5025 -20615
rect -4911 -20729 -4910 -20615
rect -5026 -20730 -4910 -20729
rect -2310 -20532 -2309 -20418
rect -2195 -20532 -2194 -20418
rect -2310 -20533 -2194 -20532
rect -12501 -21164 -12373 -21118
rect -16402 -21435 -16342 -21365
rect -16272 -21435 -16239 -21365
rect -16402 -21476 -16239 -21435
rect -18248 -22352 -18093 -22268
rect -18009 -22352 -17860 -22268
rect -24936 -23713 -24666 -22513
rect -24936 -23819 -24830 -23713
rect -24724 -23819 -24666 -23713
rect -18248 -23670 -17860 -22352
rect -12501 -22533 -12375 -21164
rect -12501 -22575 -12373 -22533
rect -18248 -23754 -18095 -23670
rect -18011 -23754 -17860 -23670
rect -24936 -24060 -24666 -23819
rect -18248 -25050 -17860 -23754
rect -12501 -23697 -12471 -22575
rect -12399 -23697 -12373 -22575
rect 5006 -22982 5318 -18832
rect 5581 -19274 6823 -19241
rect 5581 -19283 6502 -19274
rect 5581 -19302 6062 -19283
rect 5581 -19574 5624 -19302
rect 5896 -19555 6062 -19302
rect 6334 -19546 6502 -19283
rect 6774 -19546 6823 -19274
rect 6334 -19555 6823 -19546
rect 5896 -19574 6823 -19555
rect 5581 -19608 6823 -19574
rect 12121 -19756 12450 -19604
rect 13576 -19756 13912 -18816
rect 12121 -19766 13912 -19756
rect 12121 -19784 12193 -19766
rect 11317 -19998 12193 -19784
rect 12425 -19998 13912 -19766
rect 11317 -20092 13912 -19998
rect 11317 -20113 12450 -20092
rect 7156 -20877 11207 -20853
rect 7156 -20878 9982 -20877
rect 7156 -21150 7180 -20878
rect 7452 -21150 8115 -20878
rect 8387 -21150 9051 -20878
rect 9323 -21149 9982 -20878
rect 10254 -20878 11207 -20877
rect 10254 -21149 10909 -20878
rect 9323 -21150 10909 -21149
rect 11181 -21150 11207 -20878
rect 7156 -21174 11207 -21150
rect 11317 -21806 11646 -20113
rect 12414 -21344 12821 -21232
rect 12128 -21348 12821 -21344
rect 12128 -21359 13042 -21348
rect 12128 -21631 12157 -21359
rect 12429 -21374 13042 -21359
rect 12429 -21400 13186 -21374
rect 12429 -21631 12884 -21400
rect 12128 -21661 12884 -21631
rect 12467 -21672 12884 -21661
rect 13156 -21672 13186 -21400
rect 11317 -22135 11889 -21806
rect 12467 -21820 13186 -21672
rect 12796 -21853 13186 -21820
rect 11560 -22399 11889 -22135
rect 11560 -22468 12159 -22399
rect 11560 -22720 11889 -22468
rect 12141 -22544 12159 -22468
rect 13576 -22544 13912 -20092
rect 12141 -22720 13912 -22544
rect 11560 -22768 13912 -22720
rect 11814 -22880 13912 -22768
rect 5006 -23294 6904 -22982
rect -12501 -23743 -12373 -23697
rect -18248 -25134 -18089 -25050
rect -18005 -25134 -17860 -25050
rect -18248 -25311 -17860 -25134
rect -12501 -25301 -12375 -23743
rect -12501 -25343 -12373 -25301
rect -12501 -26465 -12471 -25343
rect -12399 -26465 -12373 -25343
rect -12501 -26511 -12373 -26465
rect -12501 -27934 -12375 -26511
rect 5006 -27658 5318 -23294
rect 5581 -23802 6823 -23769
rect 5581 -23811 6502 -23802
rect 5581 -23830 6062 -23811
rect 5581 -24102 5624 -23830
rect 5896 -24083 6062 -23830
rect 6334 -24074 6502 -23811
rect 6774 -24074 6823 -23802
rect 6334 -24083 6823 -24074
rect 5896 -24102 6823 -24083
rect 5581 -24136 6823 -24102
rect 12121 -24278 12450 -24132
rect 13576 -24278 13912 -22880
rect 12121 -24294 13912 -24278
rect 12121 -24312 12193 -24294
rect 11317 -24526 12193 -24312
rect 12425 -24526 13912 -24294
rect 11317 -24614 13912 -24526
rect 11317 -24641 12450 -24614
rect 7156 -25405 11207 -25381
rect 7156 -25406 9982 -25405
rect 7156 -25678 7180 -25406
rect 7452 -25678 8115 -25406
rect 8387 -25678 9051 -25406
rect 9323 -25677 9982 -25406
rect 10254 -25406 11207 -25405
rect 10254 -25677 10909 -25406
rect 9323 -25678 10909 -25677
rect 11181 -25678 11207 -25406
rect 7156 -25702 11207 -25678
rect 11317 -26334 11646 -24641
rect 12414 -25872 12821 -25760
rect 12128 -25876 12821 -25872
rect 12128 -25887 13042 -25876
rect 12128 -26159 12157 -25887
rect 12429 -25902 13042 -25887
rect 12429 -25928 13186 -25902
rect 12429 -26159 12884 -25928
rect 12128 -26189 12884 -26159
rect 12467 -26200 12884 -26189
rect 13156 -26200 13186 -25928
rect 11317 -26663 11889 -26334
rect 12467 -26348 13186 -26200
rect 12796 -26381 13186 -26348
rect 11560 -26858 11889 -26663
rect 13576 -26858 13912 -24614
rect 11560 -26996 13912 -26858
rect 11560 -27248 11889 -26996
rect 12141 -27194 13912 -26996
rect 12141 -27248 12159 -27194
rect 11560 -27296 12159 -27248
rect -12501 -27976 -12373 -27934
rect -12501 -29098 -12471 -27976
rect -12399 -29098 -12373 -27976
rect 5006 -27970 6774 -27658
rect -12501 -29144 -12373 -29098
rect -12501 -30543 -12375 -29144
rect -12501 -30585 -12373 -30543
rect -12501 -31707 -12471 -30585
rect -12399 -31707 -12373 -30585
rect -12501 -31753 -12373 -31707
rect -12501 -33205 -12375 -31753
rect 5006 -32178 5318 -27970
rect 5581 -28330 6823 -28297
rect 5581 -28339 6502 -28330
rect 5581 -28358 6062 -28339
rect 5581 -28630 5624 -28358
rect 5896 -28611 6062 -28358
rect 6334 -28602 6502 -28339
rect 6774 -28602 6823 -28330
rect 6334 -28611 6823 -28602
rect 5896 -28630 6823 -28611
rect 5581 -28664 6823 -28630
rect 12121 -28748 12450 -28660
rect 13576 -28748 13912 -27194
rect 12120 -28822 13912 -28748
rect 12120 -28840 12193 -28822
rect 11317 -29054 12193 -28840
rect 12425 -29054 13912 -28822
rect 11317 -29084 13912 -29054
rect 11317 -29169 12450 -29084
rect 7156 -29933 11207 -29909
rect 7156 -29934 9982 -29933
rect 7156 -30206 7180 -29934
rect 7452 -30206 8115 -29934
rect 8387 -30206 9051 -29934
rect 9323 -30205 9982 -29934
rect 10254 -29934 11207 -29933
rect 10254 -30205 10909 -29934
rect 9323 -30206 10909 -30205
rect 11181 -30206 11207 -29934
rect 7156 -30230 11207 -30206
rect 11317 -30862 11646 -29169
rect 12414 -30400 12821 -30288
rect 12128 -30404 12821 -30400
rect 12128 -30415 13042 -30404
rect 12128 -30687 12157 -30415
rect 12429 -30430 13042 -30415
rect 12429 -30456 13186 -30430
rect 12429 -30687 12884 -30456
rect 12128 -30717 12884 -30687
rect 12467 -30728 12884 -30717
rect 13156 -30728 13186 -30456
rect 11317 -31191 11889 -30862
rect 12467 -30876 13186 -30728
rect 12796 -30909 13186 -30876
rect 11560 -31455 11889 -31191
rect 11560 -31524 12159 -31455
rect 11560 -31776 11889 -31524
rect 12141 -31544 12159 -31524
rect 13576 -31544 13912 -29084
rect 12141 -31776 13912 -31544
rect 11560 -31824 13912 -31776
rect 11824 -31880 13912 -31824
rect 5006 -32490 6962 -32178
rect 5006 -32698 5318 -32490
rect 5581 -32858 6823 -32825
rect 5581 -32867 6502 -32858
rect 5581 -32886 6062 -32867
rect 5581 -33158 5624 -32886
rect 5896 -33139 6062 -32886
rect 6334 -33130 6502 -32867
rect 6774 -33130 6823 -32858
rect 6334 -33139 6823 -33130
rect 5896 -33158 6823 -33139
rect 5581 -33192 6823 -33158
rect -12501 -34327 -12473 -33205
rect -12401 -34327 -12375 -33205
rect 12121 -33282 12450 -33188
rect 13576 -33282 13912 -31880
rect 12121 -33350 14308 -33282
rect 12121 -33368 12193 -33350
rect 11317 -33582 12193 -33368
rect 12425 -33582 14308 -33350
rect 11317 -33618 14308 -33582
rect 11317 -33697 12450 -33618
rect -12501 -34373 -12375 -34327
rect 7156 -34461 11207 -34437
rect 7156 -34462 9982 -34461
rect 7156 -34734 7180 -34462
rect 7452 -34734 8115 -34462
rect 8387 -34734 9051 -34462
rect 9323 -34733 9982 -34462
rect 10254 -34462 11207 -34461
rect 10254 -34733 10909 -34462
rect 9323 -34734 10909 -34733
rect 11181 -34734 11207 -34462
rect 7156 -34758 11207 -34734
rect 11317 -35390 11646 -33697
rect 12414 -34928 12821 -34816
rect 12128 -34932 12821 -34928
rect 12128 -34943 13042 -34932
rect 12128 -35215 12157 -34943
rect 12429 -34958 13042 -34943
rect 12429 -34984 13186 -34958
rect 12429 -35215 12884 -34984
rect 12128 -35245 12884 -35215
rect 12467 -35256 12884 -35245
rect 13156 -35256 13186 -34984
rect 11317 -35719 11889 -35390
rect 12467 -35404 13186 -35256
rect 12796 -35437 13186 -35404
rect 11560 -35983 11889 -35719
rect 13972 -35856 14308 -33618
rect 11560 -36052 12159 -35983
rect 11560 -36304 11889 -36052
rect 12141 -36304 12254 -36052
rect 13480 -35954 14308 -35856
rect 13480 -36068 13553 -35954
rect 13667 -36068 14308 -35954
rect 13480 -36192 14308 -36068
rect 11560 -36352 12254 -36304
rect 13972 -36352 14308 -36192
rect 11918 -36688 14308 -36352
<< via4 >>
rect 2195 4854 2467 4955
rect 2195 4784 2296 4854
rect 2296 4784 2366 4854
rect 2366 4784 2467 4854
rect 2195 4683 2467 4784
rect 3801 4854 4073 4955
rect 3801 4784 3902 4854
rect 3902 4784 3972 4854
rect 3972 4784 4073 4854
rect 3801 4683 4073 4784
rect 5505 4852 5777 4953
rect 5505 4782 5606 4852
rect 5606 4782 5676 4852
rect 5676 4782 5777 4852
rect 5505 4681 5777 4782
rect -23504 3130 -23232 3231
rect -23504 3060 -23403 3130
rect -23403 3060 -23333 3130
rect -23333 3060 -23232 3130
rect -23504 2959 -23232 3060
rect -20213 3130 -19941 3231
rect -20213 3060 -20112 3130
rect -20112 3060 -20042 3130
rect -20042 3060 -19941 3130
rect -20213 2959 -19941 3060
rect -16922 3130 -16650 3231
rect -16922 3060 -16821 3130
rect -16821 3060 -16751 3130
rect -16751 3060 -16650 3130
rect -16922 2959 -16650 3060
rect -13631 3130 -13359 3231
rect -13631 3060 -13530 3130
rect -13530 3060 -13460 3130
rect -13460 3060 -13359 3130
rect -13631 2959 -13359 3060
rect -10340 3130 -10068 3231
rect -10340 3060 -10239 3130
rect -10239 3060 -10169 3130
rect -10169 3060 -10068 3130
rect -10340 2959 -10068 3060
rect -7050 3130 -6778 3231
rect -7050 3060 -6949 3130
rect -6949 3060 -6879 3130
rect -6879 3060 -6778 3130
rect -7050 2959 -6778 3060
rect -3759 3130 -3487 3231
rect -3759 3060 -3658 3130
rect -3658 3060 -3588 3130
rect -3588 3060 -3487 3130
rect -3759 2959 -3487 3060
rect -468 3130 -196 3231
rect -468 3060 -367 3130
rect -367 3060 -297 3130
rect -297 3060 -196 3130
rect -468 2959 -196 3060
rect -24316 1346 -24044 1447
rect -24316 1276 -24215 1346
rect -24215 1276 -24145 1346
rect -24145 1276 -24044 1346
rect -24316 1175 -24044 1276
rect -22757 1346 -22485 1447
rect -22757 1276 -22656 1346
rect -22656 1276 -22586 1346
rect -22586 1276 -22485 1346
rect -22757 1175 -22485 1276
rect -21025 1346 -20753 1447
rect -21025 1276 -20924 1346
rect -20924 1276 -20854 1346
rect -20854 1276 -20753 1346
rect -21025 1175 -20753 1276
rect -19466 1346 -19194 1447
rect -19466 1276 -19365 1346
rect -19365 1276 -19295 1346
rect -19295 1276 -19194 1346
rect -19466 1175 -19194 1276
rect -17734 1346 -17462 1447
rect -17734 1276 -17633 1346
rect -17633 1276 -17563 1346
rect -17563 1276 -17462 1346
rect -17734 1175 -17462 1276
rect -16175 1346 -15903 1447
rect -16175 1276 -16074 1346
rect -16074 1276 -16004 1346
rect -16004 1276 -15903 1346
rect -16175 1175 -15903 1276
rect -14443 1346 -14171 1447
rect -14443 1276 -14342 1346
rect -14342 1276 -14272 1346
rect -14272 1276 -14171 1346
rect -14443 1175 -14171 1276
rect -12884 1346 -12612 1447
rect -12884 1276 -12783 1346
rect -12783 1276 -12713 1346
rect -12713 1276 -12612 1346
rect -12884 1175 -12612 1276
rect -11152 1346 -10880 1447
rect -11152 1276 -11051 1346
rect -11051 1276 -10981 1346
rect -10981 1276 -10880 1346
rect -11152 1175 -10880 1276
rect -9593 1346 -9321 1447
rect -9593 1276 -9492 1346
rect -9492 1276 -9422 1346
rect -9422 1276 -9321 1346
rect -9593 1175 -9321 1276
rect -7862 1346 -7590 1447
rect -7862 1276 -7761 1346
rect -7761 1276 -7691 1346
rect -7691 1276 -7590 1346
rect -7862 1175 -7590 1276
rect -6303 1346 -6031 1447
rect -6303 1276 -6202 1346
rect -6202 1276 -6132 1346
rect -6132 1276 -6031 1346
rect -6303 1175 -6031 1276
rect -4571 1346 -4299 1447
rect -4571 1276 -4470 1346
rect -4470 1276 -4400 1346
rect -4400 1276 -4299 1346
rect -4571 1175 -4299 1276
rect -3012 1346 -2740 1447
rect -3012 1276 -2911 1346
rect -2911 1276 -2841 1346
rect -2841 1276 -2740 1346
rect -3012 1175 -2740 1276
rect -1280 1346 -1008 1447
rect -1280 1276 -1179 1346
rect -1179 1276 -1109 1346
rect -1109 1276 -1008 1346
rect -1280 1175 -1008 1276
rect 279 1346 551 1447
rect 279 1276 380 1346
rect 380 1276 450 1346
rect 450 1276 551 1346
rect 279 1175 551 1276
rect -24336 267 -24001 457
rect -24336 221 -24001 267
rect -23205 255 -22933 355
rect -23205 183 -23105 255
rect -23105 183 -23033 255
rect -23033 183 -22933 255
rect -23205 83 -22933 183
rect -22343 230 -22071 333
rect -22343 164 -22240 230
rect -22240 164 -22174 230
rect -22174 164 -22071 230
rect -21045 267 -20710 457
rect -21045 221 -20710 267
rect -22343 61 -22071 164
rect -19914 255 -19642 355
rect -19914 183 -19814 255
rect -19814 183 -19742 255
rect -19742 183 -19642 255
rect -19914 83 -19642 183
rect -19052 230 -18780 333
rect -19052 164 -18949 230
rect -18949 164 -18883 230
rect -18883 164 -18780 230
rect -17754 267 -17419 457
rect -17754 221 -17419 267
rect -16623 255 -16351 355
rect -19052 61 -18780 164
rect -16623 183 -16523 255
rect -16523 183 -16451 255
rect -16451 183 -16351 255
rect -16623 83 -16351 183
rect -15761 230 -15489 333
rect -15761 164 -15658 230
rect -15658 164 -15592 230
rect -15592 164 -15489 230
rect -14463 267 -14128 457
rect -14463 221 -14128 267
rect -13332 255 -13060 355
rect -15761 61 -15489 164
rect -13332 183 -13232 255
rect -13232 183 -13160 255
rect -13160 183 -13060 255
rect -13332 83 -13060 183
rect -12470 230 -12198 333
rect -12470 164 -12367 230
rect -12367 164 -12301 230
rect -12301 164 -12198 230
rect -11172 267 -10837 457
rect -11172 221 -10837 267
rect -10041 255 -9769 355
rect -12470 61 -12198 164
rect -10041 183 -9941 255
rect -9941 183 -9869 255
rect -9869 183 -9769 255
rect -10041 83 -9769 183
rect -9179 230 -8907 333
rect -9179 164 -9076 230
rect -9076 164 -9010 230
rect -9010 164 -8907 230
rect -7882 267 -7547 457
rect -7882 221 -7547 267
rect -6751 255 -6479 355
rect -9179 61 -8907 164
rect -6751 183 -6651 255
rect -6651 183 -6579 255
rect -6579 183 -6479 255
rect -6751 83 -6479 183
rect -5889 230 -5617 333
rect -5889 164 -5786 230
rect -5786 164 -5720 230
rect -5720 164 -5617 230
rect -4591 267 -4256 457
rect -4591 221 -4256 267
rect -3460 255 -3188 355
rect -5889 61 -5617 164
rect -3460 183 -3360 255
rect -3360 183 -3288 255
rect -3288 183 -3188 255
rect -3460 83 -3188 183
rect -2598 230 -2326 333
rect -2598 164 -2495 230
rect -2495 164 -2429 230
rect -2429 164 -2326 230
rect -1300 267 -965 457
rect -1300 221 -965 267
rect -169 255 103 355
rect -2598 61 -2326 164
rect -169 183 -69 255
rect -69 183 3 255
rect 3 183 103 255
rect -169 83 103 183
rect 693 230 965 333
rect 693 164 796 230
rect 796 164 862 230
rect 862 164 965 230
rect 693 61 965 164
rect 5624 3235 5896 3338
rect 5624 3169 5727 3235
rect 5727 3169 5793 3235
rect 5793 3169 5896 3235
rect 5624 3066 5896 3169
rect 6062 3254 6334 3357
rect 6062 3188 6165 3254
rect 6165 3188 6231 3254
rect 6231 3188 6334 3254
rect 6062 3085 6334 3188
rect 6502 3263 6774 3366
rect 6502 3197 6605 3263
rect 6605 3197 6671 3263
rect 6671 3197 6774 3263
rect 6502 3094 6774 3197
rect 7180 1720 7452 1762
rect 7180 1532 7222 1720
rect 7222 1532 7410 1720
rect 7410 1532 7452 1720
rect 7180 1490 7452 1532
rect 8115 1720 8387 1762
rect 8115 1532 8157 1720
rect 8157 1532 8345 1720
rect 8345 1532 8387 1720
rect 8115 1490 8387 1532
rect 9051 1720 9323 1762
rect 9051 1532 9093 1720
rect 9093 1532 9281 1720
rect 9281 1532 9323 1720
rect 9051 1490 9323 1532
rect 9982 1720 10254 1763
rect 9982 1533 10024 1720
rect 10024 1533 10211 1720
rect 10211 1533 10254 1720
rect 9982 1491 10254 1533
rect 10909 1720 11181 1762
rect 10909 1532 10951 1720
rect 10951 1532 11139 1720
rect 11139 1532 11181 1720
rect 10909 1490 11181 1532
rect 12157 1209 12429 1281
rect 12157 1080 12228 1209
rect 12228 1080 12357 1209
rect 12357 1080 12429 1209
rect 12157 1009 12429 1080
rect 12884 1168 13156 1240
rect 12884 1039 12955 1168
rect 12955 1039 13084 1168
rect 13084 1039 13156 1168
rect 12884 968 13156 1039
rect 5624 -1293 5896 -1190
rect 5624 -1359 5727 -1293
rect 5727 -1359 5793 -1293
rect 5793 -1359 5896 -1293
rect 5624 -1462 5896 -1359
rect 6062 -1274 6334 -1171
rect 6062 -1340 6165 -1274
rect 6165 -1340 6231 -1274
rect 6231 -1340 6334 -1274
rect 6062 -1443 6334 -1340
rect 6502 -1265 6774 -1162
rect 6502 -1331 6605 -1265
rect 6605 -1331 6671 -1265
rect 6671 -1331 6774 -1265
rect 6502 -1434 6774 -1331
rect -23987 -2974 -23601 -2883
rect -23601 -2974 -23452 -2883
rect -23452 -2974 -21717 -2883
rect -23987 -2983 -21717 -2974
rect -23987 -3057 -23844 -2983
rect -23844 -3057 -22147 -2983
rect -22147 -3057 -21807 -2983
rect -21807 -3057 -21717 -2983
rect -23987 -3191 -21717 -3057
rect -20247 -2974 -19840 -2914
rect -19840 -2974 -19691 -2914
rect -19691 -2974 -18061 -2914
rect -18061 -2974 -17977 -2914
rect -20247 -2983 -17977 -2974
rect -20247 -3057 -20077 -2983
rect -20077 -3057 -18657 -2983
rect -18657 -3057 -18317 -2983
rect -18317 -3057 -17977 -2983
rect -20247 -3222 -17977 -3057
rect -24007 -4690 -21737 -4612
rect -24007 -4786 -23557 -4690
rect -23557 -4786 -23408 -4690
rect -23408 -4786 -21819 -4690
rect -21819 -4786 -21737 -4690
rect -24007 -4795 -21737 -4786
rect -24007 -4869 -23793 -4795
rect -23793 -4869 -22397 -4795
rect -22397 -4869 -22057 -4795
rect -22057 -4869 -21737 -4795
rect -24007 -4920 -21737 -4869
rect -20249 -5214 -19977 -5113
rect -20249 -5284 -20148 -5214
rect -20148 -5284 -20078 -5214
rect -20078 -5284 -19977 -5214
rect -20249 -5385 -19977 -5284
rect -18690 -5214 -18418 -5113
rect -18690 -5284 -18589 -5214
rect -18589 -5284 -18519 -5214
rect -18519 -5284 -18418 -5214
rect -18690 -5385 -18418 -5284
rect -16958 -5214 -16686 -5113
rect -16958 -5284 -16857 -5214
rect -16857 -5284 -16787 -5214
rect -16787 -5284 -16686 -5214
rect -16958 -5385 -16686 -5284
rect -15399 -5214 -15127 -5113
rect -15399 -5284 -15298 -5214
rect -15298 -5284 -15228 -5214
rect -15228 -5284 -15127 -5214
rect -15399 -5385 -15127 -5284
rect -13667 -5214 -13395 -5113
rect -13667 -5284 -13566 -5214
rect -13566 -5284 -13496 -5214
rect -13496 -5284 -13395 -5214
rect -13667 -5385 -13395 -5284
rect -12108 -5214 -11836 -5113
rect -12108 -5284 -12007 -5214
rect -12007 -5284 -11937 -5214
rect -11937 -5284 -11836 -5214
rect -12108 -5385 -11836 -5284
rect -10376 -5214 -10104 -5113
rect -10376 -5284 -10275 -5214
rect -10275 -5284 -10205 -5214
rect -10205 -5284 -10104 -5214
rect -10376 -5385 -10104 -5284
rect 7180 -2808 7452 -2766
rect 7180 -2996 7222 -2808
rect 7222 -2996 7410 -2808
rect 7410 -2996 7452 -2808
rect 7180 -3038 7452 -2996
rect 8115 -2808 8387 -2766
rect 8115 -2996 8157 -2808
rect 8157 -2996 8345 -2808
rect 8345 -2996 8387 -2808
rect 8115 -3038 8387 -2996
rect 9051 -2808 9323 -2766
rect 9051 -2996 9093 -2808
rect 9093 -2996 9281 -2808
rect 9281 -2996 9323 -2808
rect 9051 -3038 9323 -2996
rect 9982 -2808 10254 -2765
rect 9982 -2995 10024 -2808
rect 10024 -2995 10211 -2808
rect 10211 -2995 10254 -2808
rect 9982 -3037 10254 -2995
rect 10909 -2808 11181 -2766
rect 10909 -2996 10951 -2808
rect 10951 -2996 11139 -2808
rect 11139 -2996 11181 -2808
rect 10909 -3038 11181 -2996
rect 12157 -3319 12429 -3247
rect 12157 -3448 12228 -3319
rect 12228 -3448 12357 -3319
rect 12357 -3448 12429 -3319
rect 12157 -3519 12429 -3448
rect 12884 -3360 13156 -3288
rect 12884 -3489 12955 -3360
rect 12955 -3489 13084 -3360
rect 13084 -3489 13156 -3360
rect 12884 -3560 13156 -3489
rect -8817 -5214 -8545 -5113
rect -8817 -5284 -8716 -5214
rect -8716 -5284 -8646 -5214
rect -8646 -5284 -8545 -5214
rect -8817 -5385 -8545 -5284
rect -24008 -5982 -21738 -5976
rect -24008 -6078 -23559 -5982
rect -23559 -6078 -23410 -5982
rect -23410 -6078 -21825 -5982
rect -21825 -6078 -21738 -5982
rect -24008 -6087 -21738 -6078
rect -24008 -6161 -23793 -6087
rect -23793 -6161 -22397 -6087
rect -22397 -6161 -22057 -6087
rect -22057 -6161 -21738 -6087
rect -24008 -6284 -21738 -6161
rect -20269 -6293 -19934 -6103
rect -20269 -6339 -19934 -6293
rect -19138 -6305 -18866 -6205
rect -19138 -6377 -19038 -6305
rect -19038 -6377 -18966 -6305
rect -18966 -6377 -18866 -6305
rect -19138 -6477 -18866 -6377
rect -18276 -6330 -18004 -6227
rect -18276 -6396 -18173 -6330
rect -18173 -6396 -18107 -6330
rect -18107 -6396 -18004 -6330
rect -18276 -6499 -18004 -6396
rect -16978 -6293 -16643 -6103
rect -16978 -6339 -16643 -6293
rect -15847 -6305 -15575 -6205
rect -15847 -6377 -15747 -6305
rect -15747 -6377 -15675 -6305
rect -15675 -6377 -15575 -6305
rect -15847 -6477 -15575 -6377
rect -14985 -6330 -14713 -6227
rect -14985 -6396 -14882 -6330
rect -14882 -6396 -14816 -6330
rect -14816 -6396 -14713 -6330
rect -14985 -6499 -14713 -6396
rect -13687 -6293 -13352 -6103
rect -13687 -6339 -13352 -6293
rect -12556 -6305 -12284 -6205
rect -12556 -6377 -12456 -6305
rect -12456 -6377 -12384 -6305
rect -12384 -6377 -12284 -6305
rect -12556 -6477 -12284 -6377
rect -11694 -6330 -11422 -6227
rect -11694 -6396 -11591 -6330
rect -11591 -6396 -11525 -6330
rect -11525 -6396 -11422 -6330
rect -11694 -6499 -11422 -6396
rect -10396 -6293 -10061 -6103
rect -10396 -6339 -10061 -6293
rect -9265 -6305 -8993 -6205
rect -9265 -6377 -9165 -6305
rect -9165 -6377 -9093 -6305
rect -9093 -6377 -8993 -6305
rect -9265 -6477 -8993 -6377
rect -8403 -6330 -8131 -6227
rect -8403 -6396 -8300 -6330
rect -8300 -6396 -8234 -6330
rect -8234 -6396 -8131 -6330
rect -8403 -6499 -8131 -6396
rect -24046 -7955 -21776 -7870
rect -24046 -8051 -23558 -7955
rect -23558 -8051 -23409 -7955
rect -23409 -8051 -21823 -7955
rect -21823 -8051 -21776 -7955
rect -24046 -8060 -21776 -8051
rect -24046 -8134 -23793 -8060
rect -23793 -8134 -22396 -8060
rect -22396 -8134 -22056 -8060
rect -22056 -8134 -21776 -8060
rect -24046 -8178 -21776 -8134
rect -20249 -8479 -19977 -8378
rect -20249 -8549 -20148 -8479
rect -20148 -8549 -20078 -8479
rect -20078 -8549 -19977 -8479
rect -20249 -8650 -19977 -8549
rect -18690 -8479 -18418 -8378
rect -18690 -8549 -18589 -8479
rect -18589 -8549 -18519 -8479
rect -18519 -8549 -18418 -8479
rect -18690 -8650 -18418 -8549
rect -16958 -8479 -16686 -8378
rect -16958 -8549 -16857 -8479
rect -16857 -8549 -16787 -8479
rect -16787 -8549 -16686 -8479
rect -16958 -8650 -16686 -8549
rect -15399 -8479 -15127 -8378
rect -15399 -8549 -15298 -8479
rect -15298 -8549 -15228 -8479
rect -15228 -8549 -15127 -8479
rect -15399 -8650 -15127 -8549
rect -13667 -8479 -13395 -8378
rect -13667 -8549 -13566 -8479
rect -13566 -8549 -13496 -8479
rect -13496 -8549 -13395 -8479
rect -13667 -8650 -13395 -8549
rect -12108 -8479 -11836 -8378
rect -12108 -8549 -12007 -8479
rect -12007 -8549 -11937 -8479
rect -11937 -8549 -11836 -8479
rect -12108 -8650 -11836 -8549
rect -10376 -8479 -10104 -8378
rect -10376 -8549 -10275 -8479
rect -10275 -8549 -10205 -8479
rect -10205 -8549 -10104 -8479
rect -10376 -8650 -10104 -8549
rect -8817 -8479 -8545 -8378
rect -8817 -8549 -8716 -8479
rect -8716 -8549 -8646 -8479
rect -8646 -8549 -8545 -8479
rect -8817 -8650 -8545 -8549
rect -24060 -9343 -23556 -9248
rect -23556 -9343 -23407 -9248
rect -23407 -9343 -21819 -9248
rect -21819 -9343 -21790 -9248
rect -24060 -9352 -21790 -9343
rect -24060 -9426 -23793 -9352
rect -23793 -9426 -22397 -9352
rect -22397 -9426 -22057 -9352
rect -22057 -9426 -21790 -9352
rect -24060 -9556 -21790 -9426
rect -20269 -9558 -19934 -9368
rect -20269 -9604 -19934 -9558
rect -19138 -9570 -18866 -9470
rect -19138 -9642 -19038 -9570
rect -19038 -9642 -18966 -9570
rect -18966 -9642 -18866 -9570
rect -19138 -9742 -18866 -9642
rect -18276 -9595 -18004 -9492
rect -18276 -9661 -18173 -9595
rect -18173 -9661 -18107 -9595
rect -18107 -9661 -18004 -9595
rect -18276 -9764 -18004 -9661
rect -16978 -9558 -16643 -9368
rect -16978 -9604 -16643 -9558
rect -15847 -9570 -15575 -9470
rect -15847 -9642 -15747 -9570
rect -15747 -9642 -15675 -9570
rect -15675 -9642 -15575 -9570
rect -15847 -9742 -15575 -9642
rect -14985 -9595 -14713 -9492
rect -14985 -9661 -14882 -9595
rect -14882 -9661 -14816 -9595
rect -14816 -9661 -14713 -9595
rect -14985 -9764 -14713 -9661
rect -13687 -9558 -13352 -9368
rect -13687 -9604 -13352 -9558
rect -12556 -9570 -12284 -9470
rect -12556 -9642 -12456 -9570
rect -12456 -9642 -12384 -9570
rect -12384 -9642 -12284 -9570
rect -12556 -9742 -12284 -9642
rect -11694 -9595 -11422 -9492
rect -11694 -9661 -11591 -9595
rect -11591 -9661 -11525 -9595
rect -11525 -9661 -11422 -9595
rect -11694 -9764 -11422 -9661
rect -10396 -9558 -10061 -9368
rect 5624 -5721 5896 -5618
rect 5624 -5787 5727 -5721
rect 5727 -5787 5793 -5721
rect 5793 -5787 5896 -5721
rect 5624 -5890 5896 -5787
rect 6062 -5702 6334 -5599
rect 6062 -5768 6165 -5702
rect 6165 -5768 6231 -5702
rect 6231 -5768 6334 -5702
rect 6062 -5871 6334 -5768
rect 6502 -5693 6774 -5590
rect 6502 -5759 6605 -5693
rect 6605 -5759 6671 -5693
rect 6671 -5759 6774 -5693
rect 6502 -5862 6774 -5759
rect 7180 -7236 7452 -7194
rect 7180 -7424 7222 -7236
rect 7222 -7424 7410 -7236
rect 7410 -7424 7452 -7236
rect 7180 -7466 7452 -7424
rect 8115 -7236 8387 -7194
rect 8115 -7424 8157 -7236
rect 8157 -7424 8345 -7236
rect 8345 -7424 8387 -7236
rect 8115 -7466 8387 -7424
rect 9051 -7236 9323 -7194
rect 9051 -7424 9093 -7236
rect 9093 -7424 9281 -7236
rect 9281 -7424 9323 -7236
rect 9051 -7466 9323 -7424
rect 9982 -7236 10254 -7193
rect 9982 -7423 10024 -7236
rect 10024 -7423 10211 -7236
rect 10211 -7423 10254 -7236
rect 9982 -7465 10254 -7423
rect 10909 -7236 11181 -7194
rect 10909 -7424 10951 -7236
rect 10951 -7424 11139 -7236
rect 11139 -7424 11181 -7236
rect 10909 -7466 11181 -7424
rect 12157 -7747 12429 -7675
rect 12157 -7876 12228 -7747
rect 12228 -7876 12357 -7747
rect 12357 -7876 12429 -7747
rect 12157 -7947 12429 -7876
rect 12884 -7788 13156 -7716
rect 12884 -7917 12955 -7788
rect 12955 -7917 13084 -7788
rect 13084 -7917 13156 -7788
rect 12884 -7988 13156 -7917
rect -10396 -9604 -10061 -9558
rect -9265 -9570 -8993 -9470
rect -9265 -9642 -9165 -9570
rect -9165 -9642 -9093 -9570
rect -9093 -9642 -8993 -9570
rect -9265 -9742 -8993 -9642
rect -8403 -9595 -8131 -9492
rect -8403 -9661 -8300 -9595
rect -8300 -9661 -8234 -9595
rect -8234 -9661 -8131 -9595
rect -8403 -9764 -8131 -9661
rect -24018 -11219 -21748 -11202
rect -24018 -11315 -23556 -11219
rect -23556 -11315 -23407 -11219
rect -23407 -11315 -21823 -11219
rect -21823 -11315 -21748 -11219
rect -24018 -11324 -21748 -11315
rect -24018 -11398 -23793 -11324
rect -23793 -11398 -22396 -11324
rect -22396 -11398 -22056 -11324
rect -22056 -11398 -21748 -11324
rect -24018 -11510 -21748 -11398
rect -20249 -11743 -19977 -11642
rect -20249 -11813 -20148 -11743
rect -20148 -11813 -20078 -11743
rect -20078 -11813 -19977 -11743
rect -20249 -11914 -19977 -11813
rect -18690 -11743 -18418 -11642
rect -18690 -11813 -18589 -11743
rect -18589 -11813 -18519 -11743
rect -18519 -11813 -18418 -11743
rect -18690 -11914 -18418 -11813
rect -16958 -11743 -16686 -11642
rect -16958 -11813 -16857 -11743
rect -16857 -11813 -16787 -11743
rect -16787 -11813 -16686 -11743
rect -16958 -11914 -16686 -11813
rect -15399 -11743 -15127 -11642
rect -15399 -11813 -15298 -11743
rect -15298 -11813 -15228 -11743
rect -15228 -11813 -15127 -11743
rect -15399 -11914 -15127 -11813
rect -13667 -11743 -13395 -11642
rect -13667 -11813 -13566 -11743
rect -13566 -11813 -13496 -11743
rect -13496 -11813 -13395 -11743
rect -13667 -11914 -13395 -11813
rect -12108 -11743 -11836 -11642
rect -12108 -11813 -12007 -11743
rect -12007 -11813 -11937 -11743
rect -11937 -11813 -11836 -11743
rect -12108 -11914 -11836 -11813
rect -10376 -11743 -10104 -11642
rect -10376 -11813 -10275 -11743
rect -10275 -11813 -10205 -11743
rect -10205 -11813 -10104 -11743
rect -10376 -11914 -10104 -11813
rect -8817 -11743 -8545 -11642
rect -8817 -11813 -8716 -11743
rect -8716 -11813 -8646 -11743
rect -8646 -11813 -8545 -11743
rect -8817 -11914 -8545 -11813
rect -24029 -12607 -23556 -12535
rect -23556 -12607 -23407 -12535
rect -23407 -12607 -21827 -12535
rect -21827 -12607 -21759 -12535
rect -24029 -12616 -21759 -12607
rect -24029 -12690 -23793 -12616
rect -23793 -12690 -22396 -12616
rect -22396 -12690 -22056 -12616
rect -22056 -12690 -21759 -12616
rect -24029 -12843 -21759 -12690
rect -23531 -15070 -23211 -14965
rect -23531 -15181 -23426 -15070
rect -23426 -15181 -23315 -15070
rect -23315 -15181 -23211 -15070
rect -23531 -15285 -23211 -15181
rect -20269 -12822 -19934 -12632
rect -20269 -12868 -19934 -12822
rect -19138 -12834 -18866 -12734
rect -19138 -12906 -19038 -12834
rect -19038 -12906 -18966 -12834
rect -18966 -12906 -18866 -12834
rect -19138 -13006 -18866 -12906
rect -18276 -12859 -18004 -12756
rect -18276 -12925 -18173 -12859
rect -18173 -12925 -18107 -12859
rect -18107 -12925 -18004 -12859
rect -16978 -12822 -16643 -12632
rect -16978 -12868 -16643 -12822
rect -15847 -12834 -15575 -12734
rect -18276 -13028 -18004 -12925
rect -15847 -12906 -15747 -12834
rect -15747 -12906 -15675 -12834
rect -15675 -12906 -15575 -12834
rect -15847 -13006 -15575 -12906
rect -14985 -12859 -14713 -12756
rect -14985 -12925 -14882 -12859
rect -14882 -12925 -14816 -12859
rect -14816 -12925 -14713 -12859
rect -13687 -12822 -13352 -12632
rect -13687 -12868 -13352 -12822
rect -12556 -12834 -12284 -12734
rect -14985 -13028 -14713 -12925
rect -12556 -12906 -12456 -12834
rect -12456 -12906 -12384 -12834
rect -12384 -12906 -12284 -12834
rect -12556 -13006 -12284 -12906
rect -11694 -12859 -11422 -12756
rect -11694 -12925 -11591 -12859
rect -11591 -12925 -11525 -12859
rect -11525 -12925 -11422 -12859
rect -10396 -12822 -10061 -12632
rect -10396 -12868 -10061 -12822
rect -9265 -12834 -8993 -12734
rect -11694 -13028 -11422 -12925
rect -9265 -12906 -9165 -12834
rect -9165 -12906 -9093 -12834
rect -9093 -12906 -8993 -12834
rect -9265 -13006 -8993 -12906
rect -8403 -12859 -8131 -12756
rect -8403 -12925 -8300 -12859
rect -8300 -12925 -8234 -12859
rect -8234 -12925 -8131 -12859
rect -8403 -13028 -8131 -12925
rect -17039 -15321 -16719 -15196
rect -17039 -15391 -16914 -15321
rect -16914 -15391 -16844 -15321
rect -16844 -15391 -16719 -15321
rect -17039 -15516 -16719 -15391
rect 5624 -10349 5896 -10246
rect 5624 -10415 5727 -10349
rect 5727 -10415 5793 -10349
rect 5793 -10415 5896 -10349
rect 5624 -10518 5896 -10415
rect 6062 -10330 6334 -10227
rect 6062 -10396 6165 -10330
rect 6165 -10396 6231 -10330
rect 6231 -10396 6334 -10330
rect 6062 -10499 6334 -10396
rect 6502 -10321 6774 -10218
rect 6502 -10387 6605 -10321
rect 6605 -10387 6671 -10321
rect 6671 -10387 6774 -10321
rect 6502 -10490 6774 -10387
rect 7180 -11864 7452 -11822
rect 7180 -12052 7222 -11864
rect 7222 -12052 7410 -11864
rect 7410 -12052 7452 -11864
rect 7180 -12094 7452 -12052
rect 8115 -11864 8387 -11822
rect 8115 -12052 8157 -11864
rect 8157 -12052 8345 -11864
rect 8345 -12052 8387 -11864
rect 8115 -12094 8387 -12052
rect 9051 -11864 9323 -11822
rect 9051 -12052 9093 -11864
rect 9093 -12052 9281 -11864
rect 9281 -12052 9323 -11864
rect 9051 -12094 9323 -12052
rect 9982 -11864 10254 -11821
rect 9982 -12051 10024 -11864
rect 10024 -12051 10211 -11864
rect 10211 -12051 10254 -11864
rect 9982 -12093 10254 -12051
rect 10909 -11864 11181 -11822
rect 10909 -12052 10951 -11864
rect 10951 -12052 11139 -11864
rect 11139 -12052 11181 -11864
rect 10909 -12094 11181 -12052
rect 12157 -12375 12429 -12303
rect 12157 -12504 12228 -12375
rect 12228 -12504 12357 -12375
rect 12357 -12504 12429 -12375
rect 12157 -12575 12429 -12504
rect 12884 -12416 13156 -12344
rect 12884 -12545 12955 -12416
rect 12955 -12545 13084 -12416
rect 13084 -12545 13156 -12416
rect 12884 -12616 13156 -12545
rect -4092 -14245 -3820 -14163
rect -4092 -14352 -4009 -14245
rect -4009 -14352 -3902 -14245
rect -3902 -14352 -3820 -14245
rect -4092 -14435 -3820 -14352
rect -11187 -14820 -10915 -14719
rect -11187 -14890 -11086 -14820
rect -11086 -14890 -11016 -14820
rect -11016 -14890 -10915 -14820
rect -11187 -14991 -10915 -14890
rect -1376 -14069 -1104 -13986
rect -1376 -14176 -1293 -14069
rect -1293 -14176 -1186 -14069
rect -1186 -14176 -1104 -14069
rect -1376 -14258 -1104 -14176
rect -7320 -15392 -7000 -15281
rect -7320 -15491 -7209 -15392
rect -7209 -15491 -7110 -15392
rect -7110 -15491 -7000 -15392
rect -7320 -15601 -7000 -15491
rect -4092 -14878 -3820 -14796
rect -4092 -14985 -4009 -14878
rect -4009 -14985 -3902 -14878
rect -3902 -14985 -3820 -14878
rect -4092 -15068 -3820 -14985
rect -23488 -16266 -23168 -16161
rect -23488 -16377 -23383 -16266
rect -23383 -16377 -23272 -16266
rect -23272 -16377 -23168 -16266
rect -23488 -16481 -23168 -16377
rect -23479 -17478 -23159 -17373
rect -23479 -17589 -23374 -17478
rect -23374 -17589 -23263 -17478
rect -23263 -17589 -23159 -17478
rect -23479 -17693 -23159 -17589
rect -7327 -15885 -7007 -15774
rect -7327 -15984 -7216 -15885
rect -7216 -15984 -7117 -15885
rect -7117 -15984 -7007 -15885
rect -7327 -16094 -7007 -15984
rect -23471 -18619 -23151 -18514
rect -23471 -18730 -23366 -18619
rect -23366 -18730 -23255 -18619
rect -23255 -18730 -23151 -18619
rect -23471 -18834 -23151 -18730
rect -20759 -18080 -20439 -17969
rect -20759 -18179 -20648 -18080
rect -20648 -18179 -20549 -18080
rect -20549 -18179 -20439 -18080
rect -20759 -18289 -20439 -18179
rect -17039 -16727 -16719 -16602
rect -17039 -16797 -16914 -16727
rect -16914 -16797 -16844 -16727
rect -16844 -16797 -16719 -16727
rect -17039 -16922 -16719 -16797
rect -7328 -16371 -7008 -16260
rect -7328 -16470 -7217 -16371
rect -7217 -16470 -7118 -16371
rect -7118 -16470 -7008 -16371
rect -7328 -16580 -7008 -16470
rect -4092 -15697 -3820 -15615
rect -4092 -15804 -4009 -15697
rect -4009 -15804 -3902 -15697
rect -3902 -15804 -3820 -15697
rect -4092 -15887 -3820 -15804
rect -1376 -14888 -1104 -14805
rect -1376 -14995 -1293 -14888
rect -1293 -14995 -1186 -14888
rect -1186 -14995 -1104 -14888
rect -1376 -15077 -1104 -14995
rect -20766 -18573 -20446 -18462
rect -20766 -18672 -20655 -18573
rect -20655 -18672 -20556 -18573
rect -20556 -18672 -20446 -18573
rect -20766 -18782 -20446 -18672
rect -20767 -19059 -20447 -18948
rect -20767 -19158 -20656 -19059
rect -20656 -19158 -20557 -19059
rect -20557 -19158 -20447 -19059
rect -20767 -19268 -20447 -19158
rect -23448 -19791 -23128 -19686
rect -23448 -19902 -23343 -19791
rect -23343 -19902 -23232 -19791
rect -23232 -19902 -23128 -19791
rect -23448 -20006 -23128 -19902
rect -20771 -19566 -20451 -19455
rect -20771 -19665 -20660 -19566
rect -20660 -19665 -20561 -19566
rect -20561 -19665 -20451 -19566
rect -20771 -19775 -20451 -19665
rect -17170 -18158 -16850 -18033
rect -17170 -18228 -17045 -18158
rect -17045 -18228 -16975 -18158
rect -16975 -18228 -16850 -18158
rect -17170 -18353 -16850 -18228
rect -15168 -17951 -14848 -17840
rect -15168 -18050 -15057 -17951
rect -15057 -18050 -14958 -17951
rect -14958 -18050 -14848 -17951
rect -15168 -18160 -14848 -18050
rect -7332 -16878 -7012 -16767
rect -7332 -16977 -7221 -16878
rect -7221 -16977 -7122 -16878
rect -7122 -16977 -7012 -16878
rect -7332 -17087 -7012 -16977
rect -11185 -17636 -10913 -17535
rect -11185 -17706 -11084 -17636
rect -11084 -17706 -11014 -17636
rect -11014 -17706 -10913 -17636
rect -11185 -17807 -10913 -17706
rect -7331 -17353 -7011 -17242
rect -7331 -17452 -7220 -17353
rect -7220 -17452 -7121 -17353
rect -7121 -17452 -7011 -17353
rect -7331 -17562 -7011 -17452
rect -4092 -16516 -3820 -16434
rect -4092 -16623 -4009 -16516
rect -4009 -16623 -3902 -16516
rect -3902 -16623 -3820 -16516
rect -4092 -16706 -3820 -16623
rect -1376 -15707 -1104 -15624
rect -1376 -15814 -1293 -15707
rect -1293 -15814 -1186 -15707
rect -1186 -15814 -1104 -15707
rect -1376 -15896 -1104 -15814
rect -15175 -18444 -14855 -18333
rect -15175 -18543 -15064 -18444
rect -15064 -18543 -14965 -18444
rect -14965 -18543 -14855 -18444
rect -15175 -18653 -14855 -18543
rect -20770 -20041 -20450 -19930
rect -20770 -20140 -20659 -20041
rect -20659 -20140 -20560 -20041
rect -20560 -20140 -20450 -20041
rect -20770 -20250 -20450 -20140
rect -17055 -19613 -16735 -19488
rect -17055 -19683 -16930 -19613
rect -16930 -19683 -16860 -19613
rect -16860 -19683 -16735 -19613
rect -17055 -19808 -16735 -19683
rect -15176 -18930 -14856 -18819
rect -15176 -19029 -15065 -18930
rect -15065 -19029 -14966 -18930
rect -14966 -19029 -14856 -18930
rect -15176 -19139 -14856 -19029
rect -15180 -19437 -14860 -19326
rect -15180 -19536 -15069 -19437
rect -15069 -19536 -14970 -19437
rect -14970 -19536 -14860 -19437
rect -15180 -19646 -14860 -19536
rect -15179 -19912 -14859 -19801
rect -15179 -20011 -15068 -19912
rect -15068 -20011 -14969 -19912
rect -14969 -20011 -14859 -19912
rect -15179 -20121 -14859 -20011
rect -7326 -17805 -7006 -17694
rect -7326 -17904 -7215 -17805
rect -7215 -17904 -7116 -17805
rect -7116 -17904 -7006 -17805
rect -7326 -18014 -7006 -17904
rect -7326 -18247 -7006 -18136
rect -7326 -18346 -7215 -18247
rect -7215 -18346 -7116 -18247
rect -7116 -18346 -7006 -18247
rect -7326 -18456 -7006 -18346
rect -4092 -17335 -3820 -17253
rect -4092 -17442 -4009 -17335
rect -4009 -17442 -3902 -17335
rect -3902 -17442 -3820 -17335
rect -4092 -17525 -3820 -17442
rect -1376 -16526 -1104 -16443
rect -1376 -16633 -1293 -16526
rect -1293 -16633 -1186 -16526
rect -1186 -16633 -1104 -16526
rect -1376 -16715 -1104 -16633
rect -7332 -18728 -7012 -18617
rect -7332 -18827 -7221 -18728
rect -7221 -18827 -7122 -18728
rect -7122 -18827 -7012 -18728
rect -7332 -18937 -7012 -18827
rect -4092 -18154 -3820 -18072
rect -4092 -18261 -4009 -18154
rect -4009 -18261 -3902 -18154
rect -3902 -18261 -3820 -18154
rect -4092 -18344 -3820 -18261
rect -1376 -17345 -1104 -17262
rect -1376 -17452 -1293 -17345
rect -1293 -17452 -1186 -17345
rect -1186 -17452 -1104 -17345
rect -1376 -17534 -1104 -17452
rect -4092 -18973 -3820 -18891
rect -4092 -19080 -4009 -18973
rect -4009 -19080 -3902 -18973
rect -3902 -19080 -3820 -18973
rect -4092 -19163 -3820 -19080
rect -1376 -18164 -1104 -18081
rect -1376 -18271 -1293 -18164
rect -1293 -18271 -1186 -18164
rect -1186 -18271 -1104 -18164
rect -1376 -18353 -1104 -18271
rect 5624 -14877 5896 -14774
rect 5624 -14943 5727 -14877
rect 5727 -14943 5793 -14877
rect 5793 -14943 5896 -14877
rect 5624 -15046 5896 -14943
rect 6062 -14858 6334 -14755
rect 6062 -14924 6165 -14858
rect 6165 -14924 6231 -14858
rect 6231 -14924 6334 -14858
rect 6062 -15027 6334 -14924
rect 6502 -14849 6774 -14746
rect 6502 -14915 6605 -14849
rect 6605 -14915 6671 -14849
rect 6671 -14915 6774 -14849
rect 6502 -15018 6774 -14915
rect 7180 -16392 7452 -16350
rect 7180 -16580 7222 -16392
rect 7222 -16580 7410 -16392
rect 7410 -16580 7452 -16392
rect 7180 -16622 7452 -16580
rect 8115 -16392 8387 -16350
rect 8115 -16580 8157 -16392
rect 8157 -16580 8345 -16392
rect 8345 -16580 8387 -16392
rect 8115 -16622 8387 -16580
rect 9051 -16392 9323 -16350
rect 9051 -16580 9093 -16392
rect 9093 -16580 9281 -16392
rect 9281 -16580 9323 -16392
rect 9051 -16622 9323 -16580
rect 9982 -16392 10254 -16349
rect 9982 -16579 10024 -16392
rect 10024 -16579 10211 -16392
rect 10211 -16579 10254 -16392
rect 9982 -16621 10254 -16579
rect 10909 -16392 11181 -16350
rect 10909 -16580 10951 -16392
rect 10951 -16580 11139 -16392
rect 11139 -16580 11181 -16392
rect 10909 -16622 11181 -16580
rect 12157 -16903 12429 -16831
rect 12157 -17032 12228 -16903
rect 12228 -17032 12357 -16903
rect 12357 -17032 12429 -16903
rect 12157 -17103 12429 -17032
rect 12884 -16944 13156 -16872
rect 12884 -17073 12955 -16944
rect 12955 -17073 13084 -16944
rect 13084 -17073 13156 -16944
rect 12884 -17144 13156 -17073
rect 16278 -16732 16550 -16730
rect 16278 -17000 16280 -16732
rect 16280 -17000 16548 -16732
rect 16548 -17000 16550 -16732
rect 16278 -17002 16550 -17000
rect -23439 -20989 -23119 -20884
rect -23439 -21100 -23334 -20989
rect -23334 -21100 -23223 -20989
rect -23223 -21100 -23119 -20989
rect -23439 -21204 -23119 -21100
rect -20765 -20493 -20445 -20382
rect -20765 -20592 -20654 -20493
rect -20654 -20592 -20555 -20493
rect -20555 -20592 -20445 -20493
rect -20765 -20702 -20445 -20592
rect -20765 -20935 -20445 -20824
rect -20765 -21034 -20654 -20935
rect -20654 -21034 -20555 -20935
rect -20555 -21034 -20445 -20935
rect -20765 -21144 -20445 -21034
rect -15174 -20364 -14854 -20253
rect -15174 -20463 -15063 -20364
rect -15063 -20463 -14964 -20364
rect -14964 -20463 -14854 -20364
rect -15174 -20573 -14854 -20463
rect -20771 -21416 -20451 -21305
rect -20771 -21515 -20660 -21416
rect -20660 -21515 -20561 -21416
rect -20561 -21515 -20451 -21416
rect -20771 -21625 -20451 -21515
rect -23442 -22283 -23122 -22178
rect -23442 -22394 -23337 -22283
rect -23337 -22394 -23226 -22283
rect -23226 -22394 -23122 -22283
rect -23442 -22498 -23122 -22394
rect -17045 -21008 -16725 -20884
rect -17045 -21080 -16921 -21008
rect -16921 -21080 -16849 -21008
rect -16849 -21080 -16725 -21008
rect -17045 -21204 -16725 -21080
rect -15174 -20806 -14854 -20695
rect -15174 -20905 -15063 -20806
rect -15063 -20905 -14964 -20806
rect -14964 -20905 -14854 -20806
rect -15174 -21015 -14854 -20905
rect -11185 -20593 -10913 -20492
rect -11185 -20663 -11084 -20593
rect -11084 -20663 -11014 -20593
rect -11014 -20663 -10913 -20593
rect -11185 -20764 -10913 -20663
rect -4092 -19792 -3820 -19710
rect -4092 -19899 -4009 -19792
rect -4009 -19899 -3902 -19792
rect -3902 -19899 -3820 -19792
rect -4092 -19982 -3820 -19899
rect -1376 -18983 -1104 -18900
rect -1376 -19090 -1293 -18983
rect -1293 -19090 -1186 -18983
rect -1186 -19090 -1104 -18983
rect -1376 -19172 -1104 -19090
rect -1376 -19802 -1104 -19719
rect -1376 -19909 -1293 -19802
rect -1293 -19909 -1186 -19802
rect -1186 -19909 -1104 -19802
rect -1376 -19991 -1104 -19909
rect -4092 -20611 -3820 -20529
rect -1376 -20435 -1104 -20352
rect -4092 -20718 -4009 -20611
rect -4009 -20718 -3902 -20611
rect -3902 -20718 -3820 -20611
rect -1376 -20542 -1293 -20435
rect -1293 -20542 -1186 -20435
rect -1186 -20542 -1104 -20435
rect -1376 -20624 -1104 -20542
rect -4092 -20801 -3820 -20718
rect -15180 -21287 -14860 -21176
rect -15180 -21386 -15069 -21287
rect -15069 -21386 -14970 -21287
rect -14970 -21386 -14860 -21287
rect -15180 -21496 -14860 -21386
rect -16854 -21978 -16534 -21855
rect -16854 -22052 -16731 -21978
rect -16731 -22052 -16657 -21978
rect -16657 -22052 -16534 -21978
rect -16854 -22175 -16534 -22052
rect -23482 -23599 -23162 -23494
rect -23482 -23710 -23377 -23599
rect -23377 -23710 -23266 -23599
rect -23266 -23710 -23162 -23599
rect -23482 -23814 -23162 -23710
rect -16809 -23362 -16489 -23246
rect -16809 -23450 -16693 -23362
rect -16693 -23450 -16605 -23362
rect -16605 -23450 -16489 -23362
rect -16809 -23566 -16489 -23450
rect 5624 -19405 5896 -19302
rect 5624 -19471 5727 -19405
rect 5727 -19471 5793 -19405
rect 5793 -19471 5896 -19405
rect 5624 -19574 5896 -19471
rect 6062 -19386 6334 -19283
rect 6062 -19452 6165 -19386
rect 6165 -19452 6231 -19386
rect 6231 -19452 6334 -19386
rect 6062 -19555 6334 -19452
rect 6502 -19377 6774 -19274
rect 6502 -19443 6605 -19377
rect 6605 -19443 6671 -19377
rect 6671 -19443 6774 -19377
rect 6502 -19546 6774 -19443
rect 17877 -18864 18149 -18768
rect 17877 -18945 17972 -18864
rect 17972 -18945 18053 -18864
rect 18053 -18945 18149 -18864
rect 17877 -19040 18149 -18945
rect 7180 -20920 7452 -20878
rect 7180 -21108 7222 -20920
rect 7222 -21108 7410 -20920
rect 7410 -21108 7452 -20920
rect 7180 -21150 7452 -21108
rect 8115 -20920 8387 -20878
rect 8115 -21108 8157 -20920
rect 8157 -21108 8345 -20920
rect 8345 -21108 8387 -20920
rect 8115 -21150 8387 -21108
rect 9051 -20920 9323 -20878
rect 9051 -21108 9093 -20920
rect 9093 -21108 9281 -20920
rect 9281 -21108 9323 -20920
rect 9051 -21150 9323 -21108
rect 9982 -20920 10254 -20877
rect 9982 -21107 10024 -20920
rect 10024 -21107 10211 -20920
rect 10211 -21107 10254 -20920
rect 9982 -21149 10254 -21107
rect 10909 -20920 11181 -20878
rect 10909 -21108 10951 -20920
rect 10951 -21108 11139 -20920
rect 11139 -21108 11181 -20920
rect 10909 -21150 11181 -21108
rect 12157 -21431 12429 -21359
rect 12157 -21560 12228 -21431
rect 12228 -21560 12357 -21431
rect 12357 -21560 12429 -21431
rect 12157 -21631 12429 -21560
rect 12884 -21472 13156 -21400
rect 12884 -21601 12955 -21472
rect 12955 -21601 13084 -21472
rect 13084 -21601 13156 -21472
rect 12884 -21672 13156 -21601
rect 16220 -20172 16492 -20170
rect 16220 -20441 16226 -20172
rect 16226 -20441 16485 -20172
rect 16485 -20441 16492 -20172
rect 16220 -20442 16492 -20441
rect -11185 -23172 -10913 -23071
rect -11185 -23242 -11084 -23172
rect -11084 -23242 -11014 -23172
rect -11014 -23242 -10913 -23172
rect -11185 -23343 -10913 -23242
rect -16811 -24770 -16491 -24652
rect -16811 -24854 -16693 -24770
rect -16693 -24854 -16609 -24770
rect -16609 -24854 -16491 -24770
rect -16811 -24972 -16491 -24854
rect -11185 -25940 -10913 -25839
rect -11185 -26010 -11084 -25940
rect -11084 -26010 -11014 -25940
rect -11014 -26010 -10913 -25940
rect -11185 -26111 -10913 -26010
rect 5624 -23933 5896 -23830
rect 5624 -23999 5727 -23933
rect 5727 -23999 5793 -23933
rect 5793 -23999 5896 -23933
rect 5624 -24102 5896 -23999
rect 6062 -23914 6334 -23811
rect 6062 -23980 6165 -23914
rect 6165 -23980 6231 -23914
rect 6231 -23980 6334 -23914
rect 6062 -24083 6334 -23980
rect 6502 -23905 6774 -23802
rect 6502 -23971 6605 -23905
rect 6605 -23971 6671 -23905
rect 6671 -23971 6774 -23905
rect 6502 -24074 6774 -23971
rect 7180 -25448 7452 -25406
rect 7180 -25636 7222 -25448
rect 7222 -25636 7410 -25448
rect 7410 -25636 7452 -25448
rect 7180 -25678 7452 -25636
rect 8115 -25448 8387 -25406
rect 8115 -25636 8157 -25448
rect 8157 -25636 8345 -25448
rect 8345 -25636 8387 -25448
rect 8115 -25678 8387 -25636
rect 9051 -25448 9323 -25406
rect 9051 -25636 9093 -25448
rect 9093 -25636 9281 -25448
rect 9281 -25636 9323 -25448
rect 9051 -25678 9323 -25636
rect 9982 -25448 10254 -25405
rect 9982 -25635 10024 -25448
rect 10024 -25635 10211 -25448
rect 10211 -25635 10254 -25448
rect 9982 -25677 10254 -25635
rect 10909 -25448 11181 -25406
rect 10909 -25636 10951 -25448
rect 10951 -25636 11139 -25448
rect 11139 -25636 11181 -25448
rect 10909 -25678 11181 -25636
rect 12157 -25959 12429 -25887
rect 12157 -26088 12228 -25959
rect 12228 -26088 12357 -25959
rect 12357 -26088 12429 -25959
rect 12157 -26159 12429 -26088
rect 12884 -26000 13156 -25928
rect 12884 -26129 12955 -26000
rect 12955 -26129 13084 -26000
rect 13084 -26129 13156 -26000
rect 12884 -26200 13156 -26129
rect -11185 -28573 -10913 -28472
rect -11185 -28643 -11084 -28573
rect -11084 -28643 -11014 -28573
rect -11014 -28643 -10913 -28573
rect -11185 -28744 -10913 -28643
rect -11185 -31182 -10913 -31081
rect -11185 -31252 -11084 -31182
rect -11084 -31252 -11014 -31182
rect -11014 -31252 -10913 -31182
rect -11185 -31353 -10913 -31252
rect 5624 -28461 5896 -28358
rect 5624 -28527 5727 -28461
rect 5727 -28527 5793 -28461
rect 5793 -28527 5896 -28461
rect 5624 -28630 5896 -28527
rect 6062 -28442 6334 -28339
rect 6062 -28508 6165 -28442
rect 6165 -28508 6231 -28442
rect 6231 -28508 6334 -28442
rect 6062 -28611 6334 -28508
rect 6502 -28433 6774 -28330
rect 6502 -28499 6605 -28433
rect 6605 -28499 6671 -28433
rect 6671 -28499 6774 -28433
rect 6502 -28602 6774 -28499
rect 7180 -29976 7452 -29934
rect 7180 -30164 7222 -29976
rect 7222 -30164 7410 -29976
rect 7410 -30164 7452 -29976
rect 7180 -30206 7452 -30164
rect 8115 -29976 8387 -29934
rect 8115 -30164 8157 -29976
rect 8157 -30164 8345 -29976
rect 8345 -30164 8387 -29976
rect 8115 -30206 8387 -30164
rect 9051 -29976 9323 -29934
rect 9051 -30164 9093 -29976
rect 9093 -30164 9281 -29976
rect 9281 -30164 9323 -29976
rect 9051 -30206 9323 -30164
rect 9982 -29976 10254 -29933
rect 9982 -30163 10024 -29976
rect 10024 -30163 10211 -29976
rect 10211 -30163 10254 -29976
rect 9982 -30205 10254 -30163
rect 10909 -29976 11181 -29934
rect 10909 -30164 10951 -29976
rect 10951 -30164 11139 -29976
rect 11139 -30164 11181 -29976
rect 10909 -30206 11181 -30164
rect 12157 -30487 12429 -30415
rect 12157 -30616 12228 -30487
rect 12228 -30616 12357 -30487
rect 12357 -30616 12429 -30487
rect 12157 -30687 12429 -30616
rect 12884 -30528 13156 -30456
rect 12884 -30657 12955 -30528
rect 12955 -30657 13084 -30528
rect 13084 -30657 13156 -30528
rect 12884 -30728 13156 -30657
rect 5624 -32989 5896 -32886
rect 5624 -33055 5727 -32989
rect 5727 -33055 5793 -32989
rect 5793 -33055 5896 -32989
rect 5624 -33158 5896 -33055
rect 6062 -32970 6334 -32867
rect 6062 -33036 6165 -32970
rect 6165 -33036 6231 -32970
rect 6231 -33036 6334 -32970
rect 6062 -33139 6334 -33036
rect 6502 -32961 6774 -32858
rect 6502 -33027 6605 -32961
rect 6605 -33027 6671 -32961
rect 6671 -33027 6774 -32961
rect 6502 -33130 6774 -33027
rect -11187 -33802 -10915 -33701
rect -11187 -33872 -11086 -33802
rect -11086 -33872 -11016 -33802
rect -11016 -33872 -10915 -33802
rect -11187 -33973 -10915 -33872
rect 7180 -34504 7452 -34462
rect 7180 -34692 7222 -34504
rect 7222 -34692 7410 -34504
rect 7410 -34692 7452 -34504
rect 7180 -34734 7452 -34692
rect 8115 -34504 8387 -34462
rect 8115 -34692 8157 -34504
rect 8157 -34692 8345 -34504
rect 8345 -34692 8387 -34504
rect 8115 -34734 8387 -34692
rect 9051 -34504 9323 -34462
rect 9051 -34692 9093 -34504
rect 9093 -34692 9281 -34504
rect 9281 -34692 9323 -34504
rect 9051 -34734 9323 -34692
rect 9982 -34504 10254 -34461
rect 9982 -34691 10024 -34504
rect 10024 -34691 10211 -34504
rect 10211 -34691 10254 -34504
rect 9982 -34733 10254 -34691
rect 10909 -34504 11181 -34462
rect 10909 -34692 10951 -34504
rect 10951 -34692 11139 -34504
rect 11139 -34692 11181 -34504
rect 10909 -34734 11181 -34692
rect 12157 -35015 12429 -34943
rect 12157 -35144 12228 -35015
rect 12228 -35144 12357 -35015
rect 12357 -35144 12429 -35015
rect 12157 -35215 12429 -35144
rect 12884 -35056 13156 -34984
rect 12884 -35185 12955 -35056
rect 12955 -35185 13084 -35056
rect 13084 -35185 13156 -35056
rect 12884 -35256 13156 -35185
rect 12462 -35950 12734 -35868
rect 12462 -36057 12544 -35950
rect 12544 -36057 12651 -35950
rect 12651 -36057 12734 -35950
rect 12462 -36140 12734 -36057
<< metal5 >>
rect -27804 4955 20350 6916
rect -27804 4683 2195 4955
rect 2467 4683 3801 4955
rect 4073 4953 20350 4955
rect 4073 4683 5505 4953
rect -27804 4681 5505 4683
rect 5777 4681 20350 4953
rect -27804 3366 20350 4681
rect -27804 3357 6502 3366
rect -27804 3338 6062 3357
rect -27804 3231 5624 3338
rect -27804 2959 -23504 3231
rect -23232 2959 -20213 3231
rect -19941 2959 -16922 3231
rect -16650 2959 -13631 3231
rect -13359 2959 -10340 3231
rect -10068 2959 -7050 3231
rect -6778 2959 -3759 3231
rect -3487 2959 -468 3231
rect -196 3066 5624 3231
rect 5896 3085 6062 3338
rect 6334 3094 6502 3357
rect 6774 3094 20350 3366
rect 6334 3085 20350 3094
rect 5896 3066 20350 3085
rect -196 2959 20350 3066
rect -27804 1763 20350 2959
rect -27804 1762 9982 1763
rect -27804 1490 7180 1762
rect 7452 1490 8115 1762
rect 8387 1490 9051 1762
rect 9323 1491 9982 1762
rect 10254 1762 20350 1763
rect 10254 1491 10909 1762
rect 9323 1490 10909 1491
rect 11181 1490 20350 1762
rect -27804 1447 20350 1490
rect -27804 1175 -24316 1447
rect -24044 1175 -22757 1447
rect -22485 1175 -21025 1447
rect -20753 1175 -19466 1447
rect -19194 1175 -17734 1447
rect -17462 1175 -16175 1447
rect -15903 1175 -14443 1447
rect -14171 1175 -12884 1447
rect -12612 1175 -11152 1447
rect -10880 1175 -9593 1447
rect -9321 1175 -7862 1447
rect -7590 1175 -6303 1447
rect -6031 1175 -4571 1447
rect -4299 1175 -3012 1447
rect -2740 1175 -1280 1447
rect -1008 1175 279 1447
rect 551 1281 20350 1447
rect 551 1175 12157 1281
rect -27804 1009 12157 1175
rect 12429 1240 20350 1281
rect 12429 1009 12884 1240
rect -27804 968 12884 1009
rect 13156 968 20350 1240
rect -27804 457 20350 968
rect -27804 221 -24336 457
rect -24001 355 -21045 457
rect -24001 221 -23205 355
rect -27804 83 -23205 221
rect -22933 333 -21045 355
rect -22933 83 -22343 333
rect -27804 61 -22343 83
rect -22071 221 -21045 333
rect -20710 355 -17754 457
rect -20710 221 -19914 355
rect -22071 83 -19914 221
rect -19642 333 -17754 355
rect -19642 83 -19052 333
rect -22071 61 -19052 83
rect -18780 221 -17754 333
rect -17419 355 -14463 457
rect -17419 221 -16623 355
rect -18780 83 -16623 221
rect -16351 333 -14463 355
rect -16351 83 -15761 333
rect -18780 61 -15761 83
rect -15489 221 -14463 333
rect -14128 355 -11172 457
rect -14128 221 -13332 355
rect -15489 83 -13332 221
rect -13060 333 -11172 355
rect -13060 83 -12470 333
rect -15489 61 -12470 83
rect -12198 221 -11172 333
rect -10837 355 -7882 457
rect -10837 221 -10041 355
rect -12198 83 -10041 221
rect -9769 333 -7882 355
rect -9769 83 -9179 333
rect -12198 61 -9179 83
rect -8907 221 -7882 333
rect -7547 355 -4591 457
rect -7547 221 -6751 355
rect -8907 83 -6751 221
rect -6479 333 -4591 355
rect -6479 83 -5889 333
rect -8907 61 -5889 83
rect -5617 221 -4591 333
rect -4256 355 -1300 457
rect -4256 221 -3460 355
rect -5617 83 -3460 221
rect -3188 333 -1300 355
rect -3188 83 -2598 333
rect -5617 61 -2598 83
rect -2326 221 -1300 333
rect -965 355 20350 457
rect -965 221 -169 355
rect -2326 83 -169 221
rect 103 333 20350 355
rect 103 83 693 333
rect -2326 61 693 83
rect 965 61 20350 333
rect -27804 -1162 20350 61
rect -27804 -1171 6502 -1162
rect -27804 -1190 6062 -1171
rect -27804 -1462 5624 -1190
rect 5896 -1443 6062 -1190
rect 6334 -1434 6502 -1171
rect 6774 -1434 20350 -1162
rect 6334 -1443 20350 -1434
rect 5896 -1462 20350 -1443
rect -27804 -2765 20350 -1462
rect -27804 -2766 9982 -2765
rect -27804 -2883 7180 -2766
rect -27804 -3191 -23987 -2883
rect -21717 -2914 7180 -2883
rect -21717 -3191 -20247 -2914
rect -27804 -3222 -20247 -3191
rect -17977 -3038 7180 -2914
rect 7452 -3038 8115 -2766
rect 8387 -3038 9051 -2766
rect 9323 -3037 9982 -2766
rect 10254 -2766 20350 -2765
rect 10254 -3037 10909 -2766
rect 9323 -3038 10909 -3037
rect 11181 -3038 20350 -2766
rect -17977 -3222 20350 -3038
rect -27804 -3247 20350 -3222
rect -27804 -3519 12157 -3247
rect 12429 -3288 20350 -3247
rect 12429 -3519 12884 -3288
rect -27804 -3560 12884 -3519
rect 13156 -3560 20350 -3288
rect -27804 -4612 20350 -3560
rect -27804 -4920 -24007 -4612
rect -21737 -4920 20350 -4612
rect -27804 -5113 20350 -4920
rect -27804 -5385 -20249 -5113
rect -19977 -5385 -18690 -5113
rect -18418 -5385 -16958 -5113
rect -16686 -5385 -15399 -5113
rect -15127 -5385 -13667 -5113
rect -13395 -5385 -12108 -5113
rect -11836 -5385 -10376 -5113
rect -10104 -5385 -8817 -5113
rect -8545 -5385 20350 -5113
rect -27804 -5590 20350 -5385
rect -27804 -5599 6502 -5590
rect -27804 -5618 6062 -5599
rect -27804 -5890 5624 -5618
rect 5896 -5871 6062 -5618
rect 6334 -5862 6502 -5599
rect 6774 -5862 20350 -5590
rect 6334 -5871 20350 -5862
rect 5896 -5890 20350 -5871
rect -27804 -5976 20350 -5890
rect -27804 -6284 -24008 -5976
rect -21738 -6103 20350 -5976
rect -21738 -6284 -20269 -6103
rect -27804 -6339 -20269 -6284
rect -19934 -6205 -16978 -6103
rect -19934 -6339 -19138 -6205
rect -27804 -6477 -19138 -6339
rect -18866 -6227 -16978 -6205
rect -18866 -6477 -18276 -6227
rect -27804 -6499 -18276 -6477
rect -18004 -6339 -16978 -6227
rect -16643 -6205 -13687 -6103
rect -16643 -6339 -15847 -6205
rect -18004 -6477 -15847 -6339
rect -15575 -6227 -13687 -6205
rect -15575 -6477 -14985 -6227
rect -18004 -6499 -14985 -6477
rect -14713 -6339 -13687 -6227
rect -13352 -6205 -10396 -6103
rect -13352 -6339 -12556 -6205
rect -14713 -6477 -12556 -6339
rect -12284 -6227 -10396 -6205
rect -12284 -6477 -11694 -6227
rect -14713 -6499 -11694 -6477
rect -11422 -6339 -10396 -6227
rect -10061 -6205 20350 -6103
rect -10061 -6339 -9265 -6205
rect -11422 -6477 -9265 -6339
rect -8993 -6227 20350 -6205
rect -8993 -6477 -8403 -6227
rect -11422 -6499 -8403 -6477
rect -8131 -6499 20350 -6227
rect -27804 -7193 20350 -6499
rect -27804 -7194 9982 -7193
rect -27804 -7466 7180 -7194
rect 7452 -7466 8115 -7194
rect 8387 -7466 9051 -7194
rect 9323 -7465 9982 -7194
rect 10254 -7194 20350 -7193
rect 10254 -7465 10909 -7194
rect 9323 -7466 10909 -7465
rect 11181 -7466 20350 -7194
rect -27804 -7675 20350 -7466
rect -27804 -7870 12157 -7675
rect -27804 -8178 -24046 -7870
rect -21776 -7947 12157 -7870
rect 12429 -7716 20350 -7675
rect 12429 -7947 12884 -7716
rect -21776 -7988 12884 -7947
rect 13156 -7988 20350 -7716
rect -21776 -8178 20350 -7988
rect -27804 -8378 20350 -8178
rect -27804 -8650 -20249 -8378
rect -19977 -8650 -18690 -8378
rect -18418 -8650 -16958 -8378
rect -16686 -8650 -15399 -8378
rect -15127 -8650 -13667 -8378
rect -13395 -8650 -12108 -8378
rect -11836 -8650 -10376 -8378
rect -10104 -8650 -8817 -8378
rect -8545 -8650 20350 -8378
rect -27804 -9248 20350 -8650
rect -27804 -9556 -24060 -9248
rect -21790 -9368 20350 -9248
rect -21790 -9556 -20269 -9368
rect -27804 -9604 -20269 -9556
rect -19934 -9470 -16978 -9368
rect -19934 -9604 -19138 -9470
rect -27804 -9742 -19138 -9604
rect -18866 -9492 -16978 -9470
rect -18866 -9742 -18276 -9492
rect -27804 -9764 -18276 -9742
rect -18004 -9604 -16978 -9492
rect -16643 -9470 -13687 -9368
rect -16643 -9604 -15847 -9470
rect -18004 -9742 -15847 -9604
rect -15575 -9492 -13687 -9470
rect -15575 -9742 -14985 -9492
rect -18004 -9764 -14985 -9742
rect -14713 -9604 -13687 -9492
rect -13352 -9470 -10396 -9368
rect -13352 -9604 -12556 -9470
rect -14713 -9742 -12556 -9604
rect -12284 -9492 -10396 -9470
rect -12284 -9742 -11694 -9492
rect -14713 -9764 -11694 -9742
rect -11422 -9604 -10396 -9492
rect -10061 -9470 20350 -9368
rect -10061 -9604 -9265 -9470
rect -11422 -9742 -9265 -9604
rect -8993 -9492 20350 -9470
rect -8993 -9742 -8403 -9492
rect -11422 -9764 -8403 -9742
rect -8131 -9764 20350 -9492
rect -27804 -10218 20350 -9764
rect -27804 -10227 6502 -10218
rect -27804 -10246 6062 -10227
rect -27804 -10518 5624 -10246
rect 5896 -10499 6062 -10246
rect 6334 -10490 6502 -10227
rect 6774 -10490 20350 -10218
rect 6334 -10499 20350 -10490
rect 5896 -10518 20350 -10499
rect -27804 -11202 20350 -10518
rect -27804 -11510 -24018 -11202
rect -21748 -11510 20350 -11202
rect -27804 -11642 20350 -11510
rect -27804 -11914 -20249 -11642
rect -19977 -11914 -18690 -11642
rect -18418 -11914 -16958 -11642
rect -16686 -11914 -15399 -11642
rect -15127 -11914 -13667 -11642
rect -13395 -11914 -12108 -11642
rect -11836 -11914 -10376 -11642
rect -10104 -11914 -8817 -11642
rect -8545 -11821 20350 -11642
rect -8545 -11822 9982 -11821
rect -8545 -11914 7180 -11822
rect -27804 -12094 7180 -11914
rect 7452 -12094 8115 -11822
rect 8387 -12094 9051 -11822
rect 9323 -12093 9982 -11822
rect 10254 -11822 20350 -11821
rect 10254 -12093 10909 -11822
rect 9323 -12094 10909 -12093
rect 11181 -12094 20350 -11822
rect -27804 -12303 20350 -12094
rect -27804 -12535 12157 -12303
rect -27804 -12843 -24029 -12535
rect -21759 -12575 12157 -12535
rect 12429 -12344 20350 -12303
rect 12429 -12575 12884 -12344
rect -21759 -12616 12884 -12575
rect 13156 -12616 20350 -12344
rect -21759 -12632 20350 -12616
rect -21759 -12843 -20269 -12632
rect -27804 -12868 -20269 -12843
rect -19934 -12734 -16978 -12632
rect -19934 -12868 -19138 -12734
rect -27804 -13006 -19138 -12868
rect -18866 -12756 -16978 -12734
rect -18866 -13006 -18276 -12756
rect -27804 -13028 -18276 -13006
rect -18004 -12868 -16978 -12756
rect -16643 -12734 -13687 -12632
rect -16643 -12868 -15847 -12734
rect -18004 -13006 -15847 -12868
rect -15575 -12756 -13687 -12734
rect -15575 -13006 -14985 -12756
rect -18004 -13028 -14985 -13006
rect -14713 -12868 -13687 -12756
rect -13352 -12734 -10396 -12632
rect -13352 -12868 -12556 -12734
rect -14713 -13006 -12556 -12868
rect -12284 -12756 -10396 -12734
rect -12284 -13006 -11694 -12756
rect -14713 -13028 -11694 -13006
rect -11422 -12868 -10396 -12756
rect -10061 -12734 20350 -12632
rect -10061 -12868 -9265 -12734
rect -11422 -13006 -9265 -12868
rect -8993 -12756 20350 -12734
rect -8993 -13006 -8403 -12756
rect -11422 -13028 -8403 -13006
rect -8131 -13028 20350 -12756
rect -27804 -13986 20350 -13028
rect -27804 -14163 -1376 -13986
rect -27804 -14435 -4092 -14163
rect -3820 -14258 -1376 -14163
rect -1104 -14258 20350 -13986
rect -3820 -14435 20350 -14258
rect -27804 -14719 20350 -14435
rect -27804 -14965 -11187 -14719
rect -27804 -15285 -23531 -14965
rect -23211 -14991 -11187 -14965
rect -10915 -14746 20350 -14719
rect -10915 -14755 6502 -14746
rect -10915 -14774 6062 -14755
rect -10915 -14796 5624 -14774
rect -10915 -14991 -4092 -14796
rect -23211 -15068 -4092 -14991
rect -3820 -14805 5624 -14796
rect -3820 -15068 -1376 -14805
rect -23211 -15077 -1376 -15068
rect -1104 -15046 5624 -14805
rect 5896 -15027 6062 -14774
rect 6334 -15018 6502 -14755
rect 6774 -15018 20350 -14746
rect 6334 -15027 20350 -15018
rect 5896 -15046 20350 -15027
rect -1104 -15077 20350 -15046
rect -23211 -15196 20350 -15077
rect -23211 -15285 -17039 -15196
rect -27804 -15516 -17039 -15285
rect -16719 -15281 20350 -15196
rect -16719 -15516 -7320 -15281
rect -27804 -15601 -7320 -15516
rect -7000 -15601 20350 -15281
rect -27804 -15615 20350 -15601
rect -27804 -15774 -4092 -15615
rect -27804 -16094 -7327 -15774
rect -7007 -15887 -4092 -15774
rect -3820 -15624 20350 -15615
rect -3820 -15887 -1376 -15624
rect -7007 -15896 -1376 -15887
rect -1104 -15896 20350 -15624
rect -7007 -16094 20350 -15896
rect -27804 -16161 20350 -16094
rect -27804 -16481 -23488 -16161
rect -23168 -16260 20350 -16161
rect -23168 -16481 -7328 -16260
rect -27804 -16580 -7328 -16481
rect -7008 -16349 20350 -16260
rect -7008 -16350 9982 -16349
rect -7008 -16434 7180 -16350
rect -7008 -16580 -4092 -16434
rect -27804 -16602 -4092 -16580
rect -27804 -16922 -17039 -16602
rect -16719 -16706 -4092 -16602
rect -3820 -16443 7180 -16434
rect -3820 -16706 -1376 -16443
rect -16719 -16715 -1376 -16706
rect -1104 -16622 7180 -16443
rect 7452 -16622 8115 -16350
rect 8387 -16622 9051 -16350
rect 9323 -16621 9982 -16350
rect 10254 -16350 20350 -16349
rect 10254 -16621 10909 -16350
rect 9323 -16622 10909 -16621
rect 11181 -16622 20350 -16350
rect -1104 -16715 20350 -16622
rect -16719 -16730 20350 -16715
rect -16719 -16767 16278 -16730
rect -16719 -16922 -7332 -16767
rect -27804 -17087 -7332 -16922
rect -7012 -16831 16278 -16767
rect -7012 -17087 12157 -16831
rect -27804 -17103 12157 -17087
rect 12429 -16872 16278 -16831
rect 12429 -17103 12884 -16872
rect -27804 -17144 12884 -17103
rect 13156 -17002 16278 -16872
rect 16550 -17002 20350 -16730
rect 13156 -17144 20350 -17002
rect -27804 -17242 20350 -17144
rect -27804 -17373 -7331 -17242
rect -27804 -17693 -23479 -17373
rect -23159 -17535 -7331 -17373
rect -23159 -17693 -11185 -17535
rect -27804 -17807 -11185 -17693
rect -10913 -17562 -7331 -17535
rect -7011 -17253 20350 -17242
rect -7011 -17525 -4092 -17253
rect -3820 -17262 20350 -17253
rect -3820 -17525 -1376 -17262
rect -7011 -17534 -1376 -17525
rect -1104 -17534 20350 -17262
rect -7011 -17562 20350 -17534
rect -10913 -17694 20350 -17562
rect -10913 -17807 -7326 -17694
rect -27804 -17840 -7326 -17807
rect -27804 -17969 -15168 -17840
rect -27804 -18289 -20759 -17969
rect -20439 -18033 -15168 -17969
rect -20439 -18289 -17170 -18033
rect -27804 -18353 -17170 -18289
rect -16850 -18160 -15168 -18033
rect -14848 -18014 -7326 -17840
rect -7006 -18014 20350 -17694
rect -14848 -18072 20350 -18014
rect -14848 -18136 -4092 -18072
rect -14848 -18160 -7326 -18136
rect -16850 -18333 -7326 -18160
rect -16850 -18353 -15175 -18333
rect -27804 -18462 -15175 -18353
rect -27804 -18514 -20766 -18462
rect -27804 -18834 -23471 -18514
rect -23151 -18782 -20766 -18514
rect -20446 -18653 -15175 -18462
rect -14855 -18456 -7326 -18333
rect -7006 -18344 -4092 -18136
rect -3820 -18081 20350 -18072
rect -3820 -18344 -1376 -18081
rect -7006 -18353 -1376 -18344
rect -1104 -18353 20350 -18081
rect -7006 -18456 20350 -18353
rect -14855 -18617 20350 -18456
rect -14855 -18653 -7332 -18617
rect -20446 -18782 -7332 -18653
rect -23151 -18819 -7332 -18782
rect -23151 -18834 -15176 -18819
rect -27804 -18948 -15176 -18834
rect -27804 -19268 -20767 -18948
rect -20447 -19139 -15176 -18948
rect -14856 -18937 -7332 -18819
rect -7012 -18768 20350 -18617
rect -7012 -18891 17877 -18768
rect -7012 -18937 -4092 -18891
rect -14856 -19139 -4092 -18937
rect -20447 -19163 -4092 -19139
rect -3820 -18900 17877 -18891
rect -3820 -19163 -1376 -18900
rect -20447 -19172 -1376 -19163
rect -1104 -19040 17877 -18900
rect 18149 -19040 20350 -18768
rect -1104 -19172 20350 -19040
rect -20447 -19268 20350 -19172
rect -27804 -19274 20350 -19268
rect -27804 -19283 6502 -19274
rect -27804 -19302 6062 -19283
rect -27804 -19326 5624 -19302
rect -27804 -19455 -15180 -19326
rect -27804 -19686 -20771 -19455
rect -27804 -20006 -23448 -19686
rect -23128 -19775 -20771 -19686
rect -20451 -19488 -15180 -19455
rect -20451 -19775 -17055 -19488
rect -23128 -19808 -17055 -19775
rect -16735 -19646 -15180 -19488
rect -14860 -19574 5624 -19326
rect 5896 -19555 6062 -19302
rect 6334 -19546 6502 -19283
rect 6774 -19546 20350 -19274
rect 6334 -19555 20350 -19546
rect 5896 -19574 20350 -19555
rect -14860 -19646 20350 -19574
rect -16735 -19710 20350 -19646
rect -16735 -19801 -4092 -19710
rect -16735 -19808 -15179 -19801
rect -23128 -19930 -15179 -19808
rect -23128 -20006 -20770 -19930
rect -27804 -20250 -20770 -20006
rect -20450 -20121 -15179 -19930
rect -14859 -19982 -4092 -19801
rect -3820 -19719 20350 -19710
rect -3820 -19982 -1376 -19719
rect -14859 -19991 -1376 -19982
rect -1104 -19991 20350 -19719
rect -14859 -20121 20350 -19991
rect -20450 -20170 20350 -20121
rect -20450 -20250 16220 -20170
rect -27804 -20253 16220 -20250
rect -27804 -20382 -15174 -20253
rect -27804 -20702 -20765 -20382
rect -20445 -20573 -15174 -20382
rect -14854 -20352 16220 -20253
rect -14854 -20492 -1376 -20352
rect -14854 -20573 -11185 -20492
rect -20445 -20695 -11185 -20573
rect -20445 -20702 -15174 -20695
rect -27804 -20824 -15174 -20702
rect -27804 -20884 -20765 -20824
rect -27804 -21204 -23439 -20884
rect -23119 -21144 -20765 -20884
rect -20445 -20884 -15174 -20824
rect -20445 -21144 -17045 -20884
rect -23119 -21204 -17045 -21144
rect -16725 -21015 -15174 -20884
rect -14854 -20764 -11185 -20695
rect -10913 -20529 -1376 -20492
rect -10913 -20764 -4092 -20529
rect -14854 -20801 -4092 -20764
rect -3820 -20624 -1376 -20529
rect -1104 -20442 16220 -20352
rect 16492 -20442 20350 -20170
rect -1104 -20624 20350 -20442
rect -3820 -20801 20350 -20624
rect -14854 -20877 20350 -20801
rect -14854 -20878 9982 -20877
rect -14854 -21015 7180 -20878
rect -16725 -21150 7180 -21015
rect 7452 -21150 8115 -20878
rect 8387 -21150 9051 -20878
rect 9323 -21149 9982 -20878
rect 10254 -20878 20350 -20877
rect 10254 -21149 10909 -20878
rect 9323 -21150 10909 -21149
rect 11181 -21150 20350 -20878
rect -16725 -21176 20350 -21150
rect -16725 -21204 -15180 -21176
rect -27804 -21305 -15180 -21204
rect -27804 -21625 -20771 -21305
rect -20451 -21496 -15180 -21305
rect -14860 -21359 20350 -21176
rect -14860 -21496 12157 -21359
rect -20451 -21625 12157 -21496
rect -27804 -21631 12157 -21625
rect 12429 -21400 20350 -21359
rect 12429 -21631 12884 -21400
rect -27804 -21672 12884 -21631
rect 13156 -21672 20350 -21400
rect -27804 -21855 20350 -21672
rect -27804 -22175 -16854 -21855
rect -16534 -22175 20350 -21855
rect -27804 -22178 20350 -22175
rect -27804 -22498 -23442 -22178
rect -23122 -22498 20350 -22178
rect -27804 -23071 20350 -22498
rect -27804 -23246 -11185 -23071
rect -27804 -23494 -16809 -23246
rect -27804 -23814 -23482 -23494
rect -23162 -23566 -16809 -23494
rect -16489 -23343 -11185 -23246
rect -10913 -23343 20350 -23071
rect -16489 -23566 20350 -23343
rect -23162 -23802 20350 -23566
rect -23162 -23811 6502 -23802
rect -23162 -23814 6062 -23811
rect -27804 -23830 6062 -23814
rect -27804 -24102 5624 -23830
rect 5896 -24083 6062 -23830
rect 6334 -24074 6502 -23811
rect 6774 -24074 20350 -23802
rect 6334 -24083 20350 -24074
rect 5896 -24102 20350 -24083
rect -27804 -24652 20350 -24102
rect -27804 -24972 -16811 -24652
rect -16491 -24972 20350 -24652
rect -27804 -25405 20350 -24972
rect -27804 -25406 9982 -25405
rect -27804 -25678 7180 -25406
rect 7452 -25678 8115 -25406
rect 8387 -25678 9051 -25406
rect 9323 -25677 9982 -25406
rect 10254 -25406 20350 -25405
rect 10254 -25677 10909 -25406
rect 9323 -25678 10909 -25677
rect 11181 -25678 20350 -25406
rect -27804 -25839 20350 -25678
rect -27804 -26111 -11185 -25839
rect -10913 -25887 20350 -25839
rect -10913 -26111 12157 -25887
rect -27804 -26159 12157 -26111
rect 12429 -25928 20350 -25887
rect 12429 -26159 12884 -25928
rect -27804 -26200 12884 -26159
rect 13156 -26200 20350 -25928
rect -27804 -28330 20350 -26200
rect -27804 -28339 6502 -28330
rect -27804 -28358 6062 -28339
rect -27804 -28472 5624 -28358
rect -27804 -28744 -11185 -28472
rect -10913 -28630 5624 -28472
rect 5896 -28611 6062 -28358
rect 6334 -28602 6502 -28339
rect 6774 -28602 20350 -28330
rect 6334 -28611 20350 -28602
rect 5896 -28630 20350 -28611
rect -10913 -28744 20350 -28630
rect -27804 -29933 20350 -28744
rect -27804 -29934 9982 -29933
rect -27804 -30206 7180 -29934
rect 7452 -30206 8115 -29934
rect 8387 -30206 9051 -29934
rect 9323 -30205 9982 -29934
rect 10254 -29934 20350 -29933
rect 10254 -30205 10909 -29934
rect 9323 -30206 10909 -30205
rect 11181 -30206 20350 -29934
rect -27804 -30415 20350 -30206
rect -27804 -30687 12157 -30415
rect 12429 -30456 20350 -30415
rect 12429 -30687 12884 -30456
rect -27804 -30728 12884 -30687
rect 13156 -30728 20350 -30456
rect -27804 -31081 20350 -30728
rect -27804 -31353 -11185 -31081
rect -10913 -31353 20350 -31081
rect -27804 -32858 20350 -31353
rect -27804 -32867 6502 -32858
rect -27804 -32886 6062 -32867
rect -27804 -33158 5624 -32886
rect 5896 -33139 6062 -32886
rect 6334 -33130 6502 -32867
rect 6774 -33130 20350 -32858
rect 6334 -33139 20350 -33130
rect 5896 -33158 20350 -33139
rect -27804 -33701 20350 -33158
rect -27804 -33973 -11187 -33701
rect -10915 -33973 20350 -33701
rect -27804 -34461 20350 -33973
rect -27804 -34462 9982 -34461
rect -27804 -34734 7180 -34462
rect 7452 -34734 8115 -34462
rect 8387 -34734 9051 -34462
rect 9323 -34733 9982 -34462
rect 10254 -34462 20350 -34461
rect 10254 -34733 10909 -34462
rect 9323 -34734 10909 -34733
rect 11181 -34734 20350 -34462
rect -27804 -34943 20350 -34734
rect -27804 -35215 12157 -34943
rect 12429 -34984 20350 -34943
rect 12429 -35215 12884 -34984
rect -27804 -35256 12884 -35215
rect 13156 -35256 20350 -34984
rect -27804 -35868 20350 -35256
rect -27804 -36140 12462 -35868
rect 12734 -36140 20350 -35868
rect -27804 -37316 20350 -36140
<< labels >>
flabel metal3 -24908 -15649 -24849 -15604 0 FreeSans 800 0 0 0 B0
port 0 nsew
flabel metal3 -24899 -16827 -24840 -16782 0 FreeSans 800 0 0 0 B1
port 1 nsew
flabel metal3 -24910 -18036 -24851 -17991 0 FreeSans 800 0 0 0 B2
port 2 nsew
flabel metal3 -24840 -19162 -24781 -19117 0 FreeSans 800 0 0 0 B3
port 3 nsew
flabel metal3 -24887 -20352 -24828 -20307 0 FreeSans 800 0 0 0 B4
port 4 nsew
flabel metal3 -24879 -21556 -24820 -21511 0 FreeSans 800 0 0 0 B5
port 5 nsew
flabel metal3 -24879 -22857 -24820 -22812 0 FreeSans 800 0 0 0 B6
port 6 nsew
flabel metal3 -24878 -15812 -24819 -15767 0 FreeSans 800 0 0 0 A0
port 8 nsew
flabel metal3 -24898 -16988 -24839 -16943 0 FreeSans 800 0 0 0 A1
port 9 nsew
flabel metal3 -24905 -18196 -24846 -18151 0 FreeSans 800 0 0 0 A2
port 10 nsew
flabel metal3 -24846 -19319 -24787 -19274 0 FreeSans 800 0 0 0 A3
port 11 nsew
flabel metal3 -24884 -20512 -24825 -20467 0 FreeSans 800 0 0 0 A4
port 12 nsew
flabel metal3 -24902 -21706 -24843 -21661 0 FreeSans 800 0 0 0 A5
port 13 nsew
flabel metal3 -24888 -23019 -24829 -22974 0 FreeSans 800 0 0 0 A6
port 15 nsew
flabel metal3 -24885 -24327 -24826 -24282 0 FreeSans 800 0 0 0 A7
port 16 nsew
flabel metal1 13169 -3047 13216 -2964 0 FreeSans 800 0 0 0 Y0
port 17 nsew
flabel metal1 13172 -7413 13219 -7330 0 FreeSans 800 0 0 0 Y1
port 18 nsew
flabel metal1 13183 -12104 13230 -12021 0 FreeSans 800 0 0 0 Y2
port 20 nsew
flabel metal1 13178 -16546 13225 -16463 0 FreeSans 800 0 0 0 Y3
port 21 nsew
flabel metal1 13181 -21117 13228 -21034 0 FreeSans 800 0 0 0 Y4
port 22 nsew
flabel metal1 13179 -25614 13226 -25531 0 FreeSans 800 0 0 0 Y5
port 23 nsew
flabel metal1 13178 -30106 13225 -30058 0 FreeSans 800 0 0 0 Y6
port 24 nsew
flabel metal1 13035 -36363 13082 -36280 0 FreeSans 800 0 0 0 S
port 26 nsew
flabel metal1 18354 -18573 18391 -18471 0 FreeSans 800 0 0 0 Z
port 27 nsew
flabel metal1 13152 1469 13208 1558 0 FreeSans 800 0 0 0 C
port 28 nsew
flabel metal1 8026 5020 8106 5116 0 FreeSans 1600 0 0 0 V
port 29 nsew
flabel metal5 8982 4290 9670 4732 0 FreeSans 1600 0 0 0 VSS
port 32 nsew
flabel metal1 13172 -34752 13202 -34724 0 FreeSans 1600 0 0 0 Y7
port 34 nsew
flabel metal3 -25060 -24176 -24986 -24108 0 FreeSans 1600 0 0 0 B7
port 36 nsew
flabel metal2 6442 4066 6500 4126 0 FreeSans 160 0 0 0 SEL0
port 39 nsew
flabel metal2 6010 4070 6050 4099 0 FreeSans 160 0 0 0 SEL1
port 40 nsew
flabel metal2 5574 4072 5614 4099 0 FreeSans 160 0 0 0 SEL2
port 41 nsew
flabel metal2 5360 4068 5400 4114 0 FreeSans 160 0 0 0 SEL3
port 42 nsew
flabel metal4 5770 4214 6082 4324 0 FreeSans 1600 0 0 0 VDD
port 43 nsew
flabel metal1 -17948 -25417 -17920 -25375 0 FreeSans 160 0 0 0 OR8_0.A7
flabel metal1 -17952 -24045 -17924 -24003 0 FreeSans 160 0 0 0 OR8_0.A6
flabel metal1 -17944 -22655 -17916 -22613 0 FreeSans 160 0 0 0 OR8_0.A5
flabel metal1 -17948 -21233 -17920 -21191 0 FreeSans 160 0 0 0 OR8_0.A4
flabel metal1 -17944 -19837 -17916 -19795 0 FreeSans 160 0 0 0 OR8_0.A3
flabel metal1 -17944 -18449 -17916 -18407 0 FreeSans 160 0 0 0 OR8_0.A2
flabel metal1 -17950 -17041 -17922 -16999 0 FreeSans 160 0 0 0 OR8_0.A1
flabel metal1 -17948 -15645 -17920 -15603 0 FreeSans 160 0 0 0 OR8_0.A0
flabel metal1 -17950 -15779 -17922 -15737 0 FreeSans 160 0 0 0 OR8_0.B0
flabel metal1 -17950 -17171 -17922 -17129 0 FreeSans 160 0 0 0 OR8_0.B1
flabel metal1 -17944 -18569 -17916 -18527 0 FreeSans 160 0 0 0 OR8_0.B2
flabel metal1 -17944 -19951 -17916 -19909 0 FreeSans 160 0 0 0 OR8_0.B3
flabel metal1 -17948 -21327 -17920 -21285 0 FreeSans 160 0 0 0 OR8_0.B4
flabel metal1 -17944 -22761 -17916 -22719 0 FreeSans 160 0 0 0 OR8_0.B5
flabel metal1 -17952 -24153 -17924 -24111 0 FreeSans 160 0 0 0 OR8_0.B6
flabel metal1 -17948 -25531 -17920 -25489 0 FreeSans 160 0 0 0 OR8_0.B7
flabel metal1 -14796 -17849 -14764 -17815 0 FreeSans 160 0 0 0 OR8_0.S0
flabel metal1 -14794 -18349 -14762 -18315 0 FreeSans 160 0 0 0 OR8_0.S1
flabel metal1 -14796 -18829 -14764 -18795 0 FreeSans 160 0 0 0 OR8_0.S2
flabel metal1 -14796 -19329 -14764 -19295 0 FreeSans 160 0 0 0 OR8_0.S3
flabel metal1 -14796 -19809 -14764 -19775 0 FreeSans 160 0 0 0 OR8_0.S4
flabel metal1 -14796 -20269 -14764 -20235 0 FreeSans 160 0 0 0 OR8_0.S5
flabel metal1 -14796 -20729 -14764 -20695 0 FreeSans 160 0 0 0 OR8_0.S6
flabel metal1 -14796 -21209 -14764 -21175 0 FreeSans 160 0 0 0 OR8_0.S7
flabel metal4 -18090 -25135 -18004 -25051 0 FreeSans 1600 0 0 0 OR8_0.VDD
flabel metal5 -15070 -21387 -14968 -21287 0 FreeSans 1600 0 0 0 OR8_0.VSS
rlabel metal1 -14797 -17851 -14764 -17816 7 OR8_0.NOT8_0.S0
rlabel metal1 -14804 -18350 -14771 -18315 7 OR8_0.NOT8_0.S1
rlabel metal1 -14797 -18829 -14764 -18794 7 OR8_0.NOT8_0.S2
rlabel metal1 -14796 -19329 -14763 -19294 7 OR8_0.NOT8_0.S3
rlabel metal1 -14796 -19809 -14763 -19774 7 OR8_0.NOT8_0.S4
rlabel metal1 -14796 -20268 -14763 -20233 7 OR8_0.NOT8_0.S5
rlabel metal1 -14796 -20729 -14763 -20694 7 OR8_0.NOT8_0.S6
rlabel metal1 -14797 -21209 -14764 -21174 7 OR8_0.NOT8_0.S7
rlabel metal1 -16394 -18210 -16347 -18159 3 OR8_0.NOT8_0.A0
rlabel metal1 -16396 -18710 -16349 -18659 3 OR8_0.NOT8_0.A1
rlabel metal1 -16397 -19191 -16350 -19140 3 OR8_0.NOT8_0.A2
rlabel metal1 -16396 -19690 -16349 -19639 3 OR8_0.NOT8_0.A3
rlabel metal1 -16395 -20171 -16348 -20120 3 OR8_0.NOT8_0.A4
rlabel metal1 -16394 -20631 -16347 -20580 3 OR8_0.NOT8_0.A5
rlabel metal1 -16397 -21090 -16350 -21039 3 OR8_0.NOT8_0.A6
rlabel metal1 -16397 -21571 -16350 -21520 3 OR8_0.NOT8_0.A7
flabel metal4 -16385 -19395 -16315 -19297 0 FreeSans 160 0 0 0 OR8_0.NOT8_0.VDD
flabel metal5 -14847 -19245 -14777 -19147 0 FreeSans 160 0 0 0 OR8_0.NOT8_0.VSS
rlabel metal1 -15723 -18219 -15723 -18219 1 OR8_0.NOT8_0.inv_7.A
rlabel metal1 -15334 -18021 -15334 -18021 3 OR8_0.NOT8_0.inv_7.VSS
rlabel metal1 -16131 -18009 -16131 -18009 3 OR8_0.NOT8_0.inv_7.VDD
rlabel metal1 -15723 -17807 -15723 -17807 1 OR8_0.NOT8_0.inv_7.Y
rlabel metal1 -15722 -18719 -15722 -18719 1 OR8_0.NOT8_0.inv_6.A
rlabel metal1 -15333 -18521 -15333 -18521 3 OR8_0.NOT8_0.inv_6.VSS
rlabel metal1 -16130 -18509 -16130 -18509 3 OR8_0.NOT8_0.inv_6.VDD
rlabel metal1 -15722 -18307 -15722 -18307 1 OR8_0.NOT8_0.inv_6.Y
rlabel metal1 -15723 -19199 -15723 -19199 1 OR8_0.NOT8_0.inv_5.A
rlabel metal1 -15334 -19001 -15334 -19001 3 OR8_0.NOT8_0.inv_5.VSS
rlabel metal1 -16131 -18989 -16131 -18989 3 OR8_0.NOT8_0.inv_5.VDD
rlabel metal1 -15723 -18787 -15723 -18787 1 OR8_0.NOT8_0.inv_5.Y
rlabel metal1 -15723 -20179 -15723 -20179 1 OR8_0.NOT8_0.inv_4.A
rlabel metal1 -15334 -19981 -15334 -19981 3 OR8_0.NOT8_0.inv_4.VSS
rlabel metal1 -16131 -19969 -16131 -19969 3 OR8_0.NOT8_0.inv_4.VDD
rlabel metal1 -15723 -19767 -15723 -19767 1 OR8_0.NOT8_0.inv_4.Y
rlabel metal1 -15723 -20639 -15723 -20639 1 OR8_0.NOT8_0.inv_3.A
rlabel metal1 -15334 -20441 -15334 -20441 3 OR8_0.NOT8_0.inv_3.VSS
rlabel metal1 -16131 -20429 -16131 -20429 3 OR8_0.NOT8_0.inv_3.VDD
rlabel metal1 -15723 -20227 -15723 -20227 1 OR8_0.NOT8_0.inv_3.Y
rlabel metal1 -15737 -21099 -15737 -21099 1 OR8_0.NOT8_0.inv_2.A
rlabel metal1 -15348 -20901 -15348 -20901 3 OR8_0.NOT8_0.inv_2.VSS
rlabel metal1 -16145 -20889 -16145 -20889 3 OR8_0.NOT8_0.inv_2.VDD
rlabel metal1 -15737 -20687 -15737 -20687 1 OR8_0.NOT8_0.inv_2.Y
rlabel metal1 -15735 -21579 -15735 -21579 1 OR8_0.NOT8_0.inv_1.A
rlabel metal1 -15346 -21381 -15346 -21381 3 OR8_0.NOT8_0.inv_1.VSS
rlabel metal1 -16143 -21369 -16143 -21369 3 OR8_0.NOT8_0.inv_1.VDD
rlabel metal1 -15735 -21167 -15735 -21167 1 OR8_0.NOT8_0.inv_1.Y
rlabel metal1 -15723 -19699 -15723 -19699 1 OR8_0.NOT8_0.inv_0.A
rlabel metal1 -15334 -19501 -15334 -19501 3 OR8_0.NOT8_0.inv_0.VSS
rlabel metal1 -16131 -19489 -16131 -19489 3 OR8_0.NOT8_0.inv_0.VDD
rlabel metal1 -15723 -19287 -15723 -19287 1 OR8_0.NOT8_0.inv_0.Y
flabel metal1 -17380 -16946 -17328 -16869 7 FreeSerif 320 0 0 0 OR8_0.nor2_7.A
rlabel metal1 -17828 -16700 -17828 -16700 3 OR8_0.nor2_7.VDD
flabel metal1 -17274 -16945 -17222 -16868 7 FreeSerif 320 0 0 0 OR8_0.nor2_7.B
flabel metal1 -17268 -15941 -17216 -15864 7 FreeSerif 320 0 0 0 OR8_0.nor2_7.Y
rlabel metal1 -16850 -16404 -16850 -16404 3 OR8_0.nor2_7.VSS
flabel metal1 -17380 -18346 -17328 -18269 7 FreeSerif 320 0 0 0 OR8_0.nor2_6.A
rlabel metal1 -17828 -18100 -17828 -18100 3 OR8_0.nor2_6.VDD
flabel metal1 -17274 -18345 -17222 -18268 7 FreeSerif 320 0 0 0 OR8_0.nor2_6.B
flabel metal1 -17268 -17341 -17216 -17264 7 FreeSerif 320 0 0 0 OR8_0.nor2_6.Y
rlabel metal1 -16850 -17804 -16850 -17804 3 OR8_0.nor2_6.VSS
flabel metal1 -17380 -19746 -17328 -19669 7 FreeSerif 320 0 0 0 OR8_0.nor2_5.A
rlabel metal1 -17828 -19500 -17828 -19500 3 OR8_0.nor2_5.VDD
flabel metal1 -17274 -19745 -17222 -19668 7 FreeSerif 320 0 0 0 OR8_0.nor2_5.B
flabel metal1 -17268 -18741 -17216 -18664 7 FreeSerif 320 0 0 0 OR8_0.nor2_5.Y
rlabel metal1 -16850 -19204 -16850 -19204 3 OR8_0.nor2_5.VSS
flabel metal1 -17380 -21146 -17328 -21069 7 FreeSerif 320 0 0 0 OR8_0.nor2_4.A
rlabel metal1 -17828 -20900 -17828 -20900 3 OR8_0.nor2_4.VDD
flabel metal1 -17274 -21145 -17222 -21068 7 FreeSerif 320 0 0 0 OR8_0.nor2_4.B
flabel metal1 -17268 -20141 -17216 -20064 7 FreeSerif 320 0 0 0 OR8_0.nor2_4.Y
rlabel metal1 -16850 -20604 -16850 -20604 3 OR8_0.nor2_4.VSS
flabel metal1 -17380 -22546 -17328 -22469 7 FreeSerif 320 0 0 0 OR8_0.nor2_3.A
rlabel metal1 -17828 -22300 -17828 -22300 3 OR8_0.nor2_3.VDD
flabel metal1 -17274 -22545 -17222 -22468 7 FreeSerif 320 0 0 0 OR8_0.nor2_3.B
flabel metal1 -17268 -21541 -17216 -21464 7 FreeSerif 320 0 0 0 OR8_0.nor2_3.Y
rlabel metal1 -16850 -22004 -16850 -22004 3 OR8_0.nor2_3.VSS
flabel metal1 -17380 -23946 -17328 -23869 7 FreeSerif 320 0 0 0 OR8_0.nor2_2.A
rlabel metal1 -17828 -23700 -17828 -23700 3 OR8_0.nor2_2.VDD
flabel metal1 -17274 -23945 -17222 -23868 7 FreeSerif 320 0 0 0 OR8_0.nor2_2.B
flabel metal1 -17268 -22941 -17216 -22864 7 FreeSerif 320 0 0 0 OR8_0.nor2_2.Y
rlabel metal1 -16850 -23404 -16850 -23404 3 OR8_0.nor2_2.VSS
flabel metal1 -17380 -25346 -17328 -25269 7 FreeSerif 320 0 0 0 OR8_0.nor2_1.A
rlabel metal1 -17828 -25100 -17828 -25100 3 OR8_0.nor2_1.VDD
flabel metal1 -17274 -25345 -17222 -25268 7 FreeSerif 320 0 0 0 OR8_0.nor2_1.B
flabel metal1 -17268 -24341 -17216 -24264 7 FreeSerif 320 0 0 0 OR8_0.nor2_1.Y
rlabel metal1 -16850 -24804 -16850 -24804 3 OR8_0.nor2_1.VSS
flabel metal1 -17380 -15546 -17328 -15469 7 FreeSerif 320 0 0 0 OR8_0.nor2_0.A
rlabel metal1 -17828 -15300 -17828 -15300 3 OR8_0.nor2_0.VDD
flabel metal1 -17274 -15545 -17222 -15468 7 FreeSerif 320 0 0 0 OR8_0.nor2_0.B
flabel metal1 -17268 -14541 -17216 -14464 7 FreeSerif 320 0 0 0 OR8_0.nor2_0.Y
rlabel metal1 -16850 -15004 -16850 -15004 3 OR8_0.nor2_0.VSS
flabel metal1 -24917 -24332 -24855 -24296 0 FreeSans 160 0 0 0 AND8_0.A7
flabel metal1 -24925 -24162 -24863 -24126 0 FreeSans 160 0 0 0 AND8_0.B7
flabel metal1 -24917 -23012 -24855 -22976 0 FreeSans 160 0 0 0 AND8_0.A6
flabel metal1 -24921 -22848 -24859 -22812 0 FreeSans 160 0 0 0 AND8_0.B6
flabel metal1 -24921 -21716 -24859 -21680 0 FreeSans 160 0 0 0 AND8_0.A5
flabel metal1 -24921 -21550 -24859 -21514 0 FreeSans 160 0 0 0 AND8_0.B5
flabel metal1 -24917 -20506 -24855 -20470 0 FreeSans 160 0 0 0 AND8_0.A4
flabel metal1 -24923 -20344 -24861 -20308 0 FreeSans 160 0 0 0 AND8_0.B4
flabel metal1 -24923 -19318 -24861 -19282 0 FreeSans 160 0 0 0 AND8_0.A3
flabel metal1 -24921 -19156 -24859 -19120 0 FreeSans 160 0 0 0 AND8_0.B3
flabel metal1 -24919 -18192 -24857 -18156 0 FreeSans 160 0 0 0 AND8_0.A2
flabel metal1 -24923 -18038 -24861 -18002 0 FreeSans 160 0 0 0 AND8_0.B2
flabel metal1 -24923 -16984 -24861 -16948 0 FreeSans 160 0 0 0 AND8_0.A1
flabel metal1 -24923 -16826 -24861 -16790 0 FreeSans 160 0 0 0 AND8_0.B1
flabel metal1 -24919 -15802 -24857 -15766 0 FreeSans 160 0 0 0 AND8_0.A0
flabel metal1 -24919 -15640 -24857 -15604 0 FreeSans 160 0 0 0 AND8_0.B0
flabel metal1 -20379 -17972 -20361 -17952 0 FreeSans 160 0 0 0 AND8_0.S0
flabel metal1 -20381 -18468 -20363 -18448 0 FreeSans 160 0 0 0 AND8_0.S1
flabel metal1 -20379 -18950 -20361 -18930 0 FreeSans 160 0 0 0 AND8_0.S2
flabel metal1 -20381 -19448 -20363 -19428 0 FreeSans 160 0 0 0 AND8_0.S3
flabel metal1 -20381 -19926 -20363 -19906 0 FreeSans 160 0 0 0 AND8_0.S4
flabel metal1 -20381 -20390 -20363 -20370 0 FreeSans 160 0 0 0 AND8_0.S5
flabel metal1 -20383 -20850 -20365 -20830 0 FreeSans 160 0 0 0 AND8_0.S6
flabel metal1 -20381 -21334 -20363 -21314 0 FreeSans 160 0 0 0 AND8_0.S7
rlabel metal1 -20388 -17980 -20355 -17945 7 AND8_0.NOT8_0.S0
rlabel metal1 -20395 -18479 -20362 -18444 7 AND8_0.NOT8_0.S1
rlabel metal1 -20388 -18958 -20355 -18923 7 AND8_0.NOT8_0.S2
rlabel metal1 -20387 -19458 -20354 -19423 7 AND8_0.NOT8_0.S3
rlabel metal1 -20387 -19938 -20354 -19903 7 AND8_0.NOT8_0.S4
rlabel metal1 -20387 -20397 -20354 -20362 7 AND8_0.NOT8_0.S5
rlabel metal1 -20387 -20858 -20354 -20823 7 AND8_0.NOT8_0.S6
rlabel metal1 -20388 -21338 -20355 -21303 7 AND8_0.NOT8_0.S7
rlabel metal1 -21985 -18339 -21938 -18288 3 AND8_0.NOT8_0.A0
rlabel metal1 -21987 -18839 -21940 -18788 3 AND8_0.NOT8_0.A1
rlabel metal1 -21988 -19320 -21941 -19269 3 AND8_0.NOT8_0.A2
rlabel metal1 -21987 -19819 -21940 -19768 3 AND8_0.NOT8_0.A3
rlabel metal1 -21986 -20300 -21939 -20249 3 AND8_0.NOT8_0.A4
rlabel metal1 -21985 -20760 -21938 -20709 3 AND8_0.NOT8_0.A5
rlabel metal1 -21988 -21219 -21941 -21168 3 AND8_0.NOT8_0.A6
rlabel metal1 -21988 -21700 -21941 -21649 3 AND8_0.NOT8_0.A7
flabel metal4 -21976 -19524 -21906 -19426 0 FreeSans 160 0 0 0 AND8_0.NOT8_0.VDD
flabel metal5 -20438 -19374 -20368 -19276 0 FreeSans 160 0 0 0 AND8_0.NOT8_0.VSS
rlabel metal1 -21314 -18348 -21314 -18348 1 AND8_0.NOT8_0.inv_7.A
rlabel metal1 -20925 -18150 -20925 -18150 3 AND8_0.NOT8_0.inv_7.VSS
rlabel metal1 -21722 -18138 -21722 -18138 3 AND8_0.NOT8_0.inv_7.VDD
rlabel metal1 -21314 -17936 -21314 -17936 1 AND8_0.NOT8_0.inv_7.Y
rlabel metal1 -21313 -18848 -21313 -18848 1 AND8_0.NOT8_0.inv_6.A
rlabel metal1 -20924 -18650 -20924 -18650 3 AND8_0.NOT8_0.inv_6.VSS
rlabel metal1 -21721 -18638 -21721 -18638 3 AND8_0.NOT8_0.inv_6.VDD
rlabel metal1 -21313 -18436 -21313 -18436 1 AND8_0.NOT8_0.inv_6.Y
rlabel metal1 -21314 -19328 -21314 -19328 1 AND8_0.NOT8_0.inv_5.A
rlabel metal1 -20925 -19130 -20925 -19130 3 AND8_0.NOT8_0.inv_5.VSS
rlabel metal1 -21722 -19118 -21722 -19118 3 AND8_0.NOT8_0.inv_5.VDD
rlabel metal1 -21314 -18916 -21314 -18916 1 AND8_0.NOT8_0.inv_5.Y
rlabel metal1 -21314 -20308 -21314 -20308 1 AND8_0.NOT8_0.inv_4.A
rlabel metal1 -20925 -20110 -20925 -20110 3 AND8_0.NOT8_0.inv_4.VSS
rlabel metal1 -21722 -20098 -21722 -20098 3 AND8_0.NOT8_0.inv_4.VDD
rlabel metal1 -21314 -19896 -21314 -19896 1 AND8_0.NOT8_0.inv_4.Y
rlabel metal1 -21314 -20768 -21314 -20768 1 AND8_0.NOT8_0.inv_3.A
rlabel metal1 -20925 -20570 -20925 -20570 3 AND8_0.NOT8_0.inv_3.VSS
rlabel metal1 -21722 -20558 -21722 -20558 3 AND8_0.NOT8_0.inv_3.VDD
rlabel metal1 -21314 -20356 -21314 -20356 1 AND8_0.NOT8_0.inv_3.Y
rlabel metal1 -21328 -21228 -21328 -21228 1 AND8_0.NOT8_0.inv_2.A
rlabel metal1 -20939 -21030 -20939 -21030 3 AND8_0.NOT8_0.inv_2.VSS
rlabel metal1 -21736 -21018 -21736 -21018 3 AND8_0.NOT8_0.inv_2.VDD
rlabel metal1 -21328 -20816 -21328 -20816 1 AND8_0.NOT8_0.inv_2.Y
rlabel metal1 -21326 -21708 -21326 -21708 1 AND8_0.NOT8_0.inv_1.A
rlabel metal1 -20937 -21510 -20937 -21510 3 AND8_0.NOT8_0.inv_1.VSS
rlabel metal1 -21734 -21498 -21734 -21498 3 AND8_0.NOT8_0.inv_1.VDD
rlabel metal1 -21326 -21296 -21326 -21296 1 AND8_0.NOT8_0.inv_1.Y
rlabel metal1 -21314 -19828 -21314 -19828 1 AND8_0.NOT8_0.inv_0.A
rlabel metal1 -20925 -19630 -20925 -19630 3 AND8_0.NOT8_0.inv_0.VSS
rlabel metal1 -21722 -19618 -21722 -19618 3 AND8_0.NOT8_0.inv_0.VDD
rlabel metal1 -21314 -19416 -21314 -19416 1 AND8_0.NOT8_0.inv_0.Y
rlabel metal1 -24928 -24341 -24871 -24274 7 AND8_0.NAND8_0.A0
rlabel metal1 -24928 -24172 -24871 -24116 7 AND8_0.NAND8_0.B0
rlabel metal1 -24930 -23035 -24866 -22960 7 AND8_0.NAND8_0.A1
rlabel metal1 -24929 -22860 -24866 -22806 7 AND8_0.NAND8_0.B1
rlabel metal1 -24928 -21731 -24872 -21662 7 AND8_0.NAND8_0.A2
rlabel metal1 -24927 -21559 -24872 -21503 7 AND8_0.NAND8_0.B2
rlabel metal1 -24927 -20525 -24859 -20452 7 AND8_0.NAND8_0.A3
rlabel metal1 -24927 -20355 -24860 -20299 7 AND8_0.NAND8_0.B3
rlabel metal1 -24929 -19337 -24860 -19265 7 AND8_0.NAND8_0.A4
rlabel metal1 -24929 -19170 -24860 -19108 7 AND8_0.NAND8_0.B4
rlabel metal1 -24930 -18211 -24849 -18137 7 AND8_0.NAND8_0.A5
rlabel metal1 -24930 -18045 -24852 -17991 7 AND8_0.NAND8_0.B5
rlabel metal1 -24931 -17008 -24848 -16929 7 AND8_0.NAND8_0.A6
rlabel metal1 -24930 -16834 -24848 -16774 7 AND8_0.NAND8_0.B6
rlabel metal1 -24928 -15822 -24846 -15748 7 AND8_0.NAND8_0.A7
rlabel metal1 -24927 -15651 -24846 -15592 7 AND8_0.NAND8_0.B7
rlabel metal1 -23079 -23334 -23010 -23269 3 AND8_0.NAND8_0.P0
rlabel metal1 -23080 -22028 -23011 -21963 3 AND8_0.NAND8_0.P1
rlabel metal1 -23079 -20727 -23010 -20662 3 AND8_0.NAND8_0.P2
rlabel metal1 -23078 -19528 -23009 -19463 3 AND8_0.NAND8_0.P3
rlabel metal1 -23079 -18338 -23010 -18273 3 AND8_0.NAND8_0.P4
rlabel metal1 -23078 -17236 -23009 -17171 3 AND8_0.NAND8_0.P5
rlabel metal1 -23079 -16033 -23010 -15968 3 AND8_0.NAND8_0.P6
rlabel metal1 -23079 -14837 -23010 -14772 3 AND8_0.NAND8_0.P7
rlabel metal1 -24088 -21497 -24088 -21497 5 AND8_0.NAND8_0.NAND2_9.A
rlabel metal1 -23920 -21497 -23920 -21497 5 AND8_0.NAND8_0.NAND2_9.B
rlabel metal1 -23801 -21027 -23801 -21027 3 AND8_0.NAND8_0.NAND2_9.VSS
rlabel metal1 -24431 -21144 -24431 -21144 7 AND8_0.NAND8_0.NAND2_9.VDD
rlabel metal1 -24198 -20791 -24198 -20791 1 AND8_0.NAND8_0.NAND2_9.Y
rlabel metal1 -24089 -22800 -24089 -22800 5 AND8_0.NAND8_0.NAND2_8.A
rlabel metal1 -23921 -22800 -23921 -22800 5 AND8_0.NAND8_0.NAND2_8.B
rlabel metal1 -23802 -22330 -23802 -22330 3 AND8_0.NAND8_0.NAND2_8.VSS
rlabel metal1 -24432 -22447 -24432 -22447 7 AND8_0.NAND8_0.NAND2_8.VDD
rlabel metal1 -24199 -22094 -24199 -22094 1 AND8_0.NAND8_0.NAND2_8.Y
rlabel metal1 -24141 -16771 -24141 -16771 5 AND8_0.NAND8_0.NAND2_7.A
rlabel metal1 -23973 -16771 -23973 -16771 5 AND8_0.NAND8_0.NAND2_7.B
rlabel metal1 -23854 -16301 -23854 -16301 3 AND8_0.NAND8_0.NAND2_7.VSS
rlabel metal1 -24484 -16418 -24484 -16418 7 AND8_0.NAND8_0.NAND2_7.VDD
rlabel metal1 -24251 -16065 -24251 -16065 1 AND8_0.NAND8_0.NAND2_7.Y
rlabel metal1 -24136 -17984 -24136 -17984 5 AND8_0.NAND8_0.NAND2_6.A
rlabel metal1 -23968 -17984 -23968 -17984 5 AND8_0.NAND8_0.NAND2_6.B
rlabel metal1 -23849 -17514 -23849 -17514 3 AND8_0.NAND8_0.NAND2_6.VSS
rlabel metal1 -24479 -17631 -24479 -17631 7 AND8_0.NAND8_0.NAND2_6.VDD
rlabel metal1 -24246 -17278 -24246 -17278 1 AND8_0.NAND8_0.NAND2_6.Y
rlabel metal1 -24089 -24109 -24089 -24109 5 AND8_0.NAND8_0.NAND2_4.A
rlabel metal1 -23921 -24109 -23921 -24109 5 AND8_0.NAND8_0.NAND2_4.B
rlabel metal1 -23802 -23639 -23802 -23639 3 AND8_0.NAND8_0.NAND2_4.VSS
rlabel metal1 -24432 -23756 -24432 -23756 7 AND8_0.NAND8_0.NAND2_4.VDD
rlabel metal1 -24199 -23403 -24199 -23403 1 AND8_0.NAND8_0.NAND2_4.Y
rlabel metal1 -24119 -20297 -24119 -20297 5 AND8_0.NAND8_0.NAND2_2.A
rlabel metal1 -23951 -20297 -23951 -20297 5 AND8_0.NAND8_0.NAND2_2.B
rlabel metal1 -23832 -19827 -23832 -19827 3 AND8_0.NAND8_0.NAND2_2.VSS
rlabel metal1 -24462 -19944 -24462 -19944 7 AND8_0.NAND8_0.NAND2_2.VDD
rlabel metal1 -24229 -19591 -24229 -19591 1 AND8_0.NAND8_0.NAND2_2.Y
rlabel metal1 -24121 -19103 -24121 -19103 5 AND8_0.NAND8_0.NAND2_1.A
rlabel metal1 -23953 -19103 -23953 -19103 5 AND8_0.NAND8_0.NAND2_1.B
rlabel metal1 -23834 -18633 -23834 -18633 3 AND8_0.NAND8_0.NAND2_1.VSS
rlabel metal1 -24464 -18750 -24464 -18750 7 AND8_0.NAND8_0.NAND2_1.VDD
rlabel metal1 -24231 -18397 -24231 -18397 1 AND8_0.NAND8_0.NAND2_1.Y
rlabel metal1 -24142 -15586 -24142 -15586 5 AND8_0.NAND8_0.NAND2_0.A
rlabel metal1 -23974 -15586 -23974 -15586 5 AND8_0.NAND8_0.NAND2_0.B
rlabel metal1 -23855 -15116 -23855 -15116 3 AND8_0.NAND8_0.NAND2_0.VSS
rlabel metal1 -24485 -15233 -24485 -15233 7 AND8_0.NAND8_0.NAND2_0.VDD
rlabel metal1 -24252 -14880 -24252 -14880 1 AND8_0.NAND8_0.NAND2_0.Y
flabel metal1 -12607 -34754 -12545 -34675 0 FreeSans 160 0 0 0 XOR8_0.B7
flabel metal1 -12598 -34572 -12552 -34515 0 FreeSans 160 0 0 0 XOR8_0.A7
flabel metal1 -12606 -31990 -12560 -31933 0 FreeSans 160 0 0 0 XOR8_0.A6
flabel metal1 -12600 -29449 -12554 -29392 0 FreeSans 160 0 0 0 XOR8_0.A5
flabel metal1 -12598 -26817 -12552 -26760 0 FreeSans 160 0 0 0 XOR8_0.A4
flabel metal1 -12604 -24024 -12558 -23967 0 FreeSans 160 0 0 0 XOR8_0.A3
flabel metal1 -12603 -21438 -12557 -21381 0 FreeSans 160 0 0 0 XOR8_0.A2
flabel metal1 -12602 -18468 -12556 -18411 0 FreeSans 160 0 0 0 XOR8_0.A1
flabel metal1 -12601 -15660 -12555 -15603 0 FreeSans 160 0 0 0 XOR8_0.A0
flabel metal1 -12600 -15816 -12554 -15759 0 FreeSans 160 0 0 0 XOR8_0.B0
flabel metal1 -12604 -18635 -12558 -18578 0 FreeSans 160 0 0 0 XOR8_0.B1
flabel metal1 -12601 -21563 -12555 -21506 0 FreeSans 160 0 0 0 XOR8_0.B2
flabel metal1 -12606 -24149 -12560 -24092 0 FreeSans 160 0 0 0 XOR8_0.B3
flabel metal1 -12600 -26994 -12554 -26937 0 FreeSans 160 0 0 0 XOR8_0.B4
flabel metal1 -12601 -29598 -12555 -29541 0 FreeSans 160 0 0 0 XOR8_0.B5
flabel metal1 -12604 -32120 -12558 -32063 0 FreeSans 160 0 0 0 XOR8_0.B6
flabel metal1 -10837 -32994 -10791 -32937 0 FreeSans 160 0 0 0 XOR8_0.S7
flabel metal1 -10839 -30313 -10793 -30256 0 FreeSans 160 0 0 0 XOR8_0.S6
flabel metal1 -10832 -27745 -10786 -27688 0 FreeSans 160 0 0 0 XOR8_0.S5
flabel metal1 -10835 -25055 -10789 -24998 0 FreeSans 160 0 0 0 XOR8_0.S4
flabel metal1 -10832 -22319 -10786 -22262 0 FreeSans 160 0 0 0 XOR8_0.S3
flabel metal1 -10839 -19695 -10793 -19638 0 FreeSans 160 0 0 0 XOR8_0.S2
flabel metal1 -10834 -16756 -10788 -16699 0 FreeSans 160 0 0 0 XOR8_0.S1
flabel metal1 -10836 -13961 -10790 -13904 0 FreeSans 160 0 0 0 XOR8_0.S0
rlabel poly -11549 -18316 -11509 -18292 5 XOR8_0.XOR2_7.A
rlabel metal1 -11405 -18338 -11365 -18314 5 XOR8_0.XOR2_7.B
rlabel via1 -12447 -17806 -12421 -17712 3 XOR8_0.XOR2_7.VDD
rlabel metal1 -11471 -16948 -11393 -16896 3 XOR8_0.XOR2_7.Y
rlabel metal1 -11059 -17876 -11033 -17782 3 XOR8_0.XOR2_7.VSS
rlabel poly -11549 -21273 -11509 -21249 5 XOR8_0.XOR2_6.A
rlabel metal1 -11405 -21295 -11365 -21271 5 XOR8_0.XOR2_6.B
rlabel via1 -12447 -20763 -12421 -20669 3 XOR8_0.XOR2_6.VDD
rlabel metal1 -11471 -19905 -11393 -19853 3 XOR8_0.XOR2_6.Y
rlabel metal1 -11059 -20833 -11033 -20739 3 XOR8_0.XOR2_6.VSS
rlabel poly -11549 -23852 -11509 -23828 5 XOR8_0.XOR2_5.A
rlabel metal1 -11405 -23874 -11365 -23850 5 XOR8_0.XOR2_5.B
rlabel via1 -12447 -23342 -12421 -23248 3 XOR8_0.XOR2_5.VDD
rlabel metal1 -11471 -22484 -11393 -22432 3 XOR8_0.XOR2_5.Y
rlabel metal1 -11059 -23412 -11033 -23318 3 XOR8_0.XOR2_5.VSS
rlabel poly -11549 -26620 -11509 -26596 5 XOR8_0.XOR2_4.A
rlabel metal1 -11405 -26642 -11365 -26618 5 XOR8_0.XOR2_4.B
rlabel via1 -12447 -26110 -12421 -26016 3 XOR8_0.XOR2_4.VDD
rlabel metal1 -11471 -25252 -11393 -25200 3 XOR8_0.XOR2_4.Y
rlabel metal1 -11059 -26180 -11033 -26086 3 XOR8_0.XOR2_4.VSS
rlabel poly -11549 -29253 -11509 -29229 5 XOR8_0.XOR2_3.A
rlabel metal1 -11405 -29275 -11365 -29251 5 XOR8_0.XOR2_3.B
rlabel via1 -12447 -28743 -12421 -28649 3 XOR8_0.XOR2_3.VDD
rlabel metal1 -11471 -27885 -11393 -27833 3 XOR8_0.XOR2_3.Y
rlabel metal1 -11059 -28813 -11033 -28719 3 XOR8_0.XOR2_3.VSS
rlabel poly -11549 -31862 -11509 -31838 5 XOR8_0.XOR2_2.A
rlabel metal1 -11405 -31884 -11365 -31860 5 XOR8_0.XOR2_2.B
rlabel via1 -12447 -31352 -12421 -31258 3 XOR8_0.XOR2_2.VDD
rlabel metal1 -11471 -30494 -11393 -30442 3 XOR8_0.XOR2_2.Y
rlabel metal1 -11059 -31422 -11033 -31328 3 XOR8_0.XOR2_2.VSS
rlabel poly -11551 -34482 -11511 -34458 5 XOR8_0.XOR2_1.A
rlabel metal1 -11407 -34504 -11367 -34480 5 XOR8_0.XOR2_1.B
rlabel via1 -12449 -33972 -12423 -33878 3 XOR8_0.XOR2_1.VDD
rlabel metal1 -11473 -33114 -11395 -33062 3 XOR8_0.XOR2_1.Y
rlabel metal1 -11061 -34042 -11035 -33948 3 XOR8_0.XOR2_1.VSS
rlabel poly -11551 -15500 -11511 -15476 5 XOR8_0.XOR2_0.A
rlabel metal1 -11407 -15522 -11367 -15498 5 XOR8_0.XOR2_0.B
rlabel via1 -12449 -14990 -12423 -14896 3 XOR8_0.XOR2_0.VDD
rlabel metal1 -11473 -14132 -11395 -14080 3 XOR8_0.XOR2_0.Y
rlabel metal1 -11061 -15060 -11035 -14966 3 XOR8_0.XOR2_0.VSS
rlabel metal1 -2332 -14527 -2332 -14527 3 right_shifter_0.A0
rlabel metal1 -2332 -15341 -2332 -15341 3 right_shifter_0.A1
rlabel metal1 -2332 -16155 -2332 -16155 3 right_shifter_0.A2
rlabel metal1 -2332 -16982 -2332 -16982 3 right_shifter_0.A3
rlabel metal1 -2332 -17797 -2332 -17797 3 right_shifter_0.A4
rlabel metal1 -2332 -18624 -2332 -18624 3 right_shifter_0.A5
rlabel metal1 -2332 -19442 -2332 -19442 3 right_shifter_0.A6
rlabel metal1 -2332 -20253 -2332 -20253 3 right_shifter_0.A7
rlabel metal1 -1058 -13713 -1058 -13713 3 right_shifter_0.C
rlabel metal1 -1058 -14528 -1058 -14528 3 right_shifter_0.S0
rlabel metal1 -1058 -15347 -1058 -15347 3 right_shifter_0.S1
rlabel metal1 -1058 -16175 -1058 -16175 3 right_shifter_0.S2
rlabel metal1 -1058 -16991 -1058 -16991 3 right_shifter_0.S3
rlabel metal1 -1058 -17808 -1058 -17808 3 right_shifter_0.S4
rlabel metal1 -1058 -18625 -1058 -18625 3 right_shifter_0.S5
rlabel metal1 -1058 -19444 -1058 -19444 3 right_shifter_0.S6
rlabel metal1 -1058 -20262 -1058 -20262 3 right_shifter_0.S7
rlabel metal5 -1058 -17008 -1058 -17008 3 right_shifter_0.VSS
rlabel metal4 -2310 -16982 -2310 -16982 3 right_shifter_0.VDD
rlabel metal1 -1808 -20684 -1808 -20684 1 right_shifter_0.inv_0.A
rlabel metal1 -1419 -20486 -1419 -20486 3 right_shifter_0.inv_0.VSS
rlabel metal1 -2216 -20474 -2216 -20474 3 right_shifter_0.inv_0.VDD
rlabel metal1 -1808 -20272 -1808 -20272 1 right_shifter_0.inv_0.Y
rlabel metal1 -1811 -15330 -1811 -15330 1 right_shifter_0.buffer_7.A
rlabel metal1 -1419 -14892 -1419 -14892 3 right_shifter_0.buffer_7.VSS
rlabel metal1 -1826 -14539 -1826 -14539 1 right_shifter_0.buffer_7.Y
rlabel metal1 -2216 -14879 -2216 -14879 3 right_shifter_0.buffer_7.VDD
rlabel metal1 -1808 -14951 -1808 -14951 1 right_shifter_0.buffer_7.inv_1.A
rlabel metal1 -1419 -14753 -1419 -14753 3 right_shifter_0.buffer_7.inv_1.VSS
rlabel metal1 -2216 -14741 -2216 -14741 3 right_shifter_0.buffer_7.inv_1.VDD
rlabel metal1 -1808 -14539 -1808 -14539 1 right_shifter_0.buffer_7.inv_1.Y
rlabel metal1 -1808 -15330 -1808 -15330 1 right_shifter_0.buffer_7.inv_0.A
rlabel metal1 -1419 -15132 -1419 -15132 3 right_shifter_0.buffer_7.inv_0.VSS
rlabel metal1 -2216 -15120 -2216 -15120 3 right_shifter_0.buffer_7.inv_0.VDD
rlabel metal1 -1808 -14918 -1808 -14918 1 right_shifter_0.buffer_7.inv_0.Y
rlabel metal1 -1811 -14511 -1811 -14511 1 right_shifter_0.buffer_6.A
rlabel metal1 -1419 -14073 -1419 -14073 3 right_shifter_0.buffer_6.VSS
rlabel metal1 -1826 -13720 -1826 -13720 1 right_shifter_0.buffer_6.Y
rlabel metal1 -2216 -14060 -2216 -14060 3 right_shifter_0.buffer_6.VDD
rlabel metal1 -1808 -14132 -1808 -14132 1 right_shifter_0.buffer_6.inv_1.A
rlabel metal1 -1419 -13934 -1419 -13934 3 right_shifter_0.buffer_6.inv_1.VSS
rlabel metal1 -2216 -13922 -2216 -13922 3 right_shifter_0.buffer_6.inv_1.VDD
rlabel metal1 -1808 -13720 -1808 -13720 1 right_shifter_0.buffer_6.inv_1.Y
rlabel metal1 -1808 -14511 -1808 -14511 1 right_shifter_0.buffer_6.inv_0.A
rlabel metal1 -1419 -14313 -1419 -14313 3 right_shifter_0.buffer_6.inv_0.VSS
rlabel metal1 -2216 -14301 -2216 -14301 3 right_shifter_0.buffer_6.inv_0.VDD
rlabel metal1 -1808 -14099 -1808 -14099 1 right_shifter_0.buffer_6.inv_0.Y
rlabel metal1 -1811 -16968 -1811 -16968 1 right_shifter_0.buffer_5.A
rlabel metal1 -1419 -16530 -1419 -16530 3 right_shifter_0.buffer_5.VSS
rlabel metal1 -1826 -16177 -1826 -16177 1 right_shifter_0.buffer_5.Y
rlabel metal1 -2216 -16517 -2216 -16517 3 right_shifter_0.buffer_5.VDD
rlabel metal1 -1808 -16589 -1808 -16589 1 right_shifter_0.buffer_5.inv_1.A
rlabel metal1 -1419 -16391 -1419 -16391 3 right_shifter_0.buffer_5.inv_1.VSS
rlabel metal1 -2216 -16379 -2216 -16379 3 right_shifter_0.buffer_5.inv_1.VDD
rlabel metal1 -1808 -16177 -1808 -16177 1 right_shifter_0.buffer_5.inv_1.Y
rlabel metal1 -1808 -16968 -1808 -16968 1 right_shifter_0.buffer_5.inv_0.A
rlabel metal1 -1419 -16770 -1419 -16770 3 right_shifter_0.buffer_5.inv_0.VSS
rlabel metal1 -2216 -16758 -2216 -16758 3 right_shifter_0.buffer_5.inv_0.VDD
rlabel metal1 -1808 -16556 -1808 -16556 1 right_shifter_0.buffer_5.inv_0.Y
rlabel metal1 -1811 -17787 -1811 -17787 1 right_shifter_0.buffer_4.A
rlabel metal1 -1419 -17349 -1419 -17349 3 right_shifter_0.buffer_4.VSS
rlabel metal1 -1826 -16996 -1826 -16996 1 right_shifter_0.buffer_4.Y
rlabel metal1 -2216 -17336 -2216 -17336 3 right_shifter_0.buffer_4.VDD
rlabel metal1 -1808 -17408 -1808 -17408 1 right_shifter_0.buffer_4.inv_1.A
rlabel metal1 -1419 -17210 -1419 -17210 3 right_shifter_0.buffer_4.inv_1.VSS
rlabel metal1 -2216 -17198 -2216 -17198 3 right_shifter_0.buffer_4.inv_1.VDD
rlabel metal1 -1808 -16996 -1808 -16996 1 right_shifter_0.buffer_4.inv_1.Y
rlabel metal1 -1808 -17787 -1808 -17787 1 right_shifter_0.buffer_4.inv_0.A
rlabel metal1 -1419 -17589 -1419 -17589 3 right_shifter_0.buffer_4.inv_0.VSS
rlabel metal1 -2216 -17577 -2216 -17577 3 right_shifter_0.buffer_4.inv_0.VDD
rlabel metal1 -1808 -17375 -1808 -17375 1 right_shifter_0.buffer_4.inv_0.Y
rlabel metal1 -1811 -18606 -1811 -18606 1 right_shifter_0.buffer_3.A
rlabel metal1 -1419 -18168 -1419 -18168 3 right_shifter_0.buffer_3.VSS
rlabel metal1 -1826 -17815 -1826 -17815 1 right_shifter_0.buffer_3.Y
rlabel metal1 -2216 -18155 -2216 -18155 3 right_shifter_0.buffer_3.VDD
rlabel metal1 -1808 -18227 -1808 -18227 1 right_shifter_0.buffer_3.inv_1.A
rlabel metal1 -1419 -18029 -1419 -18029 3 right_shifter_0.buffer_3.inv_1.VSS
rlabel metal1 -2216 -18017 -2216 -18017 3 right_shifter_0.buffer_3.inv_1.VDD
rlabel metal1 -1808 -17815 -1808 -17815 1 right_shifter_0.buffer_3.inv_1.Y
rlabel metal1 -1808 -18606 -1808 -18606 1 right_shifter_0.buffer_3.inv_0.A
rlabel metal1 -1419 -18408 -1419 -18408 3 right_shifter_0.buffer_3.inv_0.VSS
rlabel metal1 -2216 -18396 -2216 -18396 3 right_shifter_0.buffer_3.inv_0.VDD
rlabel metal1 -1808 -18194 -1808 -18194 1 right_shifter_0.buffer_3.inv_0.Y
rlabel metal1 -1811 -19425 -1811 -19425 1 right_shifter_0.buffer_2.A
rlabel metal1 -1419 -18987 -1419 -18987 3 right_shifter_0.buffer_2.VSS
rlabel metal1 -1826 -18634 -1826 -18634 1 right_shifter_0.buffer_2.Y
rlabel metal1 -2216 -18974 -2216 -18974 3 right_shifter_0.buffer_2.VDD
rlabel metal1 -1808 -19046 -1808 -19046 1 right_shifter_0.buffer_2.inv_1.A
rlabel metal1 -1419 -18848 -1419 -18848 3 right_shifter_0.buffer_2.inv_1.VSS
rlabel metal1 -2216 -18836 -2216 -18836 3 right_shifter_0.buffer_2.inv_1.VDD
rlabel metal1 -1808 -18634 -1808 -18634 1 right_shifter_0.buffer_2.inv_1.Y
rlabel metal1 -1808 -19425 -1808 -19425 1 right_shifter_0.buffer_2.inv_0.A
rlabel metal1 -1419 -19227 -1419 -19227 3 right_shifter_0.buffer_2.inv_0.VSS
rlabel metal1 -2216 -19215 -2216 -19215 3 right_shifter_0.buffer_2.inv_0.VDD
rlabel metal1 -1808 -19013 -1808 -19013 1 right_shifter_0.buffer_2.inv_0.Y
rlabel metal1 -1811 -20244 -1811 -20244 1 right_shifter_0.buffer_1.A
rlabel metal1 -1419 -19806 -1419 -19806 3 right_shifter_0.buffer_1.VSS
rlabel metal1 -1826 -19453 -1826 -19453 1 right_shifter_0.buffer_1.Y
rlabel metal1 -2216 -19793 -2216 -19793 3 right_shifter_0.buffer_1.VDD
rlabel metal1 -1808 -19865 -1808 -19865 1 right_shifter_0.buffer_1.inv_1.A
rlabel metal1 -1419 -19667 -1419 -19667 3 right_shifter_0.buffer_1.inv_1.VSS
rlabel metal1 -2216 -19655 -2216 -19655 3 right_shifter_0.buffer_1.inv_1.VDD
rlabel metal1 -1808 -19453 -1808 -19453 1 right_shifter_0.buffer_1.inv_1.Y
rlabel metal1 -1808 -20244 -1808 -20244 1 right_shifter_0.buffer_1.inv_0.A
rlabel metal1 -1419 -20046 -1419 -20046 3 right_shifter_0.buffer_1.inv_0.VSS
rlabel metal1 -2216 -20034 -2216 -20034 3 right_shifter_0.buffer_1.inv_0.VDD
rlabel metal1 -1808 -19832 -1808 -19832 1 right_shifter_0.buffer_1.inv_0.Y
rlabel metal1 -1811 -16149 -1811 -16149 1 right_shifter_0.buffer_0.A
rlabel metal1 -1419 -15711 -1419 -15711 3 right_shifter_0.buffer_0.VSS
rlabel metal1 -1826 -15358 -1826 -15358 1 right_shifter_0.buffer_0.Y
rlabel metal1 -2216 -15698 -2216 -15698 3 right_shifter_0.buffer_0.VDD
rlabel metal1 -1808 -15770 -1808 -15770 1 right_shifter_0.buffer_0.inv_1.A
rlabel metal1 -1419 -15572 -1419 -15572 3 right_shifter_0.buffer_0.inv_1.VSS
rlabel metal1 -2216 -15560 -2216 -15560 3 right_shifter_0.buffer_0.inv_1.VDD
rlabel metal1 -1808 -15358 -1808 -15358 1 right_shifter_0.buffer_0.inv_1.Y
rlabel metal1 -1808 -16149 -1808 -16149 1 right_shifter_0.buffer_0.inv_0.A
rlabel metal1 -1419 -15951 -1419 -15951 3 right_shifter_0.buffer_0.inv_0.VSS
rlabel metal1 -2216 -15939 -2216 -15939 3 right_shifter_0.buffer_0.inv_0.VDD
rlabel metal1 -1808 -15737 -1808 -15737 1 right_shifter_0.buffer_0.inv_0.Y
rlabel metal1 -6949 -15292 -6916 -15257 7 NOT8_0.S0
rlabel metal1 -6956 -15791 -6923 -15756 7 NOT8_0.S1
rlabel metal1 -6949 -16270 -6916 -16235 7 NOT8_0.S2
rlabel metal1 -6948 -16770 -6915 -16735 7 NOT8_0.S3
rlabel metal1 -6948 -17250 -6915 -17215 7 NOT8_0.S4
rlabel metal1 -6948 -17709 -6915 -17674 7 NOT8_0.S5
rlabel metal1 -6948 -18170 -6915 -18135 7 NOT8_0.S6
rlabel metal1 -6949 -18650 -6916 -18615 7 NOT8_0.S7
rlabel metal1 -8546 -15651 -8499 -15600 3 NOT8_0.A0
rlabel metal1 -8548 -16151 -8501 -16100 3 NOT8_0.A1
rlabel metal1 -8549 -16632 -8502 -16581 3 NOT8_0.A2
rlabel metal1 -8548 -17131 -8501 -17080 3 NOT8_0.A3
rlabel metal1 -8547 -17612 -8500 -17561 3 NOT8_0.A4
rlabel metal1 -8546 -18072 -8499 -18021 3 NOT8_0.A5
rlabel metal1 -8549 -18531 -8502 -18480 3 NOT8_0.A6
rlabel metal1 -8549 -19012 -8502 -18961 3 NOT8_0.A7
flabel metal4 -8537 -16836 -8467 -16738 0 FreeSans 160 0 0 0 NOT8_0.VDD
flabel metal5 -6999 -16686 -6929 -16588 0 FreeSans 160 0 0 0 NOT8_0.VSS
rlabel metal1 -7875 -15660 -7875 -15660 1 NOT8_0.inv_7.A
rlabel metal1 -7486 -15462 -7486 -15462 3 NOT8_0.inv_7.VSS
rlabel metal1 -8283 -15450 -8283 -15450 3 NOT8_0.inv_7.VDD
rlabel metal1 -7875 -15248 -7875 -15248 1 NOT8_0.inv_7.Y
rlabel metal1 -7874 -16160 -7874 -16160 1 NOT8_0.inv_6.A
rlabel metal1 -7485 -15962 -7485 -15962 3 NOT8_0.inv_6.VSS
rlabel metal1 -8282 -15950 -8282 -15950 3 NOT8_0.inv_6.VDD
rlabel metal1 -7874 -15748 -7874 -15748 1 NOT8_0.inv_6.Y
rlabel metal1 -7875 -16640 -7875 -16640 1 NOT8_0.inv_5.A
rlabel metal1 -7486 -16442 -7486 -16442 3 NOT8_0.inv_5.VSS
rlabel metal1 -8283 -16430 -8283 -16430 3 NOT8_0.inv_5.VDD
rlabel metal1 -7875 -16228 -7875 -16228 1 NOT8_0.inv_5.Y
rlabel metal1 -7875 -17620 -7875 -17620 1 NOT8_0.inv_4.A
rlabel metal1 -7486 -17422 -7486 -17422 3 NOT8_0.inv_4.VSS
rlabel metal1 -8283 -17410 -8283 -17410 3 NOT8_0.inv_4.VDD
rlabel metal1 -7875 -17208 -7875 -17208 1 NOT8_0.inv_4.Y
rlabel metal1 -7875 -18080 -7875 -18080 1 NOT8_0.inv_3.A
rlabel metal1 -7486 -17882 -7486 -17882 3 NOT8_0.inv_3.VSS
rlabel metal1 -8283 -17870 -8283 -17870 3 NOT8_0.inv_3.VDD
rlabel metal1 -7875 -17668 -7875 -17668 1 NOT8_0.inv_3.Y
rlabel metal1 -7889 -18540 -7889 -18540 1 NOT8_0.inv_2.A
rlabel metal1 -7500 -18342 -7500 -18342 3 NOT8_0.inv_2.VSS
rlabel metal1 -8297 -18330 -8297 -18330 3 NOT8_0.inv_2.VDD
rlabel metal1 -7889 -18128 -7889 -18128 1 NOT8_0.inv_2.Y
rlabel metal1 -7887 -19020 -7887 -19020 1 NOT8_0.inv_1.A
rlabel metal1 -7498 -18822 -7498 -18822 3 NOT8_0.inv_1.VSS
rlabel metal1 -8295 -18810 -8295 -18810 3 NOT8_0.inv_1.VDD
rlabel metal1 -7887 -18608 -7887 -18608 1 NOT8_0.inv_1.Y
rlabel metal1 -7875 -17140 -7875 -17140 1 NOT8_0.inv_0.A
rlabel metal1 -7486 -16942 -7486 -16942 3 NOT8_0.inv_0.VSS
rlabel metal1 -8283 -16930 -8283 -16930 3 NOT8_0.inv_0.VDD
rlabel metal1 -7875 -16728 -7875 -16728 1 NOT8_0.inv_0.Y
rlabel metal1 -5048 -14527 -5048 -14527 3 left_shifter_0.A0
rlabel metal1 -5048 -15349 -5048 -15349 3 left_shifter_0.A1
rlabel metal1 -5048 -16163 -5048 -16163 3 left_shifter_0.A2
rlabel metal1 -5048 -16985 -5048 -16985 3 left_shifter_0.A3
rlabel metal1 -5048 -17809 -5048 -17809 3 left_shifter_0.A4
rlabel metal1 -5048 -18628 -5048 -18628 3 left_shifter_0.A5
rlabel metal1 -5048 -19444 -5048 -19444 3 left_shifter_0.A6
rlabel metal1 -5048 -20258 -5048 -20258 3 left_shifter_0.A7
rlabel metal1 -3774 -15342 -3774 -15342 3 left_shifter_0.S1
rlabel metal1 -3774 -16159 -3774 -16159 3 left_shifter_0.S2
rlabel metal1 -3774 -16978 -3774 -16978 3 left_shifter_0.S3
rlabel metal1 -3774 -17795 -3774 -17795 3 left_shifter_0.S4
rlabel metal1 -3774 -18614 -3774 -18614 3 left_shifter_0.S5
rlabel metal1 -3774 -19451 -3774 -19451 3 left_shifter_0.S6
rlabel metal1 -3774 -20246 -3774 -20246 3 left_shifter_0.S7
rlabel metal1 -3774 -21065 -3774 -21065 3 left_shifter_0.C
rlabel metal4 -5026 -17809 -5026 -17809 3 left_shifter_0.VDD
rlabel metal5 -3774 -17812 -3774 -17812 3 left_shifter_0.VSS
rlabel metal1 -3774 -14531 -3774 -14531 3 left_shifter_0.S0
rlabel metal1 -4524 -14103 -4524 -14103 5 left_shifter_0.inv_0.A
rlabel metal1 -4135 -14301 -4135 -14301 3 left_shifter_0.inv_0.VSS
rlabel metal1 -4932 -14313 -4932 -14313 3 left_shifter_0.inv_0.VDD
rlabel metal1 -4524 -14515 -4524 -14515 5 left_shifter_0.inv_0.Y
rlabel metal1 -4527 -15362 -4527 -15362 5 left_shifter_0.buffer_7.A
rlabel metal1 -4135 -15800 -4135 -15800 3 left_shifter_0.buffer_7.VSS
rlabel metal1 -4542 -16153 -4542 -16153 5 left_shifter_0.buffer_7.Y
rlabel metal1 -4932 -15813 -4932 -15813 3 left_shifter_0.buffer_7.VDD
rlabel metal1 -4524 -15741 -4524 -15741 5 left_shifter_0.buffer_7.inv_1.A
rlabel metal1 -4135 -15939 -4135 -15939 3 left_shifter_0.buffer_7.inv_1.VSS
rlabel metal1 -4932 -15951 -4932 -15951 3 left_shifter_0.buffer_7.inv_1.VDD
rlabel metal1 -4524 -16153 -4524 -16153 5 left_shifter_0.buffer_7.inv_1.Y
rlabel metal1 -4524 -15362 -4524 -15362 5 left_shifter_0.buffer_7.inv_0.A
rlabel metal1 -4135 -15560 -4135 -15560 3 left_shifter_0.buffer_7.inv_0.VSS
rlabel metal1 -4932 -15572 -4932 -15572 3 left_shifter_0.buffer_7.inv_0.VDD
rlabel metal1 -4524 -15774 -4524 -15774 5 left_shifter_0.buffer_7.inv_0.Y
rlabel metal1 -4527 -14543 -4527 -14543 5 left_shifter_0.buffer_6.A
rlabel metal1 -4135 -14981 -4135 -14981 3 left_shifter_0.buffer_6.VSS
rlabel metal1 -4542 -15334 -4542 -15334 5 left_shifter_0.buffer_6.Y
rlabel metal1 -4932 -14994 -4932 -14994 3 left_shifter_0.buffer_6.VDD
rlabel metal1 -4524 -14922 -4524 -14922 5 left_shifter_0.buffer_6.inv_1.A
rlabel metal1 -4135 -15120 -4135 -15120 3 left_shifter_0.buffer_6.inv_1.VSS
rlabel metal1 -4932 -15132 -4932 -15132 3 left_shifter_0.buffer_6.inv_1.VDD
rlabel metal1 -4524 -15334 -4524 -15334 5 left_shifter_0.buffer_6.inv_1.Y
rlabel metal1 -4524 -14543 -4524 -14543 5 left_shifter_0.buffer_6.inv_0.A
rlabel metal1 -4135 -14741 -4135 -14741 3 left_shifter_0.buffer_6.inv_0.VSS
rlabel metal1 -4932 -14753 -4932 -14753 3 left_shifter_0.buffer_6.inv_0.VDD
rlabel metal1 -4524 -14955 -4524 -14955 5 left_shifter_0.buffer_6.inv_0.Y
rlabel metal1 -4527 -17000 -4527 -17000 5 left_shifter_0.buffer_5.A
rlabel metal1 -4135 -17438 -4135 -17438 3 left_shifter_0.buffer_5.VSS
rlabel metal1 -4542 -17791 -4542 -17791 5 left_shifter_0.buffer_5.Y
rlabel metal1 -4932 -17451 -4932 -17451 3 left_shifter_0.buffer_5.VDD
rlabel metal1 -4524 -17379 -4524 -17379 5 left_shifter_0.buffer_5.inv_1.A
rlabel metal1 -4135 -17577 -4135 -17577 3 left_shifter_0.buffer_5.inv_1.VSS
rlabel metal1 -4932 -17589 -4932 -17589 3 left_shifter_0.buffer_5.inv_1.VDD
rlabel metal1 -4524 -17791 -4524 -17791 5 left_shifter_0.buffer_5.inv_1.Y
rlabel metal1 -4524 -17000 -4524 -17000 5 left_shifter_0.buffer_5.inv_0.A
rlabel metal1 -4135 -17198 -4135 -17198 3 left_shifter_0.buffer_5.inv_0.VSS
rlabel metal1 -4932 -17210 -4932 -17210 3 left_shifter_0.buffer_5.inv_0.VDD
rlabel metal1 -4524 -17412 -4524 -17412 5 left_shifter_0.buffer_5.inv_0.Y
rlabel metal1 -4527 -17819 -4527 -17819 5 left_shifter_0.buffer_4.A
rlabel metal1 -4135 -18257 -4135 -18257 3 left_shifter_0.buffer_4.VSS
rlabel metal1 -4542 -18610 -4542 -18610 5 left_shifter_0.buffer_4.Y
rlabel metal1 -4932 -18270 -4932 -18270 3 left_shifter_0.buffer_4.VDD
rlabel metal1 -4524 -18198 -4524 -18198 5 left_shifter_0.buffer_4.inv_1.A
rlabel metal1 -4135 -18396 -4135 -18396 3 left_shifter_0.buffer_4.inv_1.VSS
rlabel metal1 -4932 -18408 -4932 -18408 3 left_shifter_0.buffer_4.inv_1.VDD
rlabel metal1 -4524 -18610 -4524 -18610 5 left_shifter_0.buffer_4.inv_1.Y
rlabel metal1 -4524 -17819 -4524 -17819 5 left_shifter_0.buffer_4.inv_0.A
rlabel metal1 -4135 -18017 -4135 -18017 3 left_shifter_0.buffer_4.inv_0.VSS
rlabel metal1 -4932 -18029 -4932 -18029 3 left_shifter_0.buffer_4.inv_0.VDD
rlabel metal1 -4524 -18231 -4524 -18231 5 left_shifter_0.buffer_4.inv_0.Y
rlabel metal1 -4527 -18638 -4527 -18638 5 left_shifter_0.buffer_3.A
rlabel metal1 -4135 -19076 -4135 -19076 3 left_shifter_0.buffer_3.VSS
rlabel metal1 -4542 -19429 -4542 -19429 5 left_shifter_0.buffer_3.Y
rlabel metal1 -4932 -19089 -4932 -19089 3 left_shifter_0.buffer_3.VDD
rlabel metal1 -4524 -19017 -4524 -19017 5 left_shifter_0.buffer_3.inv_1.A
rlabel metal1 -4135 -19215 -4135 -19215 3 left_shifter_0.buffer_3.inv_1.VSS
rlabel metal1 -4932 -19227 -4932 -19227 3 left_shifter_0.buffer_3.inv_1.VDD
rlabel metal1 -4524 -19429 -4524 -19429 5 left_shifter_0.buffer_3.inv_1.Y
rlabel metal1 -4524 -18638 -4524 -18638 5 left_shifter_0.buffer_3.inv_0.A
rlabel metal1 -4135 -18836 -4135 -18836 3 left_shifter_0.buffer_3.inv_0.VSS
rlabel metal1 -4932 -18848 -4932 -18848 3 left_shifter_0.buffer_3.inv_0.VDD
rlabel metal1 -4524 -19050 -4524 -19050 5 left_shifter_0.buffer_3.inv_0.Y
rlabel metal1 -4527 -19457 -4527 -19457 5 left_shifter_0.buffer_2.A
rlabel metal1 -4135 -19895 -4135 -19895 3 left_shifter_0.buffer_2.VSS
rlabel metal1 -4542 -20248 -4542 -20248 5 left_shifter_0.buffer_2.Y
rlabel metal1 -4932 -19908 -4932 -19908 3 left_shifter_0.buffer_2.VDD
rlabel metal1 -4524 -19836 -4524 -19836 5 left_shifter_0.buffer_2.inv_1.A
rlabel metal1 -4135 -20034 -4135 -20034 3 left_shifter_0.buffer_2.inv_1.VSS
rlabel metal1 -4932 -20046 -4932 -20046 3 left_shifter_0.buffer_2.inv_1.VDD
rlabel metal1 -4524 -20248 -4524 -20248 5 left_shifter_0.buffer_2.inv_1.Y
rlabel metal1 -4524 -19457 -4524 -19457 5 left_shifter_0.buffer_2.inv_0.A
rlabel metal1 -4135 -19655 -4135 -19655 3 left_shifter_0.buffer_2.inv_0.VSS
rlabel metal1 -4932 -19667 -4932 -19667 3 left_shifter_0.buffer_2.inv_0.VDD
rlabel metal1 -4524 -19869 -4524 -19869 5 left_shifter_0.buffer_2.inv_0.Y
rlabel metal1 -4527 -20276 -4527 -20276 5 left_shifter_0.buffer_1.A
rlabel metal1 -4135 -20714 -4135 -20714 3 left_shifter_0.buffer_1.VSS
rlabel metal1 -4542 -21067 -4542 -21067 5 left_shifter_0.buffer_1.Y
rlabel metal1 -4932 -20727 -4932 -20727 3 left_shifter_0.buffer_1.VDD
rlabel metal1 -4524 -20655 -4524 -20655 5 left_shifter_0.buffer_1.inv_1.A
rlabel metal1 -4135 -20853 -4135 -20853 3 left_shifter_0.buffer_1.inv_1.VSS
rlabel metal1 -4932 -20865 -4932 -20865 3 left_shifter_0.buffer_1.inv_1.VDD
rlabel metal1 -4524 -21067 -4524 -21067 5 left_shifter_0.buffer_1.inv_1.Y
rlabel metal1 -4524 -20276 -4524 -20276 5 left_shifter_0.buffer_1.inv_0.A
rlabel metal1 -4135 -20474 -4135 -20474 3 left_shifter_0.buffer_1.inv_0.VSS
rlabel metal1 -4932 -20486 -4932 -20486 3 left_shifter_0.buffer_1.inv_0.VDD
rlabel metal1 -4524 -20688 -4524 -20688 5 left_shifter_0.buffer_1.inv_0.Y
rlabel metal1 -4527 -16181 -4527 -16181 5 left_shifter_0.buffer_0.A
rlabel metal1 -4135 -16619 -4135 -16619 3 left_shifter_0.buffer_0.VSS
rlabel metal1 -4542 -16972 -4542 -16972 5 left_shifter_0.buffer_0.Y
rlabel metal1 -4932 -16632 -4932 -16632 3 left_shifter_0.buffer_0.VDD
rlabel metal1 -4524 -16560 -4524 -16560 5 left_shifter_0.buffer_0.inv_1.A
rlabel metal1 -4135 -16758 -4135 -16758 3 left_shifter_0.buffer_0.inv_1.VSS
rlabel metal1 -4932 -16770 -4932 -16770 3 left_shifter_0.buffer_0.inv_1.VDD
rlabel metal1 -4524 -16972 -4524 -16972 5 left_shifter_0.buffer_0.inv_1.Y
rlabel metal1 -4524 -16181 -4524 -16181 5 left_shifter_0.buffer_0.inv_0.A
rlabel metal1 -4135 -16379 -4135 -16379 3 left_shifter_0.buffer_0.inv_0.VSS
rlabel metal1 -4932 -16391 -4932 -16391 3 left_shifter_0.buffer_0.inv_0.VDD
rlabel metal1 -4524 -16593 -4524 -16593 5 left_shifter_0.buffer_0.inv_0.Y
flabel space 9272 -28311 9338 -28245 0 FreeSans 1600 0 0 0 mux8_8.000
flabel space 10238 -28318 10245 -28316 0 FreeSans 1600 0 0 0 mux8_8.001
flabel space 7382 -28312 7385 -28312 0 FreeSans 1600 0 0 0 mux8_8.010
flabel space 8270 -28307 8594 -28248 0 FreeSans 1600 0 0 0 mux8_8.011
flabel space 9211 -32023 9637 -31966 0 FreeSans 1600 0 0 0 mux8_8.100
flabel space 10193 -32045 10471 -31886 0 FreeSans 1600 0 0 0 mux8_8.101
flabel space 7299 -32096 7617 -31921 0 FreeSans 1600 0 0 0 mux8_8.110
flabel space 8304 -32074 8622 -31899 0 FreeSans 1600 0 0 0 mux8_8.111
flabel metal2 5740 -29238 5792 -29186 0 FreeSans 160 0 0 0 mux8_8.A0
flabel metal2 5743 -29333 5795 -29281 0 FreeSans 160 0 0 0 mux8_8.A1
flabel metal2 5746 -29439 5798 -29387 0 FreeSans 160 0 0 0 mux8_8.A2
flabel metal2 5741 -29545 5793 -29493 0 FreeSans 160 0 0 0 mux8_8.A3
flabel metal2 5744 -30643 5796 -30591 0 FreeSans 160 0 0 0 mux8_8.A4
flabel metal2 5746 -30767 5798 -30715 0 FreeSans 160 0 0 0 mux8_8.A5
flabel metal2 5743 -30863 5795 -30811 0 FreeSans 160 0 0 0 mux8_8.A6
flabel metal2 5739 -30984 5791 -30932 0 FreeSans 160 0 0 0 mux8_8.A7
flabel metal1 12377 -28599 12429 -28547 0 FreeSans 160 0 0 0 mux8_8.VDD
flabel metal1 13159 -30239 13211 -30187 0 FreeSans 160 0 0 0 mux8_8.Y
flabel metal5 12955 -30886 13007 -30834 0 FreeSans 160 0 0 0 mux8_8.VSS
flabel metal2 6448 -27615 6493 -27576 0 FreeSans 160 0 0 0 mux8_8.SEL0
flabel metal2 6007 -27624 6052 -27585 0 FreeSans 160 0 0 0 mux8_8.SEL1
flabel metal2 5569 -27624 5614 -27585 0 FreeSans 160 0 0 0 mux8_8.SEL2
flabel metal1 8057 -29172 8091 -29123 0 FreeSans 160 0 0 0 mux8_8.NAND4F_2.A
flabel metal1 8060 -29072 8094 -29023 0 FreeSans 160 0 0 0 mux8_8.NAND4F_2.B
flabel metal1 8061 -28984 8095 -28935 0 FreeSans 160 0 0 0 mux8_8.NAND4F_2.C
flabel metal1 8062 -28891 8096 -28842 0 FreeSans 160 0 0 0 mux8_8.NAND4F_2.D
flabel metal1 8199 -29990 8233 -29941 0 FreeSans 160 0 0 0 mux8_8.NAND4F_2.VSS
flabel nwell 8462 -28429 8496 -28380 0 FreeSans 160 0 0 0 mux8_8.NAND4F_2.VDD
flabel metal1 8895 -29109 8929 -29060 0 FreeSans 160 0 0 0 mux8_8.NAND4F_2.Y
flabel metal1 7109 -29172 7143 -29123 0 FreeSans 160 0 0 0 mux8_8.NAND4F_4.A
flabel metal1 7112 -29072 7146 -29023 0 FreeSans 160 0 0 0 mux8_8.NAND4F_4.B
flabel metal1 7113 -28984 7147 -28935 0 FreeSans 160 0 0 0 mux8_8.NAND4F_4.C
flabel metal1 7114 -28891 7148 -28842 0 FreeSans 160 0 0 0 mux8_8.NAND4F_4.D
flabel metal1 7251 -29990 7285 -29941 0 FreeSans 160 0 0 0 mux8_8.NAND4F_4.VSS
flabel nwell 7514 -28429 7548 -28380 0 FreeSans 160 0 0 0 mux8_8.NAND4F_4.VDD
flabel metal1 7947 -29109 7981 -29060 0 FreeSans 160 0 0 0 mux8_8.NAND4F_4.Y
flabel metal1 7109 -31017 7143 -30968 0 FreeSans 160 0 0 0 mux8_8.NAND4F_5.A
flabel metal1 7112 -31117 7146 -31068 0 FreeSans 160 0 0 0 mux8_8.NAND4F_5.B
flabel metal1 7113 -31205 7147 -31156 0 FreeSans 160 0 0 0 mux8_8.NAND4F_5.C
flabel metal1 7114 -31298 7148 -31249 0 FreeSans 160 0 0 0 mux8_8.NAND4F_5.D
flabel metal1 7251 -30199 7285 -30150 0 FreeSans 160 0 0 0 mux8_8.NAND4F_5.VSS
flabel nwell 7514 -31760 7548 -31711 0 FreeSans 160 0 0 0 mux8_8.NAND4F_5.VDD
flabel metal1 7947 -31080 7981 -31031 0 FreeSans 160 0 0 0 mux8_8.NAND4F_5.Y
flabel metal1 8057 -31017 8091 -30968 0 FreeSans 160 0 0 0 mux8_8.NAND4F_6.A
flabel metal1 8060 -31117 8094 -31068 0 FreeSans 160 0 0 0 mux8_8.NAND4F_6.B
flabel metal1 8061 -31205 8095 -31156 0 FreeSans 160 0 0 0 mux8_8.NAND4F_6.C
flabel metal1 8062 -31298 8096 -31249 0 FreeSans 160 0 0 0 mux8_8.NAND4F_6.D
flabel metal1 8199 -30199 8233 -30150 0 FreeSans 160 0 0 0 mux8_8.NAND4F_6.VSS
flabel nwell 8462 -31760 8496 -31711 0 FreeSans 160 0 0 0 mux8_8.NAND4F_6.VDD
flabel metal1 8895 -31080 8929 -31031 0 FreeSans 160 0 0 0 mux8_8.NAND4F_6.Y
flabel metal1 9924 -29172 9958 -29123 0 FreeSans 160 0 0 0 mux8_8.NAND4F_0.A
flabel metal1 9927 -29072 9961 -29023 0 FreeSans 160 0 0 0 mux8_8.NAND4F_0.B
flabel metal1 9928 -28984 9962 -28935 0 FreeSans 160 0 0 0 mux8_8.NAND4F_0.C
flabel metal1 9929 -28891 9963 -28842 0 FreeSans 160 0 0 0 mux8_8.NAND4F_0.D
flabel metal1 10066 -29990 10100 -29941 0 FreeSans 160 0 0 0 mux8_8.NAND4F_0.VSS
flabel nwell 10329 -28429 10363 -28380 0 FreeSans 160 0 0 0 mux8_8.NAND4F_0.VDD
flabel metal1 10762 -29109 10796 -29060 0 FreeSans 160 0 0 0 mux8_8.NAND4F_0.Y
flabel metal1 8993 -31017 9027 -30968 0 FreeSans 160 0 0 0 mux8_8.NAND4F_1.A
flabel metal1 8996 -31117 9030 -31068 0 FreeSans 160 0 0 0 mux8_8.NAND4F_1.B
flabel metal1 8997 -31205 9031 -31156 0 FreeSans 160 0 0 0 mux8_8.NAND4F_1.C
flabel metal1 8998 -31298 9032 -31249 0 FreeSans 160 0 0 0 mux8_8.NAND4F_1.D
flabel metal1 9135 -30199 9169 -30150 0 FreeSans 160 0 0 0 mux8_8.NAND4F_1.VSS
flabel nwell 9398 -31760 9432 -31711 0 FreeSans 160 0 0 0 mux8_8.NAND4F_1.VDD
flabel metal1 9831 -31080 9865 -31031 0 FreeSans 160 0 0 0 mux8_8.NAND4F_1.Y
flabel metal1 8993 -29172 9027 -29123 0 FreeSans 160 0 0 0 mux8_8.NAND4F_3.A
flabel metal1 8996 -29072 9030 -29023 0 FreeSans 160 0 0 0 mux8_8.NAND4F_3.B
flabel metal1 8997 -28984 9031 -28935 0 FreeSans 160 0 0 0 mux8_8.NAND4F_3.C
flabel metal1 8998 -28891 9032 -28842 0 FreeSans 160 0 0 0 mux8_8.NAND4F_3.D
flabel metal1 9135 -29990 9169 -29941 0 FreeSans 160 0 0 0 mux8_8.NAND4F_3.VSS
flabel nwell 9398 -28429 9432 -28380 0 FreeSans 160 0 0 0 mux8_8.NAND4F_3.VDD
flabel metal1 9831 -29109 9865 -29060 0 FreeSans 160 0 0 0 mux8_8.NAND4F_3.Y
flabel metal1 9924 -31016 9958 -30967 0 FreeSans 160 0 0 0 mux8_8.NAND4F_7.A
flabel metal1 9927 -31116 9961 -31067 0 FreeSans 160 0 0 0 mux8_8.NAND4F_7.B
flabel metal1 9928 -31204 9962 -31155 0 FreeSans 160 0 0 0 mux8_8.NAND4F_7.C
flabel metal1 9929 -31297 9963 -31248 0 FreeSans 160 0 0 0 mux8_8.NAND4F_7.D
flabel metal1 10066 -30198 10100 -30149 0 FreeSans 160 0 0 0 mux8_8.NAND4F_7.VSS
flabel nwell 10329 -31759 10363 -31710 0 FreeSans 160 0 0 0 mux8_8.NAND4F_7.VDD
flabel metal1 10762 -31079 10796 -31030 0 FreeSans 160 0 0 0 mux8_8.NAND4F_7.Y
flabel metal1 10851 -29172 10885 -29123 0 FreeSans 160 0 0 0 mux8_8.NAND4F_8.A
flabel metal1 10854 -29072 10888 -29023 0 FreeSans 160 0 0 0 mux8_8.NAND4F_8.B
flabel metal1 10855 -28984 10889 -28935 0 FreeSans 160 0 0 0 mux8_8.NAND4F_8.C
flabel metal1 10856 -28891 10890 -28842 0 FreeSans 160 0 0 0 mux8_8.NAND4F_8.D
flabel metal1 10993 -29990 11027 -29941 0 FreeSans 160 0 0 0 mux8_8.NAND4F_8.VSS
flabel nwell 11256 -28429 11290 -28380 0 FreeSans 160 0 0 0 mux8_8.NAND4F_8.VDD
flabel metal1 11689 -29109 11723 -29060 0 FreeSans 160 0 0 0 mux8_8.NAND4F_8.Y
flabel metal1 10851 -31017 10885 -30968 0 FreeSans 160 0 0 0 mux8_8.NAND4F_9.A
flabel metal1 10854 -31117 10888 -31068 0 FreeSans 160 0 0 0 mux8_8.NAND4F_9.B
flabel metal1 10855 -31205 10889 -31156 0 FreeSans 160 0 0 0 mux8_8.NAND4F_9.C
flabel metal1 10856 -31298 10890 -31249 0 FreeSans 160 0 0 0 mux8_8.NAND4F_9.D
flabel metal1 10993 -30199 11027 -30150 0 FreeSans 160 0 0 0 mux8_8.NAND4F_9.VSS
flabel nwell 11256 -31760 11290 -31711 0 FreeSans 160 0 0 0 mux8_8.NAND4F_9.VDD
flabel metal1 11689 -31080 11723 -31031 0 FreeSans 160 0 0 0 mux8_8.NAND4F_9.Y
rlabel metal1 12823 -30095 12823 -30095 3 mux8_8.inv_0.A
rlabel metal1 13021 -30484 13021 -30484 5 mux8_8.inv_0.VSS
rlabel metal1 13033 -29687 13033 -29687 5 mux8_8.inv_0.VDD
rlabel metal1 13235 -30095 13235 -30095 3 mux8_8.inv_0.Y
flabel metal1 11744 -30036 11821 -29984 1 FreeSerif 320 0 0 0 mux8_8.nor2_0.A
rlabel metal1 11990 -29536 11990 -29536 5 mux8_8.nor2_0.VDD
flabel metal1 11745 -30142 11822 -30090 1 FreeSerif 320 0 0 0 mux8_8.nor2_0.B
flabel metal1 12749 -30148 12826 -30096 1 FreeSerif 320 0 0 0 mux8_8.nor2_0.Y
rlabel metal1 12286 -30514 12286 -30514 5 mux8_8.nor2_0.VSS
rlabel metal1 5998 -28077 5998 -28077 3 mux8_8.inv_1.A
rlabel metal1 6196 -28466 6196 -28466 5 mux8_8.inv_1.VSS
rlabel metal1 6208 -27669 6208 -27669 5 mux8_8.inv_1.VDD
rlabel metal1 6410 -28077 6410 -28077 3 mux8_8.inv_1.Y
rlabel metal1 6438 -28077 6438 -28077 3 mux8_8.inv_2.A
rlabel metal1 6636 -28466 6636 -28466 5 mux8_8.inv_2.VSS
rlabel metal1 6648 -27669 6648 -27669 5 mux8_8.inv_2.VDD
rlabel metal1 6850 -28077 6850 -28077 3 mux8_8.inv_2.Y
rlabel metal1 5558 -28077 5558 -28077 3 mux8_8.inv_3.A
rlabel metal1 5756 -28466 5756 -28466 5 mux8_8.inv_3.VSS
rlabel metal1 5768 -27669 5768 -27669 5 mux8_8.inv_3.VDD
rlabel metal1 5970 -28077 5970 -28077 3 mux8_8.inv_3.Y
flabel space 9272 -23783 9338 -23717 0 FreeSans 1600 0 0 0 mux8_7.000
flabel space 10238 -23790 10245 -23788 0 FreeSans 1600 0 0 0 mux8_7.001
flabel space 7382 -23784 7385 -23784 0 FreeSans 1600 0 0 0 mux8_7.010
flabel space 8270 -23779 8594 -23720 0 FreeSans 1600 0 0 0 mux8_7.011
flabel space 9211 -27495 9637 -27438 0 FreeSans 1600 0 0 0 mux8_7.100
flabel space 10193 -27517 10471 -27358 0 FreeSans 1600 0 0 0 mux8_7.101
flabel space 7299 -27568 7617 -27393 0 FreeSans 1600 0 0 0 mux8_7.110
flabel space 8304 -27546 8622 -27371 0 FreeSans 1600 0 0 0 mux8_7.111
flabel metal2 5740 -24710 5792 -24658 0 FreeSans 160 0 0 0 mux8_7.A0
flabel metal2 5743 -24805 5795 -24753 0 FreeSans 160 0 0 0 mux8_7.A1
flabel metal2 5746 -24911 5798 -24859 0 FreeSans 160 0 0 0 mux8_7.A2
flabel metal2 5741 -25017 5793 -24965 0 FreeSans 160 0 0 0 mux8_7.A3
flabel metal2 5744 -26115 5796 -26063 0 FreeSans 160 0 0 0 mux8_7.A4
flabel metal2 5746 -26239 5798 -26187 0 FreeSans 160 0 0 0 mux8_7.A5
flabel metal2 5743 -26335 5795 -26283 0 FreeSans 160 0 0 0 mux8_7.A6
flabel metal2 5739 -26456 5791 -26404 0 FreeSans 160 0 0 0 mux8_7.A7
flabel metal1 12377 -24071 12429 -24019 0 FreeSans 160 0 0 0 mux8_7.VDD
flabel metal1 13159 -25711 13211 -25659 0 FreeSans 160 0 0 0 mux8_7.Y
flabel metal5 12955 -26358 13007 -26306 0 FreeSans 160 0 0 0 mux8_7.VSS
flabel metal2 6448 -23087 6493 -23048 0 FreeSans 160 0 0 0 mux8_7.SEL0
flabel metal2 6007 -23096 6052 -23057 0 FreeSans 160 0 0 0 mux8_7.SEL1
flabel metal2 5569 -23096 5614 -23057 0 FreeSans 160 0 0 0 mux8_7.SEL2
flabel metal1 8057 -24644 8091 -24595 0 FreeSans 160 0 0 0 mux8_7.NAND4F_2.A
flabel metal1 8060 -24544 8094 -24495 0 FreeSans 160 0 0 0 mux8_7.NAND4F_2.B
flabel metal1 8061 -24456 8095 -24407 0 FreeSans 160 0 0 0 mux8_7.NAND4F_2.C
flabel metal1 8062 -24363 8096 -24314 0 FreeSans 160 0 0 0 mux8_7.NAND4F_2.D
flabel metal1 8199 -25462 8233 -25413 0 FreeSans 160 0 0 0 mux8_7.NAND4F_2.VSS
flabel nwell 8462 -23901 8496 -23852 0 FreeSans 160 0 0 0 mux8_7.NAND4F_2.VDD
flabel metal1 8895 -24581 8929 -24532 0 FreeSans 160 0 0 0 mux8_7.NAND4F_2.Y
flabel metal1 7109 -24644 7143 -24595 0 FreeSans 160 0 0 0 mux8_7.NAND4F_4.A
flabel metal1 7112 -24544 7146 -24495 0 FreeSans 160 0 0 0 mux8_7.NAND4F_4.B
flabel metal1 7113 -24456 7147 -24407 0 FreeSans 160 0 0 0 mux8_7.NAND4F_4.C
flabel metal1 7114 -24363 7148 -24314 0 FreeSans 160 0 0 0 mux8_7.NAND4F_4.D
flabel metal1 7251 -25462 7285 -25413 0 FreeSans 160 0 0 0 mux8_7.NAND4F_4.VSS
flabel nwell 7514 -23901 7548 -23852 0 FreeSans 160 0 0 0 mux8_7.NAND4F_4.VDD
flabel metal1 7947 -24581 7981 -24532 0 FreeSans 160 0 0 0 mux8_7.NAND4F_4.Y
flabel metal1 7109 -26489 7143 -26440 0 FreeSans 160 0 0 0 mux8_7.NAND4F_5.A
flabel metal1 7112 -26589 7146 -26540 0 FreeSans 160 0 0 0 mux8_7.NAND4F_5.B
flabel metal1 7113 -26677 7147 -26628 0 FreeSans 160 0 0 0 mux8_7.NAND4F_5.C
flabel metal1 7114 -26770 7148 -26721 0 FreeSans 160 0 0 0 mux8_7.NAND4F_5.D
flabel metal1 7251 -25671 7285 -25622 0 FreeSans 160 0 0 0 mux8_7.NAND4F_5.VSS
flabel nwell 7514 -27232 7548 -27183 0 FreeSans 160 0 0 0 mux8_7.NAND4F_5.VDD
flabel metal1 7947 -26552 7981 -26503 0 FreeSans 160 0 0 0 mux8_7.NAND4F_5.Y
flabel metal1 8057 -26489 8091 -26440 0 FreeSans 160 0 0 0 mux8_7.NAND4F_6.A
flabel metal1 8060 -26589 8094 -26540 0 FreeSans 160 0 0 0 mux8_7.NAND4F_6.B
flabel metal1 8061 -26677 8095 -26628 0 FreeSans 160 0 0 0 mux8_7.NAND4F_6.C
flabel metal1 8062 -26770 8096 -26721 0 FreeSans 160 0 0 0 mux8_7.NAND4F_6.D
flabel metal1 8199 -25671 8233 -25622 0 FreeSans 160 0 0 0 mux8_7.NAND4F_6.VSS
flabel nwell 8462 -27232 8496 -27183 0 FreeSans 160 0 0 0 mux8_7.NAND4F_6.VDD
flabel metal1 8895 -26552 8929 -26503 0 FreeSans 160 0 0 0 mux8_7.NAND4F_6.Y
flabel metal1 9924 -24644 9958 -24595 0 FreeSans 160 0 0 0 mux8_7.NAND4F_0.A
flabel metal1 9927 -24544 9961 -24495 0 FreeSans 160 0 0 0 mux8_7.NAND4F_0.B
flabel metal1 9928 -24456 9962 -24407 0 FreeSans 160 0 0 0 mux8_7.NAND4F_0.C
flabel metal1 9929 -24363 9963 -24314 0 FreeSans 160 0 0 0 mux8_7.NAND4F_0.D
flabel metal1 10066 -25462 10100 -25413 0 FreeSans 160 0 0 0 mux8_7.NAND4F_0.VSS
flabel nwell 10329 -23901 10363 -23852 0 FreeSans 160 0 0 0 mux8_7.NAND4F_0.VDD
flabel metal1 10762 -24581 10796 -24532 0 FreeSans 160 0 0 0 mux8_7.NAND4F_0.Y
flabel metal1 8993 -26489 9027 -26440 0 FreeSans 160 0 0 0 mux8_7.NAND4F_1.A
flabel metal1 8996 -26589 9030 -26540 0 FreeSans 160 0 0 0 mux8_7.NAND4F_1.B
flabel metal1 8997 -26677 9031 -26628 0 FreeSans 160 0 0 0 mux8_7.NAND4F_1.C
flabel metal1 8998 -26770 9032 -26721 0 FreeSans 160 0 0 0 mux8_7.NAND4F_1.D
flabel metal1 9135 -25671 9169 -25622 0 FreeSans 160 0 0 0 mux8_7.NAND4F_1.VSS
flabel nwell 9398 -27232 9432 -27183 0 FreeSans 160 0 0 0 mux8_7.NAND4F_1.VDD
flabel metal1 9831 -26552 9865 -26503 0 FreeSans 160 0 0 0 mux8_7.NAND4F_1.Y
flabel metal1 8993 -24644 9027 -24595 0 FreeSans 160 0 0 0 mux8_7.NAND4F_3.A
flabel metal1 8996 -24544 9030 -24495 0 FreeSans 160 0 0 0 mux8_7.NAND4F_3.B
flabel metal1 8997 -24456 9031 -24407 0 FreeSans 160 0 0 0 mux8_7.NAND4F_3.C
flabel metal1 8998 -24363 9032 -24314 0 FreeSans 160 0 0 0 mux8_7.NAND4F_3.D
flabel metal1 9135 -25462 9169 -25413 0 FreeSans 160 0 0 0 mux8_7.NAND4F_3.VSS
flabel nwell 9398 -23901 9432 -23852 0 FreeSans 160 0 0 0 mux8_7.NAND4F_3.VDD
flabel metal1 9831 -24581 9865 -24532 0 FreeSans 160 0 0 0 mux8_7.NAND4F_3.Y
flabel metal1 9924 -26488 9958 -26439 0 FreeSans 160 0 0 0 mux8_7.NAND4F_7.A
flabel metal1 9927 -26588 9961 -26539 0 FreeSans 160 0 0 0 mux8_7.NAND4F_7.B
flabel metal1 9928 -26676 9962 -26627 0 FreeSans 160 0 0 0 mux8_7.NAND4F_7.C
flabel metal1 9929 -26769 9963 -26720 0 FreeSans 160 0 0 0 mux8_7.NAND4F_7.D
flabel metal1 10066 -25670 10100 -25621 0 FreeSans 160 0 0 0 mux8_7.NAND4F_7.VSS
flabel nwell 10329 -27231 10363 -27182 0 FreeSans 160 0 0 0 mux8_7.NAND4F_7.VDD
flabel metal1 10762 -26551 10796 -26502 0 FreeSans 160 0 0 0 mux8_7.NAND4F_7.Y
flabel metal1 10851 -24644 10885 -24595 0 FreeSans 160 0 0 0 mux8_7.NAND4F_8.A
flabel metal1 10854 -24544 10888 -24495 0 FreeSans 160 0 0 0 mux8_7.NAND4F_8.B
flabel metal1 10855 -24456 10889 -24407 0 FreeSans 160 0 0 0 mux8_7.NAND4F_8.C
flabel metal1 10856 -24363 10890 -24314 0 FreeSans 160 0 0 0 mux8_7.NAND4F_8.D
flabel metal1 10993 -25462 11027 -25413 0 FreeSans 160 0 0 0 mux8_7.NAND4F_8.VSS
flabel nwell 11256 -23901 11290 -23852 0 FreeSans 160 0 0 0 mux8_7.NAND4F_8.VDD
flabel metal1 11689 -24581 11723 -24532 0 FreeSans 160 0 0 0 mux8_7.NAND4F_8.Y
flabel metal1 10851 -26489 10885 -26440 0 FreeSans 160 0 0 0 mux8_7.NAND4F_9.A
flabel metal1 10854 -26589 10888 -26540 0 FreeSans 160 0 0 0 mux8_7.NAND4F_9.B
flabel metal1 10855 -26677 10889 -26628 0 FreeSans 160 0 0 0 mux8_7.NAND4F_9.C
flabel metal1 10856 -26770 10890 -26721 0 FreeSans 160 0 0 0 mux8_7.NAND4F_9.D
flabel metal1 10993 -25671 11027 -25622 0 FreeSans 160 0 0 0 mux8_7.NAND4F_9.VSS
flabel nwell 11256 -27232 11290 -27183 0 FreeSans 160 0 0 0 mux8_7.NAND4F_9.VDD
flabel metal1 11689 -26552 11723 -26503 0 FreeSans 160 0 0 0 mux8_7.NAND4F_9.Y
rlabel metal1 12823 -25567 12823 -25567 3 mux8_7.inv_0.A
rlabel metal1 13021 -25956 13021 -25956 5 mux8_7.inv_0.VSS
rlabel metal1 13033 -25159 13033 -25159 5 mux8_7.inv_0.VDD
rlabel metal1 13235 -25567 13235 -25567 3 mux8_7.inv_0.Y
flabel metal1 11744 -25508 11821 -25456 1 FreeSerif 320 0 0 0 mux8_7.nor2_0.A
rlabel metal1 11990 -25008 11990 -25008 5 mux8_7.nor2_0.VDD
flabel metal1 11745 -25614 11822 -25562 1 FreeSerif 320 0 0 0 mux8_7.nor2_0.B
flabel metal1 12749 -25620 12826 -25568 1 FreeSerif 320 0 0 0 mux8_7.nor2_0.Y
rlabel metal1 12286 -25986 12286 -25986 5 mux8_7.nor2_0.VSS
rlabel metal1 5998 -23549 5998 -23549 3 mux8_7.inv_1.A
rlabel metal1 6196 -23938 6196 -23938 5 mux8_7.inv_1.VSS
rlabel metal1 6208 -23141 6208 -23141 5 mux8_7.inv_1.VDD
rlabel metal1 6410 -23549 6410 -23549 3 mux8_7.inv_1.Y
rlabel metal1 6438 -23549 6438 -23549 3 mux8_7.inv_2.A
rlabel metal1 6636 -23938 6636 -23938 5 mux8_7.inv_2.VSS
rlabel metal1 6648 -23141 6648 -23141 5 mux8_7.inv_2.VDD
rlabel metal1 6850 -23549 6850 -23549 3 mux8_7.inv_2.Y
rlabel metal1 5558 -23549 5558 -23549 3 mux8_7.inv_3.A
rlabel metal1 5756 -23938 5756 -23938 5 mux8_7.inv_3.VSS
rlabel metal1 5768 -23141 5768 -23141 5 mux8_7.inv_3.VDD
rlabel metal1 5970 -23549 5970 -23549 3 mux8_7.inv_3.Y
flabel space 9272 -32839 9338 -32773 0 FreeSans 1600 0 0 0 mux8_6.000
flabel space 10238 -32846 10245 -32844 0 FreeSans 1600 0 0 0 mux8_6.001
flabel space 7382 -32840 7385 -32840 0 FreeSans 1600 0 0 0 mux8_6.010
flabel space 8270 -32835 8594 -32776 0 FreeSans 1600 0 0 0 mux8_6.011
flabel space 9211 -36551 9637 -36494 0 FreeSans 1600 0 0 0 mux8_6.100
flabel space 10193 -36573 10471 -36414 0 FreeSans 1600 0 0 0 mux8_6.101
flabel space 7299 -36624 7617 -36449 0 FreeSans 1600 0 0 0 mux8_6.110
flabel space 8304 -36602 8622 -36427 0 FreeSans 1600 0 0 0 mux8_6.111
flabel metal2 5740 -33766 5792 -33714 0 FreeSans 160 0 0 0 mux8_6.A0
flabel metal2 5743 -33861 5795 -33809 0 FreeSans 160 0 0 0 mux8_6.A1
flabel metal2 5746 -33967 5798 -33915 0 FreeSans 160 0 0 0 mux8_6.A2
flabel metal2 5741 -34073 5793 -34021 0 FreeSans 160 0 0 0 mux8_6.A3
flabel metal2 5744 -35171 5796 -35119 0 FreeSans 160 0 0 0 mux8_6.A4
flabel metal2 5746 -35295 5798 -35243 0 FreeSans 160 0 0 0 mux8_6.A5
flabel metal2 5743 -35391 5795 -35339 0 FreeSans 160 0 0 0 mux8_6.A6
flabel metal2 5739 -35512 5791 -35460 0 FreeSans 160 0 0 0 mux8_6.A7
flabel metal1 12377 -33127 12429 -33075 0 FreeSans 160 0 0 0 mux8_6.VDD
flabel metal1 13159 -34767 13211 -34715 0 FreeSans 160 0 0 0 mux8_6.Y
flabel metal5 12955 -35414 13007 -35362 0 FreeSans 160 0 0 0 mux8_6.VSS
flabel metal2 6448 -32143 6493 -32104 0 FreeSans 160 0 0 0 mux8_6.SEL0
flabel metal2 6007 -32152 6052 -32113 0 FreeSans 160 0 0 0 mux8_6.SEL1
flabel metal2 5569 -32152 5614 -32113 0 FreeSans 160 0 0 0 mux8_6.SEL2
flabel metal1 8057 -33700 8091 -33651 0 FreeSans 160 0 0 0 mux8_6.NAND4F_2.A
flabel metal1 8060 -33600 8094 -33551 0 FreeSans 160 0 0 0 mux8_6.NAND4F_2.B
flabel metal1 8061 -33512 8095 -33463 0 FreeSans 160 0 0 0 mux8_6.NAND4F_2.C
flabel metal1 8062 -33419 8096 -33370 0 FreeSans 160 0 0 0 mux8_6.NAND4F_2.D
flabel metal1 8199 -34518 8233 -34469 0 FreeSans 160 0 0 0 mux8_6.NAND4F_2.VSS
flabel nwell 8462 -32957 8496 -32908 0 FreeSans 160 0 0 0 mux8_6.NAND4F_2.VDD
flabel metal1 8895 -33637 8929 -33588 0 FreeSans 160 0 0 0 mux8_6.NAND4F_2.Y
flabel metal1 7109 -33700 7143 -33651 0 FreeSans 160 0 0 0 mux8_6.NAND4F_4.A
flabel metal1 7112 -33600 7146 -33551 0 FreeSans 160 0 0 0 mux8_6.NAND4F_4.B
flabel metal1 7113 -33512 7147 -33463 0 FreeSans 160 0 0 0 mux8_6.NAND4F_4.C
flabel metal1 7114 -33419 7148 -33370 0 FreeSans 160 0 0 0 mux8_6.NAND4F_4.D
flabel metal1 7251 -34518 7285 -34469 0 FreeSans 160 0 0 0 mux8_6.NAND4F_4.VSS
flabel nwell 7514 -32957 7548 -32908 0 FreeSans 160 0 0 0 mux8_6.NAND4F_4.VDD
flabel metal1 7947 -33637 7981 -33588 0 FreeSans 160 0 0 0 mux8_6.NAND4F_4.Y
flabel metal1 7109 -35545 7143 -35496 0 FreeSans 160 0 0 0 mux8_6.NAND4F_5.A
flabel metal1 7112 -35645 7146 -35596 0 FreeSans 160 0 0 0 mux8_6.NAND4F_5.B
flabel metal1 7113 -35733 7147 -35684 0 FreeSans 160 0 0 0 mux8_6.NAND4F_5.C
flabel metal1 7114 -35826 7148 -35777 0 FreeSans 160 0 0 0 mux8_6.NAND4F_5.D
flabel metal1 7251 -34727 7285 -34678 0 FreeSans 160 0 0 0 mux8_6.NAND4F_5.VSS
flabel nwell 7514 -36288 7548 -36239 0 FreeSans 160 0 0 0 mux8_6.NAND4F_5.VDD
flabel metal1 7947 -35608 7981 -35559 0 FreeSans 160 0 0 0 mux8_6.NAND4F_5.Y
flabel metal1 8057 -35545 8091 -35496 0 FreeSans 160 0 0 0 mux8_6.NAND4F_6.A
flabel metal1 8060 -35645 8094 -35596 0 FreeSans 160 0 0 0 mux8_6.NAND4F_6.B
flabel metal1 8061 -35733 8095 -35684 0 FreeSans 160 0 0 0 mux8_6.NAND4F_6.C
flabel metal1 8062 -35826 8096 -35777 0 FreeSans 160 0 0 0 mux8_6.NAND4F_6.D
flabel metal1 8199 -34727 8233 -34678 0 FreeSans 160 0 0 0 mux8_6.NAND4F_6.VSS
flabel nwell 8462 -36288 8496 -36239 0 FreeSans 160 0 0 0 mux8_6.NAND4F_6.VDD
flabel metal1 8895 -35608 8929 -35559 0 FreeSans 160 0 0 0 mux8_6.NAND4F_6.Y
flabel metal1 9924 -33700 9958 -33651 0 FreeSans 160 0 0 0 mux8_6.NAND4F_0.A
flabel metal1 9927 -33600 9961 -33551 0 FreeSans 160 0 0 0 mux8_6.NAND4F_0.B
flabel metal1 9928 -33512 9962 -33463 0 FreeSans 160 0 0 0 mux8_6.NAND4F_0.C
flabel metal1 9929 -33419 9963 -33370 0 FreeSans 160 0 0 0 mux8_6.NAND4F_0.D
flabel metal1 10066 -34518 10100 -34469 0 FreeSans 160 0 0 0 mux8_6.NAND4F_0.VSS
flabel nwell 10329 -32957 10363 -32908 0 FreeSans 160 0 0 0 mux8_6.NAND4F_0.VDD
flabel metal1 10762 -33637 10796 -33588 0 FreeSans 160 0 0 0 mux8_6.NAND4F_0.Y
flabel metal1 8993 -35545 9027 -35496 0 FreeSans 160 0 0 0 mux8_6.NAND4F_1.A
flabel metal1 8996 -35645 9030 -35596 0 FreeSans 160 0 0 0 mux8_6.NAND4F_1.B
flabel metal1 8997 -35733 9031 -35684 0 FreeSans 160 0 0 0 mux8_6.NAND4F_1.C
flabel metal1 8998 -35826 9032 -35777 0 FreeSans 160 0 0 0 mux8_6.NAND4F_1.D
flabel metal1 9135 -34727 9169 -34678 0 FreeSans 160 0 0 0 mux8_6.NAND4F_1.VSS
flabel nwell 9398 -36288 9432 -36239 0 FreeSans 160 0 0 0 mux8_6.NAND4F_1.VDD
flabel metal1 9831 -35608 9865 -35559 0 FreeSans 160 0 0 0 mux8_6.NAND4F_1.Y
flabel metal1 8993 -33700 9027 -33651 0 FreeSans 160 0 0 0 mux8_6.NAND4F_3.A
flabel metal1 8996 -33600 9030 -33551 0 FreeSans 160 0 0 0 mux8_6.NAND4F_3.B
flabel metal1 8997 -33512 9031 -33463 0 FreeSans 160 0 0 0 mux8_6.NAND4F_3.C
flabel metal1 8998 -33419 9032 -33370 0 FreeSans 160 0 0 0 mux8_6.NAND4F_3.D
flabel metal1 9135 -34518 9169 -34469 0 FreeSans 160 0 0 0 mux8_6.NAND4F_3.VSS
flabel nwell 9398 -32957 9432 -32908 0 FreeSans 160 0 0 0 mux8_6.NAND4F_3.VDD
flabel metal1 9831 -33637 9865 -33588 0 FreeSans 160 0 0 0 mux8_6.NAND4F_3.Y
flabel metal1 9924 -35544 9958 -35495 0 FreeSans 160 0 0 0 mux8_6.NAND4F_7.A
flabel metal1 9927 -35644 9961 -35595 0 FreeSans 160 0 0 0 mux8_6.NAND4F_7.B
flabel metal1 9928 -35732 9962 -35683 0 FreeSans 160 0 0 0 mux8_6.NAND4F_7.C
flabel metal1 9929 -35825 9963 -35776 0 FreeSans 160 0 0 0 mux8_6.NAND4F_7.D
flabel metal1 10066 -34726 10100 -34677 0 FreeSans 160 0 0 0 mux8_6.NAND4F_7.VSS
flabel nwell 10329 -36287 10363 -36238 0 FreeSans 160 0 0 0 mux8_6.NAND4F_7.VDD
flabel metal1 10762 -35607 10796 -35558 0 FreeSans 160 0 0 0 mux8_6.NAND4F_7.Y
flabel metal1 10851 -33700 10885 -33651 0 FreeSans 160 0 0 0 mux8_6.NAND4F_8.A
flabel metal1 10854 -33600 10888 -33551 0 FreeSans 160 0 0 0 mux8_6.NAND4F_8.B
flabel metal1 10855 -33512 10889 -33463 0 FreeSans 160 0 0 0 mux8_6.NAND4F_8.C
flabel metal1 10856 -33419 10890 -33370 0 FreeSans 160 0 0 0 mux8_6.NAND4F_8.D
flabel metal1 10993 -34518 11027 -34469 0 FreeSans 160 0 0 0 mux8_6.NAND4F_8.VSS
flabel nwell 11256 -32957 11290 -32908 0 FreeSans 160 0 0 0 mux8_6.NAND4F_8.VDD
flabel metal1 11689 -33637 11723 -33588 0 FreeSans 160 0 0 0 mux8_6.NAND4F_8.Y
flabel metal1 10851 -35545 10885 -35496 0 FreeSans 160 0 0 0 mux8_6.NAND4F_9.A
flabel metal1 10854 -35645 10888 -35596 0 FreeSans 160 0 0 0 mux8_6.NAND4F_9.B
flabel metal1 10855 -35733 10889 -35684 0 FreeSans 160 0 0 0 mux8_6.NAND4F_9.C
flabel metal1 10856 -35826 10890 -35777 0 FreeSans 160 0 0 0 mux8_6.NAND4F_9.D
flabel metal1 10993 -34727 11027 -34678 0 FreeSans 160 0 0 0 mux8_6.NAND4F_9.VSS
flabel nwell 11256 -36288 11290 -36239 0 FreeSans 160 0 0 0 mux8_6.NAND4F_9.VDD
flabel metal1 11689 -35608 11723 -35559 0 FreeSans 160 0 0 0 mux8_6.NAND4F_9.Y
rlabel metal1 12823 -34623 12823 -34623 3 mux8_6.inv_0.A
rlabel metal1 13021 -35012 13021 -35012 5 mux8_6.inv_0.VSS
rlabel metal1 13033 -34215 13033 -34215 5 mux8_6.inv_0.VDD
rlabel metal1 13235 -34623 13235 -34623 3 mux8_6.inv_0.Y
flabel metal1 11744 -34564 11821 -34512 1 FreeSerif 320 0 0 0 mux8_6.nor2_0.A
rlabel metal1 11990 -34064 11990 -34064 5 mux8_6.nor2_0.VDD
flabel metal1 11745 -34670 11822 -34618 1 FreeSerif 320 0 0 0 mux8_6.nor2_0.B
flabel metal1 12749 -34676 12826 -34624 1 FreeSerif 320 0 0 0 mux8_6.nor2_0.Y
rlabel metal1 12286 -35042 12286 -35042 5 mux8_6.nor2_0.VSS
rlabel metal1 5998 -32605 5998 -32605 3 mux8_6.inv_1.A
rlabel metal1 6196 -32994 6196 -32994 5 mux8_6.inv_1.VSS
rlabel metal1 6208 -32197 6208 -32197 5 mux8_6.inv_1.VDD
rlabel metal1 6410 -32605 6410 -32605 3 mux8_6.inv_1.Y
rlabel metal1 6438 -32605 6438 -32605 3 mux8_6.inv_2.A
rlabel metal1 6636 -32994 6636 -32994 5 mux8_6.inv_2.VSS
rlabel metal1 6648 -32197 6648 -32197 5 mux8_6.inv_2.VDD
rlabel metal1 6850 -32605 6850 -32605 3 mux8_6.inv_2.Y
rlabel metal1 5558 -32605 5558 -32605 3 mux8_6.inv_3.A
rlabel metal1 5756 -32994 5756 -32994 5 mux8_6.inv_3.VSS
rlabel metal1 5768 -32197 5768 -32197 5 mux8_6.inv_3.VDD
rlabel metal1 5970 -32605 5970 -32605 3 mux8_6.inv_3.Y
flabel space 9272 -19255 9338 -19189 0 FreeSans 1600 0 0 0 mux8_5.000
flabel space 10238 -19262 10245 -19260 0 FreeSans 1600 0 0 0 mux8_5.001
flabel space 7382 -19256 7385 -19256 0 FreeSans 1600 0 0 0 mux8_5.010
flabel space 8270 -19251 8594 -19192 0 FreeSans 1600 0 0 0 mux8_5.011
flabel space 9211 -22967 9637 -22910 0 FreeSans 1600 0 0 0 mux8_5.100
flabel space 10193 -22989 10471 -22830 0 FreeSans 1600 0 0 0 mux8_5.101
flabel space 7299 -23040 7617 -22865 0 FreeSans 1600 0 0 0 mux8_5.110
flabel space 8304 -23018 8622 -22843 0 FreeSans 1600 0 0 0 mux8_5.111
flabel metal2 5740 -20182 5792 -20130 0 FreeSans 160 0 0 0 mux8_5.A0
flabel metal2 5743 -20277 5795 -20225 0 FreeSans 160 0 0 0 mux8_5.A1
flabel metal2 5746 -20383 5798 -20331 0 FreeSans 160 0 0 0 mux8_5.A2
flabel metal2 5741 -20489 5793 -20437 0 FreeSans 160 0 0 0 mux8_5.A3
flabel metal2 5744 -21587 5796 -21535 0 FreeSans 160 0 0 0 mux8_5.A4
flabel metal2 5746 -21711 5798 -21659 0 FreeSans 160 0 0 0 mux8_5.A5
flabel metal2 5743 -21807 5795 -21755 0 FreeSans 160 0 0 0 mux8_5.A6
flabel metal2 5739 -21928 5791 -21876 0 FreeSans 160 0 0 0 mux8_5.A7
flabel metal1 12377 -19543 12429 -19491 0 FreeSans 160 0 0 0 mux8_5.VDD
flabel metal1 13159 -21183 13211 -21131 0 FreeSans 160 0 0 0 mux8_5.Y
flabel metal5 12955 -21830 13007 -21778 0 FreeSans 160 0 0 0 mux8_5.VSS
flabel metal2 6448 -18559 6493 -18520 0 FreeSans 160 0 0 0 mux8_5.SEL0
flabel metal2 6007 -18568 6052 -18529 0 FreeSans 160 0 0 0 mux8_5.SEL1
flabel metal2 5569 -18568 5614 -18529 0 FreeSans 160 0 0 0 mux8_5.SEL2
flabel metal1 8057 -20116 8091 -20067 0 FreeSans 160 0 0 0 mux8_5.NAND4F_2.A
flabel metal1 8060 -20016 8094 -19967 0 FreeSans 160 0 0 0 mux8_5.NAND4F_2.B
flabel metal1 8061 -19928 8095 -19879 0 FreeSans 160 0 0 0 mux8_5.NAND4F_2.C
flabel metal1 8062 -19835 8096 -19786 0 FreeSans 160 0 0 0 mux8_5.NAND4F_2.D
flabel metal1 8199 -20934 8233 -20885 0 FreeSans 160 0 0 0 mux8_5.NAND4F_2.VSS
flabel nwell 8462 -19373 8496 -19324 0 FreeSans 160 0 0 0 mux8_5.NAND4F_2.VDD
flabel metal1 8895 -20053 8929 -20004 0 FreeSans 160 0 0 0 mux8_5.NAND4F_2.Y
flabel metal1 7109 -20116 7143 -20067 0 FreeSans 160 0 0 0 mux8_5.NAND4F_4.A
flabel metal1 7112 -20016 7146 -19967 0 FreeSans 160 0 0 0 mux8_5.NAND4F_4.B
flabel metal1 7113 -19928 7147 -19879 0 FreeSans 160 0 0 0 mux8_5.NAND4F_4.C
flabel metal1 7114 -19835 7148 -19786 0 FreeSans 160 0 0 0 mux8_5.NAND4F_4.D
flabel metal1 7251 -20934 7285 -20885 0 FreeSans 160 0 0 0 mux8_5.NAND4F_4.VSS
flabel nwell 7514 -19373 7548 -19324 0 FreeSans 160 0 0 0 mux8_5.NAND4F_4.VDD
flabel metal1 7947 -20053 7981 -20004 0 FreeSans 160 0 0 0 mux8_5.NAND4F_4.Y
flabel metal1 7109 -21961 7143 -21912 0 FreeSans 160 0 0 0 mux8_5.NAND4F_5.A
flabel metal1 7112 -22061 7146 -22012 0 FreeSans 160 0 0 0 mux8_5.NAND4F_5.B
flabel metal1 7113 -22149 7147 -22100 0 FreeSans 160 0 0 0 mux8_5.NAND4F_5.C
flabel metal1 7114 -22242 7148 -22193 0 FreeSans 160 0 0 0 mux8_5.NAND4F_5.D
flabel metal1 7251 -21143 7285 -21094 0 FreeSans 160 0 0 0 mux8_5.NAND4F_5.VSS
flabel nwell 7514 -22704 7548 -22655 0 FreeSans 160 0 0 0 mux8_5.NAND4F_5.VDD
flabel metal1 7947 -22024 7981 -21975 0 FreeSans 160 0 0 0 mux8_5.NAND4F_5.Y
flabel metal1 8057 -21961 8091 -21912 0 FreeSans 160 0 0 0 mux8_5.NAND4F_6.A
flabel metal1 8060 -22061 8094 -22012 0 FreeSans 160 0 0 0 mux8_5.NAND4F_6.B
flabel metal1 8061 -22149 8095 -22100 0 FreeSans 160 0 0 0 mux8_5.NAND4F_6.C
flabel metal1 8062 -22242 8096 -22193 0 FreeSans 160 0 0 0 mux8_5.NAND4F_6.D
flabel metal1 8199 -21143 8233 -21094 0 FreeSans 160 0 0 0 mux8_5.NAND4F_6.VSS
flabel nwell 8462 -22704 8496 -22655 0 FreeSans 160 0 0 0 mux8_5.NAND4F_6.VDD
flabel metal1 8895 -22024 8929 -21975 0 FreeSans 160 0 0 0 mux8_5.NAND4F_6.Y
flabel metal1 9924 -20116 9958 -20067 0 FreeSans 160 0 0 0 mux8_5.NAND4F_0.A
flabel metal1 9927 -20016 9961 -19967 0 FreeSans 160 0 0 0 mux8_5.NAND4F_0.B
flabel metal1 9928 -19928 9962 -19879 0 FreeSans 160 0 0 0 mux8_5.NAND4F_0.C
flabel metal1 9929 -19835 9963 -19786 0 FreeSans 160 0 0 0 mux8_5.NAND4F_0.D
flabel metal1 10066 -20934 10100 -20885 0 FreeSans 160 0 0 0 mux8_5.NAND4F_0.VSS
flabel nwell 10329 -19373 10363 -19324 0 FreeSans 160 0 0 0 mux8_5.NAND4F_0.VDD
flabel metal1 10762 -20053 10796 -20004 0 FreeSans 160 0 0 0 mux8_5.NAND4F_0.Y
flabel metal1 8993 -21961 9027 -21912 0 FreeSans 160 0 0 0 mux8_5.NAND4F_1.A
flabel metal1 8996 -22061 9030 -22012 0 FreeSans 160 0 0 0 mux8_5.NAND4F_1.B
flabel metal1 8997 -22149 9031 -22100 0 FreeSans 160 0 0 0 mux8_5.NAND4F_1.C
flabel metal1 8998 -22242 9032 -22193 0 FreeSans 160 0 0 0 mux8_5.NAND4F_1.D
flabel metal1 9135 -21143 9169 -21094 0 FreeSans 160 0 0 0 mux8_5.NAND4F_1.VSS
flabel nwell 9398 -22704 9432 -22655 0 FreeSans 160 0 0 0 mux8_5.NAND4F_1.VDD
flabel metal1 9831 -22024 9865 -21975 0 FreeSans 160 0 0 0 mux8_5.NAND4F_1.Y
flabel metal1 8993 -20116 9027 -20067 0 FreeSans 160 0 0 0 mux8_5.NAND4F_3.A
flabel metal1 8996 -20016 9030 -19967 0 FreeSans 160 0 0 0 mux8_5.NAND4F_3.B
flabel metal1 8997 -19928 9031 -19879 0 FreeSans 160 0 0 0 mux8_5.NAND4F_3.C
flabel metal1 8998 -19835 9032 -19786 0 FreeSans 160 0 0 0 mux8_5.NAND4F_3.D
flabel metal1 9135 -20934 9169 -20885 0 FreeSans 160 0 0 0 mux8_5.NAND4F_3.VSS
flabel nwell 9398 -19373 9432 -19324 0 FreeSans 160 0 0 0 mux8_5.NAND4F_3.VDD
flabel metal1 9831 -20053 9865 -20004 0 FreeSans 160 0 0 0 mux8_5.NAND4F_3.Y
flabel metal1 9924 -21960 9958 -21911 0 FreeSans 160 0 0 0 mux8_5.NAND4F_7.A
flabel metal1 9927 -22060 9961 -22011 0 FreeSans 160 0 0 0 mux8_5.NAND4F_7.B
flabel metal1 9928 -22148 9962 -22099 0 FreeSans 160 0 0 0 mux8_5.NAND4F_7.C
flabel metal1 9929 -22241 9963 -22192 0 FreeSans 160 0 0 0 mux8_5.NAND4F_7.D
flabel metal1 10066 -21142 10100 -21093 0 FreeSans 160 0 0 0 mux8_5.NAND4F_7.VSS
flabel nwell 10329 -22703 10363 -22654 0 FreeSans 160 0 0 0 mux8_5.NAND4F_7.VDD
flabel metal1 10762 -22023 10796 -21974 0 FreeSans 160 0 0 0 mux8_5.NAND4F_7.Y
flabel metal1 10851 -20116 10885 -20067 0 FreeSans 160 0 0 0 mux8_5.NAND4F_8.A
flabel metal1 10854 -20016 10888 -19967 0 FreeSans 160 0 0 0 mux8_5.NAND4F_8.B
flabel metal1 10855 -19928 10889 -19879 0 FreeSans 160 0 0 0 mux8_5.NAND4F_8.C
flabel metal1 10856 -19835 10890 -19786 0 FreeSans 160 0 0 0 mux8_5.NAND4F_8.D
flabel metal1 10993 -20934 11027 -20885 0 FreeSans 160 0 0 0 mux8_5.NAND4F_8.VSS
flabel nwell 11256 -19373 11290 -19324 0 FreeSans 160 0 0 0 mux8_5.NAND4F_8.VDD
flabel metal1 11689 -20053 11723 -20004 0 FreeSans 160 0 0 0 mux8_5.NAND4F_8.Y
flabel metal1 10851 -21961 10885 -21912 0 FreeSans 160 0 0 0 mux8_5.NAND4F_9.A
flabel metal1 10854 -22061 10888 -22012 0 FreeSans 160 0 0 0 mux8_5.NAND4F_9.B
flabel metal1 10855 -22149 10889 -22100 0 FreeSans 160 0 0 0 mux8_5.NAND4F_9.C
flabel metal1 10856 -22242 10890 -22193 0 FreeSans 160 0 0 0 mux8_5.NAND4F_9.D
flabel metal1 10993 -21143 11027 -21094 0 FreeSans 160 0 0 0 mux8_5.NAND4F_9.VSS
flabel nwell 11256 -22704 11290 -22655 0 FreeSans 160 0 0 0 mux8_5.NAND4F_9.VDD
flabel metal1 11689 -22024 11723 -21975 0 FreeSans 160 0 0 0 mux8_5.NAND4F_9.Y
rlabel metal1 12823 -21039 12823 -21039 3 mux8_5.inv_0.A
rlabel metal1 13021 -21428 13021 -21428 5 mux8_5.inv_0.VSS
rlabel metal1 13033 -20631 13033 -20631 5 mux8_5.inv_0.VDD
rlabel metal1 13235 -21039 13235 -21039 3 mux8_5.inv_0.Y
flabel metal1 11744 -20980 11821 -20928 1 FreeSerif 320 0 0 0 mux8_5.nor2_0.A
rlabel metal1 11990 -20480 11990 -20480 5 mux8_5.nor2_0.VDD
flabel metal1 11745 -21086 11822 -21034 1 FreeSerif 320 0 0 0 mux8_5.nor2_0.B
flabel metal1 12749 -21092 12826 -21040 1 FreeSerif 320 0 0 0 mux8_5.nor2_0.Y
rlabel metal1 12286 -21458 12286 -21458 5 mux8_5.nor2_0.VSS
rlabel metal1 5998 -19021 5998 -19021 3 mux8_5.inv_1.A
rlabel metal1 6196 -19410 6196 -19410 5 mux8_5.inv_1.VSS
rlabel metal1 6208 -18613 6208 -18613 5 mux8_5.inv_1.VDD
rlabel metal1 6410 -19021 6410 -19021 3 mux8_5.inv_1.Y
rlabel metal1 6438 -19021 6438 -19021 3 mux8_5.inv_2.A
rlabel metal1 6636 -19410 6636 -19410 5 mux8_5.inv_2.VSS
rlabel metal1 6648 -18613 6648 -18613 5 mux8_5.inv_2.VDD
rlabel metal1 6850 -19021 6850 -19021 3 mux8_5.inv_2.Y
rlabel metal1 5558 -19021 5558 -19021 3 mux8_5.inv_3.A
rlabel metal1 5756 -19410 5756 -19410 5 mux8_5.inv_3.VSS
rlabel metal1 5768 -18613 5768 -18613 5 mux8_5.inv_3.VDD
rlabel metal1 5970 -19021 5970 -19021 3 mux8_5.inv_3.Y
flabel space 9272 -14727 9338 -14661 0 FreeSans 1600 0 0 0 mux8_4.000
flabel space 10238 -14734 10245 -14732 0 FreeSans 1600 0 0 0 mux8_4.001
flabel space 7382 -14728 7385 -14728 0 FreeSans 1600 0 0 0 mux8_4.010
flabel space 8270 -14723 8594 -14664 0 FreeSans 1600 0 0 0 mux8_4.011
flabel space 9211 -18439 9637 -18382 0 FreeSans 1600 0 0 0 mux8_4.100
flabel space 10193 -18461 10471 -18302 0 FreeSans 1600 0 0 0 mux8_4.101
flabel space 7299 -18512 7617 -18337 0 FreeSans 1600 0 0 0 mux8_4.110
flabel space 8304 -18490 8622 -18315 0 FreeSans 1600 0 0 0 mux8_4.111
flabel metal2 5740 -15654 5792 -15602 0 FreeSans 160 0 0 0 mux8_4.A0
flabel metal2 5743 -15749 5795 -15697 0 FreeSans 160 0 0 0 mux8_4.A1
flabel metal2 5746 -15855 5798 -15803 0 FreeSans 160 0 0 0 mux8_4.A2
flabel metal2 5741 -15961 5793 -15909 0 FreeSans 160 0 0 0 mux8_4.A3
flabel metal2 5744 -17059 5796 -17007 0 FreeSans 160 0 0 0 mux8_4.A4
flabel metal2 5746 -17183 5798 -17131 0 FreeSans 160 0 0 0 mux8_4.A5
flabel metal2 5743 -17279 5795 -17227 0 FreeSans 160 0 0 0 mux8_4.A6
flabel metal2 5739 -17400 5791 -17348 0 FreeSans 160 0 0 0 mux8_4.A7
flabel metal1 12377 -15015 12429 -14963 0 FreeSans 160 0 0 0 mux8_4.VDD
flabel metal1 13159 -16655 13211 -16603 0 FreeSans 160 0 0 0 mux8_4.Y
flabel metal5 12955 -17302 13007 -17250 0 FreeSans 160 0 0 0 mux8_4.VSS
flabel metal2 6448 -14031 6493 -13992 0 FreeSans 160 0 0 0 mux8_4.SEL0
flabel metal2 6007 -14040 6052 -14001 0 FreeSans 160 0 0 0 mux8_4.SEL1
flabel metal2 5569 -14040 5614 -14001 0 FreeSans 160 0 0 0 mux8_4.SEL2
flabel metal1 8057 -15588 8091 -15539 0 FreeSans 160 0 0 0 mux8_4.NAND4F_2.A
flabel metal1 8060 -15488 8094 -15439 0 FreeSans 160 0 0 0 mux8_4.NAND4F_2.B
flabel metal1 8061 -15400 8095 -15351 0 FreeSans 160 0 0 0 mux8_4.NAND4F_2.C
flabel metal1 8062 -15307 8096 -15258 0 FreeSans 160 0 0 0 mux8_4.NAND4F_2.D
flabel metal1 8199 -16406 8233 -16357 0 FreeSans 160 0 0 0 mux8_4.NAND4F_2.VSS
flabel nwell 8462 -14845 8496 -14796 0 FreeSans 160 0 0 0 mux8_4.NAND4F_2.VDD
flabel metal1 8895 -15525 8929 -15476 0 FreeSans 160 0 0 0 mux8_4.NAND4F_2.Y
flabel metal1 7109 -15588 7143 -15539 0 FreeSans 160 0 0 0 mux8_4.NAND4F_4.A
flabel metal1 7112 -15488 7146 -15439 0 FreeSans 160 0 0 0 mux8_4.NAND4F_4.B
flabel metal1 7113 -15400 7147 -15351 0 FreeSans 160 0 0 0 mux8_4.NAND4F_4.C
flabel metal1 7114 -15307 7148 -15258 0 FreeSans 160 0 0 0 mux8_4.NAND4F_4.D
flabel metal1 7251 -16406 7285 -16357 0 FreeSans 160 0 0 0 mux8_4.NAND4F_4.VSS
flabel nwell 7514 -14845 7548 -14796 0 FreeSans 160 0 0 0 mux8_4.NAND4F_4.VDD
flabel metal1 7947 -15525 7981 -15476 0 FreeSans 160 0 0 0 mux8_4.NAND4F_4.Y
flabel metal1 7109 -17433 7143 -17384 0 FreeSans 160 0 0 0 mux8_4.NAND4F_5.A
flabel metal1 7112 -17533 7146 -17484 0 FreeSans 160 0 0 0 mux8_4.NAND4F_5.B
flabel metal1 7113 -17621 7147 -17572 0 FreeSans 160 0 0 0 mux8_4.NAND4F_5.C
flabel metal1 7114 -17714 7148 -17665 0 FreeSans 160 0 0 0 mux8_4.NAND4F_5.D
flabel metal1 7251 -16615 7285 -16566 0 FreeSans 160 0 0 0 mux8_4.NAND4F_5.VSS
flabel nwell 7514 -18176 7548 -18127 0 FreeSans 160 0 0 0 mux8_4.NAND4F_5.VDD
flabel metal1 7947 -17496 7981 -17447 0 FreeSans 160 0 0 0 mux8_4.NAND4F_5.Y
flabel metal1 8057 -17433 8091 -17384 0 FreeSans 160 0 0 0 mux8_4.NAND4F_6.A
flabel metal1 8060 -17533 8094 -17484 0 FreeSans 160 0 0 0 mux8_4.NAND4F_6.B
flabel metal1 8061 -17621 8095 -17572 0 FreeSans 160 0 0 0 mux8_4.NAND4F_6.C
flabel metal1 8062 -17714 8096 -17665 0 FreeSans 160 0 0 0 mux8_4.NAND4F_6.D
flabel metal1 8199 -16615 8233 -16566 0 FreeSans 160 0 0 0 mux8_4.NAND4F_6.VSS
flabel nwell 8462 -18176 8496 -18127 0 FreeSans 160 0 0 0 mux8_4.NAND4F_6.VDD
flabel metal1 8895 -17496 8929 -17447 0 FreeSans 160 0 0 0 mux8_4.NAND4F_6.Y
flabel metal1 9924 -15588 9958 -15539 0 FreeSans 160 0 0 0 mux8_4.NAND4F_0.A
flabel metal1 9927 -15488 9961 -15439 0 FreeSans 160 0 0 0 mux8_4.NAND4F_0.B
flabel metal1 9928 -15400 9962 -15351 0 FreeSans 160 0 0 0 mux8_4.NAND4F_0.C
flabel metal1 9929 -15307 9963 -15258 0 FreeSans 160 0 0 0 mux8_4.NAND4F_0.D
flabel metal1 10066 -16406 10100 -16357 0 FreeSans 160 0 0 0 mux8_4.NAND4F_0.VSS
flabel nwell 10329 -14845 10363 -14796 0 FreeSans 160 0 0 0 mux8_4.NAND4F_0.VDD
flabel metal1 10762 -15525 10796 -15476 0 FreeSans 160 0 0 0 mux8_4.NAND4F_0.Y
flabel metal1 8993 -17433 9027 -17384 0 FreeSans 160 0 0 0 mux8_4.NAND4F_1.A
flabel metal1 8996 -17533 9030 -17484 0 FreeSans 160 0 0 0 mux8_4.NAND4F_1.B
flabel metal1 8997 -17621 9031 -17572 0 FreeSans 160 0 0 0 mux8_4.NAND4F_1.C
flabel metal1 8998 -17714 9032 -17665 0 FreeSans 160 0 0 0 mux8_4.NAND4F_1.D
flabel metal1 9135 -16615 9169 -16566 0 FreeSans 160 0 0 0 mux8_4.NAND4F_1.VSS
flabel nwell 9398 -18176 9432 -18127 0 FreeSans 160 0 0 0 mux8_4.NAND4F_1.VDD
flabel metal1 9831 -17496 9865 -17447 0 FreeSans 160 0 0 0 mux8_4.NAND4F_1.Y
flabel metal1 8993 -15588 9027 -15539 0 FreeSans 160 0 0 0 mux8_4.NAND4F_3.A
flabel metal1 8996 -15488 9030 -15439 0 FreeSans 160 0 0 0 mux8_4.NAND4F_3.B
flabel metal1 8997 -15400 9031 -15351 0 FreeSans 160 0 0 0 mux8_4.NAND4F_3.C
flabel metal1 8998 -15307 9032 -15258 0 FreeSans 160 0 0 0 mux8_4.NAND4F_3.D
flabel metal1 9135 -16406 9169 -16357 0 FreeSans 160 0 0 0 mux8_4.NAND4F_3.VSS
flabel nwell 9398 -14845 9432 -14796 0 FreeSans 160 0 0 0 mux8_4.NAND4F_3.VDD
flabel metal1 9831 -15525 9865 -15476 0 FreeSans 160 0 0 0 mux8_4.NAND4F_3.Y
flabel metal1 9924 -17432 9958 -17383 0 FreeSans 160 0 0 0 mux8_4.NAND4F_7.A
flabel metal1 9927 -17532 9961 -17483 0 FreeSans 160 0 0 0 mux8_4.NAND4F_7.B
flabel metal1 9928 -17620 9962 -17571 0 FreeSans 160 0 0 0 mux8_4.NAND4F_7.C
flabel metal1 9929 -17713 9963 -17664 0 FreeSans 160 0 0 0 mux8_4.NAND4F_7.D
flabel metal1 10066 -16614 10100 -16565 0 FreeSans 160 0 0 0 mux8_4.NAND4F_7.VSS
flabel nwell 10329 -18175 10363 -18126 0 FreeSans 160 0 0 0 mux8_4.NAND4F_7.VDD
flabel metal1 10762 -17495 10796 -17446 0 FreeSans 160 0 0 0 mux8_4.NAND4F_7.Y
flabel metal1 10851 -15588 10885 -15539 0 FreeSans 160 0 0 0 mux8_4.NAND4F_8.A
flabel metal1 10854 -15488 10888 -15439 0 FreeSans 160 0 0 0 mux8_4.NAND4F_8.B
flabel metal1 10855 -15400 10889 -15351 0 FreeSans 160 0 0 0 mux8_4.NAND4F_8.C
flabel metal1 10856 -15307 10890 -15258 0 FreeSans 160 0 0 0 mux8_4.NAND4F_8.D
flabel metal1 10993 -16406 11027 -16357 0 FreeSans 160 0 0 0 mux8_4.NAND4F_8.VSS
flabel nwell 11256 -14845 11290 -14796 0 FreeSans 160 0 0 0 mux8_4.NAND4F_8.VDD
flabel metal1 11689 -15525 11723 -15476 0 FreeSans 160 0 0 0 mux8_4.NAND4F_8.Y
flabel metal1 10851 -17433 10885 -17384 0 FreeSans 160 0 0 0 mux8_4.NAND4F_9.A
flabel metal1 10854 -17533 10888 -17484 0 FreeSans 160 0 0 0 mux8_4.NAND4F_9.B
flabel metal1 10855 -17621 10889 -17572 0 FreeSans 160 0 0 0 mux8_4.NAND4F_9.C
flabel metal1 10856 -17714 10890 -17665 0 FreeSans 160 0 0 0 mux8_4.NAND4F_9.D
flabel metal1 10993 -16615 11027 -16566 0 FreeSans 160 0 0 0 mux8_4.NAND4F_9.VSS
flabel nwell 11256 -18176 11290 -18127 0 FreeSans 160 0 0 0 mux8_4.NAND4F_9.VDD
flabel metal1 11689 -17496 11723 -17447 0 FreeSans 160 0 0 0 mux8_4.NAND4F_9.Y
rlabel metal1 12823 -16511 12823 -16511 3 mux8_4.inv_0.A
rlabel metal1 13021 -16900 13021 -16900 5 mux8_4.inv_0.VSS
rlabel metal1 13033 -16103 13033 -16103 5 mux8_4.inv_0.VDD
rlabel metal1 13235 -16511 13235 -16511 3 mux8_4.inv_0.Y
flabel metal1 11744 -16452 11821 -16400 1 FreeSerif 320 0 0 0 mux8_4.nor2_0.A
rlabel metal1 11990 -15952 11990 -15952 5 mux8_4.nor2_0.VDD
flabel metal1 11745 -16558 11822 -16506 1 FreeSerif 320 0 0 0 mux8_4.nor2_0.B
flabel metal1 12749 -16564 12826 -16512 1 FreeSerif 320 0 0 0 mux8_4.nor2_0.Y
rlabel metal1 12286 -16930 12286 -16930 5 mux8_4.nor2_0.VSS
rlabel metal1 5998 -14493 5998 -14493 3 mux8_4.inv_1.A
rlabel metal1 6196 -14882 6196 -14882 5 mux8_4.inv_1.VSS
rlabel metal1 6208 -14085 6208 -14085 5 mux8_4.inv_1.VDD
rlabel metal1 6410 -14493 6410 -14493 3 mux8_4.inv_1.Y
rlabel metal1 6438 -14493 6438 -14493 3 mux8_4.inv_2.A
rlabel metal1 6636 -14882 6636 -14882 5 mux8_4.inv_2.VSS
rlabel metal1 6648 -14085 6648 -14085 5 mux8_4.inv_2.VDD
rlabel metal1 6850 -14493 6850 -14493 3 mux8_4.inv_2.Y
rlabel metal1 5558 -14493 5558 -14493 3 mux8_4.inv_3.A
rlabel metal1 5756 -14882 5756 -14882 5 mux8_4.inv_3.VSS
rlabel metal1 5768 -14085 5768 -14085 5 mux8_4.inv_3.VDD
rlabel metal1 5970 -14493 5970 -14493 3 mux8_4.inv_3.Y
rlabel metal1 13169 -35615 13169 -35615 5 buffer_0.A
rlabel metal1 12777 -36053 12777 -36053 7 buffer_0.VSS
rlabel metal1 13184 -36406 13184 -36406 5 buffer_0.Y
rlabel metal1 13574 -36066 13574 -36066 7 buffer_0.VDD
rlabel metal1 13166 -35994 13166 -35994 5 buffer_0.inv_1.A
rlabel metal1 12777 -36192 12777 -36192 7 buffer_0.inv_1.VSS
rlabel metal1 13574 -36204 13574 -36204 7 buffer_0.inv_1.VDD
rlabel metal1 13166 -36406 13166 -36406 5 buffer_0.inv_1.Y
rlabel metal1 13166 -35615 13166 -35615 5 buffer_0.inv_0.A
rlabel metal1 12777 -35813 12777 -35813 7 buffer_0.inv_0.VSS
rlabel metal1 13574 -35825 13574 -35825 7 buffer_0.inv_0.VDD
rlabel metal1 13166 -36027 13166 -36027 5 buffer_0.inv_0.Y
flabel metal1 15629 -17342 15641 -17306 0 FreeSans 160 0 0 0 ZFLAG_0.A0
flabel metal1 15631 -17434 15643 -17398 0 FreeSans 160 0 0 0 ZFLAG_0.A1
flabel metal1 15631 -17528 15643 -17492 0 FreeSans 160 0 0 0 ZFLAG_0.A2
flabel metal1 15631 -17624 15643 -17588 0 FreeSans 160 0 0 0 ZFLAG_0.A3
flabel metal1 15625 -19588 15649 -19548 0 FreeSans 160 0 0 0 ZFLAG_0.A4
flabel metal1 15631 -19684 15655 -19644 0 FreeSans 160 0 0 0 ZFLAG_0.A5
flabel metal1 15629 -19780 15653 -19740 0 FreeSans 160 0 0 0 ZFLAG_0.A6
flabel metal1 15629 -19872 15653 -19832 0 FreeSans 160 0 0 0 ZFLAG_0.A7
flabel metal4 15639 -18642 15683 -18532 0 FreeSans 160 0 0 0 ZFLAG_0.VDD
flabel metal1 18357 -18653 18397 -18531 0 FreeSans 160 0 0 0 ZFLAG_0.Z
rlabel metal5 17042 -20468 17448 -20227 5 ZFLAG_0.VSS
rlabel metal1 15617 -19571 15617 -19571 3 ZFLAG_0.nor4_1.A
rlabel metal1 15617 -19663 15617 -19663 3 ZFLAG_0.nor4_1.B
rlabel metal1 15617 -19759 15617 -19759 3 ZFLAG_0.nor4_1.C
rlabel metal1 15617 -19854 15617 -19854 3 ZFLAG_0.nor4_1.D
rlabel metal1 16377 -20365 16377 -20365 5 ZFLAG_0.nor4_1.VSS
rlabel metal1 15688 -19317 15688 -19317 5 ZFLAG_0.nor4_1.VDD
rlabel metal1 17009 -19570 17009 -19570 3 ZFLAG_0.nor4_1.Y
rlabel metal1 15617 -17601 15617 -17601 3 ZFLAG_0.nor4_0.A
rlabel metal1 15617 -17509 15617 -17509 3 ZFLAG_0.nor4_0.B
rlabel metal1 15617 -17413 15617 -17413 3 ZFLAG_0.nor4_0.C
rlabel metal1 15617 -17318 15617 -17318 3 ZFLAG_0.nor4_0.D
rlabel metal1 16377 -16807 16377 -16807 1 ZFLAG_0.nor4_0.VSS
rlabel metal1 15688 -17855 15688 -17855 1 ZFLAG_0.nor4_0.VDD
rlabel metal1 17009 -17602 17009 -17602 3 ZFLAG_0.nor4_0.Y
rlabel metal1 17258 -18582 17258 -18582 7 ZFLAG_0.NAND2_0.A
rlabel metal1 17258 -18750 17258 -18750 7 ZFLAG_0.NAND2_0.B
rlabel metal1 17728 -18869 17728 -18869 5 ZFLAG_0.NAND2_0.VSS
rlabel metal1 17611 -18239 17611 -18239 1 ZFLAG_0.NAND2_0.VDD
rlabel metal1 17964 -18472 17964 -18472 3 ZFLAG_0.NAND2_0.Y
rlabel metal1 17996 -18551 17996 -18551 3 ZFLAG_0.inv_0.A
rlabel metal1 18194 -18940 18194 -18940 5 ZFLAG_0.inv_0.VSS
rlabel metal1 18206 -18143 18206 -18143 5 ZFLAG_0.inv_0.VDD
rlabel metal1 18408 -18551 18408 -18551 3 ZFLAG_0.inv_0.Y
rlabel metal4 -15250 4413 -14951 4623 5 8bit_ADDER_0.VDD
rlabel metal5 -11927 4574 -11848 4674 5 8bit_ADDER_0.VSS
rlabel metal1 -24905 1129 -24853 1190 5 8bit_ADDER_0.C
flabel metal2 -21805 200 -21730 282 0 FreeSans 160 0 0 0 8bit_ADDER_0.S7
flabel metal2 -18510 203 -18435 285 0 FreeSans 160 0 0 0 8bit_ADDER_0.S6
flabel metal2 -15222 206 -15147 288 0 FreeSans 160 0 0 0 8bit_ADDER_0.S5
flabel metal2 -11935 207 -11860 289 0 FreeSans 160 0 0 0 8bit_ADDER_0.S4
flabel metal2 -8633 204 -8558 286 0 FreeSans 160 0 0 0 8bit_ADDER_0.S3
flabel metal2 -5355 203 -5280 285 0 FreeSans 160 0 0 0 8bit_ADDER_0.S2
flabel metal2 -2056 213 -1981 295 0 FreeSans 160 0 0 0 8bit_ADDER_0.S1
flabel metal2 1234 207 1309 289 0 FreeSans 160 0 0 0 8bit_ADDER_0.S0
flabel metal1 -25107 4474 -25012 4540 0 FreeSans 160 0 0 0 8bit_ADDER_0.A7
flabel metal1 -21816 4468 -21721 4534 0 FreeSans 160 0 0 0 8bit_ADDER_0.A6
flabel metal1 -18526 4476 -18431 4542 0 FreeSans 160 0 0 0 8bit_ADDER_0.A5
flabel metal1 -15233 4478 -15138 4544 0 FreeSans 160 0 0 0 8bit_ADDER_0.A4
flabel metal1 -11943 4476 -11848 4542 0 FreeSans 160 0 0 0 8bit_ADDER_0.A3
flabel metal1 -8651 4470 -8556 4536 0 FreeSans 160 0 0 0 8bit_ADDER_0.A2
flabel metal1 -5360 4474 -5265 4540 0 FreeSans 160 0 0 0 8bit_ADDER_0.A1
flabel metal1 -2071 4480 -1976 4546 0 FreeSans 160 0 0 0 8bit_ADDER_0.A0
flabel metal1 -22626 4457 -22531 4523 0 FreeSans 160 0 0 0 8bit_ADDER_0.B7
flabel metal1 -19340 4451 -19245 4517 0 FreeSans 160 0 0 0 8bit_ADDER_0.B6
flabel metal1 -16041 4455 -15946 4521 0 FreeSans 160 0 0 0 8bit_ADDER_0.B5
flabel metal1 -12755 4448 -12660 4514 0 FreeSans 160 0 0 0 8bit_ADDER_0.B4
flabel metal1 -9450 4453 -9355 4519 0 FreeSans 160 0 0 0 8bit_ADDER_0.B3
flabel metal1 -6174 4466 -6079 4532 0 FreeSans 160 0 0 0 8bit_ADDER_0.B2
flabel metal1 -2875 4472 -2780 4538 0 FreeSans 160 0 0 0 8bit_ADDER_0.B1
flabel metal1 397 4462 492 4528 0 FreeSans 160 0 0 0 8bit_ADDER_0.B0
rlabel metal2 602 4379 774 4550 5 8bit_ADDER_0.K
rlabel metal2 -2054 3916 -2000 3988 5 8bit_ADDER_0.FULL_ADDER_XORED_7.A
rlabel metal1 426 4442 490 4544 5 8bit_ADDER_0.FULL_ADDER_XORED_7.B
rlabel metal1 670 4428 734 4530 5 8bit_ADDER_0.FULL_ADDER_XORED_7.K
rlabel metal1 -1866 1126 -1830 1196 5 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT
rlabel metal2 1228 212 1308 292 5 8bit_ADDER_0.FULL_ADDER_XORED_7.OUT
rlabel metal1 1022 1134 1172 1178 5 8bit_ADDER_0.FULL_ADDER_XORED_7.CIN
rlabel metal4 -571 4442 -170 4519 5 8bit_ADDER_0.FULL_ADDER_XORED_7.VDD
rlabel metal5 -1353 -43 -952 34 5 8bit_ADDER_0.FULL_ADDER_XORED_7.VSS
rlabel poly 289 3555 313 3595 3 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.A
rlabel metal1 311 3411 335 3451 3 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.B
rlabel via1 -291 4467 -197 4493 5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.VDD
rlabel metal1 -1107 3439 -1055 3517 5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y
rlabel metal1 -221 3079 -127 3105 5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.VSS
rlabel poly -230 1771 -206 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A
rlabel metal1 -252 1627 -228 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.B
rlabel via1 280 2683 374 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.VDD
rlabel metal1 1138 1655 1190 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.Y
rlabel metal1 210 1295 304 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.VSS
rlabel poly -1789 1771 -1765 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_0.A
rlabel metal1 -1811 1627 -1787 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_0.B
rlabel via1 -1279 2683 -1185 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_0.VDD
rlabel metal1 -421 1655 -369 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_0.Y
rlabel metal1 -1349 1295 -1255 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_0.VSS
rlabel metal1 394 568 394 568 7 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A
rlabel metal1 394 400 394 400 7 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B
rlabel metal1 864 281 864 281 5 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.VSS
rlabel metal1 747 911 747 911 1 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.VDD
rlabel metal1 1100 678 1100 678 3 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.Y
rlabel metal1 -488 568 -488 568 7 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_1.A
rlabel metal1 -488 400 -488 400 7 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_1.B
rlabel metal1 -18 281 -18 281 5 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_1.VSS
rlabel metal1 -135 911 -135 911 1 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_1.VDD
rlabel metal1 218 678 218 678 3 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_1.Y
rlabel metal1 -1597 568 -1597 568 7 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_0.A
rlabel metal1 -1597 400 -1597 400 7 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_0.B
rlabel metal1 -1127 281 -1127 281 5 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_0.VSS
rlabel metal1 -1244 911 -1244 911 1 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_0.VDD
rlabel metal1 -891 678 -891 678 3 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_0.Y
rlabel metal2 -5345 3916 -5291 3988 5 8bit_ADDER_0.FULL_ADDER_XORED_6.A
rlabel metal1 -2865 4442 -2801 4544 5 8bit_ADDER_0.FULL_ADDER_XORED_6.B
rlabel metal1 -2621 4428 -2557 4530 5 8bit_ADDER_0.FULL_ADDER_XORED_6.K
rlabel metal1 -5157 1126 -5121 1196 5 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT
rlabel metal2 -2063 212 -1983 292 5 8bit_ADDER_0.FULL_ADDER_XORED_6.OUT
rlabel metal1 -2269 1134 -2119 1178 5 8bit_ADDER_0.FULL_ADDER_XORED_6.CIN
rlabel metal4 -3862 4442 -3461 4519 5 8bit_ADDER_0.FULL_ADDER_XORED_6.VDD
rlabel metal5 -4644 -43 -4243 34 5 8bit_ADDER_0.FULL_ADDER_XORED_6.VSS
rlabel poly -3002 3555 -2978 3595 3 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.A
rlabel metal1 -2980 3411 -2956 3451 3 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.B
rlabel via1 -3582 4467 -3488 4493 5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.VDD
rlabel metal1 -4398 3439 -4346 3517 5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y
rlabel metal1 -3512 3079 -3418 3105 5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.VSS
rlabel poly -3521 1771 -3497 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A
rlabel metal1 -3543 1627 -3519 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.B
rlabel via1 -3011 2683 -2917 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.VDD
rlabel metal1 -2153 1655 -2101 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.Y
rlabel metal1 -3081 1295 -2987 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.VSS
rlabel poly -5080 1771 -5056 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_0.A
rlabel metal1 -5102 1627 -5078 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_0.B
rlabel via1 -4570 2683 -4476 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_0.VDD
rlabel metal1 -3712 1655 -3660 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_0.Y
rlabel metal1 -4640 1295 -4546 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_0.VSS
rlabel metal1 -2897 568 -2897 568 7 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A
rlabel metal1 -2897 400 -2897 400 7 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B
rlabel metal1 -2427 281 -2427 281 5 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.VSS
rlabel metal1 -2544 911 -2544 911 1 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.VDD
rlabel metal1 -2191 678 -2191 678 3 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.Y
rlabel metal1 -3779 568 -3779 568 7 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_1.A
rlabel metal1 -3779 400 -3779 400 7 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_1.B
rlabel metal1 -3309 281 -3309 281 5 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_1.VSS
rlabel metal1 -3426 911 -3426 911 1 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_1.VDD
rlabel metal1 -3073 678 -3073 678 3 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_1.Y
rlabel metal1 -4888 568 -4888 568 7 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_0.A
rlabel metal1 -4888 400 -4888 400 7 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_0.B
rlabel metal1 -4418 281 -4418 281 5 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_0.VSS
rlabel metal1 -4535 911 -4535 911 1 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_0.VDD
rlabel metal1 -4182 678 -4182 678 3 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_0.Y
rlabel metal2 -8636 3916 -8582 3988 5 8bit_ADDER_0.FULL_ADDER_XORED_5.A
rlabel metal1 -6156 4442 -6092 4544 5 8bit_ADDER_0.FULL_ADDER_XORED_5.B
rlabel metal1 -5912 4428 -5848 4530 5 8bit_ADDER_0.FULL_ADDER_XORED_5.K
rlabel metal1 -8448 1126 -8412 1196 5 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT
rlabel metal2 -5354 212 -5274 292 5 8bit_ADDER_0.FULL_ADDER_XORED_5.OUT
rlabel metal1 -5560 1134 -5410 1178 5 8bit_ADDER_0.FULL_ADDER_XORED_5.CIN
rlabel metal4 -7153 4442 -6752 4519 5 8bit_ADDER_0.FULL_ADDER_XORED_5.VDD
rlabel metal5 -7935 -43 -7534 34 5 8bit_ADDER_0.FULL_ADDER_XORED_5.VSS
rlabel poly -6293 3555 -6269 3595 3 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.A
rlabel metal1 -6271 3411 -6247 3451 3 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.B
rlabel via1 -6873 4467 -6779 4493 5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.VDD
rlabel metal1 -7689 3439 -7637 3517 5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y
rlabel metal1 -6803 3079 -6709 3105 5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.VSS
rlabel poly -6812 1771 -6788 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A
rlabel metal1 -6834 1627 -6810 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.B
rlabel via1 -6302 2683 -6208 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.VDD
rlabel metal1 -5444 1655 -5392 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.Y
rlabel metal1 -6372 1295 -6278 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.VSS
rlabel poly -8371 1771 -8347 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_0.A
rlabel metal1 -8393 1627 -8369 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_0.B
rlabel via1 -7861 2683 -7767 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_0.VDD
rlabel metal1 -7003 1655 -6951 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_0.Y
rlabel metal1 -7931 1295 -7837 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_0.VSS
rlabel metal1 -6188 568 -6188 568 7 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A
rlabel metal1 -6188 400 -6188 400 7 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B
rlabel metal1 -5718 281 -5718 281 5 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.VSS
rlabel metal1 -5835 911 -5835 911 1 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.VDD
rlabel metal1 -5482 678 -5482 678 3 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.Y
rlabel metal1 -7070 568 -7070 568 7 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_1.A
rlabel metal1 -7070 400 -7070 400 7 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_1.B
rlabel metal1 -6600 281 -6600 281 5 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_1.VSS
rlabel metal1 -6717 911 -6717 911 1 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_1.VDD
rlabel metal1 -6364 678 -6364 678 3 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_1.Y
rlabel metal1 -8179 568 -8179 568 7 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_0.A
rlabel metal1 -8179 400 -8179 400 7 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_0.B
rlabel metal1 -7709 281 -7709 281 5 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_0.VSS
rlabel metal1 -7826 911 -7826 911 1 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_0.VDD
rlabel metal1 -7473 678 -7473 678 3 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_0.Y
rlabel metal2 -11926 3916 -11872 3988 5 8bit_ADDER_0.FULL_ADDER_XORED_4.A
rlabel metal1 -9446 4442 -9382 4544 5 8bit_ADDER_0.FULL_ADDER_XORED_4.B
rlabel metal1 -9202 4428 -9138 4530 5 8bit_ADDER_0.FULL_ADDER_XORED_4.K
rlabel metal1 -11738 1126 -11702 1196 5 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT
rlabel metal2 -8644 212 -8564 292 5 8bit_ADDER_0.FULL_ADDER_XORED_4.OUT
rlabel metal1 -8850 1134 -8700 1178 5 8bit_ADDER_0.FULL_ADDER_XORED_4.CIN
rlabel metal4 -10443 4442 -10042 4519 5 8bit_ADDER_0.FULL_ADDER_XORED_4.VDD
rlabel metal5 -11225 -43 -10824 34 5 8bit_ADDER_0.FULL_ADDER_XORED_4.VSS
rlabel poly -9583 3555 -9559 3595 3 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.A
rlabel metal1 -9561 3411 -9537 3451 3 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.B
rlabel via1 -10163 4467 -10069 4493 5 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.VDD
rlabel metal1 -10979 3439 -10927 3517 5 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y
rlabel metal1 -10093 3079 -9999 3105 5 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.VSS
rlabel poly -10102 1771 -10078 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A
rlabel metal1 -10124 1627 -10100 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.B
rlabel via1 -9592 2683 -9498 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.VDD
rlabel metal1 -8734 1655 -8682 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.Y
rlabel metal1 -9662 1295 -9568 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.VSS
rlabel poly -11661 1771 -11637 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_0.A
rlabel metal1 -11683 1627 -11659 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_0.B
rlabel via1 -11151 2683 -11057 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_0.VDD
rlabel metal1 -10293 1655 -10241 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_0.Y
rlabel metal1 -11221 1295 -11127 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_0.VSS
rlabel metal1 -9478 568 -9478 568 7 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A
rlabel metal1 -9478 400 -9478 400 7 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B
rlabel metal1 -9008 281 -9008 281 5 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.VSS
rlabel metal1 -9125 911 -9125 911 1 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.VDD
rlabel metal1 -8772 678 -8772 678 3 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.Y
rlabel metal1 -10360 568 -10360 568 7 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_1.A
rlabel metal1 -10360 400 -10360 400 7 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_1.B
rlabel metal1 -9890 281 -9890 281 5 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_1.VSS
rlabel metal1 -10007 911 -10007 911 1 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_1.VDD
rlabel metal1 -9654 678 -9654 678 3 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_1.Y
rlabel metal1 -11469 568 -11469 568 7 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_0.A
rlabel metal1 -11469 400 -11469 400 7 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_0.B
rlabel metal1 -10999 281 -10999 281 5 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_0.VSS
rlabel metal1 -11116 911 -11116 911 1 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_0.VDD
rlabel metal1 -10763 678 -10763 678 3 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_0.Y
rlabel metal2 -15217 3916 -15163 3988 5 8bit_ADDER_0.FULL_ADDER_XORED_3.A
rlabel metal1 -12737 4442 -12673 4544 5 8bit_ADDER_0.FULL_ADDER_XORED_3.B
rlabel metal1 -12493 4428 -12429 4530 5 8bit_ADDER_0.FULL_ADDER_XORED_3.K
rlabel metal1 -15029 1126 -14993 1196 5 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT
rlabel metal2 -11935 212 -11855 292 5 8bit_ADDER_0.FULL_ADDER_XORED_3.OUT
rlabel metal1 -12141 1134 -11991 1178 5 8bit_ADDER_0.FULL_ADDER_XORED_3.CIN
rlabel metal4 -13734 4442 -13333 4519 5 8bit_ADDER_0.FULL_ADDER_XORED_3.VDD
rlabel metal5 -14516 -43 -14115 34 5 8bit_ADDER_0.FULL_ADDER_XORED_3.VSS
rlabel poly -12874 3555 -12850 3595 3 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.A
rlabel metal1 -12852 3411 -12828 3451 3 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.B
rlabel via1 -13454 4467 -13360 4493 5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.VDD
rlabel metal1 -14270 3439 -14218 3517 5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y
rlabel metal1 -13384 3079 -13290 3105 5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.VSS
rlabel poly -13393 1771 -13369 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A
rlabel metal1 -13415 1627 -13391 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.B
rlabel via1 -12883 2683 -12789 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.VDD
rlabel metal1 -12025 1655 -11973 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.Y
rlabel metal1 -12953 1295 -12859 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.VSS
rlabel poly -14952 1771 -14928 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_0.A
rlabel metal1 -14974 1627 -14950 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_0.B
rlabel via1 -14442 2683 -14348 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_0.VDD
rlabel metal1 -13584 1655 -13532 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_0.Y
rlabel metal1 -14512 1295 -14418 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_0.VSS
rlabel metal1 -12769 568 -12769 568 7 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A
rlabel metal1 -12769 400 -12769 400 7 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B
rlabel metal1 -12299 281 -12299 281 5 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.VSS
rlabel metal1 -12416 911 -12416 911 1 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.VDD
rlabel metal1 -12063 678 -12063 678 3 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.Y
rlabel metal1 -13651 568 -13651 568 7 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_1.A
rlabel metal1 -13651 400 -13651 400 7 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_1.B
rlabel metal1 -13181 281 -13181 281 5 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_1.VSS
rlabel metal1 -13298 911 -13298 911 1 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_1.VDD
rlabel metal1 -12945 678 -12945 678 3 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_1.Y
rlabel metal1 -14760 568 -14760 568 7 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_0.A
rlabel metal1 -14760 400 -14760 400 7 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_0.B
rlabel metal1 -14290 281 -14290 281 5 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_0.VSS
rlabel metal1 -14407 911 -14407 911 1 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_0.VDD
rlabel metal1 -14054 678 -14054 678 3 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_0.Y
rlabel metal2 -18508 3916 -18454 3988 5 8bit_ADDER_0.FULL_ADDER_XORED_2.A
rlabel metal1 -16028 4442 -15964 4544 5 8bit_ADDER_0.FULL_ADDER_XORED_2.B
rlabel metal1 -15784 4428 -15720 4530 5 8bit_ADDER_0.FULL_ADDER_XORED_2.K
rlabel metal1 -18320 1126 -18284 1196 5 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT
rlabel metal2 -15226 212 -15146 292 5 8bit_ADDER_0.FULL_ADDER_XORED_2.OUT
rlabel metal1 -15432 1134 -15282 1178 5 8bit_ADDER_0.FULL_ADDER_XORED_2.CIN
rlabel metal4 -17025 4442 -16624 4519 5 8bit_ADDER_0.FULL_ADDER_XORED_2.VDD
rlabel metal5 -17807 -43 -17406 34 5 8bit_ADDER_0.FULL_ADDER_XORED_2.VSS
rlabel poly -16165 3555 -16141 3595 3 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.A
rlabel metal1 -16143 3411 -16119 3451 3 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.B
rlabel via1 -16745 4467 -16651 4493 5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.VDD
rlabel metal1 -17561 3439 -17509 3517 5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y
rlabel metal1 -16675 3079 -16581 3105 5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.VSS
rlabel poly -16684 1771 -16660 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A
rlabel metal1 -16706 1627 -16682 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.B
rlabel via1 -16174 2683 -16080 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.VDD
rlabel metal1 -15316 1655 -15264 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.Y
rlabel metal1 -16244 1295 -16150 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.VSS
rlabel poly -18243 1771 -18219 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_0.A
rlabel metal1 -18265 1627 -18241 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_0.B
rlabel via1 -17733 2683 -17639 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_0.VDD
rlabel metal1 -16875 1655 -16823 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_0.Y
rlabel metal1 -17803 1295 -17709 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_0.VSS
rlabel metal1 -16060 568 -16060 568 7 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A
rlabel metal1 -16060 400 -16060 400 7 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B
rlabel metal1 -15590 281 -15590 281 5 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.VSS
rlabel metal1 -15707 911 -15707 911 1 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.VDD
rlabel metal1 -15354 678 -15354 678 3 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.Y
rlabel metal1 -16942 568 -16942 568 7 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_1.A
rlabel metal1 -16942 400 -16942 400 7 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_1.B
rlabel metal1 -16472 281 -16472 281 5 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_1.VSS
rlabel metal1 -16589 911 -16589 911 1 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_1.VDD
rlabel metal1 -16236 678 -16236 678 3 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_1.Y
rlabel metal1 -18051 568 -18051 568 7 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_0.A
rlabel metal1 -18051 400 -18051 400 7 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_0.B
rlabel metal1 -17581 281 -17581 281 5 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_0.VSS
rlabel metal1 -17698 911 -17698 911 1 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_0.VDD
rlabel metal1 -17345 678 -17345 678 3 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_0.Y
rlabel metal2 -21799 3916 -21745 3988 5 8bit_ADDER_0.FULL_ADDER_XORED_1.A
rlabel metal1 -19319 4442 -19255 4544 5 8bit_ADDER_0.FULL_ADDER_XORED_1.B
rlabel metal1 -19075 4428 -19011 4530 5 8bit_ADDER_0.FULL_ADDER_XORED_1.K
rlabel metal1 -21611 1126 -21575 1196 5 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT
rlabel metal2 -18517 212 -18437 292 5 8bit_ADDER_0.FULL_ADDER_XORED_1.OUT
rlabel metal1 -18723 1134 -18573 1178 5 8bit_ADDER_0.FULL_ADDER_XORED_1.CIN
rlabel metal4 -20316 4442 -19915 4519 5 8bit_ADDER_0.FULL_ADDER_XORED_1.VDD
rlabel metal5 -21098 -43 -20697 34 5 8bit_ADDER_0.FULL_ADDER_XORED_1.VSS
rlabel poly -19456 3555 -19432 3595 3 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.A
rlabel metal1 -19434 3411 -19410 3451 3 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.B
rlabel via1 -20036 4467 -19942 4493 5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.VDD
rlabel metal1 -20852 3439 -20800 3517 5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y
rlabel metal1 -19966 3079 -19872 3105 5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.VSS
rlabel poly -19975 1771 -19951 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A
rlabel metal1 -19997 1627 -19973 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.B
rlabel via1 -19465 2683 -19371 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.VDD
rlabel metal1 -18607 1655 -18555 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.Y
rlabel metal1 -19535 1295 -19441 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.VSS
rlabel poly -21534 1771 -21510 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_0.A
rlabel metal1 -21556 1627 -21532 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_0.B
rlabel via1 -21024 2683 -20930 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_0.VDD
rlabel metal1 -20166 1655 -20114 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_0.Y
rlabel metal1 -21094 1295 -21000 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_0.VSS
rlabel metal1 -19351 568 -19351 568 7 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A
rlabel metal1 -19351 400 -19351 400 7 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B
rlabel metal1 -18881 281 -18881 281 5 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.VSS
rlabel metal1 -18998 911 -18998 911 1 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.VDD
rlabel metal1 -18645 678 -18645 678 3 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.Y
rlabel metal1 -20233 568 -20233 568 7 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_1.A
rlabel metal1 -20233 400 -20233 400 7 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_1.B
rlabel metal1 -19763 281 -19763 281 5 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_1.VSS
rlabel metal1 -19880 911 -19880 911 1 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_1.VDD
rlabel metal1 -19527 678 -19527 678 3 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_1.Y
rlabel metal1 -21342 568 -21342 568 7 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_0.A
rlabel metal1 -21342 400 -21342 400 7 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_0.B
rlabel metal1 -20872 281 -20872 281 5 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_0.VSS
rlabel metal1 -20989 911 -20989 911 1 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_0.VDD
rlabel metal1 -20636 678 -20636 678 3 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_0.Y
rlabel metal2 -25090 3916 -25036 3988 5 8bit_ADDER_0.FULL_ADDER_XORED_0.A
rlabel metal1 -22610 4442 -22546 4544 5 8bit_ADDER_0.FULL_ADDER_XORED_0.B
rlabel metal1 -22366 4428 -22302 4530 5 8bit_ADDER_0.FULL_ADDER_XORED_0.K
rlabel metal1 -24902 1126 -24866 1196 5 8bit_ADDER_0.FULL_ADDER_XORED_0.COUT
rlabel metal2 -21808 212 -21728 292 5 8bit_ADDER_0.FULL_ADDER_XORED_0.OUT
rlabel metal1 -22014 1134 -21864 1178 5 8bit_ADDER_0.FULL_ADDER_XORED_0.CIN
rlabel metal4 -23607 4442 -23206 4519 5 8bit_ADDER_0.FULL_ADDER_XORED_0.VDD
rlabel metal5 -24389 -43 -23988 34 5 8bit_ADDER_0.FULL_ADDER_XORED_0.VSS
rlabel poly -22747 3555 -22723 3595 3 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.A
rlabel metal1 -22725 3411 -22701 3451 3 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.B
rlabel via1 -23327 4467 -23233 4493 5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.VDD
rlabel metal1 -24143 3439 -24091 3517 5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y
rlabel metal1 -23257 3079 -23163 3105 5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.VSS
rlabel poly -23266 1771 -23242 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A
rlabel metal1 -23288 1627 -23264 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.B
rlabel via1 -22756 2683 -22662 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.VDD
rlabel metal1 -21898 1655 -21846 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.Y
rlabel metal1 -22826 1295 -22732 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.VSS
rlabel poly -24825 1771 -24801 1811 7 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_0.A
rlabel metal1 -24847 1627 -24823 1667 7 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_0.B
rlabel via1 -24315 2683 -24221 2709 5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_0.VDD
rlabel metal1 -23457 1655 -23405 1733 5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_0.Y
rlabel metal1 -24385 1295 -24291 1321 5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_0.VSS
rlabel metal1 -22642 568 -22642 568 7 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A
rlabel metal1 -22642 400 -22642 400 7 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B
rlabel metal1 -22172 281 -22172 281 5 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.VSS
rlabel metal1 -22289 911 -22289 911 1 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.VDD
rlabel metal1 -21936 678 -21936 678 3 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.Y
rlabel metal1 -23524 568 -23524 568 7 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_1.A
rlabel metal1 -23524 400 -23524 400 7 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_1.B
rlabel metal1 -23054 281 -23054 281 5 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_1.VSS
rlabel metal1 -23171 911 -23171 911 1 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_1.VDD
rlabel metal1 -22818 678 -22818 678 3 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_1.Y
rlabel metal1 -24633 568 -24633 568 7 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_0.A
rlabel metal1 -24633 400 -24633 400 7 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_0.B
rlabel metal1 -24163 281 -24163 281 5 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_0.VSS
rlabel metal1 -24280 911 -24280 911 1 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_0.VDD
rlabel metal1 -23927 678 -23927 678 3 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_0.Y
flabel metal2 -24272 -8421 -24152 -8301 1 FreeSerif 160 0 0 0 MULT_0.B2
flabel metal2 -24264 -11683 -24144 -11563 1 FreeSerif 160 0 0 0 MULT_0.B3
flabel metal2 -23996 -6807 -23876 -6687 1 FreeSerif 160 0 0 0 MULT_0.A1
flabel metal2 -8224 -3177 -8104 -3057 1 FreeSerif 160 0 0 0 MULT_0.SO
flabel metal3 -23190 -6433 -23070 -6313 1 FreeSerif 160 0 0 0 MULT_0.A2
flabel metal1 -24838 -4585 -24718 -4465 1 FreeSerif 160 0 0 0 MULT_0.A0
flabel metal3 -24234 -3553 -24114 -3433 1 FreeSerif 160 0 0 0 MULT_0.A3
flabel metal2 -24628 -2345 -24508 -2225 1 FreeSerif 160 0 0 0 MULT_0.B0
flabel metal2 -20990 -12959 -20894 -12873 1 FreeSerif 160 0 0 0 MULT_0.S7
flabel metal2 -7862 -12895 -7766 -12809 1 FreeSerif 160 0 0 0 MULT_0.S3
flabel metal2 -11166 -12901 -11070 -12815 1 FreeSerif 160 0 0 0 MULT_0.S4
flabel metal2 -14458 -12899 -14362 -12813 1 FreeSerif 160 0 0 0 MULT_0.S5
flabel metal2 -7862 -9625 -7766 -9539 1 FreeSerif 160 0 0 0 MULT_0.S2
flabel metal2 -7878 -6263 -7782 -6177 1 FreeSerif 160 0 0 0 MULT_0.S1
flabel metal2 -17750 -12895 -17654 -12809 1 FreeSerif 160 0 0 0 MULT_0.S6
flabel metal5 -15068 -13179 -12970 -11583 0 FreeSans 160 0 0 0 MULT_0.VSS
flabel metal4 -14354 -3907 -14222 -3813 0 FreeSans 160 0 0 0 MULT_0.VDD
flabel metal2 -24606 -5123 -24492 -5005 0 FreeSans 160 0 0 0 MULT_0.B1
rlabel metal1 -22695 -12353 -22695 -12353 7 MULT_0.NAND2_15.A
rlabel metal1 -22695 -12521 -22695 -12521 7 MULT_0.NAND2_15.B
rlabel metal1 -22225 -12640 -22225 -12640 5 MULT_0.NAND2_15.VSS
rlabel metal1 -22342 -12010 -22342 -12010 1 MULT_0.NAND2_15.VDD
rlabel metal1 -21989 -12243 -21989 -12243 3 MULT_0.NAND2_15.Y
rlabel metal1 -24432 -12353 -24432 -12353 7 MULT_0.NAND2_9.A
rlabel metal1 -24432 -12521 -24432 -12521 7 MULT_0.NAND2_9.B
rlabel metal1 -23962 -12640 -23962 -12640 5 MULT_0.NAND2_9.VSS
rlabel metal1 -24079 -12010 -24079 -12010 1 MULT_0.NAND2_9.VDD
rlabel metal1 -23726 -12243 -23726 -12243 3 MULT_0.NAND2_9.Y
rlabel metal1 -21954 -12244 -21954 -12244 3 MULT_0.inv_15.A
rlabel metal1 -21756 -12633 -21756 -12633 5 MULT_0.inv_15.VSS
rlabel metal1 -21744 -11836 -21744 -11836 5 MULT_0.inv_15.VDD
rlabel metal1 -21542 -12244 -21542 -12244 3 MULT_0.inv_15.Y
rlabel metal1 -23683 -12244 -23683 -12244 3 MULT_0.inv_9.A
rlabel metal1 -23485 -12633 -23485 -12633 5 MULT_0.inv_9.VSS
rlabel metal1 -23473 -11836 -23473 -11836 5 MULT_0.inv_9.VDD
rlabel metal1 -23271 -12244 -23271 -12244 3 MULT_0.inv_9.Y
rlabel metal1 -22695 -11061 -22695 -11061 7 MULT_0.NAND2_14.A
rlabel metal1 -22695 -11229 -22695 -11229 7 MULT_0.NAND2_14.B
rlabel metal1 -22225 -11348 -22225 -11348 5 MULT_0.NAND2_14.VSS
rlabel metal1 -22342 -10718 -22342 -10718 1 MULT_0.NAND2_14.VDD
rlabel metal1 -21989 -10951 -21989 -10951 3 MULT_0.NAND2_14.Y
rlabel metal1 -24432 -11061 -24432 -11061 7 MULT_0.NAND2_8.A
rlabel metal1 -24432 -11229 -24432 -11229 7 MULT_0.NAND2_8.B
rlabel metal1 -23962 -11348 -23962 -11348 5 MULT_0.NAND2_8.VSS
rlabel metal1 -24079 -10718 -24079 -10718 1 MULT_0.NAND2_8.VDD
rlabel metal1 -23726 -10951 -23726 -10951 3 MULT_0.NAND2_8.Y
rlabel metal1 -21950 -10952 -21950 -10952 3 MULT_0.inv_14.A
rlabel metal1 -21752 -11341 -21752 -11341 5 MULT_0.inv_14.VSS
rlabel metal1 -21740 -10544 -21740 -10544 5 MULT_0.inv_14.VDD
rlabel metal1 -21538 -10952 -21538 -10952 3 MULT_0.inv_14.Y
rlabel metal1 -23683 -10952 -23683 -10952 3 MULT_0.inv_8.A
rlabel metal1 -23485 -11341 -23485 -11341 5 MULT_0.inv_8.VSS
rlabel metal1 -23473 -10544 -23473 -10544 5 MULT_0.inv_8.VDD
rlabel metal1 -23271 -10952 -23271 -10952 3 MULT_0.inv_8.Y
flabel metal2 -21031 -10351 -20961 -10291 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.A3
flabel metal2 -17735 -10371 -17665 -10311 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.A2
flabel metal2 -14447 -10373 -14377 -10313 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.A1
flabel metal2 -11155 -10357 -11085 -10297 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.A0
flabel metal2 -10977 -10357 -10907 -10297 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.B0
flabel metal2 -14267 -10373 -14197 -10313 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.B1
flabel metal2 -17561 -10371 -17491 -10311 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.B2
flabel metal2 -20847 -10351 -20777 -10291 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.B3
flabel metal1 -7765 -11959 -7693 -11889 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.C
flabel metal2 -7865 -12881 -7793 -12811 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.S0
flabel metal2 -11159 -12877 -11081 -12797 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.S1
flabel metal2 -14451 -12877 -14373 -12797 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.S2
flabel metal2 -17741 -12877 -17663 -12797 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.S3
flabel metal2 -21025 -13025 -20887 -12913 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.Cout
flabel metal5 -15355 -13199 -15217 -13087 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.VSS
flabel metal4 -15387 -10443 -15249 -10331 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_2.VDD
rlabel metal1 -10962 -11963 -10926 -11893 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT
rlabel metal2 -7868 -12877 -7788 -12797 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.OUT
rlabel metal1 -8074 -11955 -7924 -11911 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.CIN
rlabel metal5 -10449 -13132 -10048 -13055 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.VSS
rlabel metal2 -11161 -10341 -11081 -10282 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.A
rlabel metal2 -10984 -10341 -10904 -10282 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.B
rlabel metal4 -9527 -10428 -9272 -10326 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.VDD
rlabel poly -9326 -11318 -9302 -11278 7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A
rlabel metal1 -9348 -11462 -9324 -11422 7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.B
rlabel via1 -8816 -10406 -8722 -10380 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.VDD
rlabel metal1 -7958 -11434 -7906 -11356 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.Y
rlabel metal1 -8886 -11794 -8792 -11768 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.VSS
rlabel poly -10885 -11318 -10861 -11278 7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_0.A
rlabel metal1 -10907 -11462 -10883 -11422 7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_0.B
rlabel via1 -10375 -10406 -10281 -10380 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_0.VDD
rlabel metal1 -9517 -11434 -9465 -11356 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_0.Y
rlabel metal1 -10445 -11794 -10351 -11768 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_0.VSS
rlabel metal1 -8702 -12521 -8702 -12521 7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A
rlabel metal1 -8702 -12689 -8702 -12689 7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B
rlabel metal1 -8232 -12808 -8232 -12808 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.VSS
rlabel metal1 -8349 -12178 -8349 -12178 1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.VDD
rlabel metal1 -7996 -12411 -7996 -12411 3 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.Y
rlabel metal1 -9584 -12521 -9584 -12521 7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_1.A
rlabel metal1 -9584 -12689 -9584 -12689 7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_1.B
rlabel metal1 -9114 -12808 -9114 -12808 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_1.VSS
rlabel metal1 -9231 -12178 -9231 -12178 1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_1.VDD
rlabel metal1 -8878 -12411 -8878 -12411 3 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_1.Y
rlabel metal1 -10693 -12521 -10693 -12521 7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_0.A
rlabel metal1 -10693 -12689 -10693 -12689 7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_0.B
rlabel metal1 -10223 -12808 -10223 -12808 5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_0.VSS
rlabel metal1 -10340 -12178 -10340 -12178 1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_0.VDD
rlabel metal1 -9987 -12411 -9987 -12411 3 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_0.Y
rlabel metal1 -14253 -11963 -14217 -11893 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT
rlabel metal2 -11159 -12877 -11079 -12797 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.OUT
rlabel metal1 -11365 -11955 -11215 -11911 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.CIN
rlabel metal5 -13740 -13132 -13339 -13055 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.VSS
rlabel metal2 -14452 -10341 -14372 -10282 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.A
rlabel metal2 -14275 -10341 -14195 -10282 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.B
rlabel metal4 -12818 -10428 -12563 -10326 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.VDD
rlabel poly -12617 -11318 -12593 -11278 7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A
rlabel metal1 -12639 -11462 -12615 -11422 7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.B
rlabel via1 -12107 -10406 -12013 -10380 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.VDD
rlabel metal1 -11249 -11434 -11197 -11356 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.Y
rlabel metal1 -12177 -11794 -12083 -11768 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.VSS
rlabel poly -14176 -11318 -14152 -11278 7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_0.A
rlabel metal1 -14198 -11462 -14174 -11422 7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_0.B
rlabel via1 -13666 -10406 -13572 -10380 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_0.VDD
rlabel metal1 -12808 -11434 -12756 -11356 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_0.Y
rlabel metal1 -13736 -11794 -13642 -11768 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_0.VSS
rlabel metal1 -11993 -12521 -11993 -12521 7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A
rlabel metal1 -11993 -12689 -11993 -12689 7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B
rlabel metal1 -11523 -12808 -11523 -12808 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.VSS
rlabel metal1 -11640 -12178 -11640 -12178 1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.VDD
rlabel metal1 -11287 -12411 -11287 -12411 3 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.Y
rlabel metal1 -12875 -12521 -12875 -12521 7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_1.A
rlabel metal1 -12875 -12689 -12875 -12689 7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_1.B
rlabel metal1 -12405 -12808 -12405 -12808 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_1.VSS
rlabel metal1 -12522 -12178 -12522 -12178 1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_1.VDD
rlabel metal1 -12169 -12411 -12169 -12411 3 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_1.Y
rlabel metal1 -13984 -12521 -13984 -12521 7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_0.A
rlabel metal1 -13984 -12689 -13984 -12689 7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_0.B
rlabel metal1 -13514 -12808 -13514 -12808 5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_0.VSS
rlabel metal1 -13631 -12178 -13631 -12178 1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_0.VDD
rlabel metal1 -13278 -12411 -13278 -12411 3 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_0.Y
rlabel metal1 -17544 -11963 -17508 -11893 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT
rlabel metal2 -14450 -12877 -14370 -12797 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.OUT
rlabel metal1 -14656 -11955 -14506 -11911 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.CIN
rlabel metal5 -17031 -13132 -16630 -13055 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.VSS
rlabel metal2 -17743 -10341 -17663 -10282 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.A
rlabel metal2 -17566 -10341 -17486 -10282 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.B
rlabel metal4 -16109 -10428 -15854 -10326 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.VDD
rlabel poly -15908 -11318 -15884 -11278 7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A
rlabel metal1 -15930 -11462 -15906 -11422 7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.B
rlabel via1 -15398 -10406 -15304 -10380 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.VDD
rlabel metal1 -14540 -11434 -14488 -11356 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.Y
rlabel metal1 -15468 -11794 -15374 -11768 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.VSS
rlabel poly -17467 -11318 -17443 -11278 7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_0.A
rlabel metal1 -17489 -11462 -17465 -11422 7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_0.B
rlabel via1 -16957 -10406 -16863 -10380 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_0.VDD
rlabel metal1 -16099 -11434 -16047 -11356 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_0.Y
rlabel metal1 -17027 -11794 -16933 -11768 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_0.VSS
rlabel metal1 -15284 -12521 -15284 -12521 7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A
rlabel metal1 -15284 -12689 -15284 -12689 7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B
rlabel metal1 -14814 -12808 -14814 -12808 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.VSS
rlabel metal1 -14931 -12178 -14931 -12178 1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.VDD
rlabel metal1 -14578 -12411 -14578 -12411 3 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.Y
rlabel metal1 -16166 -12521 -16166 -12521 7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_1.A
rlabel metal1 -16166 -12689 -16166 -12689 7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_1.B
rlabel metal1 -15696 -12808 -15696 -12808 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_1.VSS
rlabel metal1 -15813 -12178 -15813 -12178 1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_1.VDD
rlabel metal1 -15460 -12411 -15460 -12411 3 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_1.Y
rlabel metal1 -17275 -12521 -17275 -12521 7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_0.A
rlabel metal1 -17275 -12689 -17275 -12689 7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_0.B
rlabel metal1 -16805 -12808 -16805 -12808 5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_0.VSS
rlabel metal1 -16922 -12178 -16922 -12178 1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_0.VDD
rlabel metal1 -16569 -12411 -16569 -12411 3 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_0.Y
rlabel metal1 -20835 -11963 -20799 -11893 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.COUT
rlabel metal2 -17741 -12877 -17661 -12797 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.OUT
rlabel metal1 -17947 -11955 -17797 -11911 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.CIN
rlabel metal5 -20322 -13132 -19921 -13055 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.VSS
rlabel metal2 -21034 -10341 -20954 -10282 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.A
rlabel metal2 -20857 -10341 -20777 -10282 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.B
rlabel metal4 -19400 -10428 -19145 -10326 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.VDD
rlabel poly -19199 -11318 -19175 -11278 7 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A
rlabel metal1 -19221 -11462 -19197 -11422 7 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.B
rlabel via1 -18689 -10406 -18595 -10380 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.VDD
rlabel metal1 -17831 -11434 -17779 -11356 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.Y
rlabel metal1 -18759 -11794 -18665 -11768 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.VSS
rlabel poly -20758 -11318 -20734 -11278 7 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_0.A
rlabel metal1 -20780 -11462 -20756 -11422 7 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_0.B
rlabel via1 -20248 -10406 -20154 -10380 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_0.VDD
rlabel metal1 -19390 -11434 -19338 -11356 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_0.Y
rlabel metal1 -20318 -11794 -20224 -11768 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_0.VSS
rlabel metal1 -18575 -12521 -18575 -12521 7 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A
rlabel metal1 -18575 -12689 -18575 -12689 7 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B
rlabel metal1 -18105 -12808 -18105 -12808 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.VSS
rlabel metal1 -18222 -12178 -18222 -12178 1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.VDD
rlabel metal1 -17869 -12411 -17869 -12411 3 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.Y
rlabel metal1 -19457 -12521 -19457 -12521 7 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_1.A
rlabel metal1 -19457 -12689 -19457 -12689 7 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_1.B
rlabel metal1 -18987 -12808 -18987 -12808 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_1.VSS
rlabel metal1 -19104 -12178 -19104 -12178 1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_1.VDD
rlabel metal1 -18751 -12411 -18751 -12411 3 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_1.Y
rlabel metal1 -20566 -12521 -20566 -12521 7 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_0.A
rlabel metal1 -20566 -12689 -20566 -12689 7 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_0.B
rlabel metal1 -20096 -12808 -20096 -12808 5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_0.VSS
rlabel metal1 -20213 -12178 -20213 -12178 1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_0.VDD
rlabel metal1 -19860 -12411 -19860 -12411 3 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_0.Y
flabel metal2 -21031 -7087 -20961 -7027 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.A3
flabel metal2 -17735 -7107 -17665 -7047 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.A2
flabel metal2 -14447 -7109 -14377 -7049 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.A1
flabel metal2 -11155 -7093 -11085 -7033 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.A0
flabel metal2 -10977 -7093 -10907 -7033 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.B0
flabel metal2 -14267 -7109 -14197 -7049 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.B1
flabel metal2 -17561 -7107 -17491 -7047 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.B2
flabel metal2 -20847 -7087 -20777 -7027 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.B3
flabel metal1 -7765 -8695 -7693 -8625 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.C
flabel metal2 -7865 -9617 -7793 -9547 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.S0
flabel metal2 -11159 -9613 -11081 -9533 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.S1
flabel metal2 -14451 -9613 -14373 -9533 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.S2
flabel metal2 -17741 -9613 -17663 -9533 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.S3
flabel metal2 -21025 -9761 -20887 -9649 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.Cout
flabel metal5 -15355 -9935 -15217 -9823 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.VSS
flabel metal4 -15387 -7179 -15249 -7067 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_1.VDD
rlabel metal1 -10962 -8699 -10926 -8629 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT
rlabel metal2 -7868 -9613 -7788 -9533 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.OUT
rlabel metal1 -8074 -8691 -7924 -8647 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.CIN
rlabel metal5 -10449 -9868 -10048 -9791 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.VSS
rlabel metal2 -11161 -7077 -11081 -7018 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.A
rlabel metal2 -10984 -7077 -10904 -7018 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.B
rlabel metal4 -9527 -7164 -9272 -7062 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.VDD
rlabel poly -9326 -8054 -9302 -8014 7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A
rlabel metal1 -9348 -8198 -9324 -8158 7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.B
rlabel via1 -8816 -7142 -8722 -7116 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.VDD
rlabel metal1 -7958 -8170 -7906 -8092 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.Y
rlabel metal1 -8886 -8530 -8792 -8504 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.VSS
rlabel poly -10885 -8054 -10861 -8014 7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_0.A
rlabel metal1 -10907 -8198 -10883 -8158 7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_0.B
rlabel via1 -10375 -7142 -10281 -7116 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_0.VDD
rlabel metal1 -9517 -8170 -9465 -8092 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_0.Y
rlabel metal1 -10445 -8530 -10351 -8504 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_0.VSS
rlabel metal1 -8702 -9257 -8702 -9257 7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A
rlabel metal1 -8702 -9425 -8702 -9425 7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B
rlabel metal1 -8232 -9544 -8232 -9544 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.VSS
rlabel metal1 -8349 -8914 -8349 -8914 1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.VDD
rlabel metal1 -7996 -9147 -7996 -9147 3 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.Y
rlabel metal1 -9584 -9257 -9584 -9257 7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_1.A
rlabel metal1 -9584 -9425 -9584 -9425 7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_1.B
rlabel metal1 -9114 -9544 -9114 -9544 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_1.VSS
rlabel metal1 -9231 -8914 -9231 -8914 1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_1.VDD
rlabel metal1 -8878 -9147 -8878 -9147 3 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_1.Y
rlabel metal1 -10693 -9257 -10693 -9257 7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_0.A
rlabel metal1 -10693 -9425 -10693 -9425 7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_0.B
rlabel metal1 -10223 -9544 -10223 -9544 5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_0.VSS
rlabel metal1 -10340 -8914 -10340 -8914 1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_0.VDD
rlabel metal1 -9987 -9147 -9987 -9147 3 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_0.Y
rlabel metal1 -14253 -8699 -14217 -8629 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT
rlabel metal2 -11159 -9613 -11079 -9533 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.OUT
rlabel metal1 -11365 -8691 -11215 -8647 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.CIN
rlabel metal5 -13740 -9868 -13339 -9791 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.VSS
rlabel metal2 -14452 -7077 -14372 -7018 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.A
rlabel metal2 -14275 -7077 -14195 -7018 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.B
rlabel metal4 -12818 -7164 -12563 -7062 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.VDD
rlabel poly -12617 -8054 -12593 -8014 7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A
rlabel metal1 -12639 -8198 -12615 -8158 7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.B
rlabel via1 -12107 -7142 -12013 -7116 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.VDD
rlabel metal1 -11249 -8170 -11197 -8092 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.Y
rlabel metal1 -12177 -8530 -12083 -8504 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.VSS
rlabel poly -14176 -8054 -14152 -8014 7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_0.A
rlabel metal1 -14198 -8198 -14174 -8158 7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_0.B
rlabel via1 -13666 -7142 -13572 -7116 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_0.VDD
rlabel metal1 -12808 -8170 -12756 -8092 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_0.Y
rlabel metal1 -13736 -8530 -13642 -8504 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_0.VSS
rlabel metal1 -11993 -9257 -11993 -9257 7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A
rlabel metal1 -11993 -9425 -11993 -9425 7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B
rlabel metal1 -11523 -9544 -11523 -9544 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.VSS
rlabel metal1 -11640 -8914 -11640 -8914 1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.VDD
rlabel metal1 -11287 -9147 -11287 -9147 3 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.Y
rlabel metal1 -12875 -9257 -12875 -9257 7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_1.A
rlabel metal1 -12875 -9425 -12875 -9425 7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_1.B
rlabel metal1 -12405 -9544 -12405 -9544 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_1.VSS
rlabel metal1 -12522 -8914 -12522 -8914 1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_1.VDD
rlabel metal1 -12169 -9147 -12169 -9147 3 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_1.Y
rlabel metal1 -13984 -9257 -13984 -9257 7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_0.A
rlabel metal1 -13984 -9425 -13984 -9425 7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_0.B
rlabel metal1 -13514 -9544 -13514 -9544 5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_0.VSS
rlabel metal1 -13631 -8914 -13631 -8914 1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_0.VDD
rlabel metal1 -13278 -9147 -13278 -9147 3 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_0.Y
rlabel metal1 -17544 -8699 -17508 -8629 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT
rlabel metal2 -14450 -9613 -14370 -9533 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.OUT
rlabel metal1 -14656 -8691 -14506 -8647 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.CIN
rlabel metal5 -17031 -9868 -16630 -9791 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.VSS
rlabel metal2 -17743 -7077 -17663 -7018 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.A
rlabel metal2 -17566 -7077 -17486 -7018 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.B
rlabel metal4 -16109 -7164 -15854 -7062 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.VDD
rlabel poly -15908 -8054 -15884 -8014 7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A
rlabel metal1 -15930 -8198 -15906 -8158 7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.B
rlabel via1 -15398 -7142 -15304 -7116 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.VDD
rlabel metal1 -14540 -8170 -14488 -8092 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.Y
rlabel metal1 -15468 -8530 -15374 -8504 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.VSS
rlabel poly -17467 -8054 -17443 -8014 7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_0.A
rlabel metal1 -17489 -8198 -17465 -8158 7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_0.B
rlabel via1 -16957 -7142 -16863 -7116 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_0.VDD
rlabel metal1 -16099 -8170 -16047 -8092 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_0.Y
rlabel metal1 -17027 -8530 -16933 -8504 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_0.VSS
rlabel metal1 -15284 -9257 -15284 -9257 7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A
rlabel metal1 -15284 -9425 -15284 -9425 7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B
rlabel metal1 -14814 -9544 -14814 -9544 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.VSS
rlabel metal1 -14931 -8914 -14931 -8914 1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.VDD
rlabel metal1 -14578 -9147 -14578 -9147 3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.Y
rlabel metal1 -16166 -9257 -16166 -9257 7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_1.A
rlabel metal1 -16166 -9425 -16166 -9425 7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_1.B
rlabel metal1 -15696 -9544 -15696 -9544 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_1.VSS
rlabel metal1 -15813 -8914 -15813 -8914 1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_1.VDD
rlabel metal1 -15460 -9147 -15460 -9147 3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_1.Y
rlabel metal1 -17275 -9257 -17275 -9257 7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_0.A
rlabel metal1 -17275 -9425 -17275 -9425 7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_0.B
rlabel metal1 -16805 -9544 -16805 -9544 5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_0.VSS
rlabel metal1 -16922 -8914 -16922 -8914 1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_0.VDD
rlabel metal1 -16569 -9147 -16569 -9147 3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_0.Y
rlabel metal1 -20835 -8699 -20799 -8629 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.COUT
rlabel metal2 -17741 -9613 -17661 -9533 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.OUT
rlabel metal1 -17947 -8691 -17797 -8647 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.CIN
rlabel metal5 -20322 -9868 -19921 -9791 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.VSS
rlabel metal2 -21034 -7077 -20954 -7018 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.A
rlabel metal2 -20857 -7077 -20777 -7018 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.B
rlabel metal4 -19400 -7164 -19145 -7062 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.VDD
rlabel poly -19199 -8054 -19175 -8014 7 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A
rlabel metal1 -19221 -8198 -19197 -8158 7 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.B
rlabel via1 -18689 -7142 -18595 -7116 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.VDD
rlabel metal1 -17831 -8170 -17779 -8092 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.Y
rlabel metal1 -18759 -8530 -18665 -8504 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.VSS
rlabel poly -20758 -8054 -20734 -8014 7 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_0.A
rlabel metal1 -20780 -8198 -20756 -8158 7 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_0.B
rlabel via1 -20248 -7142 -20154 -7116 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_0.VDD
rlabel metal1 -19390 -8170 -19338 -8092 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_0.Y
rlabel metal1 -20318 -8530 -20224 -8504 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_0.VSS
rlabel metal1 -18575 -9257 -18575 -9257 7 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A
rlabel metal1 -18575 -9425 -18575 -9425 7 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B
rlabel metal1 -18105 -9544 -18105 -9544 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.VSS
rlabel metal1 -18222 -8914 -18222 -8914 1 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.VDD
rlabel metal1 -17869 -9147 -17869 -9147 3 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.Y
rlabel metal1 -19457 -9257 -19457 -9257 7 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_1.A
rlabel metal1 -19457 -9425 -19457 -9425 7 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_1.B
rlabel metal1 -18987 -9544 -18987 -9544 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_1.VSS
rlabel metal1 -19104 -8914 -19104 -8914 1 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_1.VDD
rlabel metal1 -18751 -9147 -18751 -9147 3 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_1.Y
rlabel metal1 -20566 -9257 -20566 -9257 7 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_0.A
rlabel metal1 -20566 -9425 -20566 -9425 7 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_0.B
rlabel metal1 -20096 -9544 -20096 -9544 5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_0.VSS
rlabel metal1 -20213 -8914 -20213 -8914 1 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_0.VDD
rlabel metal1 -19860 -9147 -19860 -9147 3 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_0.Y
flabel metal2 -21031 -3822 -20961 -3762 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.A3
flabel metal2 -17735 -3842 -17665 -3782 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.A2
flabel metal2 -14447 -3844 -14377 -3784 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.A1
flabel metal2 -11155 -3828 -11085 -3768 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.A0
flabel metal2 -10977 -3828 -10907 -3768 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.B0
flabel metal2 -14267 -3844 -14197 -3784 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.B1
flabel metal2 -17561 -3842 -17491 -3782 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.B2
flabel metal2 -20847 -3822 -20777 -3762 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.B3
flabel metal1 -7765 -5430 -7693 -5360 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.C
flabel metal2 -7865 -6352 -7793 -6282 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.S0
flabel metal2 -11159 -6348 -11081 -6268 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.S1
flabel metal2 -14451 -6348 -14373 -6268 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.S2
flabel metal2 -17741 -6348 -17663 -6268 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.S3
flabel metal2 -21025 -6496 -20887 -6384 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.Cout
flabel metal5 -15355 -6670 -15217 -6558 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.VSS
flabel metal4 -15387 -3914 -15249 -3802 0 FreeSans 160 0 0 0 MULT_0.4bit_ADDER_0.VDD
rlabel metal1 -10962 -5434 -10926 -5364 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT
rlabel metal2 -7868 -6348 -7788 -6268 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.OUT
rlabel metal1 -8074 -5426 -7924 -5382 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.CIN
rlabel metal5 -10449 -6603 -10048 -6526 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.VSS
rlabel metal2 -11161 -3812 -11081 -3753 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.A
rlabel metal2 -10984 -3812 -10904 -3753 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.B
rlabel metal4 -9527 -3899 -9272 -3797 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.VDD
rlabel poly -9326 -4789 -9302 -4749 7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A
rlabel metal1 -9348 -4933 -9324 -4893 7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.B
rlabel via1 -8816 -3877 -8722 -3851 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.VDD
rlabel metal1 -7958 -4905 -7906 -4827 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.Y
rlabel metal1 -8886 -5265 -8792 -5239 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.VSS
rlabel poly -10885 -4789 -10861 -4749 7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_0.A
rlabel metal1 -10907 -4933 -10883 -4893 7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_0.B
rlabel via1 -10375 -3877 -10281 -3851 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_0.VDD
rlabel metal1 -9517 -4905 -9465 -4827 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_0.Y
rlabel metal1 -10445 -5265 -10351 -5239 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_0.VSS
rlabel metal1 -8702 -5992 -8702 -5992 7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A
rlabel metal1 -8702 -6160 -8702 -6160 7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B
rlabel metal1 -8232 -6279 -8232 -6279 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.VSS
rlabel metal1 -8349 -5649 -8349 -5649 1 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.VDD
rlabel metal1 -7996 -5882 -7996 -5882 3 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.Y
rlabel metal1 -9584 -5992 -9584 -5992 7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_1.A
rlabel metal1 -9584 -6160 -9584 -6160 7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_1.B
rlabel metal1 -9114 -6279 -9114 -6279 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_1.VSS
rlabel metal1 -9231 -5649 -9231 -5649 1 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_1.VDD
rlabel metal1 -8878 -5882 -8878 -5882 3 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_1.Y
rlabel metal1 -10693 -5992 -10693 -5992 7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_0.A
rlabel metal1 -10693 -6160 -10693 -6160 7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_0.B
rlabel metal1 -10223 -6279 -10223 -6279 5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_0.VSS
rlabel metal1 -10340 -5649 -10340 -5649 1 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_0.VDD
rlabel metal1 -9987 -5882 -9987 -5882 3 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_0.Y
rlabel metal1 -14253 -5434 -14217 -5364 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT
rlabel metal2 -11159 -6348 -11079 -6268 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.OUT
rlabel metal1 -11365 -5426 -11215 -5382 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.CIN
rlabel metal5 -13740 -6603 -13339 -6526 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.VSS
rlabel metal2 -14452 -3812 -14372 -3753 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.A
rlabel metal2 -14275 -3812 -14195 -3753 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.B
rlabel metal4 -12818 -3899 -12563 -3797 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.VDD
rlabel poly -12617 -4789 -12593 -4749 7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A
rlabel metal1 -12639 -4933 -12615 -4893 7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.B
rlabel via1 -12107 -3877 -12013 -3851 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.VDD
rlabel metal1 -11249 -4905 -11197 -4827 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.Y
rlabel metal1 -12177 -5265 -12083 -5239 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.VSS
rlabel poly -14176 -4789 -14152 -4749 7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_0.A
rlabel metal1 -14198 -4933 -14174 -4893 7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_0.B
rlabel via1 -13666 -3877 -13572 -3851 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_0.VDD
rlabel metal1 -12808 -4905 -12756 -4827 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_0.Y
rlabel metal1 -13736 -5265 -13642 -5239 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_0.VSS
rlabel metal1 -11993 -5992 -11993 -5992 7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A
rlabel metal1 -11993 -6160 -11993 -6160 7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B
rlabel metal1 -11523 -6279 -11523 -6279 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.VSS
rlabel metal1 -11640 -5649 -11640 -5649 1 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.VDD
rlabel metal1 -11287 -5882 -11287 -5882 3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.Y
rlabel metal1 -12875 -5992 -12875 -5992 7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_1.A
rlabel metal1 -12875 -6160 -12875 -6160 7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_1.B
rlabel metal1 -12405 -6279 -12405 -6279 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_1.VSS
rlabel metal1 -12522 -5649 -12522 -5649 1 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_1.VDD
rlabel metal1 -12169 -5882 -12169 -5882 3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_1.Y
rlabel metal1 -13984 -5992 -13984 -5992 7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_0.A
rlabel metal1 -13984 -6160 -13984 -6160 7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_0.B
rlabel metal1 -13514 -6279 -13514 -6279 5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_0.VSS
rlabel metal1 -13631 -5649 -13631 -5649 1 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_0.VDD
rlabel metal1 -13278 -5882 -13278 -5882 3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_0.Y
rlabel metal1 -17544 -5434 -17508 -5364 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT
rlabel metal2 -14450 -6348 -14370 -6268 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.OUT
rlabel metal1 -14656 -5426 -14506 -5382 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.CIN
rlabel metal5 -17031 -6603 -16630 -6526 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.VSS
rlabel metal2 -17743 -3812 -17663 -3753 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.A
rlabel metal2 -17566 -3812 -17486 -3753 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.B
rlabel metal4 -16109 -3899 -15854 -3797 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.VDD
rlabel poly -15908 -4789 -15884 -4749 7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A
rlabel metal1 -15930 -4933 -15906 -4893 7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.B
rlabel via1 -15398 -3877 -15304 -3851 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.VDD
rlabel metal1 -14540 -4905 -14488 -4827 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.Y
rlabel metal1 -15468 -5265 -15374 -5239 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.VSS
rlabel poly -17467 -4789 -17443 -4749 7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_0.A
rlabel metal1 -17489 -4933 -17465 -4893 7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_0.B
rlabel via1 -16957 -3877 -16863 -3851 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_0.VDD
rlabel metal1 -16099 -4905 -16047 -4827 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_0.Y
rlabel metal1 -17027 -5265 -16933 -5239 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_0.VSS
rlabel metal1 -15284 -5992 -15284 -5992 7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A
rlabel metal1 -15284 -6160 -15284 -6160 7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B
rlabel metal1 -14814 -6279 -14814 -6279 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.VSS
rlabel metal1 -14931 -5649 -14931 -5649 1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.VDD
rlabel metal1 -14578 -5882 -14578 -5882 3 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.Y
rlabel metal1 -16166 -5992 -16166 -5992 7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_1.A
rlabel metal1 -16166 -6160 -16166 -6160 7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_1.B
rlabel metal1 -15696 -6279 -15696 -6279 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_1.VSS
rlabel metal1 -15813 -5649 -15813 -5649 1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_1.VDD
rlabel metal1 -15460 -5882 -15460 -5882 3 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_1.Y
rlabel metal1 -17275 -5992 -17275 -5992 7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_0.A
rlabel metal1 -17275 -6160 -17275 -6160 7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_0.B
rlabel metal1 -16805 -6279 -16805 -6279 5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_0.VSS
rlabel metal1 -16922 -5649 -16922 -5649 1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_0.VDD
rlabel metal1 -16569 -5882 -16569 -5882 3 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_0.Y
rlabel metal1 -20835 -5434 -20799 -5364 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.COUT
rlabel metal2 -17741 -6348 -17661 -6268 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.OUT
rlabel metal1 -17947 -5426 -17797 -5382 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.CIN
rlabel metal5 -20322 -6603 -19921 -6526 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.VSS
rlabel metal2 -21034 -3812 -20954 -3753 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.A
rlabel metal2 -20857 -3812 -20777 -3753 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.B
rlabel metal4 -19400 -3899 -19145 -3797 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.VDD
rlabel poly -19199 -4789 -19175 -4749 7 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A
rlabel metal1 -19221 -4933 -19197 -4893 7 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.B
rlabel via1 -18689 -3877 -18595 -3851 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.VDD
rlabel metal1 -17831 -4905 -17779 -4827 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.Y
rlabel metal1 -18759 -5265 -18665 -5239 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.VSS
rlabel poly -20758 -4789 -20734 -4749 7 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_0.A
rlabel metal1 -20780 -4933 -20756 -4893 7 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_0.B
rlabel via1 -20248 -3877 -20154 -3851 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_0.VDD
rlabel metal1 -19390 -4905 -19338 -4827 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_0.Y
rlabel metal1 -20318 -5265 -20224 -5239 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_0.VSS
rlabel metal1 -18575 -5992 -18575 -5992 7 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A
rlabel metal1 -18575 -6160 -18575 -6160 7 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B
rlabel metal1 -18105 -6279 -18105 -6279 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.VSS
rlabel metal1 -18222 -5649 -18222 -5649 1 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.VDD
rlabel metal1 -17869 -5882 -17869 -5882 3 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.Y
rlabel metal1 -19457 -5992 -19457 -5992 7 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_1.A
rlabel metal1 -19457 -6160 -19457 -6160 7 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_1.B
rlabel metal1 -18987 -6279 -18987 -6279 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_1.VSS
rlabel metal1 -19104 -5649 -19104 -5649 1 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_1.VDD
rlabel metal1 -18751 -5882 -18751 -5882 3 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_1.Y
rlabel metal1 -20566 -5992 -20566 -5992 7 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_0.A
rlabel metal1 -20566 -6160 -20566 -6160 7 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_0.B
rlabel metal1 -20096 -6279 -20096 -6279 5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_0.VSS
rlabel metal1 -20213 -5649 -20213 -5649 1 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_0.VDD
rlabel metal1 -19860 -5882 -19860 -5882 3 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_0.Y
rlabel metal1 -23684 -7688 -23684 -7688 3 MULT_0.inv_6.A
rlabel metal1 -23486 -8077 -23486 -8077 5 MULT_0.inv_6.VSS
rlabel metal1 -23474 -7280 -23474 -7280 5 MULT_0.inv_6.VDD
rlabel metal1 -23272 -7688 -23272 -7688 3 MULT_0.inv_6.Y
rlabel metal1 -23683 -8980 -23683 -8980 3 MULT_0.inv_7.A
rlabel metal1 -23485 -9369 -23485 -9369 5 MULT_0.inv_7.VSS
rlabel metal1 -23473 -8572 -23473 -8572 5 MULT_0.inv_7.VDD
rlabel metal1 -23271 -8980 -23271 -8980 3 MULT_0.inv_7.Y
rlabel metal1 -21950 -7688 -21950 -7688 3 MULT_0.inv_12.A
rlabel metal1 -21752 -8077 -21752 -8077 5 MULT_0.inv_12.VSS
rlabel metal1 -21740 -7280 -21740 -7280 5 MULT_0.inv_12.VDD
rlabel metal1 -21538 -7688 -21538 -7688 3 MULT_0.inv_12.Y
rlabel metal1 -21946 -8980 -21946 -8980 3 MULT_0.inv_13.A
rlabel metal1 -21748 -9369 -21748 -9369 5 MULT_0.inv_13.VSS
rlabel metal1 -21736 -8572 -21736 -8572 5 MULT_0.inv_13.VDD
rlabel metal1 -21534 -8980 -21534 -8980 3 MULT_0.inv_13.Y
rlabel metal1 -24432 -7797 -24432 -7797 7 MULT_0.NAND2_6.A
rlabel metal1 -24432 -7965 -24432 -7965 7 MULT_0.NAND2_6.B
rlabel metal1 -23962 -8084 -23962 -8084 5 MULT_0.NAND2_6.VSS
rlabel metal1 -24079 -7454 -24079 -7454 1 MULT_0.NAND2_6.VDD
rlabel metal1 -23726 -7687 -23726 -7687 3 MULT_0.NAND2_6.Y
rlabel metal1 -24432 -9089 -24432 -9089 7 MULT_0.NAND2_7.A
rlabel metal1 -24432 -9257 -24432 -9257 7 MULT_0.NAND2_7.B
rlabel metal1 -23962 -9376 -23962 -9376 5 MULT_0.NAND2_7.VSS
rlabel metal1 -24079 -8746 -24079 -8746 1 MULT_0.NAND2_7.VDD
rlabel metal1 -23726 -8979 -23726 -8979 3 MULT_0.NAND2_7.Y
rlabel metal1 -22695 -7797 -22695 -7797 7 MULT_0.NAND2_12.A
rlabel metal1 -22695 -7965 -22695 -7965 7 MULT_0.NAND2_12.B
rlabel metal1 -22225 -8084 -22225 -8084 5 MULT_0.NAND2_12.VSS
rlabel metal1 -22342 -7454 -22342 -7454 1 MULT_0.NAND2_12.VDD
rlabel metal1 -21989 -7687 -21989 -7687 3 MULT_0.NAND2_12.Y
rlabel metal1 -22696 -9089 -22696 -9089 7 MULT_0.NAND2_13.A
rlabel metal1 -22696 -9257 -22696 -9257 7 MULT_0.NAND2_13.B
rlabel metal1 -22226 -9376 -22226 -9376 5 MULT_0.NAND2_13.VSS
rlabel metal1 -22343 -8746 -22343 -8746 1 MULT_0.NAND2_13.VDD
rlabel metal1 -21990 -8979 -21990 -8979 3 MULT_0.NAND2_13.Y
rlabel metal1 -24432 -5824 -24432 -5824 7 MULT_0.NAND2_5.A
rlabel metal1 -24432 -5992 -24432 -5992 7 MULT_0.NAND2_5.B
rlabel metal1 -23962 -6111 -23962 -6111 5 MULT_0.NAND2_5.VSS
rlabel metal1 -24079 -5481 -24079 -5481 1 MULT_0.NAND2_5.VDD
rlabel metal1 -23726 -5714 -23726 -5714 3 MULT_0.NAND2_5.Y
rlabel metal1 -24432 -4532 -24432 -4532 7 MULT_0.NAND2_4.A
rlabel metal1 -24432 -4700 -24432 -4700 7 MULT_0.NAND2_4.B
rlabel metal1 -23962 -4819 -23962 -4819 5 MULT_0.NAND2_4.VSS
rlabel metal1 -24079 -4189 -24079 -4189 1 MULT_0.NAND2_4.VDD
rlabel metal1 -23726 -4422 -23726 -4422 3 MULT_0.NAND2_4.Y
rlabel metal1 -24483 -2720 -24483 -2720 7 MULT_0.NAND2_0.A
rlabel metal1 -24483 -2888 -24483 -2888 7 MULT_0.NAND2_0.B
rlabel metal1 -24013 -3007 -24013 -3007 5 MULT_0.NAND2_0.VSS
rlabel metal1 -24130 -2377 -24130 -2377 1 MULT_0.NAND2_0.VDD
rlabel metal1 -23777 -2610 -23777 -2610 3 MULT_0.NAND2_0.Y
rlabel metal1 -23684 -4423 -23684 -4423 3 MULT_0.inv_5.A
rlabel metal1 -23486 -4812 -23486 -4812 5 MULT_0.inv_5.VSS
rlabel metal1 -23474 -4015 -23474 -4015 5 MULT_0.inv_5.VDD
rlabel metal1 -23272 -4423 -23272 -4423 3 MULT_0.inv_5.Y
rlabel metal1 -23686 -5715 -23686 -5715 3 MULT_0.inv_4.A
rlabel metal1 -23488 -6104 -23488 -6104 5 MULT_0.inv_4.VSS
rlabel metal1 -23476 -5307 -23476 -5307 5 MULT_0.inv_4.VDD
rlabel metal1 -23274 -5715 -23274 -5715 3 MULT_0.inv_4.Y
rlabel metal1 -22696 -5824 -22696 -5824 7 MULT_0.NAND2_11.A
rlabel metal1 -22696 -5992 -22696 -5992 7 MULT_0.NAND2_11.B
rlabel metal1 -22226 -6111 -22226 -6111 5 MULT_0.NAND2_11.VSS
rlabel metal1 -22343 -5481 -22343 -5481 1 MULT_0.NAND2_11.VDD
rlabel metal1 -21990 -5714 -21990 -5714 3 MULT_0.NAND2_11.Y
rlabel metal1 -22696 -4532 -22696 -4532 7 MULT_0.NAND2_10.A
rlabel metal1 -22696 -4700 -22696 -4700 7 MULT_0.NAND2_10.B
rlabel metal1 -22226 -4819 -22226 -4819 5 MULT_0.NAND2_10.VSS
rlabel metal1 -22343 -4189 -22343 -4189 1 MULT_0.NAND2_10.VDD
rlabel metal1 -21990 -4422 -21990 -4422 3 MULT_0.NAND2_10.Y
rlabel metal1 -22446 -2720 -22446 -2720 7 MULT_0.NAND2_1.A
rlabel metal1 -22446 -2888 -22446 -2888 7 MULT_0.NAND2_1.B
rlabel metal1 -21976 -3007 -21976 -3007 5 MULT_0.NAND2_1.VSS
rlabel metal1 -22093 -2377 -22093 -2377 1 MULT_0.NAND2_1.VDD
rlabel metal1 -21740 -2610 -21740 -2610 3 MULT_0.NAND2_1.Y
rlabel metal1 -21952 -5715 -21952 -5715 3 MULT_0.inv_11.A
rlabel metal1 -21754 -6104 -21754 -6104 5 MULT_0.inv_11.VSS
rlabel metal1 -21742 -5307 -21742 -5307 5 MULT_0.inv_11.VDD
rlabel metal1 -21540 -5715 -21540 -5715 3 MULT_0.inv_11.Y
rlabel metal1 -21946 -4423 -21946 -4423 3 MULT_0.inv_10.A
rlabel metal1 -21748 -4812 -21748 -4812 5 MULT_0.inv_10.VSS
rlabel metal1 -21736 -4015 -21736 -4015 5 MULT_0.inv_10.VDD
rlabel metal1 -21534 -4423 -21534 -4423 3 MULT_0.inv_10.Y
rlabel metal1 -20716 -2720 -20716 -2720 7 MULT_0.NAND2_2.A
rlabel metal1 -20716 -2888 -20716 -2888 7 MULT_0.NAND2_2.B
rlabel metal1 -20246 -3007 -20246 -3007 5 MULT_0.NAND2_2.VSS
rlabel metal1 -20363 -2377 -20363 -2377 1 MULT_0.NAND2_2.VDD
rlabel metal1 -20010 -2610 -20010 -2610 3 MULT_0.NAND2_2.Y
rlabel metal1 -18956 -2720 -18956 -2720 7 MULT_0.NAND2_3.A
rlabel metal1 -18956 -2888 -18956 -2888 7 MULT_0.NAND2_3.B
rlabel metal1 -18486 -3007 -18486 -3007 5 MULT_0.NAND2_3.VSS
rlabel metal1 -18603 -2377 -18603 -2377 1 MULT_0.NAND2_3.VDD
rlabel metal1 -18250 -2610 -18250 -2610 3 MULT_0.NAND2_3.Y
rlabel metal1 -23728 -2611 -23728 -2611 3 MULT_0.inv_0.A
rlabel metal1 -23530 -3000 -23530 -3000 5 MULT_0.inv_0.VSS
rlabel metal1 -23518 -2203 -23518 -2203 5 MULT_0.inv_0.VDD
rlabel metal1 -23316 -2611 -23316 -2611 3 MULT_0.inv_0.Y
rlabel metal1 -21708 -2611 -21708 -2611 3 MULT_0.inv_1.A
rlabel metal1 -21510 -3000 -21510 -3000 5 MULT_0.inv_1.VSS
rlabel metal1 -21498 -2203 -21498 -2203 5 MULT_0.inv_1.VDD
rlabel metal1 -21296 -2611 -21296 -2611 3 MULT_0.inv_1.Y
rlabel metal1 -19967 -2611 -19967 -2611 3 MULT_0.inv_2.A
rlabel metal1 -19769 -3000 -19769 -3000 5 MULT_0.inv_2.VSS
rlabel metal1 -19757 -2203 -19757 -2203 5 MULT_0.inv_2.VDD
rlabel metal1 -19555 -2611 -19555 -2611 3 MULT_0.inv_2.Y
rlabel metal1 -18188 -2611 -18188 -2611 3 MULT_0.inv_3.A
rlabel metal1 -17990 -3000 -17990 -3000 5 MULT_0.inv_3.VSS
rlabel metal1 -17978 -2203 -17978 -2203 5 MULT_0.inv_3.VDD
rlabel metal1 -17776 -2611 -17776 -2611 3 MULT_0.inv_3.Y
flabel space 9272 3385 9338 3451 0 FreeSans 1600 0 0 0 mux8_0.000
flabel space 10238 3378 10245 3380 0 FreeSans 1600 0 0 0 mux8_0.001
flabel space 7382 3384 7385 3384 0 FreeSans 1600 0 0 0 mux8_0.010
flabel space 8270 3389 8594 3448 0 FreeSans 1600 0 0 0 mux8_0.011
flabel space 9211 -327 9637 -270 0 FreeSans 1600 0 0 0 mux8_0.100
flabel space 10193 -349 10471 -190 0 FreeSans 1600 0 0 0 mux8_0.101
flabel space 7299 -400 7617 -225 0 FreeSans 1600 0 0 0 mux8_0.110
flabel space 8304 -378 8622 -203 0 FreeSans 1600 0 0 0 mux8_0.111
flabel metal2 5740 2458 5792 2510 0 FreeSans 160 0 0 0 mux8_0.A0
flabel metal2 5743 2363 5795 2415 0 FreeSans 160 0 0 0 mux8_0.A1
flabel metal2 5746 2257 5798 2309 0 FreeSans 160 0 0 0 mux8_0.A2
flabel metal2 5741 2151 5793 2203 0 FreeSans 160 0 0 0 mux8_0.A3
flabel metal2 5744 1053 5796 1105 0 FreeSans 160 0 0 0 mux8_0.A4
flabel metal2 5746 929 5798 981 0 FreeSans 160 0 0 0 mux8_0.A5
flabel metal2 5743 833 5795 885 0 FreeSans 160 0 0 0 mux8_0.A6
flabel metal2 5739 712 5791 764 0 FreeSans 160 0 0 0 mux8_0.A7
flabel metal1 12377 3097 12429 3149 0 FreeSans 160 0 0 0 mux8_0.VDD
flabel metal1 13159 1457 13211 1509 0 FreeSans 160 0 0 0 mux8_0.Y
flabel metal5 12955 810 13007 862 0 FreeSans 160 0 0 0 mux8_0.VSS
flabel metal2 6448 4081 6493 4120 0 FreeSans 160 0 0 0 mux8_0.SEL0
flabel metal2 6007 4072 6052 4111 0 FreeSans 160 0 0 0 mux8_0.SEL1
flabel metal2 5569 4072 5614 4111 0 FreeSans 160 0 0 0 mux8_0.SEL2
flabel metal1 8057 2524 8091 2573 0 FreeSans 160 0 0 0 mux8_0.NAND4F_2.A
flabel metal1 8060 2624 8094 2673 0 FreeSans 160 0 0 0 mux8_0.NAND4F_2.B
flabel metal1 8061 2712 8095 2761 0 FreeSans 160 0 0 0 mux8_0.NAND4F_2.C
flabel metal1 8062 2805 8096 2854 0 FreeSans 160 0 0 0 mux8_0.NAND4F_2.D
flabel metal1 8199 1706 8233 1755 0 FreeSans 160 0 0 0 mux8_0.NAND4F_2.VSS
flabel nwell 8462 3267 8496 3316 0 FreeSans 160 0 0 0 mux8_0.NAND4F_2.VDD
flabel metal1 8895 2587 8929 2636 0 FreeSans 160 0 0 0 mux8_0.NAND4F_2.Y
flabel metal1 7109 2524 7143 2573 0 FreeSans 160 0 0 0 mux8_0.NAND4F_4.A
flabel metal1 7112 2624 7146 2673 0 FreeSans 160 0 0 0 mux8_0.NAND4F_4.B
flabel metal1 7113 2712 7147 2761 0 FreeSans 160 0 0 0 mux8_0.NAND4F_4.C
flabel metal1 7114 2805 7148 2854 0 FreeSans 160 0 0 0 mux8_0.NAND4F_4.D
flabel metal1 7251 1706 7285 1755 0 FreeSans 160 0 0 0 mux8_0.NAND4F_4.VSS
flabel nwell 7514 3267 7548 3316 0 FreeSans 160 0 0 0 mux8_0.NAND4F_4.VDD
flabel metal1 7947 2587 7981 2636 0 FreeSans 160 0 0 0 mux8_0.NAND4F_4.Y
flabel metal1 7109 679 7143 728 0 FreeSans 160 0 0 0 mux8_0.NAND4F_5.A
flabel metal1 7112 579 7146 628 0 FreeSans 160 0 0 0 mux8_0.NAND4F_5.B
flabel metal1 7113 491 7147 540 0 FreeSans 160 0 0 0 mux8_0.NAND4F_5.C
flabel metal1 7114 398 7148 447 0 FreeSans 160 0 0 0 mux8_0.NAND4F_5.D
flabel metal1 7251 1497 7285 1546 0 FreeSans 160 0 0 0 mux8_0.NAND4F_5.VSS
flabel nwell 7514 -64 7548 -15 0 FreeSans 160 0 0 0 mux8_0.NAND4F_5.VDD
flabel metal1 7947 616 7981 665 0 FreeSans 160 0 0 0 mux8_0.NAND4F_5.Y
flabel metal1 8057 679 8091 728 0 FreeSans 160 0 0 0 mux8_0.NAND4F_6.A
flabel metal1 8060 579 8094 628 0 FreeSans 160 0 0 0 mux8_0.NAND4F_6.B
flabel metal1 8061 491 8095 540 0 FreeSans 160 0 0 0 mux8_0.NAND4F_6.C
flabel metal1 8062 398 8096 447 0 FreeSans 160 0 0 0 mux8_0.NAND4F_6.D
flabel metal1 8199 1497 8233 1546 0 FreeSans 160 0 0 0 mux8_0.NAND4F_6.VSS
flabel nwell 8462 -64 8496 -15 0 FreeSans 160 0 0 0 mux8_0.NAND4F_6.VDD
flabel metal1 8895 616 8929 665 0 FreeSans 160 0 0 0 mux8_0.NAND4F_6.Y
flabel metal1 9924 2524 9958 2573 0 FreeSans 160 0 0 0 mux8_0.NAND4F_0.A
flabel metal1 9927 2624 9961 2673 0 FreeSans 160 0 0 0 mux8_0.NAND4F_0.B
flabel metal1 9928 2712 9962 2761 0 FreeSans 160 0 0 0 mux8_0.NAND4F_0.C
flabel metal1 9929 2805 9963 2854 0 FreeSans 160 0 0 0 mux8_0.NAND4F_0.D
flabel metal1 10066 1706 10100 1755 0 FreeSans 160 0 0 0 mux8_0.NAND4F_0.VSS
flabel nwell 10329 3267 10363 3316 0 FreeSans 160 0 0 0 mux8_0.NAND4F_0.VDD
flabel metal1 10762 2587 10796 2636 0 FreeSans 160 0 0 0 mux8_0.NAND4F_0.Y
flabel metal1 8993 679 9027 728 0 FreeSans 160 0 0 0 mux8_0.NAND4F_1.A
flabel metal1 8996 579 9030 628 0 FreeSans 160 0 0 0 mux8_0.NAND4F_1.B
flabel metal1 8997 491 9031 540 0 FreeSans 160 0 0 0 mux8_0.NAND4F_1.C
flabel metal1 8998 398 9032 447 0 FreeSans 160 0 0 0 mux8_0.NAND4F_1.D
flabel metal1 9135 1497 9169 1546 0 FreeSans 160 0 0 0 mux8_0.NAND4F_1.VSS
flabel nwell 9398 -64 9432 -15 0 FreeSans 160 0 0 0 mux8_0.NAND4F_1.VDD
flabel metal1 9831 616 9865 665 0 FreeSans 160 0 0 0 mux8_0.NAND4F_1.Y
flabel metal1 8993 2524 9027 2573 0 FreeSans 160 0 0 0 mux8_0.NAND4F_3.A
flabel metal1 8996 2624 9030 2673 0 FreeSans 160 0 0 0 mux8_0.NAND4F_3.B
flabel metal1 8997 2712 9031 2761 0 FreeSans 160 0 0 0 mux8_0.NAND4F_3.C
flabel metal1 8998 2805 9032 2854 0 FreeSans 160 0 0 0 mux8_0.NAND4F_3.D
flabel metal1 9135 1706 9169 1755 0 FreeSans 160 0 0 0 mux8_0.NAND4F_3.VSS
flabel nwell 9398 3267 9432 3316 0 FreeSans 160 0 0 0 mux8_0.NAND4F_3.VDD
flabel metal1 9831 2587 9865 2636 0 FreeSans 160 0 0 0 mux8_0.NAND4F_3.Y
flabel metal1 9924 680 9958 729 0 FreeSans 160 0 0 0 mux8_0.NAND4F_7.A
flabel metal1 9927 580 9961 629 0 FreeSans 160 0 0 0 mux8_0.NAND4F_7.B
flabel metal1 9928 492 9962 541 0 FreeSans 160 0 0 0 mux8_0.NAND4F_7.C
flabel metal1 9929 399 9963 448 0 FreeSans 160 0 0 0 mux8_0.NAND4F_7.D
flabel metal1 10066 1498 10100 1547 0 FreeSans 160 0 0 0 mux8_0.NAND4F_7.VSS
flabel nwell 10329 -63 10363 -14 0 FreeSans 160 0 0 0 mux8_0.NAND4F_7.VDD
flabel metal1 10762 617 10796 666 0 FreeSans 160 0 0 0 mux8_0.NAND4F_7.Y
flabel metal1 10851 2524 10885 2573 0 FreeSans 160 0 0 0 mux8_0.NAND4F_8.A
flabel metal1 10854 2624 10888 2673 0 FreeSans 160 0 0 0 mux8_0.NAND4F_8.B
flabel metal1 10855 2712 10889 2761 0 FreeSans 160 0 0 0 mux8_0.NAND4F_8.C
flabel metal1 10856 2805 10890 2854 0 FreeSans 160 0 0 0 mux8_0.NAND4F_8.D
flabel metal1 10993 1706 11027 1755 0 FreeSans 160 0 0 0 mux8_0.NAND4F_8.VSS
flabel nwell 11256 3267 11290 3316 0 FreeSans 160 0 0 0 mux8_0.NAND4F_8.VDD
flabel metal1 11689 2587 11723 2636 0 FreeSans 160 0 0 0 mux8_0.NAND4F_8.Y
flabel metal1 10851 679 10885 728 0 FreeSans 160 0 0 0 mux8_0.NAND4F_9.A
flabel metal1 10854 579 10888 628 0 FreeSans 160 0 0 0 mux8_0.NAND4F_9.B
flabel metal1 10855 491 10889 540 0 FreeSans 160 0 0 0 mux8_0.NAND4F_9.C
flabel metal1 10856 398 10890 447 0 FreeSans 160 0 0 0 mux8_0.NAND4F_9.D
flabel metal1 10993 1497 11027 1546 0 FreeSans 160 0 0 0 mux8_0.NAND4F_9.VSS
flabel nwell 11256 -64 11290 -15 0 FreeSans 160 0 0 0 mux8_0.NAND4F_9.VDD
flabel metal1 11689 616 11723 665 0 FreeSans 160 0 0 0 mux8_0.NAND4F_9.Y
rlabel metal1 12823 1601 12823 1601 3 mux8_0.inv_0.A
rlabel metal1 13021 1212 13021 1212 5 mux8_0.inv_0.VSS
rlabel metal1 13033 2009 13033 2009 5 mux8_0.inv_0.VDD
rlabel metal1 13235 1601 13235 1601 3 mux8_0.inv_0.Y
flabel metal1 11744 1660 11821 1712 1 FreeSerif 320 0 0 0 mux8_0.nor2_0.A
rlabel metal1 11990 2160 11990 2160 5 mux8_0.nor2_0.VDD
flabel metal1 11745 1554 11822 1606 1 FreeSerif 320 0 0 0 mux8_0.nor2_0.B
flabel metal1 12749 1548 12826 1600 1 FreeSerif 320 0 0 0 mux8_0.nor2_0.Y
rlabel metal1 12286 1182 12286 1182 5 mux8_0.nor2_0.VSS
rlabel metal1 5998 3619 5998 3619 3 mux8_0.inv_1.A
rlabel metal1 6196 3230 6196 3230 5 mux8_0.inv_1.VSS
rlabel metal1 6208 4027 6208 4027 5 mux8_0.inv_1.VDD
rlabel metal1 6410 3619 6410 3619 3 mux8_0.inv_1.Y
rlabel metal1 6438 3619 6438 3619 3 mux8_0.inv_2.A
rlabel metal1 6636 3230 6636 3230 5 mux8_0.inv_2.VSS
rlabel metal1 6648 4027 6648 4027 5 mux8_0.inv_2.VDD
rlabel metal1 6850 3619 6850 3619 3 mux8_0.inv_2.Y
rlabel metal1 5558 3619 5558 3619 3 mux8_0.inv_3.A
rlabel metal1 5756 3230 5756 3230 5 mux8_0.inv_3.VSS
rlabel metal1 5768 4027 5768 4027 5 mux8_0.inv_3.VDD
rlabel metal1 5970 3619 5970 3619 3 mux8_0.inv_3.Y
flabel space 9272 -1143 9338 -1077 0 FreeSans 1600 0 0 0 mux8_1.000
flabel space 10238 -1150 10245 -1148 0 FreeSans 1600 0 0 0 mux8_1.001
flabel space 7382 -1144 7385 -1144 0 FreeSans 1600 0 0 0 mux8_1.010
flabel space 8270 -1139 8594 -1080 0 FreeSans 1600 0 0 0 mux8_1.011
flabel space 9211 -4855 9637 -4798 0 FreeSans 1600 0 0 0 mux8_1.100
flabel space 10193 -4877 10471 -4718 0 FreeSans 1600 0 0 0 mux8_1.101
flabel space 7299 -4928 7617 -4753 0 FreeSans 1600 0 0 0 mux8_1.110
flabel space 8304 -4906 8622 -4731 0 FreeSans 1600 0 0 0 mux8_1.111
flabel metal2 5740 -2070 5792 -2018 0 FreeSans 160 0 0 0 mux8_1.A0
flabel metal2 5743 -2165 5795 -2113 0 FreeSans 160 0 0 0 mux8_1.A1
flabel metal2 5746 -2271 5798 -2219 0 FreeSans 160 0 0 0 mux8_1.A2
flabel metal2 5741 -2377 5793 -2325 0 FreeSans 160 0 0 0 mux8_1.A3
flabel metal2 5744 -3475 5796 -3423 0 FreeSans 160 0 0 0 mux8_1.A4
flabel metal2 5746 -3599 5798 -3547 0 FreeSans 160 0 0 0 mux8_1.A5
flabel metal2 5743 -3695 5795 -3643 0 FreeSans 160 0 0 0 mux8_1.A6
flabel metal2 5739 -3816 5791 -3764 0 FreeSans 160 0 0 0 mux8_1.A7
flabel metal1 12377 -1431 12429 -1379 0 FreeSans 160 0 0 0 mux8_1.VDD
flabel metal1 13159 -3071 13211 -3019 0 FreeSans 160 0 0 0 mux8_1.Y
flabel metal5 12955 -3718 13007 -3666 0 FreeSans 160 0 0 0 mux8_1.VSS
flabel metal2 6448 -447 6493 -408 0 FreeSans 160 0 0 0 mux8_1.SEL0
flabel metal2 6007 -456 6052 -417 0 FreeSans 160 0 0 0 mux8_1.SEL1
flabel metal2 5569 -456 5614 -417 0 FreeSans 160 0 0 0 mux8_1.SEL2
flabel metal1 8057 -2004 8091 -1955 0 FreeSans 160 0 0 0 mux8_1.NAND4F_2.A
flabel metal1 8060 -1904 8094 -1855 0 FreeSans 160 0 0 0 mux8_1.NAND4F_2.B
flabel metal1 8061 -1816 8095 -1767 0 FreeSans 160 0 0 0 mux8_1.NAND4F_2.C
flabel metal1 8062 -1723 8096 -1674 0 FreeSans 160 0 0 0 mux8_1.NAND4F_2.D
flabel metal1 8199 -2822 8233 -2773 0 FreeSans 160 0 0 0 mux8_1.NAND4F_2.VSS
flabel nwell 8462 -1261 8496 -1212 0 FreeSans 160 0 0 0 mux8_1.NAND4F_2.VDD
flabel metal1 8895 -1941 8929 -1892 0 FreeSans 160 0 0 0 mux8_1.NAND4F_2.Y
flabel metal1 7109 -2004 7143 -1955 0 FreeSans 160 0 0 0 mux8_1.NAND4F_4.A
flabel metal1 7112 -1904 7146 -1855 0 FreeSans 160 0 0 0 mux8_1.NAND4F_4.B
flabel metal1 7113 -1816 7147 -1767 0 FreeSans 160 0 0 0 mux8_1.NAND4F_4.C
flabel metal1 7114 -1723 7148 -1674 0 FreeSans 160 0 0 0 mux8_1.NAND4F_4.D
flabel metal1 7251 -2822 7285 -2773 0 FreeSans 160 0 0 0 mux8_1.NAND4F_4.VSS
flabel nwell 7514 -1261 7548 -1212 0 FreeSans 160 0 0 0 mux8_1.NAND4F_4.VDD
flabel metal1 7947 -1941 7981 -1892 0 FreeSans 160 0 0 0 mux8_1.NAND4F_4.Y
flabel metal1 7109 -3849 7143 -3800 0 FreeSans 160 0 0 0 mux8_1.NAND4F_5.A
flabel metal1 7112 -3949 7146 -3900 0 FreeSans 160 0 0 0 mux8_1.NAND4F_5.B
flabel metal1 7113 -4037 7147 -3988 0 FreeSans 160 0 0 0 mux8_1.NAND4F_5.C
flabel metal1 7114 -4130 7148 -4081 0 FreeSans 160 0 0 0 mux8_1.NAND4F_5.D
flabel metal1 7251 -3031 7285 -2982 0 FreeSans 160 0 0 0 mux8_1.NAND4F_5.VSS
flabel nwell 7514 -4592 7548 -4543 0 FreeSans 160 0 0 0 mux8_1.NAND4F_5.VDD
flabel metal1 7947 -3912 7981 -3863 0 FreeSans 160 0 0 0 mux8_1.NAND4F_5.Y
flabel metal1 8057 -3849 8091 -3800 0 FreeSans 160 0 0 0 mux8_1.NAND4F_6.A
flabel metal1 8060 -3949 8094 -3900 0 FreeSans 160 0 0 0 mux8_1.NAND4F_6.B
flabel metal1 8061 -4037 8095 -3988 0 FreeSans 160 0 0 0 mux8_1.NAND4F_6.C
flabel metal1 8062 -4130 8096 -4081 0 FreeSans 160 0 0 0 mux8_1.NAND4F_6.D
flabel metal1 8199 -3031 8233 -2982 0 FreeSans 160 0 0 0 mux8_1.NAND4F_6.VSS
flabel nwell 8462 -4592 8496 -4543 0 FreeSans 160 0 0 0 mux8_1.NAND4F_6.VDD
flabel metal1 8895 -3912 8929 -3863 0 FreeSans 160 0 0 0 mux8_1.NAND4F_6.Y
flabel metal1 9924 -2004 9958 -1955 0 FreeSans 160 0 0 0 mux8_1.NAND4F_0.A
flabel metal1 9927 -1904 9961 -1855 0 FreeSans 160 0 0 0 mux8_1.NAND4F_0.B
flabel metal1 9928 -1816 9962 -1767 0 FreeSans 160 0 0 0 mux8_1.NAND4F_0.C
flabel metal1 9929 -1723 9963 -1674 0 FreeSans 160 0 0 0 mux8_1.NAND4F_0.D
flabel metal1 10066 -2822 10100 -2773 0 FreeSans 160 0 0 0 mux8_1.NAND4F_0.VSS
flabel nwell 10329 -1261 10363 -1212 0 FreeSans 160 0 0 0 mux8_1.NAND4F_0.VDD
flabel metal1 10762 -1941 10796 -1892 0 FreeSans 160 0 0 0 mux8_1.NAND4F_0.Y
flabel metal1 8993 -3849 9027 -3800 0 FreeSans 160 0 0 0 mux8_1.NAND4F_1.A
flabel metal1 8996 -3949 9030 -3900 0 FreeSans 160 0 0 0 mux8_1.NAND4F_1.B
flabel metal1 8997 -4037 9031 -3988 0 FreeSans 160 0 0 0 mux8_1.NAND4F_1.C
flabel metal1 8998 -4130 9032 -4081 0 FreeSans 160 0 0 0 mux8_1.NAND4F_1.D
flabel metal1 9135 -3031 9169 -2982 0 FreeSans 160 0 0 0 mux8_1.NAND4F_1.VSS
flabel nwell 9398 -4592 9432 -4543 0 FreeSans 160 0 0 0 mux8_1.NAND4F_1.VDD
flabel metal1 9831 -3912 9865 -3863 0 FreeSans 160 0 0 0 mux8_1.NAND4F_1.Y
flabel metal1 8993 -2004 9027 -1955 0 FreeSans 160 0 0 0 mux8_1.NAND4F_3.A
flabel metal1 8996 -1904 9030 -1855 0 FreeSans 160 0 0 0 mux8_1.NAND4F_3.B
flabel metal1 8997 -1816 9031 -1767 0 FreeSans 160 0 0 0 mux8_1.NAND4F_3.C
flabel metal1 8998 -1723 9032 -1674 0 FreeSans 160 0 0 0 mux8_1.NAND4F_3.D
flabel metal1 9135 -2822 9169 -2773 0 FreeSans 160 0 0 0 mux8_1.NAND4F_3.VSS
flabel nwell 9398 -1261 9432 -1212 0 FreeSans 160 0 0 0 mux8_1.NAND4F_3.VDD
flabel metal1 9831 -1941 9865 -1892 0 FreeSans 160 0 0 0 mux8_1.NAND4F_3.Y
flabel metal1 9924 -3848 9958 -3799 0 FreeSans 160 0 0 0 mux8_1.NAND4F_7.A
flabel metal1 9927 -3948 9961 -3899 0 FreeSans 160 0 0 0 mux8_1.NAND4F_7.B
flabel metal1 9928 -4036 9962 -3987 0 FreeSans 160 0 0 0 mux8_1.NAND4F_7.C
flabel metal1 9929 -4129 9963 -4080 0 FreeSans 160 0 0 0 mux8_1.NAND4F_7.D
flabel metal1 10066 -3030 10100 -2981 0 FreeSans 160 0 0 0 mux8_1.NAND4F_7.VSS
flabel nwell 10329 -4591 10363 -4542 0 FreeSans 160 0 0 0 mux8_1.NAND4F_7.VDD
flabel metal1 10762 -3911 10796 -3862 0 FreeSans 160 0 0 0 mux8_1.NAND4F_7.Y
flabel metal1 10851 -2004 10885 -1955 0 FreeSans 160 0 0 0 mux8_1.NAND4F_8.A
flabel metal1 10854 -1904 10888 -1855 0 FreeSans 160 0 0 0 mux8_1.NAND4F_8.B
flabel metal1 10855 -1816 10889 -1767 0 FreeSans 160 0 0 0 mux8_1.NAND4F_8.C
flabel metal1 10856 -1723 10890 -1674 0 FreeSans 160 0 0 0 mux8_1.NAND4F_8.D
flabel metal1 10993 -2822 11027 -2773 0 FreeSans 160 0 0 0 mux8_1.NAND4F_8.VSS
flabel nwell 11256 -1261 11290 -1212 0 FreeSans 160 0 0 0 mux8_1.NAND4F_8.VDD
flabel metal1 11689 -1941 11723 -1892 0 FreeSans 160 0 0 0 mux8_1.NAND4F_8.Y
flabel metal1 10851 -3849 10885 -3800 0 FreeSans 160 0 0 0 mux8_1.NAND4F_9.A
flabel metal1 10854 -3949 10888 -3900 0 FreeSans 160 0 0 0 mux8_1.NAND4F_9.B
flabel metal1 10855 -4037 10889 -3988 0 FreeSans 160 0 0 0 mux8_1.NAND4F_9.C
flabel metal1 10856 -4130 10890 -4081 0 FreeSans 160 0 0 0 mux8_1.NAND4F_9.D
flabel metal1 10993 -3031 11027 -2982 0 FreeSans 160 0 0 0 mux8_1.NAND4F_9.VSS
flabel nwell 11256 -4592 11290 -4543 0 FreeSans 160 0 0 0 mux8_1.NAND4F_9.VDD
flabel metal1 11689 -3912 11723 -3863 0 FreeSans 160 0 0 0 mux8_1.NAND4F_9.Y
rlabel metal1 12823 -2927 12823 -2927 3 mux8_1.inv_0.A
rlabel metal1 13021 -3316 13021 -3316 5 mux8_1.inv_0.VSS
rlabel metal1 13033 -2519 13033 -2519 5 mux8_1.inv_0.VDD
rlabel metal1 13235 -2927 13235 -2927 3 mux8_1.inv_0.Y
flabel metal1 11744 -2868 11821 -2816 1 FreeSerif 320 0 0 0 mux8_1.nor2_0.A
rlabel metal1 11990 -2368 11990 -2368 5 mux8_1.nor2_0.VDD
flabel metal1 11745 -2974 11822 -2922 1 FreeSerif 320 0 0 0 mux8_1.nor2_0.B
flabel metal1 12749 -2980 12826 -2928 1 FreeSerif 320 0 0 0 mux8_1.nor2_0.Y
rlabel metal1 12286 -3346 12286 -3346 5 mux8_1.nor2_0.VSS
rlabel metal1 5998 -909 5998 -909 3 mux8_1.inv_1.A
rlabel metal1 6196 -1298 6196 -1298 5 mux8_1.inv_1.VSS
rlabel metal1 6208 -501 6208 -501 5 mux8_1.inv_1.VDD
rlabel metal1 6410 -909 6410 -909 3 mux8_1.inv_1.Y
rlabel metal1 6438 -909 6438 -909 3 mux8_1.inv_2.A
rlabel metal1 6636 -1298 6636 -1298 5 mux8_1.inv_2.VSS
rlabel metal1 6648 -501 6648 -501 5 mux8_1.inv_2.VDD
rlabel metal1 6850 -909 6850 -909 3 mux8_1.inv_2.Y
rlabel metal1 5558 -909 5558 -909 3 mux8_1.inv_3.A
rlabel metal1 5756 -1298 5756 -1298 5 mux8_1.inv_3.VSS
rlabel metal1 5768 -501 5768 -501 5 mux8_1.inv_3.VDD
rlabel metal1 5970 -909 5970 -909 3 mux8_1.inv_3.Y
flabel space 9272 -5571 9338 -5505 0 FreeSans 1600 0 0 0 mux8_2.000
flabel space 10238 -5578 10245 -5576 0 FreeSans 1600 0 0 0 mux8_2.001
flabel space 7382 -5572 7385 -5572 0 FreeSans 1600 0 0 0 mux8_2.010
flabel space 8270 -5567 8594 -5508 0 FreeSans 1600 0 0 0 mux8_2.011
flabel space 9211 -9283 9637 -9226 0 FreeSans 1600 0 0 0 mux8_2.100
flabel space 10193 -9305 10471 -9146 0 FreeSans 1600 0 0 0 mux8_2.101
flabel space 7299 -9356 7617 -9181 0 FreeSans 1600 0 0 0 mux8_2.110
flabel space 8304 -9334 8622 -9159 0 FreeSans 1600 0 0 0 mux8_2.111
flabel metal2 5740 -6498 5792 -6446 0 FreeSans 160 0 0 0 mux8_2.A0
flabel metal2 5743 -6593 5795 -6541 0 FreeSans 160 0 0 0 mux8_2.A1
flabel metal2 5746 -6699 5798 -6647 0 FreeSans 160 0 0 0 mux8_2.A2
flabel metal2 5741 -6805 5793 -6753 0 FreeSans 160 0 0 0 mux8_2.A3
flabel metal2 5744 -7903 5796 -7851 0 FreeSans 160 0 0 0 mux8_2.A4
flabel metal2 5746 -8027 5798 -7975 0 FreeSans 160 0 0 0 mux8_2.A5
flabel metal2 5743 -8123 5795 -8071 0 FreeSans 160 0 0 0 mux8_2.A6
flabel metal2 5739 -8244 5791 -8192 0 FreeSans 160 0 0 0 mux8_2.A7
flabel metal1 12377 -5859 12429 -5807 0 FreeSans 160 0 0 0 mux8_2.VDD
flabel metal1 13159 -7499 13211 -7447 0 FreeSans 160 0 0 0 mux8_2.Y
flabel metal5 12955 -8146 13007 -8094 0 FreeSans 160 0 0 0 mux8_2.VSS
flabel metal2 6448 -4875 6493 -4836 0 FreeSans 160 0 0 0 mux8_2.SEL0
flabel metal2 6007 -4884 6052 -4845 0 FreeSans 160 0 0 0 mux8_2.SEL1
flabel metal2 5569 -4884 5614 -4845 0 FreeSans 160 0 0 0 mux8_2.SEL2
flabel metal1 8057 -6432 8091 -6383 0 FreeSans 160 0 0 0 mux8_2.NAND4F_2.A
flabel metal1 8060 -6332 8094 -6283 0 FreeSans 160 0 0 0 mux8_2.NAND4F_2.B
flabel metal1 8061 -6244 8095 -6195 0 FreeSans 160 0 0 0 mux8_2.NAND4F_2.C
flabel metal1 8062 -6151 8096 -6102 0 FreeSans 160 0 0 0 mux8_2.NAND4F_2.D
flabel metal1 8199 -7250 8233 -7201 0 FreeSans 160 0 0 0 mux8_2.NAND4F_2.VSS
flabel nwell 8462 -5689 8496 -5640 0 FreeSans 160 0 0 0 mux8_2.NAND4F_2.VDD
flabel metal1 8895 -6369 8929 -6320 0 FreeSans 160 0 0 0 mux8_2.NAND4F_2.Y
flabel metal1 7109 -6432 7143 -6383 0 FreeSans 160 0 0 0 mux8_2.NAND4F_4.A
flabel metal1 7112 -6332 7146 -6283 0 FreeSans 160 0 0 0 mux8_2.NAND4F_4.B
flabel metal1 7113 -6244 7147 -6195 0 FreeSans 160 0 0 0 mux8_2.NAND4F_4.C
flabel metal1 7114 -6151 7148 -6102 0 FreeSans 160 0 0 0 mux8_2.NAND4F_4.D
flabel metal1 7251 -7250 7285 -7201 0 FreeSans 160 0 0 0 mux8_2.NAND4F_4.VSS
flabel nwell 7514 -5689 7548 -5640 0 FreeSans 160 0 0 0 mux8_2.NAND4F_4.VDD
flabel metal1 7947 -6369 7981 -6320 0 FreeSans 160 0 0 0 mux8_2.NAND4F_4.Y
flabel metal1 7109 -8277 7143 -8228 0 FreeSans 160 0 0 0 mux8_2.NAND4F_5.A
flabel metal1 7112 -8377 7146 -8328 0 FreeSans 160 0 0 0 mux8_2.NAND4F_5.B
flabel metal1 7113 -8465 7147 -8416 0 FreeSans 160 0 0 0 mux8_2.NAND4F_5.C
flabel metal1 7114 -8558 7148 -8509 0 FreeSans 160 0 0 0 mux8_2.NAND4F_5.D
flabel metal1 7251 -7459 7285 -7410 0 FreeSans 160 0 0 0 mux8_2.NAND4F_5.VSS
flabel nwell 7514 -9020 7548 -8971 0 FreeSans 160 0 0 0 mux8_2.NAND4F_5.VDD
flabel metal1 7947 -8340 7981 -8291 0 FreeSans 160 0 0 0 mux8_2.NAND4F_5.Y
flabel metal1 8057 -8277 8091 -8228 0 FreeSans 160 0 0 0 mux8_2.NAND4F_6.A
flabel metal1 8060 -8377 8094 -8328 0 FreeSans 160 0 0 0 mux8_2.NAND4F_6.B
flabel metal1 8061 -8465 8095 -8416 0 FreeSans 160 0 0 0 mux8_2.NAND4F_6.C
flabel metal1 8062 -8558 8096 -8509 0 FreeSans 160 0 0 0 mux8_2.NAND4F_6.D
flabel metal1 8199 -7459 8233 -7410 0 FreeSans 160 0 0 0 mux8_2.NAND4F_6.VSS
flabel nwell 8462 -9020 8496 -8971 0 FreeSans 160 0 0 0 mux8_2.NAND4F_6.VDD
flabel metal1 8895 -8340 8929 -8291 0 FreeSans 160 0 0 0 mux8_2.NAND4F_6.Y
flabel metal1 9924 -6432 9958 -6383 0 FreeSans 160 0 0 0 mux8_2.NAND4F_0.A
flabel metal1 9927 -6332 9961 -6283 0 FreeSans 160 0 0 0 mux8_2.NAND4F_0.B
flabel metal1 9928 -6244 9962 -6195 0 FreeSans 160 0 0 0 mux8_2.NAND4F_0.C
flabel metal1 9929 -6151 9963 -6102 0 FreeSans 160 0 0 0 mux8_2.NAND4F_0.D
flabel metal1 10066 -7250 10100 -7201 0 FreeSans 160 0 0 0 mux8_2.NAND4F_0.VSS
flabel nwell 10329 -5689 10363 -5640 0 FreeSans 160 0 0 0 mux8_2.NAND4F_0.VDD
flabel metal1 10762 -6369 10796 -6320 0 FreeSans 160 0 0 0 mux8_2.NAND4F_0.Y
flabel metal1 8993 -8277 9027 -8228 0 FreeSans 160 0 0 0 mux8_2.NAND4F_1.A
flabel metal1 8996 -8377 9030 -8328 0 FreeSans 160 0 0 0 mux8_2.NAND4F_1.B
flabel metal1 8997 -8465 9031 -8416 0 FreeSans 160 0 0 0 mux8_2.NAND4F_1.C
flabel metal1 8998 -8558 9032 -8509 0 FreeSans 160 0 0 0 mux8_2.NAND4F_1.D
flabel metal1 9135 -7459 9169 -7410 0 FreeSans 160 0 0 0 mux8_2.NAND4F_1.VSS
flabel nwell 9398 -9020 9432 -8971 0 FreeSans 160 0 0 0 mux8_2.NAND4F_1.VDD
flabel metal1 9831 -8340 9865 -8291 0 FreeSans 160 0 0 0 mux8_2.NAND4F_1.Y
flabel metal1 8993 -6432 9027 -6383 0 FreeSans 160 0 0 0 mux8_2.NAND4F_3.A
flabel metal1 8996 -6332 9030 -6283 0 FreeSans 160 0 0 0 mux8_2.NAND4F_3.B
flabel metal1 8997 -6244 9031 -6195 0 FreeSans 160 0 0 0 mux8_2.NAND4F_3.C
flabel metal1 8998 -6151 9032 -6102 0 FreeSans 160 0 0 0 mux8_2.NAND4F_3.D
flabel metal1 9135 -7250 9169 -7201 0 FreeSans 160 0 0 0 mux8_2.NAND4F_3.VSS
flabel nwell 9398 -5689 9432 -5640 0 FreeSans 160 0 0 0 mux8_2.NAND4F_3.VDD
flabel metal1 9831 -6369 9865 -6320 0 FreeSans 160 0 0 0 mux8_2.NAND4F_3.Y
flabel metal1 9924 -8276 9958 -8227 0 FreeSans 160 0 0 0 mux8_2.NAND4F_7.A
flabel metal1 9927 -8376 9961 -8327 0 FreeSans 160 0 0 0 mux8_2.NAND4F_7.B
flabel metal1 9928 -8464 9962 -8415 0 FreeSans 160 0 0 0 mux8_2.NAND4F_7.C
flabel metal1 9929 -8557 9963 -8508 0 FreeSans 160 0 0 0 mux8_2.NAND4F_7.D
flabel metal1 10066 -7458 10100 -7409 0 FreeSans 160 0 0 0 mux8_2.NAND4F_7.VSS
flabel nwell 10329 -9019 10363 -8970 0 FreeSans 160 0 0 0 mux8_2.NAND4F_7.VDD
flabel metal1 10762 -8339 10796 -8290 0 FreeSans 160 0 0 0 mux8_2.NAND4F_7.Y
flabel metal1 10851 -6432 10885 -6383 0 FreeSans 160 0 0 0 mux8_2.NAND4F_8.A
flabel metal1 10854 -6332 10888 -6283 0 FreeSans 160 0 0 0 mux8_2.NAND4F_8.B
flabel metal1 10855 -6244 10889 -6195 0 FreeSans 160 0 0 0 mux8_2.NAND4F_8.C
flabel metal1 10856 -6151 10890 -6102 0 FreeSans 160 0 0 0 mux8_2.NAND4F_8.D
flabel metal1 10993 -7250 11027 -7201 0 FreeSans 160 0 0 0 mux8_2.NAND4F_8.VSS
flabel nwell 11256 -5689 11290 -5640 0 FreeSans 160 0 0 0 mux8_2.NAND4F_8.VDD
flabel metal1 11689 -6369 11723 -6320 0 FreeSans 160 0 0 0 mux8_2.NAND4F_8.Y
flabel metal1 10851 -8277 10885 -8228 0 FreeSans 160 0 0 0 mux8_2.NAND4F_9.A
flabel metal1 10854 -8377 10888 -8328 0 FreeSans 160 0 0 0 mux8_2.NAND4F_9.B
flabel metal1 10855 -8465 10889 -8416 0 FreeSans 160 0 0 0 mux8_2.NAND4F_9.C
flabel metal1 10856 -8558 10890 -8509 0 FreeSans 160 0 0 0 mux8_2.NAND4F_9.D
flabel metal1 10993 -7459 11027 -7410 0 FreeSans 160 0 0 0 mux8_2.NAND4F_9.VSS
flabel nwell 11256 -9020 11290 -8971 0 FreeSans 160 0 0 0 mux8_2.NAND4F_9.VDD
flabel metal1 11689 -8340 11723 -8291 0 FreeSans 160 0 0 0 mux8_2.NAND4F_9.Y
rlabel metal1 12823 -7355 12823 -7355 3 mux8_2.inv_0.A
rlabel metal1 13021 -7744 13021 -7744 5 mux8_2.inv_0.VSS
rlabel metal1 13033 -6947 13033 -6947 5 mux8_2.inv_0.VDD
rlabel metal1 13235 -7355 13235 -7355 3 mux8_2.inv_0.Y
flabel metal1 11744 -7296 11821 -7244 1 FreeSerif 320 0 0 0 mux8_2.nor2_0.A
rlabel metal1 11990 -6796 11990 -6796 5 mux8_2.nor2_0.VDD
flabel metal1 11745 -7402 11822 -7350 1 FreeSerif 320 0 0 0 mux8_2.nor2_0.B
flabel metal1 12749 -7408 12826 -7356 1 FreeSerif 320 0 0 0 mux8_2.nor2_0.Y
rlabel metal1 12286 -7774 12286 -7774 5 mux8_2.nor2_0.VSS
rlabel metal1 5998 -5337 5998 -5337 3 mux8_2.inv_1.A
rlabel metal1 6196 -5726 6196 -5726 5 mux8_2.inv_1.VSS
rlabel metal1 6208 -4929 6208 -4929 5 mux8_2.inv_1.VDD
rlabel metal1 6410 -5337 6410 -5337 3 mux8_2.inv_1.Y
rlabel metal1 6438 -5337 6438 -5337 3 mux8_2.inv_2.A
rlabel metal1 6636 -5726 6636 -5726 5 mux8_2.inv_2.VSS
rlabel metal1 6648 -4929 6648 -4929 5 mux8_2.inv_2.VDD
rlabel metal1 6850 -5337 6850 -5337 3 mux8_2.inv_2.Y
rlabel metal1 5558 -5337 5558 -5337 3 mux8_2.inv_3.A
rlabel metal1 5756 -5726 5756 -5726 5 mux8_2.inv_3.VSS
rlabel metal1 5768 -4929 5768 -4929 5 mux8_2.inv_3.VDD
rlabel metal1 5970 -5337 5970 -5337 3 mux8_2.inv_3.Y
flabel space 9272 -10199 9338 -10133 0 FreeSans 1600 0 0 0 mux8_3.000
flabel space 10238 -10206 10245 -10204 0 FreeSans 1600 0 0 0 mux8_3.001
flabel space 7382 -10200 7385 -10200 0 FreeSans 1600 0 0 0 mux8_3.010
flabel space 8270 -10195 8594 -10136 0 FreeSans 1600 0 0 0 mux8_3.011
flabel space 9211 -13911 9637 -13854 0 FreeSans 1600 0 0 0 mux8_3.100
flabel space 10193 -13933 10471 -13774 0 FreeSans 1600 0 0 0 mux8_3.101
flabel space 7299 -13984 7617 -13809 0 FreeSans 1600 0 0 0 mux8_3.110
flabel space 8304 -13962 8622 -13787 0 FreeSans 1600 0 0 0 mux8_3.111
flabel metal2 5740 -11126 5792 -11074 0 FreeSans 160 0 0 0 mux8_3.A0
flabel metal2 5743 -11221 5795 -11169 0 FreeSans 160 0 0 0 mux8_3.A1
flabel metal2 5746 -11327 5798 -11275 0 FreeSans 160 0 0 0 mux8_3.A2
flabel metal2 5741 -11433 5793 -11381 0 FreeSans 160 0 0 0 mux8_3.A3
flabel metal2 5744 -12531 5796 -12479 0 FreeSans 160 0 0 0 mux8_3.A4
flabel metal2 5746 -12655 5798 -12603 0 FreeSans 160 0 0 0 mux8_3.A5
flabel metal2 5743 -12751 5795 -12699 0 FreeSans 160 0 0 0 mux8_3.A6
flabel metal2 5739 -12872 5791 -12820 0 FreeSans 160 0 0 0 mux8_3.A7
flabel metal1 12377 -10487 12429 -10435 0 FreeSans 160 0 0 0 mux8_3.VDD
flabel metal1 13159 -12127 13211 -12075 0 FreeSans 160 0 0 0 mux8_3.Y
flabel metal5 12955 -12774 13007 -12722 0 FreeSans 160 0 0 0 mux8_3.VSS
flabel metal2 6448 -9503 6493 -9464 0 FreeSans 160 0 0 0 mux8_3.SEL0
flabel metal2 6007 -9512 6052 -9473 0 FreeSans 160 0 0 0 mux8_3.SEL1
flabel metal2 5569 -9512 5614 -9473 0 FreeSans 160 0 0 0 mux8_3.SEL2
flabel metal1 8057 -11060 8091 -11011 0 FreeSans 160 0 0 0 mux8_3.NAND4F_2.A
flabel metal1 8060 -10960 8094 -10911 0 FreeSans 160 0 0 0 mux8_3.NAND4F_2.B
flabel metal1 8061 -10872 8095 -10823 0 FreeSans 160 0 0 0 mux8_3.NAND4F_2.C
flabel metal1 8062 -10779 8096 -10730 0 FreeSans 160 0 0 0 mux8_3.NAND4F_2.D
flabel metal1 8199 -11878 8233 -11829 0 FreeSans 160 0 0 0 mux8_3.NAND4F_2.VSS
flabel nwell 8462 -10317 8496 -10268 0 FreeSans 160 0 0 0 mux8_3.NAND4F_2.VDD
flabel metal1 8895 -10997 8929 -10948 0 FreeSans 160 0 0 0 mux8_3.NAND4F_2.Y
flabel metal1 7109 -11060 7143 -11011 0 FreeSans 160 0 0 0 mux8_3.NAND4F_4.A
flabel metal1 7112 -10960 7146 -10911 0 FreeSans 160 0 0 0 mux8_3.NAND4F_4.B
flabel metal1 7113 -10872 7147 -10823 0 FreeSans 160 0 0 0 mux8_3.NAND4F_4.C
flabel metal1 7114 -10779 7148 -10730 0 FreeSans 160 0 0 0 mux8_3.NAND4F_4.D
flabel metal1 7251 -11878 7285 -11829 0 FreeSans 160 0 0 0 mux8_3.NAND4F_4.VSS
flabel nwell 7514 -10317 7548 -10268 0 FreeSans 160 0 0 0 mux8_3.NAND4F_4.VDD
flabel metal1 7947 -10997 7981 -10948 0 FreeSans 160 0 0 0 mux8_3.NAND4F_4.Y
flabel metal1 7109 -12905 7143 -12856 0 FreeSans 160 0 0 0 mux8_3.NAND4F_5.A
flabel metal1 7112 -13005 7146 -12956 0 FreeSans 160 0 0 0 mux8_3.NAND4F_5.B
flabel metal1 7113 -13093 7147 -13044 0 FreeSans 160 0 0 0 mux8_3.NAND4F_5.C
flabel metal1 7114 -13186 7148 -13137 0 FreeSans 160 0 0 0 mux8_3.NAND4F_5.D
flabel metal1 7251 -12087 7285 -12038 0 FreeSans 160 0 0 0 mux8_3.NAND4F_5.VSS
flabel nwell 7514 -13648 7548 -13599 0 FreeSans 160 0 0 0 mux8_3.NAND4F_5.VDD
flabel metal1 7947 -12968 7981 -12919 0 FreeSans 160 0 0 0 mux8_3.NAND4F_5.Y
flabel metal1 8057 -12905 8091 -12856 0 FreeSans 160 0 0 0 mux8_3.NAND4F_6.A
flabel metal1 8060 -13005 8094 -12956 0 FreeSans 160 0 0 0 mux8_3.NAND4F_6.B
flabel metal1 8061 -13093 8095 -13044 0 FreeSans 160 0 0 0 mux8_3.NAND4F_6.C
flabel metal1 8062 -13186 8096 -13137 0 FreeSans 160 0 0 0 mux8_3.NAND4F_6.D
flabel metal1 8199 -12087 8233 -12038 0 FreeSans 160 0 0 0 mux8_3.NAND4F_6.VSS
flabel nwell 8462 -13648 8496 -13599 0 FreeSans 160 0 0 0 mux8_3.NAND4F_6.VDD
flabel metal1 8895 -12968 8929 -12919 0 FreeSans 160 0 0 0 mux8_3.NAND4F_6.Y
flabel metal1 9924 -11060 9958 -11011 0 FreeSans 160 0 0 0 mux8_3.NAND4F_0.A
flabel metal1 9927 -10960 9961 -10911 0 FreeSans 160 0 0 0 mux8_3.NAND4F_0.B
flabel metal1 9928 -10872 9962 -10823 0 FreeSans 160 0 0 0 mux8_3.NAND4F_0.C
flabel metal1 9929 -10779 9963 -10730 0 FreeSans 160 0 0 0 mux8_3.NAND4F_0.D
flabel metal1 10066 -11878 10100 -11829 0 FreeSans 160 0 0 0 mux8_3.NAND4F_0.VSS
flabel nwell 10329 -10317 10363 -10268 0 FreeSans 160 0 0 0 mux8_3.NAND4F_0.VDD
flabel metal1 10762 -10997 10796 -10948 0 FreeSans 160 0 0 0 mux8_3.NAND4F_0.Y
flabel metal1 8993 -12905 9027 -12856 0 FreeSans 160 0 0 0 mux8_3.NAND4F_1.A
flabel metal1 8996 -13005 9030 -12956 0 FreeSans 160 0 0 0 mux8_3.NAND4F_1.B
flabel metal1 8997 -13093 9031 -13044 0 FreeSans 160 0 0 0 mux8_3.NAND4F_1.C
flabel metal1 8998 -13186 9032 -13137 0 FreeSans 160 0 0 0 mux8_3.NAND4F_1.D
flabel metal1 9135 -12087 9169 -12038 0 FreeSans 160 0 0 0 mux8_3.NAND4F_1.VSS
flabel nwell 9398 -13648 9432 -13599 0 FreeSans 160 0 0 0 mux8_3.NAND4F_1.VDD
flabel metal1 9831 -12968 9865 -12919 0 FreeSans 160 0 0 0 mux8_3.NAND4F_1.Y
flabel metal1 8993 -11060 9027 -11011 0 FreeSans 160 0 0 0 mux8_3.NAND4F_3.A
flabel metal1 8996 -10960 9030 -10911 0 FreeSans 160 0 0 0 mux8_3.NAND4F_3.B
flabel metal1 8997 -10872 9031 -10823 0 FreeSans 160 0 0 0 mux8_3.NAND4F_3.C
flabel metal1 8998 -10779 9032 -10730 0 FreeSans 160 0 0 0 mux8_3.NAND4F_3.D
flabel metal1 9135 -11878 9169 -11829 0 FreeSans 160 0 0 0 mux8_3.NAND4F_3.VSS
flabel nwell 9398 -10317 9432 -10268 0 FreeSans 160 0 0 0 mux8_3.NAND4F_3.VDD
flabel metal1 9831 -10997 9865 -10948 0 FreeSans 160 0 0 0 mux8_3.NAND4F_3.Y
flabel metal1 9924 -12904 9958 -12855 0 FreeSans 160 0 0 0 mux8_3.NAND4F_7.A
flabel metal1 9927 -13004 9961 -12955 0 FreeSans 160 0 0 0 mux8_3.NAND4F_7.B
flabel metal1 9928 -13092 9962 -13043 0 FreeSans 160 0 0 0 mux8_3.NAND4F_7.C
flabel metal1 9929 -13185 9963 -13136 0 FreeSans 160 0 0 0 mux8_3.NAND4F_7.D
flabel metal1 10066 -12086 10100 -12037 0 FreeSans 160 0 0 0 mux8_3.NAND4F_7.VSS
flabel nwell 10329 -13647 10363 -13598 0 FreeSans 160 0 0 0 mux8_3.NAND4F_7.VDD
flabel metal1 10762 -12967 10796 -12918 0 FreeSans 160 0 0 0 mux8_3.NAND4F_7.Y
flabel metal1 10851 -11060 10885 -11011 0 FreeSans 160 0 0 0 mux8_3.NAND4F_8.A
flabel metal1 10854 -10960 10888 -10911 0 FreeSans 160 0 0 0 mux8_3.NAND4F_8.B
flabel metal1 10855 -10872 10889 -10823 0 FreeSans 160 0 0 0 mux8_3.NAND4F_8.C
flabel metal1 10856 -10779 10890 -10730 0 FreeSans 160 0 0 0 mux8_3.NAND4F_8.D
flabel metal1 10993 -11878 11027 -11829 0 FreeSans 160 0 0 0 mux8_3.NAND4F_8.VSS
flabel nwell 11256 -10317 11290 -10268 0 FreeSans 160 0 0 0 mux8_3.NAND4F_8.VDD
flabel metal1 11689 -10997 11723 -10948 0 FreeSans 160 0 0 0 mux8_3.NAND4F_8.Y
flabel metal1 10851 -12905 10885 -12856 0 FreeSans 160 0 0 0 mux8_3.NAND4F_9.A
flabel metal1 10854 -13005 10888 -12956 0 FreeSans 160 0 0 0 mux8_3.NAND4F_9.B
flabel metal1 10855 -13093 10889 -13044 0 FreeSans 160 0 0 0 mux8_3.NAND4F_9.C
flabel metal1 10856 -13186 10890 -13137 0 FreeSans 160 0 0 0 mux8_3.NAND4F_9.D
flabel metal1 10993 -12087 11027 -12038 0 FreeSans 160 0 0 0 mux8_3.NAND4F_9.VSS
flabel nwell 11256 -13648 11290 -13599 0 FreeSans 160 0 0 0 mux8_3.NAND4F_9.VDD
flabel metal1 11689 -12968 11723 -12919 0 FreeSans 160 0 0 0 mux8_3.NAND4F_9.Y
rlabel metal1 12823 -11983 12823 -11983 3 mux8_3.inv_0.A
rlabel metal1 13021 -12372 13021 -12372 5 mux8_3.inv_0.VSS
rlabel metal1 13033 -11575 13033 -11575 5 mux8_3.inv_0.VDD
rlabel metal1 13235 -11983 13235 -11983 3 mux8_3.inv_0.Y
flabel metal1 11744 -11924 11821 -11872 1 FreeSerif 320 0 0 0 mux8_3.nor2_0.A
rlabel metal1 11990 -11424 11990 -11424 5 mux8_3.nor2_0.VDD
flabel metal1 11745 -12030 11822 -11978 1 FreeSerif 320 0 0 0 mux8_3.nor2_0.B
flabel metal1 12749 -12036 12826 -11984 1 FreeSerif 320 0 0 0 mux8_3.nor2_0.Y
rlabel metal1 12286 -12402 12286 -12402 5 mux8_3.nor2_0.VSS
rlabel metal1 5998 -9965 5998 -9965 3 mux8_3.inv_1.A
rlabel metal1 6196 -10354 6196 -10354 5 mux8_3.inv_1.VSS
rlabel metal1 6208 -9557 6208 -9557 5 mux8_3.inv_1.VDD
rlabel metal1 6410 -9965 6410 -9965 3 mux8_3.inv_1.Y
rlabel metal1 6438 -9965 6438 -9965 3 mux8_3.inv_2.A
rlabel metal1 6636 -10354 6636 -10354 5 mux8_3.inv_2.VSS
rlabel metal1 6648 -9557 6648 -9557 5 mux8_3.inv_2.VDD
rlabel metal1 6850 -9965 6850 -9965 3 mux8_3.inv_2.Y
rlabel metal1 5558 -9965 5558 -9965 3 mux8_3.inv_3.A
rlabel metal1 5756 -10354 5756 -10354 5 mux8_3.inv_3.VSS
rlabel metal1 5768 -9557 5768 -9557 5 mux8_3.inv_3.VDD
rlabel metal1 5970 -9965 5970 -9965 3 mux8_3.inv_3.Y
flabel metal1 1602 6263 1649 6301 0 FreeSans 160 0 0 0 V_FLAG_0.A_MSB
flabel metal1 1407 6261 1454 6299 0 FreeSans 160 0 0 0 V_FLAG_0.B_MSB
flabel metal1 3206 6311 3253 6349 0 FreeSans 160 0 0 0 V_FLAG_0.OPCODE3
flabel metal1 4759 6303 4801 6328 0 FreeSans 160 0 0 0 V_FLAG_0.Y_MSB
flabel metal1 8048 5056 8090 5081 0 FreeSans 160 0 0 0 V_FLAG_0.V
flabel metal5 3121 4640 3295 4910 0 FreeSans 1600 0 0 0 V_FLAG_0.VSS
flabel metal4 3059 6180 3121 6252 0 FreeSans 1600 0 0 0 V_FLAG_0.VDD
rlabel poly 3292 5279 3316 5319 7 V_FLAG_0.XOR2_2.A
rlabel metal1 3270 5135 3294 5175 7 V_FLAG_0.XOR2_2.B
rlabel via1 3802 6191 3896 6217 5 V_FLAG_0.XOR2_2.VDD
rlabel metal1 4660 5163 4712 5241 5 V_FLAG_0.XOR2_2.Y
rlabel metal1 3732 4803 3826 4829 5 V_FLAG_0.XOR2_2.VSS
rlabel poly 1686 5279 1710 5319 7 V_FLAG_0.XOR2_1.A
rlabel metal1 1664 5135 1688 5175 7 V_FLAG_0.XOR2_1.B
rlabel via1 2196 6191 2290 6217 5 V_FLAG_0.XOR2_1.VDD
rlabel metal1 3054 5163 3106 5241 5 V_FLAG_0.XOR2_1.Y
rlabel metal1 2126 4803 2220 4829 5 V_FLAG_0.XOR2_1.VSS
rlabel poly 4996 5277 5020 5317 7 V_FLAG_0.XOR2_0.A
rlabel metal1 4974 5133 4998 5173 7 V_FLAG_0.XOR2_0.B
rlabel via1 5506 6189 5600 6215 5 V_FLAG_0.XOR2_0.VDD
rlabel metal1 6364 5161 6416 5239 5 V_FLAG_0.XOR2_0.Y
rlabel metal1 5436 4801 5530 4827 5 V_FLAG_0.XOR2_0.VSS
rlabel metal1 6903 5134 6903 5134 7 V_FLAG_0.NAND2_0.A
rlabel metal1 6903 4966 6903 4966 7 V_FLAG_0.NAND2_0.B
rlabel metal1 7373 4847 7373 4847 5 V_FLAG_0.NAND2_0.VSS
rlabel metal1 7256 5477 7256 5477 1 V_FLAG_0.NAND2_0.VDD
rlabel metal1 7609 5244 7609 5244 3 V_FLAG_0.NAND2_0.Y
rlabel metal1 7709 5167 7709 5167 3 V_FLAG_0.inv_0.A
rlabel metal1 7907 4778 7907 4778 5 V_FLAG_0.inv_0.VSS
rlabel metal1 7919 5575 7919 5575 5 V_FLAG_0.inv_0.VDD
rlabel metal1 8121 5167 8121 5167 3 V_FLAG_0.inv_0.Y
<< end >>
