magic
tech sky130B
magscale 1 2
timestamp 1733174445
<< error_p >>
rect -265 -73 -207 11
rect -147 -73 -89 11
rect -29 -73 29 11
rect 89 -73 147 11
rect 207 -73 265 11
<< nmos >>
rect -207 -73 -147 11
rect -89 -73 -29 11
rect 29 -73 89 11
rect 147 -73 207 11
<< ndiff >>
rect -265 -1 -207 11
rect -265 -61 -253 -1
rect -219 -61 -207 -1
rect -265 -73 -207 -61
rect -147 -1 -89 11
rect -147 -61 -135 -1
rect -101 -61 -89 -1
rect -147 -73 -89 -61
rect -29 -1 29 11
rect -29 -61 -17 -1
rect 17 -61 29 -1
rect -29 -73 29 -61
rect 89 -1 147 11
rect 89 -61 101 -1
rect 135 -61 147 -1
rect 89 -73 147 -61
rect 207 -1 265 11
rect 207 -61 219 -1
rect 253 -61 265 -1
rect 207 -73 265 -61
<< ndiffc >>
rect -253 -61 -219 -1
rect -135 -61 -101 -1
rect -17 -61 17 -1
rect 101 -61 135 -1
rect 219 -61 253 -1
<< poly >>
rect -210 83 -144 99
rect -210 49 -194 83
rect -160 49 -144 83
rect -210 33 -144 49
rect -92 83 -26 99
rect -92 49 -76 83
rect -42 49 -26 83
rect -92 33 -26 49
rect 26 83 92 99
rect 26 49 42 83
rect 76 49 92 83
rect 26 33 92 49
rect 144 83 210 99
rect 144 49 160 83
rect 194 49 210 83
rect 144 33 210 49
rect -207 11 -147 33
rect -89 11 -29 33
rect 29 11 89 33
rect 147 11 207 33
rect -207 -99 -147 -73
rect -89 -99 -29 -73
rect 29 -99 89 -73
rect 147 -99 207 -73
<< polycont >>
rect -194 49 -160 83
rect -76 49 -42 83
rect 42 49 76 83
rect 160 49 194 83
<< locali >>
rect -210 49 -194 83
rect -160 49 -144 83
rect -92 49 -76 83
rect -42 49 -26 83
rect 26 49 42 83
rect 76 49 92 83
rect 144 49 160 83
rect 194 49 210 83
rect -253 -1 -219 15
rect -253 -77 -219 -61
rect -135 -1 -101 15
rect -135 -77 -101 -61
rect -17 -1 17 15
rect -17 -77 17 -61
rect 101 -1 135 15
rect 101 -77 135 -61
rect 219 -1 253 15
rect 219 -77 253 -61
<< viali >>
rect -253 -61 -219 -1
rect -135 -61 -101 -1
rect -17 -61 17 -1
rect 101 -61 135 -1
rect 219 -61 253 -1
<< metal1 >>
rect -259 -1 -213 11
rect -259 -61 -253 -1
rect -219 -61 -213 -1
rect -259 -73 -213 -61
rect -141 -1 -95 11
rect -141 -61 -135 -1
rect -101 -61 -95 -1
rect -141 -73 -95 -61
rect -23 -1 23 11
rect -23 -61 -17 -1
rect 17 -61 23 -1
rect -23 -73 23 -61
rect 95 -1 141 11
rect 95 -61 101 -1
rect 135 -61 141 -1
rect 95 -73 141 -61
rect 213 -1 259 11
rect 213 -61 219 -1
rect 253 -61 259 -1
rect 213 -73 259 -61
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.30 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
