magic
tech sky130B
magscale 1 2
timestamp 1736600368
<< nmos >>
rect -63 -100 -33 100
rect 33 -100 63 100
<< ndiff >>
rect -125 88 -63 100
rect -125 -88 -113 88
rect -79 -88 -63 88
rect -125 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 125 100
rect 63 -88 79 88
rect 113 -88 125 88
rect 63 -100 125 -88
<< ndiffc >>
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
<< poly >>
rect -63 100 -33 126
rect 33 100 63 126
rect -63 -126 -33 -100
rect 33 -126 63 -100
<< locali >>
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
<< viali >>
rect -17 -88 17 88
<< metal1 >>
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
