magic
tech sky130B
magscale 1 2
timestamp 1734781233
<< nwell >>
rect -902 1668 1312 1671
rect -902 1199 756 1668
<< locali >>
rect -845 816 -811 1333
rect -845 95 -811 782
rect -750 440 -550 1335
rect -750 406 -667 440
rect -633 406 -550 440
rect -750 189 -550 406
rect -407 325 -373 1333
rect -407 95 -373 291
rect -312 597 -112 1316
rect 242 699 276 733
rect 144 631 178 665
rect 347 631 381 665
rect -312 563 -233 597
rect -199 563 -112 597
rect 44 563 78 597
rect -312 189 -112 563
rect 347 495 381 529
rect 151 359 185 393
rect 44 291 78 325
<< viali >>
rect -845 782 -811 816
rect -667 406 -633 440
rect -407 291 -373 325
rect 302 767 336 801
rect 144 699 178 733
rect 46 631 80 665
rect -233 563 -199 597
rect 221 563 255 597
rect 46 495 80 529
rect 144 427 178 461
rect 304 359 338 393
rect 221 291 255 325
<< metal1 >>
rect -673 1668 1312 1671
rect -764 1623 1312 1668
rect -851 821 -801 822
rect -902 816 343 821
rect -902 782 -845 816
rect -811 813 343 816
rect -811 801 344 813
rect -811 782 302 801
rect -902 776 302 782
rect 296 767 302 776
rect 336 767 344 801
rect 135 733 187 745
rect 135 699 144 733
rect 178 699 187 733
rect 40 665 88 677
rect 40 631 46 665
rect 80 631 88 665
rect -245 602 -183 603
rect 40 602 88 631
rect -245 597 88 602
rect -245 563 -233 597
rect -199 563 88 597
rect -245 558 88 563
rect -245 557 -183 558
rect 40 529 88 558
rect 40 495 46 529
rect 80 495 88 529
rect 40 483 88 495
rect 135 461 187 699
rect 135 453 144 461
rect -688 440 144 453
rect -688 406 -667 440
rect -633 427 144 440
rect 178 427 187 461
rect -633 406 187 427
rect -688 396 187 406
rect 215 597 261 610
rect 215 563 221 597
rect 255 563 261 597
rect 215 336 261 563
rect 296 393 344 767
rect 296 359 304 393
rect 338 359 344 393
rect 296 342 344 359
rect -902 325 261 336
rect -902 291 -407 325
rect -373 291 221 325
rect 255 291 261 325
rect -902 283 261 291
rect 215 279 261 283
rect -754 -15 -554 61
rect -316 -15 -116 68
rect -754 -112 54 -15
use CG4  CG4_0
timestamp 1733177410
transform 1 0 28 0 1 746
box 1 -858 1284 922
use efepmos_W107-L15-F3  efepmos_W107-L15-F3_0 ~/Documents/Dersler/VLSI/vlsi_sky130b/design/mag/inv
timestamp 1734276197
transform 0 1 -219 -1 0 1462
box -209 -207 209 169
use efepmos_W107-L15-F3  efepmos_W107-L15-F3_1
timestamp 1734276197
transform 0 1 -657 -1 0 1462
box -209 -207 209 169
use sky130_fd_pr__nfet_01v8_5D68BK  sky130_fd_pr__nfet_01v8_5D68BK_0
timestamp 1734280111
transform 0 -1 -247 1 0 128
box -73 -157 73 157
use sky130_fd_pr__nfet_01v8_BQTKEQ  sky130_fd_pr__nfet_01v8_BQTKEQ_0
timestamp 1734280111
transform 0 1 -685 -1 0 128
box -73 -157 73 157
<< labels >>
rlabel metal1 -902 317 -902 317 3 B
port 1 e
rlabel metal1 -902 797 -902 797 3 A
port 2 e
<< end >>
