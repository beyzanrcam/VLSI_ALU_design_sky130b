magic
tech sky130B
magscale 1 2
timestamp 1735230776
<< nwell >>
rect -30 403 409 644
rect 0 366 376 403
rect 101 347 104 366
rect 223 290 343 338
rect 326 288 343 290
<< psubdiff >>
rect 100 -323 301 -296
rect 100 -374 126 -323
rect 279 -374 301 -323
rect 100 -401 301 -374
<< nsubdiff >>
rect 6 513 367 585
rect 6 458 65 513
rect 283 458 367 513
rect 6 439 367 458
<< psubdiffcont >>
rect 126 -374 279 -323
<< nsubdiffcont >>
rect 65 458 283 513
<< poly >>
rect 3 -124 70 -108
rect 3 -158 19 -124
rect 53 -126 70 -124
rect 53 -156 75 -126
rect 53 -158 70 -156
rect 3 -174 70 -158
<< polycont >>
rect 19 -158 53 -124
<< locali >>
rect 49 458 65 513
rect 283 458 299 513
rect 3 -124 53 339
rect 3 -158 19 -124
rect 3 -174 53 -158
rect 110 -374 126 -323
rect 279 -374 295 -323
<< viali >>
rect 124 469 209 503
rect 19 -158 53 -124
rect 173 -361 228 -327
<< metal1 >>
rect 100 503 277 511
rect 100 469 124 503
rect 209 469 277 503
rect 100 418 277 469
rect 100 366 314 418
rect 101 347 104 366
rect 0 80 53 338
rect 223 82 376 338
rect 0 -124 69 80
rect 100 -114 376 82
rect 0 -158 19 -124
rect 53 -158 69 -124
rect 0 -175 69 -158
rect 100 -250 300 -161
rect 328 -175 376 -114
rect 150 -327 256 -250
rect 150 -361 173 -327
rect 228 -361 256 -327
rect 150 -372 256 -361
use efepmos_W107-L15-F3  efepmos_W107-L15-F3_0
timestamp 1734789349
transform 0 1 207 -1 0 209
box -209 -207 209 169
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1734789349
transform 0 1 200 -1 0 -141
box -73 -126 73 126
<< labels >>
rlabel metal1 376 -31 376 -31 3 Y
port 3 e
rlabel metal1 0 -31 0 -31 7 A
port 2 e
rlabel metal1 144 418 144 418 1 VDD
port 1 n
rlabel metal1 201 -250 201 -250 5 VSS
port 4 s
<< end >>
