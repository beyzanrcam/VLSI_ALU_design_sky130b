magic
tech sky130B
magscale 1 2
timestamp 1735982637
<< nmos >>
rect -111 -300 -81 300
rect -15 -300 15 300
rect 81 -300 111 300
<< ndiff >>
rect -173 288 -111 300
rect -173 -288 -161 288
rect -127 -288 -111 288
rect -173 -300 -111 -288
rect -81 -300 -15 300
rect 15 -300 81 300
rect 111 288 173 300
rect 111 -288 127 288
rect 161 -288 173 288
rect 111 -300 173 -288
<< ndiffc >>
rect -161 -288 -127 288
rect 127 -288 161 288
<< poly >>
rect -111 300 -81 326
rect -15 300 15 326
rect 81 300 111 326
rect -111 -326 -81 -300
rect -15 -326 15 -300
rect 81 -326 111 -300
<< locali >>
rect -161 288 -127 304
rect -161 -304 -127 -288
rect 127 288 161 304
rect 127 -304 161 -288
<< viali >>
rect -161 -288 -127 288
rect 127 -288 161 288
<< metal1 >>
rect -167 288 -121 300
rect -167 -288 -161 288
rect -127 -288 -121 288
rect -167 -300 -121 -288
rect 121 288 167 300
rect 121 -288 127 288
rect 161 -288 167 288
rect 121 -300 167 -288
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3 l 0.150 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
