magic
tech sky130B
magscale 1 2
timestamp 1734125354
<< nwell >>
rect -205 1525 789 1745
<< psubdiff >>
rect 119 219 465 240
rect 119 101 144 219
rect 420 101 465 219
rect 119 79 465 101
<< nsubdiff >>
rect -162 1694 753 1709
rect -162 1600 -135 1694
rect 78 1600 753 1694
rect -162 1582 753 1600
<< psubdiffcont >>
rect 144 101 420 219
<< nsubdiffcont >>
rect -135 1600 78 1694
<< poly >>
rect 49 799 115 814
rect 49 765 65 799
rect 99 765 115 799
rect 49 748 115 765
rect 85 661 115 748
rect 277 718 307 814
rect 259 702 325 718
rect 259 668 275 702
rect 309 668 325 702
rect 85 631 211 661
rect 259 652 325 668
rect 181 522 211 631
rect 277 522 307 652
rect 469 590 499 814
rect 373 574 499 590
rect 373 540 389 574
rect 423 560 499 574
rect 423 540 439 560
rect 373 524 439 540
rect 373 522 403 524
<< polycont >>
rect 65 765 99 799
rect 275 668 309 702
rect 389 540 423 574
<< locali >>
rect -162 1694 753 1702
rect -162 1600 -135 1694
rect 78 1600 753 1694
rect -162 1590 753 1600
rect 49 765 65 799
rect 99 765 115 799
rect 259 668 275 702
rect 309 668 325 702
rect 373 540 389 574
rect 423 540 439 574
rect 131 228 165 292
rect 323 228 357 299
rect 119 219 465 228
rect 119 101 144 219
rect 420 101 465 219
rect 119 91 465 101
<< viali >>
rect -135 1600 78 1694
rect 65 765 99 799
rect 275 668 309 702
rect 389 540 423 574
<< metal1 >>
rect -147 1694 90 1701
rect -147 1600 -135 1694
rect 78 1600 90 1694
rect -147 1593 90 1600
rect -147 1517 57 1593
rect -163 1201 75 1517
rect 221 1201 651 1517
rect -67 875 363 1171
rect 509 875 747 1171
rect -310 799 115 814
rect -310 765 65 799
rect 99 765 115 799
rect -310 747 115 765
rect -310 702 325 718
rect -310 668 275 702
rect 309 668 325 702
rect -310 652 325 668
rect -310 574 439 590
rect -310 540 389 574
rect 423 540 439 574
rect -310 524 439 540
rect 595 496 747 875
rect 221 296 747 496
use sky130_fd_pr__nfet_01v8_XGU3BH  sky130_fd_pr__nfet_01v8_XGU3BH_0
timestamp 1734121473
transform 1 0 292 0 1 396
box -173 -126 173 126
use sky130_fd_pr__pfet_01v8_KAWEF3  sky130_fd_pr__pfet_01v8_KAWEF3_0
timestamp 1734121007
transform 1 0 292 0 1 1196
box -497 -421 497 421
<< labels >>
rlabel metal1 -310 778 -310 778 7 A
port 1 w
rlabel metal1 -310 684 -310 684 7 B
port 2 w
rlabel metal1 -310 559 -310 559 3 C
port 3 e
rlabel li 246 158 246 158 1 VSS
port 4 n
rlabel metal1 -29 1648 -29 1648 5 VDD
port 5 s
rlabel metal1 676 638 676 638 3 Y
port 6 e
<< end >>
