* SPICE3 file created from nand3_x.ext - technology: sky130B

.subckt nand3 A B C VSS VDD Y
X0 a_24_224.t0 A.t0 Y.t0 VSUBS sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=0.15
X1 a_120_224.t0 B.t0 a_24_224.t1 VSUBS sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=0.15
X2 Y.t1 A.t1 VDD.t3 w_n443_743.t3 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3 VDD.t1 B.t1 Y.t7 w_n443_743.t1 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4 a_n264_224.t1 C.t0 VSS.t1 VSUBS sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.465 ps=3.62 w=1.5 l=0.15
X5 a_n168_224.t0 B.t2 a_n264_224.t0 VSUBS sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=0.15
X6 VSS.t0 C.t1 a_120_224.t1 VSUBS sky130_fd_pr__nfet_01v8 ad=0.465 pd=3.62 as=0.2475 ps=1.83 w=1.5 l=0.15
X7 VDD.t2 A.t2 Y.t2 w_n443_743.t2 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X8 Y.t4 C.t2 VDD.t4 w_n443_743.t4 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X9 VDD.t5 C.t3 Y.t5 w_n443_743.t5 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X10 Y.t6 B.t3 VDD.t0 w_n443_743.t0 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X11 Y.t3 A.t3 a_n168_224.t1 VSUBS sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=0.15
R0 A.n1 A.t0 477.18
R1 A.n0 A.t2 347.187
R2 A.n0 A.t1 329.409
R3 A.n3 A.n1 321.334
R4 A.n3 A.t3 279.49
R5 A.n6 A.n5 161.54
R6 A.n6 A.n0 161.351
R7 A.n2 A.n0 79.1168
R8 A.n4 A.n2 54.8596
R9 A.n5 A.n1 27.7155
R10 A.n4 A.n3 24.1005
R11 A.n5 A.n4 20.4855
R12 A.n2 A.n1 14.4605
R13 A A.n6 0.660513
R14 Y.n2 Y.n0 184.571
R15 Y.n2 Y.n1 184.406
R16 Y.n4 Y.n3 184.406
R17 Y Y.n5 48.7873
R18 Y.n0 Y.t5 20.1899
R19 Y.n0 Y.t4 20.1899
R20 Y.n1 Y.t7 20.1899
R21 Y.n1 Y.t6 20.1899
R22 Y.n3 Y.t2 20.1899
R23 Y.n3 Y.t1 20.1899
R24 Y.n5 Y.t0 13.2005
R25 Y.n5 Y.t3 13.2005
R26 Y.n4 Y.n2 0.164884
R27 Y Y.n4 0.0876697
R28 a_24_224.t0 a_24_224.t1 26.4005
R29 B.n0 B.t1 763.168
R30 B.n0 B.t3 763.168
R31 B.n2 B.t0 469.151
R32 B.n1 B.t2 416.19
R33 B.n2 B.n1 78.4523
R34 B.n1 B.n0 33.8878
R35 B B.n2 0.478761
R36 a_120_224.t0 a_120_224.t1 26.4005
R37 VDD.n3 VDD.t4 204.595
R38 VDD.n0 VDD.t2 204.595
R39 VDD.n5 VDD.n4 184.406
R40 VDD.n2 VDD.n1 184.406
R41 VDD.n4 VDD.t0 20.1899
R42 VDD.n4 VDD.t5 20.1899
R43 VDD.n1 VDD.t3 20.1899
R44 VDD.n1 VDD.t1 20.1899
R45 VDD.n0 VDD 0.657041
R46 VDD.n2 VDD.n0 0.115885
R47 VDD.n5 VDD.n3 0.115885
R48 VDD VDD.n2 0.0581923
R49 VDD VDD.n5 0.0581923
R50 VDD.n3 VDD 0.0179279
R51 w_n443_743.n0 w_n443_743.t4 219.835
R52 w_n443_743.t3 w_n443_743.t2 188.43
R53 w_n443_743.t1 w_n443_743.t3 188.43
R54 w_n443_743.t0 w_n443_743.t1 188.43
R55 w_n443_743.t5 w_n443_743.t0 188.43
R56 w_n443_743.t4 w_n443_743.t5 188.43
R57 C.n0 C.t1 468.93
R58 C.t0 C.n0 461.748
R59 C.n1 C.t3 329.776
R60 C.n1 C.t2 314.452
R61 C.n2 C.t0 297.443
R62 C.n3 C.n2 161.3
R63 C.n2 C.n1 88.2596
R64 C.n3 C.n0 0.743461
R65 C C.n3 0.299413
R66 VSS VSS.t0 63.3304
R67 VSS.n0 VSS.t1 62.3706
R68 VSS.n1 VSS 0.533109
R69 VSS.n1 VSS 0.185283
R70 VSS VSS.n1 0.135115
R71 VSS.n1 VSS.n0 0.0238516
R72 VSS.n0 VSS 0.0238516
R73 a_n264_224.t0 a_n264_224.t1 26.4005
R74 a_n168_224.t0 a_n168_224.t1 26.4005
C0 C B 1.65857f
C1 A VDD 0.06113f
C2 VSS Y 0.533452f
C3 B Y 0.550409f
C4 C Y 0.078409f
C5 A VSS 0.001967f
C6 A B 0.894949f
C7 A C 0.040383f
C8 A Y 0.977481f
C9 VSS VDD 6.43e-19
C10 B VDD 0.028667f
C11 C VDD 0.027842f
C12 VDD Y 1.72252f
C13 B VSS 0.007622f
C14 C VSS 1.8223f
C15 VSS VSUBS 0.696274f
C16 Y VSUBS 0.312874f
C17 VDD VSUBS 0.419562f
C18 A VSUBS 0.442732f
C19 B VSUBS 0.408572f
C20 C VSUBS 0.616474f
.ends

