* NGSPICE file created from nor2_pex.ext - technology: sky130B

.subckt nor2 A B VSS VDD Y
X0 VSS.t1 B.t0 Y.t2 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X1 Y.t4 A.t0 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X2 a_224_100.t3 A.t1 a_128_100.t0 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3 a_320_100.t1 A.t2 a_224_100.t4 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4 VDD.t12 A.t3 a_320_100.t0 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X5 a_512_100.t0 A.t4 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X6 a_704_100.t0 B.t1 a_224_100.t0 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X7 Y.t3 B.t2 a_704_100.t1 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X8 a_224_100.t5 A.t5 a_512_100.t1 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X9 a_896_100.t1 B.t3 Y.t0 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X10 a_224_100.t2 B.t4 a_896_100.t0 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X11 a_1088_100.t0 B.t5 a_224_100.t1 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X12 Y.t1 B.t6 a_1088_100.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X13 a_128_100.t1 A.t6 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
R0 B.n0 B.t6 291.829
R1 B.n5 B.t0 239.393
R2 B.n4 B.t1 221.72
R3 B.n0 B.t5 221.72
R4 B.n1 B.t4 221.72
R5 B.n2 B.t3 221.72
R6 B.n3 B.t2 221.72
R7 B B.n5 162.72
R8 B.n5 B.n4 91.5805
R9 B.n1 B.n0 70.1096
R10 B.n2 B.n1 70.1096
R11 B.n3 B.n2 70.1096
R12 B.n4 B.n3 70.1096
R13 Y.n1 Y.t1 229.641
R14 Y.n1 Y.n0 198.476
R15 Y Y.n2 66.4022
R16 Y.n0 Y.t0 30.379
R17 Y.n0 Y.t3 30.379
R18 Y.n2 Y.t2 19.8005
R19 Y.n2 Y.t4 19.8005
R20 Y Y.n1 0.411207
R21 VSS.n1 VSS.n0 585
R22 VSS.n0 VSS.t2 439.139
R23 VSS.n0 VSS.t0 387.476
R24 VSS VSS.t1 157.137
R25 VSS VSS.t3 147.976
R26 VSS.n1 VSS 10.2907
R27 VSS VSS.n1 0.376971
R28 A.n0 A.t0 388.813
R29 A.n1 A.t6 291.829
R30 A.n4 A.t4 221.72
R31 A.n0 A.t5 221.72
R32 A.n3 A.t3 221.72
R33 A.n2 A.t2 221.72
R34 A.n1 A.t1 221.72
R35 A A.n4 162.357
R36 A.n4 A.n0 70.1096
R37 A.n4 A.n3 70.1096
R38 A.n3 A.n2 70.1096
R39 A.n2 A.n1 70.1096
R40 a_128_100.t0 a_128_100.t1 60.7575
R41 a_224_100.n2 a_224_100.n1 199.335
R42 a_224_100.n2 a_224_100.n0 199.335
R43 a_224_100.n3 a_224_100.n2 198.522
R44 a_224_100.n1 a_224_100.t4 30.379
R45 a_224_100.n1 a_224_100.t3 30.379
R46 a_224_100.n0 a_224_100.t1 30.379
R47 a_224_100.n0 a_224_100.t2 30.379
R48 a_224_100.t0 a_224_100.n3 30.379
R49 a_224_100.n3 a_224_100.t5 30.379
R50 VDD.n2 VDD.n0 311.053
R51 VDD VDD.t7 304.596
R52 VDD.n2 VDD.n1 185
R53 VDD.t1 VDD.t0 158.609
R54 VDD.t2 VDD.t1 158.609
R55 VDD.t3 VDD.t2 158.609
R56 VDD.t4 VDD.t3 158.609
R57 VDD.t5 VDD.t4 158.609
R58 VDD.t8 VDD.t5 158.609
R59 VDD.t9 VDD.t8 158.609
R60 VDD.t11 VDD.t9 158.609
R61 VDD.t13 VDD.t11 158.609
R62 VDD.t14 VDD.t13 158.609
R63 VDD.n1 VDD.t6 99.1309
R64 VDD.n1 VDD.t14 59.4788
R65 VDD.n0 VDD.t10 30.379
R66 VDD.n0 VDD.t12 30.379
R67 VDD VDD.n2 0.142722
R68 a_320_100.t0 a_320_100.t1 60.7575
R69 a_512_100.t0 a_512_100.t1 60.7575
R70 a_704_100.t0 a_704_100.t1 60.7575
R71 a_896_100.t0 a_896_100.t1 60.7575
R72 a_1088_100.t0 a_1088_100.t1 60.7575
C0 B A 0.636145f
C1 B Y 0.25959f
C2 VDD A 0.216493f
C3 VDD Y 0.050776f
C4 Y A 0.018087f
C5 B VDD 0.012428f
C6 Y VSS 0.698868f
C7 B VSS 0.602316f
C8 A VSS 0.428038f
C9 VDD VSS 2.46461f
.ends

