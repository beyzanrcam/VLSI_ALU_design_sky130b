magic
tech sky130B
magscale 1 2
timestamp 1733249760
<< nwell >>
rect -530 907 1099 3113
<< nmos >>
rect 75 53 135 453
rect 193 53 253 453
rect 311 53 371 453
rect 429 53 489 453
<< pmos >>
rect -397 1047 -337 2759
rect -279 1047 -219 2759
rect -161 1047 -101 2759
rect -43 1047 17 2759
rect 75 1047 135 2759
rect 193 1047 253 2759
rect 311 1047 371 2759
rect 429 1047 489 2759
rect 547 1047 607 2759
rect 665 1047 725 2759
rect 783 1047 843 2759
rect 901 1047 961 2759
<< ndiff >>
rect 17 441 75 453
rect 17 65 29 441
rect 63 65 75 441
rect 17 53 75 65
rect 135 441 193 453
rect 135 65 147 441
rect 181 65 193 441
rect 135 53 193 65
rect 253 441 311 453
rect 253 65 265 441
rect 299 65 311 441
rect 253 53 311 65
rect 371 441 429 453
rect 371 65 383 441
rect 417 65 429 441
rect 371 53 429 65
rect 489 441 547 453
rect 489 65 501 441
rect 535 65 547 441
rect 489 53 547 65
<< pdiff >>
rect -455 2747 -397 2759
rect -455 1059 -443 2747
rect -409 1059 -397 2747
rect -455 1047 -397 1059
rect -337 2747 -279 2759
rect -337 1059 -325 2747
rect -291 1059 -279 2747
rect -337 1047 -279 1059
rect -219 2747 -161 2759
rect -219 1059 -207 2747
rect -173 1059 -161 2747
rect -219 1047 -161 1059
rect -101 2747 -43 2759
rect -101 1059 -89 2747
rect -55 1059 -43 2747
rect -101 1047 -43 1059
rect 17 2747 75 2759
rect 17 1059 29 2747
rect 63 1059 75 2747
rect 17 1047 75 1059
rect 135 2747 193 2759
rect 135 1059 147 2747
rect 181 1059 193 2747
rect 135 1047 193 1059
rect 253 2747 311 2759
rect 253 1059 265 2747
rect 299 1059 311 2747
rect 253 1047 311 1059
rect 371 2747 429 2759
rect 371 1059 383 2747
rect 417 1059 429 2747
rect 371 1047 429 1059
rect 489 2747 547 2759
rect 489 1059 501 2747
rect 535 1059 547 2747
rect 489 1047 547 1059
rect 607 2747 665 2759
rect 607 1059 619 2747
rect 653 1059 665 2747
rect 607 1047 665 1059
rect 725 2747 783 2759
rect 725 1059 737 2747
rect 771 1059 783 2747
rect 725 1047 783 1059
rect 843 2747 901 2759
rect 843 1059 855 2747
rect 889 1059 901 2747
rect 843 1047 901 1059
rect 961 2747 1019 2759
rect 961 1059 973 2747
rect 1007 1059 1019 2747
rect 961 1047 1019 1059
<< ndiffc >>
rect 29 65 63 441
rect 147 65 181 441
rect 265 65 299 441
rect 383 65 417 441
rect 501 65 535 441
<< pdiffc >>
rect -443 1059 -409 2747
rect -325 1059 -291 2747
rect -207 1059 -173 2747
rect -89 1059 -55 2747
rect 29 1059 63 2747
rect 147 1059 181 2747
rect 265 1059 299 2747
rect 383 1059 417 2747
rect 501 1059 535 2747
rect 619 1059 653 2747
rect 737 1059 771 2747
rect 855 1059 889 2747
rect 973 1059 1007 2747
<< psubdiff >>
rect 17 -69 547 -1
rect 17 -182 81 -69
rect 467 -182 547 -69
rect 17 -258 547 -182
<< nsubdiff >>
rect -457 2941 -128 2989
rect -457 2868 -412 2941
rect -199 2868 -128 2941
rect -457 2813 -128 2868
<< psubdiffcont >>
rect 81 -182 467 -69
<< nsubdiffcont >>
rect -412 2868 -199 2941
<< poly >>
rect -397 2759 -337 2785
rect -279 2759 -219 2785
rect -161 2759 -101 2785
rect -43 2759 17 2785
rect 75 2759 135 2785
rect 193 2759 253 2785
rect 311 2759 371 2785
rect 429 2759 489 2785
rect 547 2759 607 2785
rect 665 2759 725 2785
rect 783 2759 843 2785
rect 901 2759 961 2785
rect -397 1016 -337 1047
rect -279 1016 -219 1047
rect -161 1016 -101 1047
rect -43 1016 17 1047
rect 75 1016 135 1047
rect 193 1016 253 1047
rect 311 1016 371 1047
rect 429 1016 489 1047
rect 547 1016 607 1047
rect 665 1016 725 1047
rect 783 1016 843 1047
rect 901 1016 961 1047
rect -400 1000 -334 1016
rect -400 966 -384 1000
rect -350 966 -334 1000
rect -400 950 -334 966
rect -282 1000 -216 1016
rect -282 966 -266 1000
rect -232 966 -216 1000
rect -282 950 -216 966
rect -164 1000 -98 1016
rect -164 966 -148 1000
rect -114 966 -98 1000
rect -164 950 -98 966
rect -46 1000 20 1016
rect -46 966 -30 1000
rect 4 966 20 1000
rect -46 950 20 966
rect 72 1000 138 1016
rect 72 966 88 1000
rect 122 966 138 1000
rect 72 950 138 966
rect 190 1000 256 1016
rect 190 966 206 1000
rect 240 966 256 1000
rect 190 950 256 966
rect 308 1000 374 1016
rect 308 966 324 1000
rect 358 966 374 1000
rect 308 950 374 966
rect 426 1000 492 1016
rect 426 966 442 1000
rect 476 966 492 1000
rect 426 950 492 966
rect 544 1000 610 1016
rect 544 966 560 1000
rect 594 966 610 1000
rect 544 950 610 966
rect 662 1000 728 1016
rect 662 966 678 1000
rect 712 966 728 1000
rect 662 950 728 966
rect 780 1000 846 1016
rect 780 966 796 1000
rect 830 966 846 1000
rect 780 950 846 966
rect 898 1000 964 1016
rect 898 966 914 1000
rect 948 966 964 1000
rect 898 950 964 966
rect 72 525 138 541
rect 72 491 88 525
rect 122 491 138 525
rect 72 475 138 491
rect 190 525 256 541
rect 190 491 206 525
rect 240 491 256 525
rect 190 475 256 491
rect 308 525 374 541
rect 308 491 324 525
rect 358 491 374 525
rect 308 475 374 491
rect 426 525 492 541
rect 426 491 442 525
rect 476 491 492 525
rect 426 475 492 491
rect 75 453 135 475
rect 193 453 253 475
rect 311 453 371 475
rect 429 453 489 475
rect 75 27 135 53
rect 193 27 253 53
rect 311 27 371 53
rect 429 27 489 53
<< polycont >>
rect -384 966 -350 1000
rect -266 966 -232 1000
rect -148 966 -114 1000
rect -30 966 4 1000
rect 88 966 122 1000
rect 206 966 240 1000
rect 324 966 358 1000
rect 442 966 476 1000
rect 560 966 594 1000
rect 678 966 712 1000
rect 796 966 830 1000
rect 914 966 948 1000
rect 88 491 122 525
rect 206 491 240 525
rect 324 491 358 525
rect 442 491 476 525
<< locali >>
rect -457 2941 -128 2953
rect -457 2868 -412 2941
rect -199 2868 -128 2941
rect -457 2851 -128 2868
rect -443 2747 -409 2763
rect -443 1043 -409 1059
rect -325 2747 -291 2763
rect -325 1043 -291 1059
rect -207 2747 -173 2763
rect -207 1043 -173 1059
rect -89 2747 -55 2763
rect -89 1043 -55 1059
rect 29 2747 63 2763
rect 29 1043 63 1059
rect 147 2747 181 2763
rect 147 1043 181 1059
rect 265 2747 299 2763
rect 265 1043 299 1059
rect 383 2747 417 2763
rect 383 1043 417 1059
rect 501 2747 535 2763
rect 501 1043 535 1059
rect 619 2747 653 2763
rect 619 1043 653 1059
rect 737 2747 771 2763
rect 737 1043 771 1059
rect 855 2747 889 2763
rect 855 1043 889 1059
rect 973 2747 1007 2763
rect 973 1043 1007 1059
rect -400 966 -384 1000
rect -350 966 -266 1000
rect -232 966 -148 1000
rect -114 966 -98 1000
rect -46 966 -30 1000
rect 4 966 88 1000
rect 122 966 206 1000
rect 240 966 256 1000
rect 308 966 324 1000
rect 358 966 442 1000
rect 476 966 560 1000
rect 594 966 610 1000
rect 662 966 678 1000
rect 712 966 796 1000
rect 830 966 914 1000
rect 948 966 964 1000
rect -282 556 -216 966
rect 72 849 138 966
rect 426 849 492 966
rect 72 792 256 849
rect 190 671 256 792
rect 190 617 195 671
rect 247 617 256 671
rect -282 551 138 556
rect -282 497 -273 551
rect -221 525 138 551
rect -221 497 88 525
rect -282 491 88 497
rect 122 491 138 525
rect 190 525 256 617
rect 190 491 206 525
rect 240 491 256 525
rect 308 792 492 849
rect 780 911 846 966
rect 780 863 788 911
rect 839 863 846 911
rect 308 789 374 792
rect 308 735 316 789
rect 368 735 374 789
rect 308 525 374 735
rect 780 556 846 863
rect 308 491 324 525
rect 358 491 374 525
rect 426 525 846 556
rect 426 491 442 525
rect 476 491 846 525
rect 29 441 63 457
rect 29 -1 63 65
rect 147 441 181 457
rect 147 49 181 65
rect 265 441 299 457
rect 265 -1 299 65
rect 383 441 417 457
rect 383 49 417 65
rect 501 441 535 457
rect 501 -1 535 65
rect 29 -69 535 -1
rect 29 -182 81 -69
rect 467 -182 535 -69
rect 29 -230 535 -182
<< viali >>
rect -412 2868 -199 2941
rect -443 1904 -409 2747
rect -325 1059 -291 1822
rect -207 1904 -173 2747
rect -89 1059 -55 1822
rect 29 1904 63 2747
rect 147 1059 181 1822
rect 265 1904 299 2747
rect 383 1059 417 1822
rect 501 1904 535 2747
rect 619 1059 653 1822
rect 737 1904 771 2747
rect 855 1059 889 1822
rect 973 1904 1007 2747
rect 195 617 247 671
rect -273 497 -221 551
rect 788 863 839 911
rect 316 735 368 789
rect 147 243 181 441
rect 383 243 417 441
<< metal1 >>
rect -450 2941 -167 2947
rect -450 2868 -412 2941
rect -199 2868 -167 2941
rect -450 2750 -167 2868
rect -449 2747 -167 2750
rect -449 1904 -443 2747
rect -409 1904 -207 2747
rect -173 1904 -167 2747
rect -449 1892 -167 1904
rect 23 2747 541 2759
rect 23 1904 29 2747
rect 63 1904 265 2747
rect 299 1904 501 2747
rect 535 1904 541 2747
rect 23 1892 541 1904
rect 730 2747 1013 2759
rect 730 1904 737 2747
rect 771 1904 973 2747
rect 1007 1904 1013 2747
rect 730 1892 1013 1904
rect -331 1822 187 1834
rect -331 1059 -325 1822
rect -291 1059 -89 1822
rect -55 1059 147 1822
rect 181 1059 187 1822
rect -331 1047 187 1059
rect 377 1822 895 1834
rect 377 1059 383 1822
rect 417 1059 619 1822
rect 653 1059 855 1822
rect 889 1059 895 1822
rect 377 1047 895 1059
rect -600 911 851 928
rect -600 863 788 911
rect 839 863 851 911
rect -600 846 851 863
rect -600 789 374 803
rect -600 735 316 789
rect 368 735 374 789
rect -600 715 374 735
rect -600 714 -485 715
rect -601 671 258 685
rect -601 617 195 671
rect 247 617 258 671
rect -601 597 258 617
rect -602 551 -198 568
rect -602 497 -273 551
rect -221 497 -198 551
rect -602 479 -198 497
rect 924 454 1013 1892
rect 369 453 1013 454
rect 141 441 1013 453
rect 141 243 147 441
rect 181 243 383 441
rect 417 243 1013 441
rect 141 231 1013 243
<< labels >>
flabel metal1 -590 488 -523 557 1 FreeSerif 320 0 0 0 A
port 1 n
flabel metal1 -590 608 -523 677 1 FreeSerif 320 0 0 0 B
port 2 n
flabel metal1 -589 723 -522 792 1 FreeSerif 320 0 0 0 C
port 3 n
flabel metal1 -589 853 -522 922 1 FreeSerif 320 0 0 0 D
port 4 n
flabel metal1 869 297 997 427 1 FreeSerif 320 0 0 0 Y
port 5 n
flabel nwell -369 2833 -242 2945 1 FreeSerif 320 0 0 0 VDD
port 6 n
flabel psubdiffcont 218 -182 345 -70 1 FreeSerif 320 0 0 0 VSS
port 7 n
<< end >>
