* NGSPICE file created from nor4_pex.ext - technology: sky130B

.subckt nor4 A B C D VSS VDD Y
X0 a_212_1047.t2 D.t0 Y.t6 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X1 Y.t1 C.t0 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2 VSS.t7 D.t1 Y.t3 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X3 a_n364_1047.t4 A.t0 VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=1.3268 ps=9.18 w=4.28 l=0.15
X4 a_n76_1047.t2 B.t0 a_n364_1047.t1 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X5 a_212_1047.t5 C.t1 a_n76_1047.t5 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X6 VSS.t1 B.t1 Y.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X7 VDD.t2 A.t1 a_n364_1047.t3 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X8 Y.t5 D.t2 a_212_1047.t1 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X9 a_n364_1047.t2 A.t2 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X10 a_212_1047.t3 C.t2 a_n76_1047.t4 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X11 Y.t4 D.t3 a_212_1047.t0 VDD.t7 sky130_fd_pr__pfet_01v8 ad=1.3268 pd=9.18 as=0.7062 ps=4.61 w=4.28 l=0.15
X12 a_n364_1047.t5 B.t2 a_n76_1047.t1 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X13 Y.t2 A.t3 VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X14 a_n76_1047.t0 B.t3 a_n364_1047.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X15 a_n76_1047.t3 C.t3 a_212_1047.t4 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
R0 D.n0 D.t3 883.668
R1 D.n1 D.t2 729.428
R2 D.n0 D.t0 729.428
R3 D.n2 D.t1 462.137
R4 D.n2 D.n1 437.014
R5 D D.n2 163.326
R6 D.n1 D.n0 154.24
R7 Y.n1 Y.t4 148.196
R8 Y.n1 Y.n0 140.636
R9 Y.n4 Y.n2 66.4372
R10 Y.n4 Y.n3 66.3172
R11 Y.n2 Y.t0 19.8005
R12 Y.n2 Y.t2 19.8005
R13 Y.n3 Y.t3 19.8005
R14 Y.n3 Y.t1 19.8005
R15 Y.n0 Y.t6 7.59513
R16 Y.n0 Y.t5 7.59513
R17 Y.n5 Y.n4 0.594743
R18 Y Y.n5 0.0800455
R19 Y.n5 Y.n1 0.0588942
R20 a_212_1047.n2 a_212_1047.n0 140.274
R21 a_212_1047.n3 a_212_1047.n2 140.274
R22 a_212_1047.n2 a_212_1047.n1 140.21
R23 a_212_1047.n0 a_212_1047.t4 7.59513
R24 a_212_1047.n0 a_212_1047.t5 7.59513
R25 a_212_1047.n1 a_212_1047.t1 7.59513
R26 a_212_1047.n1 a_212_1047.t3 7.59513
R27 a_212_1047.n3 a_212_1047.t0 7.59513
R28 a_212_1047.t2 a_212_1047.n3 7.59513
R29 VDD.n2 VDD.t13 192.784
R30 VDD.n1 VDD.t14 148.181
R31 VDD.n1 VDD.n0 140.65
R32 VDD.t9 VDD.t7 93.539
R33 VDD.t8 VDD.t9 93.539
R34 VDD.t10 VDD.t8 93.539
R35 VDD.t11 VDD.t10 93.539
R36 VDD.t12 VDD.t11 93.539
R37 VDD.t5 VDD.t12 93.539
R38 VDD.t6 VDD.t5 93.539
R39 VDD.t0 VDD.t6 93.539
R40 VDD.t3 VDD.t0 93.539
R41 VDD.t1 VDD.t3 93.539
R42 VDD.t13 VDD.t1 93.539
R43 VDD.n0 VDD.t4 7.59513
R44 VDD.n0 VDD.t2 7.59513
R45 VDD.n2 VDD.n1 0.0243095
R46 VDD VDD.n2 0.011082
R47 C.n0 C.t2 883.668
R48 C.n1 C.t1 740.381
R49 C.n0 C.t3 729.428
R50 C.n2 C.t0 700.508
R51 C C.n2 163.012
R52 C.n1 C.n0 72.3005
R53 C.n2 C.n1 16.7975
R54 VSS.t2 VSS.t6 483.849
R55 VSS.t0 VSS.t4 483.849
R56 VSS.n0 VSS.t0 282.245
R57 VSS.n0 VSS.t2 201.605
R58 VSS.n2 VSS.t5 150.175
R59 VSS.n3 VSS.t7 149.728
R60 VSS.n2 VSS.n1 119.644
R61 VSS.n3 VSS.n0 117.001
R62 VSS.n1 VSS.t3 19.8005
R63 VSS.n1 VSS.t1 19.8005
R64 VSS VSS.n3 0.952746
R65 VSS.n3 VSS.n2 0.447662
R66 A.n2 A.t3 960.788
R67 A.n0 A.t0 883.668
R68 A.n1 A.t2 740.381
R69 A.n0 A.t1 729.428
R70 A A.n2 162.053
R71 A.n1 A.n0 72.3005
R72 A.n2 A.n1 16.7975
R73 a_n364_1047.n2 a_n364_1047.n0 140.274
R74 a_n364_1047.n3 a_n364_1047.n2 140.274
R75 a_n364_1047.n2 a_n364_1047.n1 140.21
R76 a_n364_1047.n1 a_n364_1047.t0 7.59513
R77 a_n364_1047.n1 a_n364_1047.t2 7.59513
R78 a_n364_1047.n0 a_n364_1047.t1 7.59513
R79 a_n364_1047.n0 a_n364_1047.t5 7.59513
R80 a_n364_1047.n3 a_n364_1047.t3 7.59513
R81 a_n364_1047.t4 a_n364_1047.n3 7.59513
R82 B.n0 B.t3 883.668
R83 B.n1 B.t0 740.381
R84 B.n0 B.t2 729.428
R85 B.n2 B.t1 700.508
R86 B B.n2 162.65
R87 B.n1 B.n0 72.3005
R88 B.n2 B.n1 16.7975
R89 a_n76_1047.n2 a_n76_1047.n1 140.65
R90 a_n76_1047.n2 a_n76_1047.n0 140.65
R91 a_n76_1047.n3 a_n76_1047.n2 140.587
R92 a_n76_1047.n1 a_n76_1047.t1 7.59513
R93 a_n76_1047.n1 a_n76_1047.t0 7.59513
R94 a_n76_1047.n0 a_n76_1047.t4 7.59513
R95 a_n76_1047.n0 a_n76_1047.t3 7.59513
R96 a_n76_1047.n3 a_n76_1047.t5 7.59513
R97 a_n76_1047.t2 a_n76_1047.n3 7.59513
C0 D A 0.021716f
C1 Y B 0.012947f
C2 A VDD 0.471721f
C3 D VDD 0.001869f
C4 Y A 0.006044f
C5 Y D 0.571578f
C6 B C 1.18011f
C7 Y VDD 0.023399f
C8 A C 0.016869f
C9 D C 0.982733f
C10 C VDD 0.003911f
C11 A B 0.737801f
C12 D B 0.010577f
C13 Y C 0.043552f
C14 B VDD 0.01148f
C15 Y VSS 1.39979f
C16 D VSS 0.754994f
C17 C VSS 0.428671f
C18 B VSS 0.386825f
C19 A VSS 0.560463f
C20 VDD VSS 4.36813f
.ends

