magic
tech sky130B
magscale 1 2
timestamp 1733177410
<< nwell >>
rect 2 715 1284 922
<< psubdiff >>
rect 38 -777 1248 -761
rect 38 -843 100 -777
rect 1186 -843 1248 -777
rect 38 -858 1248 -843
<< nsubdiff >>
rect 38 869 1248 886
rect 38 803 100 869
rect 1186 803 1248 869
rect 38 787 1248 803
<< psubdiffcont >>
rect 100 -843 1186 -777
<< nsubdiffcont >>
rect 100 803 1186 869
<< locali >>
rect 38 869 1248 886
rect 38 803 100 869
rect 1186 803 1248 869
rect 38 787 1248 803
rect 1 21 308 55
rect 402 -13 596 24
rect 1 -47 596 -13
rect 690 -81 884 24
rect 1 -115 884 -81
rect 978 -149 1172 24
rect 1 -183 1172 -149
rect 1 -251 1172 -217
rect 1 -319 884 -285
rect 1 -387 596 -353
rect 1 -455 308 -421
rect 402 -428 596 -387
rect 690 -424 884 -319
rect 978 -424 1172 -251
rect 38 -777 1248 -761
rect 38 -843 100 -777
rect 1186 -843 1248 -777
rect 38 -858 1248 -843
<< viali >>
rect 100 803 1186 869
rect 50 559 84 661
rect 242 559 276 661
rect 434 557 468 659
rect 626 556 660 658
rect 818 556 852 658
rect 1010 556 1044 658
rect 1202 556 1236 658
rect 146 351 180 475
rect 338 351 372 475
rect 530 351 564 475
rect 722 351 756 475
rect 914 351 948 475
rect 1106 350 1140 474
rect 50 164 84 266
rect 242 164 276 266
rect 434 158 468 260
rect 626 141 660 243
rect 818 158 852 260
rect 1010 165 1044 267
rect 1202 165 1236 267
rect 50 -557 84 -523
rect 242 -557 276 -523
rect 434 -557 468 -523
rect 626 -557 660 -523
rect 818 -557 852 -523
rect 1010 -557 1044 -523
rect 1202 -557 1236 -523
rect 146 -661 180 -627
rect 338 -661 372 -627
rect 530 -662 564 -628
rect 722 -661 756 -627
rect 914 -661 948 -627
rect 1106 -661 1140 -627
rect 100 -843 1186 -777
<< metal1 >>
rect 2 869 1284 886
rect 2 803 100 869
rect 1186 803 1284 869
rect 2 787 1284 803
rect 38 661 292 787
rect 38 559 50 661
rect 84 559 242 661
rect 276 559 292 661
rect 38 538 292 559
rect 418 659 868 685
rect 418 557 434 659
rect 468 658 868 659
rect 468 557 626 658
rect 418 556 626 557
rect 660 556 818 658
rect 852 556 868 658
rect 418 538 868 556
rect 994 658 1248 787
rect 994 556 1010 658
rect 1044 556 1202 658
rect 1236 556 1248 658
rect 994 538 1248 556
rect 130 475 1156 500
rect 130 351 146 475
rect 180 351 338 475
rect 372 351 530 475
rect 564 351 722 475
rect 756 351 914 475
rect 948 474 1156 475
rect 948 351 1106 474
rect 130 350 1106 351
rect 1140 350 1156 474
rect 130 321 1156 350
rect 38 266 292 288
rect 38 164 50 266
rect 84 164 242 266
rect 276 164 292 266
rect 38 141 292 164
rect 418 260 867 277
rect 418 158 434 260
rect 468 243 818 260
rect 468 158 626 243
rect 418 141 626 158
rect 660 158 818 243
rect 852 158 867 260
rect 660 141 867 158
rect 994 267 1249 288
rect 994 165 1010 267
rect 1044 165 1202 267
rect 1236 165 1249 267
rect 994 141 1249 165
rect 610 -148 676 141
rect 610 -251 1284 -148
rect 610 -505 676 -251
rect 38 -523 292 -505
rect 38 -557 50 -523
rect 84 -557 242 -523
rect 276 -557 292 -523
rect 38 -573 292 -557
rect 418 -523 868 -505
rect 418 -557 434 -523
rect 468 -557 626 -523
rect 660 -557 818 -523
rect 852 -557 868 -523
rect 418 -573 868 -557
rect 994 -523 1248 -505
rect 994 -557 1010 -523
rect 1044 -557 1202 -523
rect 1236 -557 1248 -523
rect 994 -573 1248 -557
rect 38 -761 100 -573
rect 130 -627 580 -615
rect 130 -661 146 -627
rect 180 -661 338 -627
rect 372 -628 580 -627
rect 372 -661 530 -628
rect 130 -662 530 -661
rect 564 -662 580 -628
rect 130 -683 580 -662
rect 706 -627 1156 -615
rect 706 -661 722 -627
rect 756 -661 914 -627
rect 948 -661 1106 -627
rect 1140 -661 1156 -627
rect 706 -683 1156 -661
rect 1186 -761 1248 -573
rect 2 -777 1284 -761
rect 2 -843 100 -777
rect 1186 -843 1284 -777
rect 2 -858 1284 -843
use nfet_3_200_15  nfet_3_200_15_0
timestamp 1733177410
transform -1 0 211 0 -1 -592
box -173 -170 173 91
use nfet_3_200_15  nfet_3_200_15_1
timestamp 1733177410
transform -1 0 499 0 -1 -592
box -173 -170 173 91
use nfet_3_200_15  nfet_3_200_15_2
timestamp 1733177410
transform -1 0 1075 0 -1 -592
box -173 -170 173 91
use nfet_3_200_15  nfet_3_200_15_3
timestamp 1733177410
transform -1 0 787 0 -1 -592
box -173 -170 173 91
use pfet_3_825_15  pfet_3_825_15_0
timestamp 1733177410
transform 1 0 211 0 1 404
box -209 -398 209 311
use pfet_3_825_15  pfet_3_825_15_1
timestamp 1733177410
transform 1 0 499 0 1 404
box -209 -398 209 311
use pfet_3_825_15  pfet_3_825_15_2
timestamp 1733177410
transform 1 0 787 0 1 404
box -209 -398 209 311
use pfet_3_825_15  pfet_3_825_15_3
timestamp 1733177410
transform 1 0 1075 0 1 404
box -209 -398 209 311
<< labels >>
flabel metal1 602 818 756 870 1 FreeSerif 80 0 0 0 VDD
port 1 n
flabel metal1 592 -835 746 -783 1 FreeSerif 80 0 0 0 VSS
port 2 n
flabel locali 13 -243 34 -223 1 FreeSerif 80 0 0 0 N1
port 3 n
flabel locali 12 -311 33 -291 1 FreeSerif 80 0 0 0 N2
port 4 n
flabel locali 12 -380 33 -360 1 FreeSerif 80 0 0 0 N3
port 5 n
flabel locali 12 -448 33 -428 1 FreeSerif 80 0 0 0 N4
port 6 n
flabel locali 13 -177 34 -157 1 FreeSerif 80 0 0 0 P1
port 7 n
flabel locali 13 -108 34 -88 1 FreeSerif 80 0 0 0 P2
port 8 n
flabel locali 13 -39 34 -19 1 FreeSerif 80 0 0 0 P3
port 9 n
flabel locali 13 28 34 48 1 FreeSerif 80 0 0 0 P4
port 10 n
flabel metal1 1183 -228 1257 -164 1 FreeSerif 80 0 0 0 OUT
port 11 n
<< end >>
