magic
tech sky130B
magscale 1 2
timestamp 1736595726
<< nwell >>
rect -1843 2757 -550 3243
rect 493 2589 3416 2590
rect 493 2013 3470 2589
rect -298 -329 3416 -328
rect -298 -904 3462 -329
<< metal1 >>
rect -1740 3153 -719 3243
rect -669 3140 -43 3243
rect -1842 3095 -1773 3101
rect -1842 3020 -1773 3026
rect -1402 3095 -1333 3101
rect -1402 3020 -1333 3026
rect -962 3095 -893 3101
rect -962 3020 -893 3026
rect -1841 2505 -1772 2751
rect -1842 2446 -1772 2505
rect -1499 2530 -1430 2751
rect -1666 2474 -1615 2493
rect -1841 2330 -1772 2446
rect -1697 2444 -1577 2474
rect -1697 2392 -1666 2444
rect -1614 2392 -1577 2444
rect -1499 2440 -1430 2461
rect -1697 2361 -1577 2392
rect -1841 2261 -1499 2330
rect -1841 2249 -1772 2261
rect -1568 -332 -1499 2261
rect -1402 1997 -1333 2751
rect -1059 2528 -990 2590
rect -1228 2499 -1177 2512
rect -1257 2463 -1137 2499
rect -1257 2411 -1228 2463
rect -1176 2411 -1137 2463
rect -1059 2446 -990 2459
rect -1257 2386 -1137 2411
rect -1408 1991 -1327 1997
rect -1408 1922 -1402 1991
rect -1333 1988 -1327 1991
rect -1333 1922 -1315 1988
rect -1408 1916 -1327 1922
rect -1402 -238 -1333 1916
rect -962 1856 -893 2587
rect -619 2537 -550 2597
rect -146 2542 -43 3140
rect 4460 2543 5009 2544
rect 5350 2543 5692 2544
rect -788 2490 -737 2521
rect -620 2506 -550 2537
rect -820 2472 -700 2490
rect -820 2420 -788 2472
rect -736 2420 -700 2472
rect -820 2377 -700 2420
rect -962 1781 -893 1787
rect -620 1894 -551 2506
rect -262 2301 3380 2542
rect 4294 2301 5692 2543
rect -294 2077 -242 2083
rect -294 2019 -242 2025
rect 3369 2016 3510 2082
rect 4460 2077 5692 2301
rect -303 1983 -232 1988
rect 705 1984 715 1986
rect -303 1931 -287 1983
rect -235 1931 -232 1983
rect 709 1932 715 1984
rect -303 1922 -232 1931
rect 705 1927 715 1932
rect 1018 1901 1099 1918
rect -620 1828 -231 1894
rect -79 1828 -73 1894
rect -7 1828 -1 1894
rect 1018 1849 1024 1901
rect 1093 1849 1099 1901
rect 1589 1888 1642 1894
rect 1589 1829 1642 1835
rect 4460 1874 4789 2077
rect 5010 1874 5692 2077
rect -620 -135 -551 1828
rect -294 1533 -228 1800
rect -294 1461 -228 1467
rect 650 1429 716 1800
rect 1586 1735 1652 1800
rect 2398 1778 2464 1784
rect 2398 1706 2464 1712
rect 1586 1651 1652 1669
rect 2517 1639 2583 1800
rect 2517 1567 2583 1573
rect 1418 1530 1484 1536
rect 1418 1458 1484 1464
rect 650 1357 716 1363
rect 4460 1359 5692 1874
rect 472 1276 538 1282
rect 4460 1272 4503 1359
rect 5326 1218 5692 1359
rect 472 1204 538 1210
rect 5632 1181 5676 1218
rect -179 753 -173 931
rect 5 753 11 931
rect 4303 733 4415 830
rect 5753 659 5823 742
rect 453 483 519 489
rect 4833 420 4952 421
rect 453 411 519 417
rect 1589 327 1655 333
rect -298 107 -232 113
rect -298 -116 -232 41
rect 1437 73 1503 79
rect 1437 1 1503 7
rect 650 -14 716 -8
rect 650 -116 716 -80
rect 1589 -116 1655 261
rect 4674 301 4833 417
rect 4952 301 5073 417
rect 5521 379 5721 435
rect 5521 357 5560 379
rect 4674 227 5073 301
rect 5523 260 5560 357
rect 5679 357 5721 379
rect 5679 260 5713 357
rect 2517 205 2583 211
rect 5523 202 5713 260
rect 2407 -21 2473 -13
rect 2407 -91 2473 -85
rect 2517 -115 2583 139
rect -626 -204 -620 -135
rect -551 -144 -545 -135
rect -551 -204 -232 -144
rect -620 -210 -232 -204
rect 3482 -210 3488 -144
rect 3554 -210 3559 -144
rect -1402 -302 -1334 -238
rect -1401 -304 -1334 -302
rect -1268 -304 -232 -238
rect -1568 -398 -459 -332
rect -393 -398 -229 -332
rect 3373 -398 3510 -332
rect -1568 -408 -1499 -398
rect -263 -857 3379 -616
rect 4483 -617 4747 -606
rect 4258 -859 4494 -617
rect 4736 -859 4747 -617
rect 4483 -870 4747 -859
<< via1 >>
rect -1842 3026 -1773 3095
rect -1402 3026 -1333 3095
rect -962 3026 -893 3095
rect -1666 2392 -1614 2444
rect -1499 2461 -1430 2530
rect -1228 2411 -1176 2463
rect -1059 2459 -990 2528
rect -1402 1922 -1333 1991
rect -788 2420 -736 2472
rect -962 1787 -893 1856
rect -294 2025 -242 2077
rect 669 2024 722 2076
rect 1602 2025 1655 2077
rect 2533 2025 2586 2077
rect -287 1931 -235 1983
rect 657 1932 709 1984
rect 1600 1927 1652 1979
rect 2535 1927 2587 1979
rect -73 1828 -7 1894
rect 1024 1849 1093 1901
rect 1589 1835 1642 1888
rect 2862 1863 2931 1932
rect 3460 1922 3526 1988
rect 3458 1828 3524 1894
rect 4789 1874 5010 2077
rect -294 1467 -228 1533
rect 1586 1669 1652 1735
rect 2398 1712 2464 1778
rect 3450 1734 3515 1800
rect 2517 1573 2583 1639
rect 1418 1464 1484 1530
rect 650 1363 716 1429
rect 472 1210 538 1276
rect -173 753 5 931
rect 762 753 940 931
rect 1698 753 1876 931
rect 2629 754 2806 931
rect 3556 753 3734 931
rect 453 417 519 483
rect 1589 261 1655 327
rect -298 41 -232 107
rect 1437 7 1503 73
rect 650 -80 716 -14
rect 4833 301 4952 420
rect 5560 260 5679 379
rect 2517 139 2583 205
rect 2407 -85 2473 -21
rect 3450 -116 3516 -50
rect -620 -204 -551 -135
rect 1001 -215 1065 -151
rect 1593 -210 1659 -144
rect 2864 -211 2924 -151
rect 3488 -210 3554 -144
rect -1334 -304 -1268 -238
rect 679 -299 731 -247
rect 1601 -304 1667 -238
rect 2537 -303 2603 -237
rect 3459 -304 3525 -238
rect -459 -398 -393 -332
rect 663 -393 728 -341
rect 1592 -393 1657 -341
rect 2551 -393 2616 -341
rect 4494 -859 4736 -617
<< metal2 >>
rect -1842 3095 -1773 3344
rect -1402 3095 -1333 3344
rect -962 3095 -893 3344
rect -1848 3026 -1842 3095
rect -1773 3026 -1767 3095
rect -1408 3026 -1402 3095
rect -1333 3026 -1327 3095
rect -968 3026 -962 3095
rect -893 3026 -887 3095
rect -1499 2641 -287 2710
rect -1499 2530 -1430 2641
rect -1697 2446 -1577 2474
rect -1499 2455 -1430 2461
rect -1242 2465 -1164 2475
rect -1697 2390 -1668 2446
rect -1612 2390 -1577 2446
rect -1242 2409 -1230 2465
rect -1174 2409 -1164 2465
rect -1065 2459 -1059 2528
rect -990 2459 -984 2528
rect -820 2474 -700 2490
rect -1242 2394 -1164 2409
rect -1697 2361 -1577 2390
rect -1059 2363 -990 2459
rect -820 2418 -790 2474
rect -734 2418 -700 2474
rect -820 2377 -700 2418
rect -1059 2295 -990 2304
rect -356 2086 -287 2641
rect -356 2077 2740 2086
rect -356 2025 -294 2077
rect -242 2076 1602 2077
rect -242 2025 669 2076
rect -356 2024 669 2025
rect 722 2025 1602 2076
rect 1655 2025 2533 2077
rect 2586 2025 2740 2077
rect 722 2024 2740 2025
rect -356 2017 2740 2024
rect 4787 2085 5031 2096
rect 4787 2077 4798 2085
rect -1408 1991 -1327 1997
rect -1408 1922 -1402 1991
rect -1333 1986 -1327 1991
rect -1333 1984 715 1986
rect -1333 1983 657 1984
rect -1333 1931 -287 1983
rect -235 1932 657 1983
rect 709 1932 715 1984
rect -235 1931 715 1932
rect -1333 1927 715 1931
rect 782 1936 1514 1989
rect 2529 1983 2600 1985
rect -1333 1922 -1327 1927
rect -1408 1916 -1327 1922
rect -79 1894 -7 1899
rect 782 1894 848 1936
rect -971 1856 -884 1865
rect -971 1787 -962 1856
rect -893 1787 -884 1856
rect -79 1828 -73 1894
rect -7 1828 848 1894
rect 1024 1901 1093 1907
rect 1461 1888 1514 1936
rect 1589 1925 1598 1981
rect 1654 1925 1663 1981
rect 2523 1927 2535 1983
rect 2591 1927 2600 1983
rect 2856 1932 2936 1938
rect 2529 1921 2593 1927
rect 1141 1856 1200 1860
rect 1093 1851 1205 1856
rect 1093 1849 1141 1851
rect -79 1822 -7 1828
rect 1024 1792 1141 1849
rect 1200 1792 1205 1851
rect 1461 1835 1589 1888
rect 1642 1835 1648 1888
rect 2856 1863 2862 1932
rect 2931 1863 2936 1932
rect 2856 1856 2936 1863
rect 3005 1922 3460 1988
rect 3526 1922 3532 1988
rect 1024 1787 1205 1792
rect -971 1778 -884 1787
rect 1141 1783 1200 1787
rect 3005 1778 3071 1922
rect -1668 1669 1586 1735
rect 1652 1669 1658 1735
rect 2392 1712 2398 1778
rect 2464 1712 3071 1778
rect 3136 1828 3458 1894
rect 3524 1828 3530 1894
rect 4787 1874 4789 2077
rect 4787 1863 4798 1874
rect 5020 1863 5041 2085
rect 4787 1852 5031 1863
rect -1668 1573 2517 1639
rect 2583 1573 2589 1639
rect -1668 1467 -294 1533
rect -228 1467 -222 1533
rect 3136 1530 3202 1828
rect 1412 1464 1418 1530
rect 1484 1464 3202 1530
rect 3259 1734 3450 1800
rect 3515 1734 3521 1800
rect -1668 1363 650 1429
rect 716 1363 722 1429
rect 3259 1276 3325 1734
rect 466 1210 472 1276
rect 538 1210 3325 1276
rect -244 931 3807 1003
rect -244 753 -173 931
rect 5 753 762 931
rect 940 753 1698 931
rect 1876 754 2629 931
rect 2806 754 3556 931
rect 1876 753 3556 754
rect 3734 753 3807 931
rect -244 682 3807 753
rect 5014 512 5421 624
rect 4728 508 5421 512
rect 447 417 453 483
rect 519 417 2721 483
rect -1668 261 1589 327
rect 1655 261 1661 327
rect 2655 205 2721 417
rect 4728 482 5642 508
rect 4728 420 5786 482
rect 4728 301 4833 420
rect 4952 379 5786 420
rect 4952 301 5560 379
rect 4728 260 5560 301
rect 5679 260 5786 379
rect -1668 139 2517 205
rect 2583 139 2589 205
rect 2655 139 3304 205
rect 4728 195 5786 260
rect -1668 41 -298 107
rect -232 41 -226 107
rect 1431 7 1437 73
rect 1503 7 3188 73
rect -1668 -80 650 -14
rect 716 -80 722 -14
rect 2401 -85 2407 -21
rect 2473 -85 3053 -21
rect 996 -116 1070 -110
rect -620 -135 -551 -129
rect -551 -188 806 -149
rect 996 -151 1005 -116
rect 1061 -151 1070 -116
rect 996 -180 1001 -151
rect -620 -210 -551 -204
rect -1334 -238 -1268 -232
rect -1268 -247 739 -238
rect -1268 -299 679 -247
rect 731 -299 739 -247
rect 767 -257 806 -188
rect 1065 -180 1070 -151
rect 1215 -210 1593 -144
rect 1659 -210 1665 -144
rect 2864 -151 2924 -145
rect 2857 -209 2864 -153
rect 2924 -209 2931 -153
rect 1001 -221 1065 -215
rect 1216 -257 1255 -210
rect 2864 -217 2924 -211
rect 767 -296 1255 -257
rect -1268 -304 739 -299
rect 1592 -304 1601 -238
rect 1667 -304 1676 -238
rect 2531 -303 2537 -237
rect 2603 -303 2612 -237
rect 2987 -238 3053 -85
rect 3122 -144 3188 7
rect 3238 -50 3304 139
rect 5067 36 5786 195
rect 5396 3 5786 36
rect 3238 -116 3450 -50
rect 3516 -116 3522 -50
rect 3122 -210 3488 -144
rect 3554 -210 3563 -144
rect 2987 -304 3459 -238
rect 3525 -304 3531 -238
rect -1334 -310 -1268 -304
rect -466 -398 -459 -332
rect -393 -341 2662 -332
rect -393 -393 663 -341
rect 728 -393 1592 -341
rect 1657 -393 2551 -341
rect 2616 -393 2662 -341
rect -393 -398 2662 -393
rect -459 -404 -393 -398
rect 4483 -617 4747 -606
rect 4483 -859 4494 -617
rect 4736 -859 4747 -617
rect 4483 -870 4747 -859
<< via2 >>
rect -1668 2444 -1612 2446
rect -1668 2392 -1666 2444
rect -1666 2392 -1614 2444
rect -1614 2392 -1612 2444
rect -1668 2390 -1612 2392
rect -1230 2463 -1174 2465
rect -1230 2411 -1228 2463
rect -1228 2411 -1176 2463
rect -1176 2411 -1174 2463
rect -1230 2409 -1174 2411
rect -790 2472 -734 2474
rect -790 2420 -788 2472
rect -788 2420 -736 2472
rect -736 2420 -734 2472
rect -790 2418 -734 2420
rect -1059 2304 -990 2363
rect 4798 2077 5020 2085
rect -962 1787 -893 1856
rect 1598 1979 1654 1981
rect 1598 1927 1600 1979
rect 1600 1927 1652 1979
rect 1652 1927 1654 1979
rect 1598 1925 1654 1927
rect 2535 1979 2591 1983
rect 2535 1927 2587 1979
rect 2587 1927 2591 1979
rect 1141 1792 1200 1851
rect 2867 1868 2926 1927
rect 4798 1874 5010 2077
rect 5010 1874 5020 2077
rect 4798 1863 5020 1874
rect -173 753 5 931
rect 762 753 940 931
rect 1698 753 1876 931
rect 2629 754 2806 931
rect 3556 753 3734 931
rect 4833 301 4952 420
rect 5560 260 5679 379
rect 1005 -151 1061 -116
rect 1005 -172 1061 -151
rect 2866 -209 2922 -153
rect 1601 -304 1667 -242
rect 2547 -303 2603 -242
rect 4494 -859 4736 -617
<< metal3 >>
rect -1693 2451 -1573 2475
rect -1693 2385 -1673 2451
rect -1607 2385 -1573 2451
rect -1693 2362 -1573 2385
rect -1256 2470 -1136 2496
rect -1256 2404 -1235 2470
rect -1169 2404 -1136 2470
rect -1256 2383 -1136 2404
rect -821 2479 -701 2497
rect -821 2413 -795 2479
rect -729 2413 -701 2479
rect -821 2384 -701 2413
rect -1064 2363 -985 2368
rect -1064 2304 -1059 2363
rect -990 2304 -985 2363
rect -1064 2299 -985 2304
rect -1058 2040 -989 2299
rect 4787 2090 5031 2096
rect -1109 1990 -988 2040
rect -1109 1983 2602 1990
rect -1109 1981 2535 1983
rect -1109 1971 1598 1981
rect -1101 1925 1598 1971
rect 1654 1927 2535 1981
rect 2591 1927 2602 1983
rect 1654 1925 2602 1927
rect -1101 1922 2602 1925
rect -1101 -237 -1035 1922
rect -827 1920 2602 1922
rect 2862 1927 2931 1932
rect 2862 1868 2867 1927
rect 2926 1868 2931 1927
rect -967 1856 -888 1861
rect 2862 1856 2931 1868
rect -967 1787 -962 1856
rect -893 1851 2931 1856
rect 4787 1858 4793 2090
rect 5025 1858 5031 2090
rect 4787 1852 5031 1858
rect -893 1792 1141 1851
rect 1200 1792 2931 1851
rect -893 1787 2931 1792
rect -967 1782 -888 1787
rect -967 1709 -893 1782
rect -960 -117 -900 1709
rect -244 936 3807 1003
rect -244 748 -178 936
rect 10 748 757 936
rect 945 748 1693 936
rect 1881 749 2624 936
rect 2811 749 3551 936
rect 1881 748 3551 749
rect 3739 748 3807 936
rect -244 682 3807 748
rect 5014 512 5421 624
rect 4728 508 5421 512
rect 4728 482 5642 508
rect 4728 425 5786 482
rect 4728 296 4828 425
rect 4957 384 5786 425
rect 4957 296 5555 384
rect 4728 255 5555 296
rect 5684 255 5786 384
rect 4728 195 5786 255
rect 5067 36 5786 195
rect 5396 3 5786 36
rect 998 -116 1071 -111
rect 998 -117 1005 -116
rect -960 -172 1005 -117
rect 1061 -117 1071 -116
rect 1061 -148 2924 -117
rect 1061 -153 2927 -148
rect 1061 -172 2866 -153
rect -960 -177 2866 -172
rect 2861 -209 2866 -177
rect 2922 -209 2927 -153
rect 2861 -214 2927 -209
rect -1101 -242 2621 -237
rect -1101 -303 1601 -242
rect 1596 -304 1601 -303
rect 1667 -303 2547 -242
rect 2603 -303 2621 -242
rect 1667 -304 1672 -303
rect 1596 -309 1672 -304
rect 2542 -308 2621 -303
rect 4483 -612 4747 -606
rect 4483 -864 4489 -612
rect 4741 -864 4747 -612
rect 4483 -870 4747 -864
<< via3 >>
rect -1673 2446 -1607 2451
rect -1673 2390 -1668 2446
rect -1668 2390 -1612 2446
rect -1612 2390 -1607 2446
rect -1673 2385 -1607 2390
rect -1235 2465 -1169 2470
rect -1235 2409 -1230 2465
rect -1230 2409 -1174 2465
rect -1174 2409 -1169 2465
rect -1235 2404 -1169 2409
rect -795 2474 -729 2479
rect -795 2418 -790 2474
rect -790 2418 -734 2474
rect -734 2418 -729 2474
rect -795 2413 -729 2418
rect 4793 2085 5025 2090
rect 4793 1863 4798 2085
rect 4798 1863 5020 2085
rect 5020 1863 5025 2085
rect 4793 1858 5025 1863
rect -178 931 10 936
rect -178 753 -173 931
rect -173 753 5 931
rect 5 753 10 931
rect -178 748 10 753
rect 757 931 945 936
rect 757 753 762 931
rect 762 753 940 931
rect 940 753 945 931
rect 757 748 945 753
rect 1693 931 1881 936
rect 1693 753 1698 931
rect 1698 753 1876 931
rect 1876 753 1881 931
rect 1693 748 1881 753
rect 2624 931 2811 936
rect 2624 754 2629 931
rect 2629 754 2806 931
rect 2806 754 2811 931
rect 2624 749 2811 754
rect 3551 931 3739 936
rect 3551 753 3556 931
rect 3556 753 3734 931
rect 3734 753 3739 931
rect 3551 748 3739 753
rect 4828 420 4957 425
rect 4828 301 4833 420
rect 4833 301 4952 420
rect 4952 301 4957 420
rect 4828 296 4957 301
rect 5555 379 5684 384
rect 5555 260 5560 379
rect 5560 260 5679 379
rect 5679 260 5684 379
rect 5555 255 5684 260
rect 4489 -617 4741 -612
rect 4489 -859 4494 -617
rect 4494 -859 4736 -617
rect 4736 -859 4741 -617
rect 4489 -864 4741 -859
<< metal4 >>
rect -1819 2582 -577 2615
rect -1819 2573 -898 2582
rect -1819 2554 -1338 2573
rect -1819 2282 -1776 2554
rect -1504 2301 -1338 2554
rect -1066 2310 -898 2573
rect -626 2310 -577 2582
rect -1066 2301 -577 2310
rect -1504 2282 -577 2301
rect -1819 2248 -577 2282
rect 4721 2090 5050 2252
rect 4721 2072 4793 2090
rect 3917 1858 4793 2072
rect 5025 1858 5050 2090
rect 3917 1743 5050 1858
rect -244 979 3807 1003
rect -244 978 2582 979
rect -244 706 -220 978
rect 52 706 715 978
rect 987 706 1651 978
rect 1923 707 2582 978
rect 2854 978 3807 979
rect 2854 707 3509 978
rect 1923 706 3509 707
rect 3781 706 3807 978
rect -244 682 3807 706
rect 3917 50 4246 1743
rect 5014 512 5421 624
rect 4728 508 5421 512
rect 4728 497 5642 508
rect 4728 225 4757 497
rect 5029 482 5642 497
rect 5029 456 5786 482
rect 5029 225 5484 456
rect 4728 195 5484 225
rect 5067 184 5484 195
rect 5756 184 5786 456
rect 3917 -279 4489 50
rect 5067 36 5786 184
rect 5396 3 5786 36
rect 4160 -543 4489 -279
rect 4160 -612 4759 -543
rect 4160 -864 4489 -612
rect 4741 -864 4759 -612
rect 4160 -912 4759 -864
<< via4 >>
rect -1776 2451 -1504 2554
rect -1776 2385 -1673 2451
rect -1673 2385 -1607 2451
rect -1607 2385 -1504 2451
rect -1776 2282 -1504 2385
rect -1338 2470 -1066 2573
rect -1338 2404 -1235 2470
rect -1235 2404 -1169 2470
rect -1169 2404 -1066 2470
rect -1338 2301 -1066 2404
rect -898 2479 -626 2582
rect -898 2413 -795 2479
rect -795 2413 -729 2479
rect -729 2413 -626 2479
rect -898 2310 -626 2413
rect -220 936 52 978
rect -220 748 -178 936
rect -178 748 10 936
rect 10 748 52 936
rect -220 706 52 748
rect 715 936 987 978
rect 715 748 757 936
rect 757 748 945 936
rect 945 748 987 936
rect 715 706 987 748
rect 1651 936 1923 978
rect 1651 748 1693 936
rect 1693 748 1881 936
rect 1881 748 1923 936
rect 1651 706 1923 748
rect 2582 936 2854 979
rect 2582 749 2624 936
rect 2624 749 2811 936
rect 2811 749 2854 936
rect 2582 707 2854 749
rect 3509 936 3781 978
rect 3509 748 3551 936
rect 3551 748 3739 936
rect 3739 748 3781 936
rect 3509 706 3781 748
rect 4757 425 5029 497
rect 4757 296 4828 425
rect 4828 296 4957 425
rect 4957 296 5029 425
rect 4757 225 5029 296
rect 5484 384 5756 456
rect 5484 255 5555 384
rect 5555 255 5684 384
rect 5684 255 5756 384
rect 5484 184 5756 255
<< metal5 >>
rect -1819 2582 -268 2615
rect -1819 2573 -898 2582
rect -1819 2554 -1338 2573
rect -1819 2282 -1776 2554
rect -1504 2301 -1338 2554
rect -1066 2310 -898 2573
rect -626 2310 -268 2582
rect -1066 2301 -268 2310
rect -1504 2282 -268 2301
rect -1819 2248 -268 2282
rect -954 1040 -268 2248
rect -954 1008 3856 1040
rect -954 1005 4503 1008
rect -954 979 4746 1005
rect -954 978 2582 979
rect -954 706 -220 978
rect 52 706 715 978
rect 987 706 1651 978
rect 1923 707 2582 978
rect 2854 978 4746 979
rect 2854 707 3509 978
rect 1923 706 3509 707
rect 3781 835 4746 978
rect 3781 706 5059 835
rect -954 681 5059 706
rect -954 637 3856 681
rect -954 635 -268 637
rect 4402 624 5059 681
rect 4402 508 5421 624
rect 4402 497 5642 508
rect 4402 225 4757 497
rect 5029 482 5642 497
rect 5029 456 5786 482
rect 5029 225 5484 456
rect 4402 195 5484 225
rect 5067 184 5484 195
rect 5756 184 5786 456
rect 5067 36 5786 184
rect 5396 3 5786 36
use inv  inv_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/inv
timestamp 1735843251
transform 1 0 5423 0 1 739
box 0 -311 412 486
use inv  inv_1
timestamp 1735843251
transform 1 0 -1402 0 1 2757
box 0 -311 412 486
use inv  inv_2
timestamp 1735843251
transform 1 0 -962 0 1 2757
box 0 -311 412 486
use inv  inv_3
timestamp 1735843251
transform 1 0 -1842 0 1 2757
box 0 -311 412 486
use NAND4F  NAND4F_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NAND/NAND4
timestamp 1736096163
transform 1 0 2507 0 1 2017
box 10 -1175 909 571
use NAND4F  NAND4F_1
timestamp 1736096163
transform 1 0 1576 0 -1 -333
box 10 -1175 909 571
use NAND4F  NAND4F_2
timestamp 1736096163
transform 1 0 640 0 1 2017
box 10 -1175 909 571
use NAND4F  NAND4F_3
timestamp 1736096163
transform 1 0 1576 0 1 2017
box 10 -1175 909 571
use NAND4F  NAND4F_4
timestamp 1736096163
transform 1 0 -308 0 1 2017
box 10 -1175 909 571
use NAND4F  NAND4F_5
timestamp 1736096163
transform 1 0 -308 0 -1 -333
box 10 -1175 909 571
use NAND4F  NAND4F_6
timestamp 1736096163
transform 1 0 640 0 -1 -333
box 10 -1175 909 571
use NAND4F  NAND4F_7
timestamp 1736096163
transform 1 0 2507 0 -1 -332
box 10 -1175 909 571
use NAND4F  NAND4F_8
timestamp 1736096163
transform 1 0 3434 0 1 2017
box 10 -1175 909 571
use NAND4F  NAND4F_9
timestamp 1736096163
transform 1 0 3434 0 -1 -333
box 10 -1175 909 571
use nor2  nor2_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NOR/NOR2
timestamp 1736020690
transform 1 0 4337 0 1 866
box 0 -480 1090 580
<< labels >>
flabel space 1872 2601 1938 2667 0 FreeSans 1600 0 0 0 000
flabel space 2838 2594 2845 2596 0 FreeSans 1600 0 0 0 001
flabel space -18 2600 -15 2600 0 FreeSans 1600 0 0 0 010
flabel space 870 2605 1194 2664 0 FreeSans 1600 0 0 0 011
flabel space 1811 -1111 2237 -1054 0 FreeSans 1600 0 0 0 100
flabel space 2793 -1133 3071 -974 0 FreeSans 1600 0 0 0 101
flabel space -101 -1184 217 -1009 0 FreeSans 1600 0 0 0 110
flabel space 904 -1162 1222 -987 0 FreeSans 1600 0 0 0 111
flabel metal2 -1660 1674 -1608 1726 0 FreeSans 160 0 0 0 A0
port 1 nsew
flabel metal2 -1657 1579 -1605 1631 0 FreeSans 160 0 0 0 A1
port 2 nsew
flabel metal2 -1654 1473 -1602 1525 0 FreeSans 160 0 0 0 A2
port 3 nsew
flabel metal2 -1659 1367 -1607 1419 0 FreeSans 160 0 0 0 A3
port 4 nsew
flabel metal2 -1656 269 -1604 321 0 FreeSans 160 0 0 0 A4
port 5 nsew
flabel metal2 -1654 145 -1602 197 0 FreeSans 160 0 0 0 A5
port 6 nsew
flabel metal2 -1657 49 -1605 101 0 FreeSans 160 0 0 0 A6
port 7 nsew
flabel metal2 -1661 -72 -1609 -20 0 FreeSans 160 0 0 0 A7
port 8 nsew
flabel metal1 4977 2313 5029 2365 0 FreeSans 160 0 0 0 VDD
port 10 nsew
flabel metal1 5759 673 5811 725 0 FreeSans 160 0 0 0 Y
port 12 nsew
flabel metal5 5555 26 5607 78 0 FreeSans 160 0 0 0 VSS
port 9 nsew
flabel metal2 -952 3297 -907 3336 0 FreeSans 160 0 0 0 SEL0
port 13 nsew
flabel metal2 -1393 3288 -1348 3327 0 FreeSans 160 0 0 0 SEL1
port 14 nsew
flabel metal2 -1831 3288 -1786 3327 0 FreeSans 160 0 0 0 SEL2
port 16 nsew
<< end >>
