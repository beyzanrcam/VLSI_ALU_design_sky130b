magic
tech sky130B
magscale 1 2
timestamp 1736600368
<< nwell >>
rect 0 459 1090 580
rect 1 396 1090 459
rect 42 350 486 396
<< psubdiff >>
rect 420 -401 670 -384
rect 420 -462 446 -401
rect 645 -462 670 -401
rect 420 -480 670 -462
<< nsubdiff >>
rect 46 502 466 544
rect 46 451 74 502
rect 431 451 466 502
rect 46 413 466 451
<< psubdiffcont >>
rect 446 -462 645 -401
<< nsubdiffcont >>
rect 74 451 431 502
<< poly >>
rect 417 19 433 53
rect 467 19 483 53
rect 482 -114 512 6
rect 578 -36 608 6
rect 560 -52 626 -36
rect 560 -86 576 -52
rect 610 -86 626 -52
rect 560 -102 626 -86
rect 578 -113 608 -102
<< polycont >>
rect 433 19 467 53
rect 576 -86 610 -52
<< locali >>
rect 46 502 466 522
rect 46 451 74 502
rect 431 451 466 502
rect 46 432 466 451
rect 48 363 82 432
rect 240 363 274 432
rect 432 363 466 432
rect 417 19 433 53
rect 467 19 483 53
rect 560 -86 576 -52
rect 610 -86 626 -52
rect 432 -390 466 -334
rect 624 -390 658 -334
rect 420 -401 670 -390
rect 420 -462 446 -401
rect 645 -462 670 -401
rect 420 -474 670 -462
<< viali >>
rect 74 451 431 502
rect 433 19 467 53
rect 576 -86 610 -52
rect 446 -462 645 -401
<< metal1 >>
rect 62 502 443 510
rect 62 451 74 502
rect 431 451 443 502
rect 62 444 443 451
rect 184 245 522 359
rect 568 245 714 359
rect 760 245 906 359
rect 88 103 426 217
rect 664 103 1090 217
rect 0 53 526 69
rect 0 19 433 53
rect 467 19 526 53
rect 0 3 526 19
rect 0 -52 626 -36
rect 0 -86 576 -52
rect 610 -86 626 -52
rect 0 -102 626 -86
rect 965 -136 1090 103
rect 568 -334 1090 -136
rect 568 -335 1088 -334
rect 568 -336 1037 -335
rect 434 -401 657 -394
rect 434 -462 446 -401
rect 645 -462 657 -401
rect 434 -468 657 -462
use sky130_fd_pr__nfet_01v8_LZEQWH  sky130_fd_pr__nfet_01v8_LZEQWH_0
timestamp 1736600368
transform -1 0 545 0 -1 -230
box -125 -126 125 126
use sky130_fd_pr__pfet_01v8_UFBY79  sky130_fd_pr__pfet_01v8_UFBY79_0
timestamp 1736600368
transform 1 0 545 0 1 231
box -545 -228 545 228
<< labels >>
flabel metal1 7 10 84 62 1 FreeSerif 320 0 0 0 A
port 1 e
rlabel metal1 253 510 253 510 5 VDD
port 4 s
flabel metal1 8 -96 85 -44 1 FreeSerif 320 0 0 0 B
port 2 e
flabel metal1 1012 -102 1089 -50 1 FreeSerif 320 0 0 0 Y
port 5 e
rlabel metal1 549 -468 549 -468 5 VSS
port 3 s
<< end >>
