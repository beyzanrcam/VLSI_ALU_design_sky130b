** sch_path: /home/erhangok/Documents/Dersler/VLSI/vlsi_sky130b/design/xschem/INV/buffer.sch
**.subckt buffer A Y
*.ipin A
*.opin Y
x1 A VSS VDD net1 inv
x2 net1 VSS VDD Y inv
**.ends

* expanding   symbol:  inv.sym # of pins=2
** sym_path: /home/erhangok/Documents/Dersler/VLSI/vlsi_sky130b/design/xschem/INV/inv.sym
** sch_path: /home/erhangok/Documents/Dersler/VLSI/vlsi_sky130b/design/xschem/INV/inv.sch
.subckt inv A VSS VDD Y
*.ipin A
*.opin Y
XM1 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.21 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
