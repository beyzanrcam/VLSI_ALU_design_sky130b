** sch_path: /foss/designs/HW3/mux_tb.sch
**.subckt mux_tb OUTPUT VDD VSS
*.opin OUTPUT
*.iopin VDD
*.iopin VSS
V1 VDD GND 1.2
V2 VSS GND 0
V4 INPUT GND pulse(0,1.2,0.01u,0 ,0,0.01u,0.02u)
x2 OUTPUT VSS VDD net1 inv
x3 OUTPUT VSS VDD net1 inv
x4 OUTPUT VSS VDD net1 inv
x5 OUTPUT VSS VDD net1 inv
x6 INPUT VSS VDD net2 inv
x1 INPUT net2 VDD VSS OUTPUT VSS VDD XOR2
**** begin user architecture code

** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt_mm




.control
set color0 = white

save all
tran 0.1p 0.03u
plot INPUT OUTPUT title 'a'

meas tran t_input when V(INPUT)=0.6 RISE=1
meas tran t_output when V(OUTPUT)=0.6 FALL=1
let tpdr = (t_output - t_input) * 1e9
echo tpdr (ns) is:
print tpdr
meas tran t_input when V(INPUT)=0.6 FALL=1
meas tran t_output when V(OUTPUT)=0.6 RISE=1
let tpdf = (t_output - t_input) * 1e9
echo tpdf (ns) is:
print tpdf
let tpd = (tpdf + tpdr)/2
echo tpd (ns) is:
print tpd

let p_n_ratio = @m.x1.xm1.msky130_fd_pr__pfet_01v8[w]/@m.x1.xm2.msky130_fd_pr__nfet_01v8[w]
print p_n_ratio
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/xschem/INV/inv.sym # of pins=2
** sym_path: /foss/designs/xschem/INV/inv.sym
** sch_path: /foss/designs/xschem/INV/inv.sch
.subckt inv A VSS VDD Y
*.ipin A
*.opin Y
XM1 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.21 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/xschem/XOR/XOR2.sym # of pins=5
** sym_path: /foss/designs/xschem/XOR/XOR2.sym
** sch_path: /foss/designs/xschem/XOR/XOR2.sch
.subckt XOR2 A !A B !B OUT VSS VDD
*.ipin A
*.ipin !A
*.ipin B
*.ipin !B
*.opin OUT
x1 VDD VSS B A !A !B B !B !A A OUT cg4_pex
.ends


* expanding   symbol:  /foss/designs/xschem/CG4/cg4.sym # of pins=9
** sym_path: /foss/designs/xschem/CG4/cg4.sym
** sch_path: /foss/designs/xschem/CG4/cg4.sch
.subckt cg4 P3 P4 P2 P1 OUT N2 N1 N4 N3 VSS VDD
*.ipin P3
*.ipin P1
*.ipin N1
*.ipin N3
*.ipin P4
*.ipin P2
*.ipin N2
*.ipin N4
*.opin OUT
XM1 OUT N1 net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT N2 net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 N3 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 N4 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 OUT P1 net3 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=8.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 OUT P2 net3 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=8.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net3 P3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=8.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net3 P4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=8.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.subckt cg4_pex VDD VSS N1 N2 N3 N4 P1 P2 P3 P4 OUT
X0 a_130_n657# N3 OUT VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 OUT N2 a_706_n657# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 a_706_n657# N1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3 a_130_n657# N4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.2015 ps=1.92 w=0.65 l=0.15
X4 OUT N3 a_130_n657# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_130_129# P4 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X6 OUT P3 a_130_129# VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X7 VDD P4 a_130_129# VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X8 OUT P3 a_130_129# VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X9 a_130_129# P3 OUT VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X10 a_130_129# P2 OUT VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X11 OUT P2 a_130_129# VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X12 VDD P1 a_130_129# VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X13 a_706_n657# N2 OUT VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X14 a_130_129# P2 OUT VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X15 a_130_129# P1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X16 VSS N1 a_706_n657# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X17 VDD P1 a_130_129# VDD sky130_fd_pr__pfet_01v8 ad=0.8525 pd=6.12 as=0.45375 ps=3.08 w=2.75 l=0.15
X18 a_130_129# P4 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.8525 ps=6.12 w=2.75 l=0.15
X19 a_706_n657# N2 OUT VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X20 VSS N1 a_706_n657# VSS sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X21 a_130_n657# N4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X22 OUT N3 a_130_n657# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X23 VSS N4 a_130_n657# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
C0 a_130_n657# N3 0.045367f
C1 P1 P4 0.001451f
C2 a_130_129# N3 3.96e-19
C3 P3 OUT 0.133874f
C4 VDD N2 9.08e-19
C5 P2 N3 5.53e-19
C6 a_130_n657# VDD 6.93e-19
C7 a_130_129# VDD 1.64045f
C8 VDD P2 0.222988f
C9 N1 P3 8.72e-19
C10 N1 OUT 0.150265f
C11 N4 N3 0.180425f
C12 P3 N2 5.72e-19
C13 OUT N2 0.202994f
C14 N3 P4 4.01e-19
C15 a_130_n657# P3 6.59e-19
C16 a_130_n657# OUT 0.226686f
C17 P1 N3 8.38e-19
C18 a_130_129# P3 0.067886f
C19 a_130_129# OUT 1.61616f
C20 VDD N4 0.001147f
C21 VDD P4 0.336708f
C22 P2 P3 0.314455f
C23 P2 OUT 0.223063f
C24 VDD P1 0.326566f
C25 N1 N2 0.441185f
C26 N3 a_706_n657# 0.00109f
C27 a_130_n657# N1 4.66e-19
C28 a_130_129# N1 2.25e-19
C29 P2 N1 8.72e-19
C30 a_130_n657# N2 0.001764f
C31 a_130_129# N2 1.8e-19
C32 N4 P3 3.9e-19
C33 N4 OUT 0.003557f
C34 a_130_n657# a_130_129# 0.006295f
C35 P4 P3 0.186817f
C36 P4 OUT 0.007562f
C37 P2 N2 0.011231f
C38 P1 P3 0.001451f
C39 P1 OUT 0.155969f
C40 a_130_n657# P2 2.59e-19
C41 a_130_129# P2 0.05964f
C42 VDD N3 7.36e-19
C43 N4 N1 0.001382f
C44 OUT a_706_n657# 0.241167f
C45 N1 P4 8.72e-19
C46 P1 N1 0.495583f
C47 N4 N2 0.00251f
C48 P4 N2 5.72e-19
C49 a_130_n657# N4 0.036845f
C50 N1 a_706_n657# 0.04127f
C51 P1 N2 8.38e-19
C52 a_130_129# N4 2.33e-19
C53 a_130_n657# P4 4.39e-19
C54 a_130_129# P4 0.053985f
C55 a_130_n657# P1 3.4e-19
C56 a_130_129# P1 0.059392f
C57 N3 P3 0.009408f
C58 N4 P2 5.53e-19
C59 N3 OUT 0.114666f
C60 P2 P4 0.002654f
C61 N2 a_706_n657# 0.037344f
C62 P1 P2 0.445343f
C63 a_130_n657# a_706_n657# 0.017f
C64 VDD P3 0.228019f
C65 VDD OUT 0.403107f
C66 N3 N1 0.001382f
C67 N4 P4 0.008118f
C68 VDD N1 0.00121f
C69 N3 N2 0.310116f
C70 N4 P1 8.38e-19
C71 N1 VSS 0.599227f
C72 N2 VSS 0.415774f
C73 N3 VSS 0.380342f
C74 N4 VSS 0.447347f
C75 OUT VSS 0.484091f
C76 P1 VSS 0.303348f
C77 P2 VSS 0.201325f
C78 P3 VSS 0.158256f
C79 P4 VSS 0.145307f
C80 VDD VSS 4.37553f
C81 a_706_n657# VSS 0.506348f
C82 a_130_n657# VSS 0.506356f
C83 a_130_129# VSS 0.227118f
.ends



.GLOBAL GND
.end
