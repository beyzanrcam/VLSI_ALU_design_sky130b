magic
tech sky130A
magscale 1 2
timestamp 1733177410
<< nwell >>
rect -209 -398 209 311
<< pmos >>
rect -111 -275 -81 275
rect -15 -275 15 275
rect 81 -275 111 275
<< pdiff >>
rect -173 263 -111 275
rect -173 -263 -161 263
rect -127 -263 -111 263
rect -173 -275 -111 -263
rect -81 263 -15 275
rect -81 -263 -65 263
rect -31 -263 -15 263
rect -81 -275 -15 -263
rect 15 263 81 275
rect 15 -263 31 263
rect 65 -263 81 263
rect 15 -275 81 -263
rect 111 263 173 275
rect 111 -263 127 263
rect 161 -263 173 263
rect 111 -275 173 -263
<< pdiffc >>
rect -161 -263 -127 263
rect -65 -263 -31 263
rect 31 -263 65 263
rect 127 -263 161 263
<< poly >>
rect -111 275 -81 306
rect -15 275 15 306
rect 81 275 111 306
rect -111 -306 -81 -275
rect -15 -306 15 -275
rect 81 -306 111 -275
rect -111 -330 111 -306
rect -111 -364 -81 -330
rect 81 -364 111 -330
rect -111 -388 111 -364
<< polycont >>
rect -81 -364 81 -330
<< locali >>
rect -161 263 -127 279
rect -161 -279 -127 -263
rect -65 263 -31 279
rect -65 -279 -31 -263
rect 31 263 65 279
rect 31 -279 65 -263
rect 127 263 161 279
rect 127 -279 161 -263
rect -97 -330 97 -314
rect -97 -364 -81 -330
rect 81 -364 97 -330
rect -97 -380 97 -364
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.75 l 0.15 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
