magic
tech sky130B
magscale 1 2
timestamp 1735575029
<< nwell >>
rect 309 632 519 736
rect -5 328 -3 334
rect 407 250 419 632
rect 785 345 786 347
<< metal1 >>
rect 305 824 475 852
rect 305 720 339 824
rect 443 736 475 824
rect 443 720 519 736
rect 305 691 519 720
rect 309 632 519 691
rect 309 616 474 632
rect -5 328 -3 334
rect 407 75 419 588
rect 785 345 786 347
rect 295 -61 519 36
rect 335 -192 432 -61
rect 335 -295 432 -289
<< via1 >>
rect 339 720 443 824
rect 335 -289 432 -192
<< metal2 >>
rect 330 720 339 824
rect 443 720 452 824
rect 326 -289 335 -192
rect 432 -289 441 -192
<< via2 >>
rect 339 720 443 824
rect 335 -289 432 -192
<< metal3 >>
rect 334 829 448 835
rect 334 709 448 715
rect 330 -187 437 -181
rect 330 -300 437 -294
<< via3 >>
rect 334 824 448 829
rect 334 720 339 824
rect 339 720 443 824
rect 443 720 448 824
rect 334 715 448 720
rect 330 -192 437 -187
rect 330 -289 335 -192
rect 335 -289 432 -192
rect 432 -289 437 -192
rect 330 -294 437 -289
<< metal4 >>
rect 333 829 449 830
rect 333 715 334 829
rect 448 715 449 829
rect 333 714 449 715
<< via4 >>
rect 248 -187 520 -104
rect 248 -294 330 -187
rect 330 -294 437 -187
rect 437 -294 520 -187
rect 248 -376 520 -294
<< metal5 >>
rect 175 -104 619 -61
rect 175 -376 248 -104
rect 520 -376 619 -104
rect 175 -422 619 -376
use inv  inv_0
timestamp 1735572721
transform 1 0 -5 0 1 250
box 0 -311 412 486
use inv  inv_1
timestamp 1735572721
transform 1 0 374 0 1 250
box 0 -311 412 486
<< labels >>
rlabel metal1 -5 331 -5 331 3 A
port 1 e
rlabel metal1 433 -61 433 -61 5 VSS
port 2 s
rlabel metal1 786 346 786 346 3 Y
port 4 e
rlabel metal1 446 736 446 736 5 VDD
port 3 s
<< end >>
