magic
tech sky130B
magscale 1 2
timestamp 1736008794
<< error_p >>
rect -545 -228 545 228
<< nwell >>
rect -545 -228 545 228
<< pmos >>
rect -447 -128 -417 128
rect -351 -128 -321 128
rect -255 -128 -225 128
rect -159 -128 -129 128
rect -63 -128 -33 128
rect 33 -128 63 128
rect 129 -128 159 128
rect 225 -128 255 128
rect 321 -128 351 128
rect 417 -128 447 128
<< pdiff >>
rect -509 116 -447 128
rect -509 -116 -497 116
rect -463 -116 -447 116
rect -509 -128 -447 -116
rect -417 116 -351 128
rect -417 -116 -401 116
rect -367 -116 -351 116
rect -417 -128 -351 -116
rect -321 116 -255 128
rect -321 -116 -305 116
rect -271 -116 -255 116
rect -321 -128 -255 -116
rect -225 116 -159 128
rect -225 -116 -209 116
rect -175 -116 -159 116
rect -225 -128 -159 -116
rect -129 116 -63 128
rect -129 -116 -113 116
rect -79 -116 -63 116
rect -129 -128 -63 -116
rect -33 116 33 128
rect -33 -116 -17 116
rect 17 -116 33 116
rect -33 -128 33 -116
rect 63 116 129 128
rect 63 -116 79 116
rect 113 -116 129 116
rect 63 -128 129 -116
rect 159 116 225 128
rect 159 -116 175 116
rect 209 -116 225 116
rect 159 -128 225 -116
rect 255 116 321 128
rect 255 -116 271 116
rect 305 -116 321 116
rect 255 -128 321 -116
rect 351 116 417 128
rect 351 -116 367 116
rect 401 -116 417 116
rect 351 -128 417 -116
rect 447 116 509 128
rect 447 -116 463 116
rect 497 -116 509 116
rect 447 -128 509 -116
<< pdiffc >>
rect -497 -116 -463 116
rect -401 -116 -367 116
rect -305 -116 -271 116
rect -209 -116 -175 116
rect -113 -116 -79 116
rect -17 -116 17 116
rect 79 -116 113 116
rect 175 -116 209 116
rect 271 -116 305 116
rect 367 -116 401 116
rect 463 -116 497 116
<< poly >>
rect -447 128 -417 154
rect -351 128 -321 154
rect -255 128 -225 154
rect -159 128 -129 154
rect -63 128 -33 154
rect 33 128 63 154
rect 129 128 159 154
rect 225 128 255 154
rect 321 128 351 154
rect 417 128 447 154
rect -447 -154 -417 -128
rect -351 -154 -321 -128
rect -255 -154 -225 -128
rect -159 -154 -129 -128
rect -63 -154 -33 -128
rect -447 -225 -33 -154
rect 33 -154 63 -128
rect 129 -154 159 -128
rect 225 -154 255 -128
rect 321 -154 351 -128
rect 417 -154 447 -128
rect 33 -225 447 -154
<< locali >>
rect -497 116 -463 132
rect -497 -132 -463 -116
rect -401 116 -367 132
rect -401 -132 -367 -116
rect -305 116 -271 132
rect -305 -132 -271 -116
rect -209 116 -175 132
rect -209 -132 -175 -116
rect -113 116 -79 132
rect -113 -132 -79 -116
rect -17 116 17 132
rect -17 -132 17 -116
rect 79 116 113 132
rect 79 -132 113 -116
rect 175 116 209 132
rect 175 -132 209 -116
rect 271 116 305 132
rect 271 -132 305 -116
rect 367 116 401 132
rect 367 -132 401 -116
rect 463 116 497 132
rect 463 -132 497 -116
<< viali >>
rect -497 -116 -463 -26
rect -401 26 -367 116
rect -305 -116 -271 -26
rect -209 26 -175 116
rect -113 -116 -79 -26
rect -17 26 17 116
rect 79 -116 113 -26
rect 175 26 209 116
rect 271 -116 305 -26
rect 367 26 401 116
rect 463 -116 497 -26
<< metal1 >>
rect -407 116 -361 128
rect -407 26 -401 116
rect -367 26 -361 116
rect -407 14 -361 26
rect -215 116 -169 128
rect -215 26 -209 116
rect -175 26 -169 116
rect -215 14 -169 26
rect -23 116 23 128
rect -23 26 -17 116
rect 17 26 23 116
rect -23 14 23 26
rect 169 116 215 128
rect 169 26 175 116
rect 209 26 215 116
rect 169 14 215 26
rect 361 116 407 128
rect 361 26 367 116
rect 401 26 407 116
rect 361 14 407 26
rect -503 -26 -457 -14
rect -503 -116 -497 -26
rect -463 -116 -457 -26
rect -503 -128 -457 -116
rect -311 -26 -265 -14
rect -311 -116 -305 -26
rect -271 -116 -265 -26
rect -311 -128 -265 -116
rect -119 -26 -73 -14
rect -119 -116 -113 -26
rect -79 -116 -73 -26
rect -119 -128 -73 -116
rect 73 -26 119 -14
rect 73 -116 79 -26
rect 113 -116 119 -26
rect 73 -128 119 -116
rect 265 -26 311 -14
rect 265 -116 271 -26
rect 305 -116 311 -26
rect 265 -128 311 -116
rect 457 -26 503 -14
rect 457 -116 463 -26
rect 497 -116 503 -26
rect 457 -128 503 -116
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.284 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
