magic
tech sky130B
magscale 1 2
timestamp 1733167563
<< nwell >>
rect -443 743 263 1227
<< nmos >>
rect -294 224 -264 524
rect -198 224 -168 524
rect -102 224 -72 524
rect -6 224 24 524
rect 90 224 120 524
rect 186 224 216 524
<< pmos >>
rect -345 843 -315 1165
rect -249 843 -219 1165
rect -153 843 -123 1165
rect -57 843 -27 1165
rect 39 843 69 1165
rect 135 843 165 1165
<< ndiff >>
rect -356 512 -294 524
rect -356 236 -344 512
rect -310 236 -294 512
rect -356 224 -294 236
rect -264 224 -198 524
rect -168 224 -102 524
rect -72 512 -6 524
rect -72 236 -56 512
rect -22 236 -6 512
rect -72 224 -6 236
rect 24 224 90 524
rect 120 224 186 524
rect 216 512 278 524
rect 216 236 232 512
rect 266 236 278 512
rect 216 224 278 236
<< pdiff >>
rect -407 1153 -345 1165
rect -407 855 -395 1153
rect -361 855 -345 1153
rect -407 843 -345 855
rect -315 1153 -249 1165
rect -315 855 -299 1153
rect -265 855 -249 1153
rect -315 843 -249 855
rect -219 1153 -153 1165
rect -219 855 -203 1153
rect -169 855 -153 1153
rect -219 843 -153 855
rect -123 1153 -57 1165
rect -123 855 -107 1153
rect -73 855 -57 1153
rect -123 843 -57 855
rect -27 1153 39 1165
rect -27 855 -11 1153
rect 23 855 39 1153
rect -27 843 39 855
rect 69 1153 135 1165
rect 69 855 85 1153
rect 119 855 135 1153
rect 69 843 135 855
rect 165 1153 227 1165
rect 165 855 181 1153
rect 215 855 227 1153
rect 165 843 227 855
<< ndiffc >>
rect -344 236 -310 512
rect -56 236 -22 512
rect 232 236 266 512
<< pdiffc >>
rect -395 855 -361 1153
rect -299 855 -265 1153
rect -203 855 -169 1153
rect -107 855 -73 1153
rect -11 855 23 1153
rect 85 855 119 1153
rect 181 855 215 1153
<< poly >>
rect -345 1165 -315 1191
rect -249 1165 -219 1191
rect -153 1165 -123 1191
rect -57 1165 -27 1191
rect 39 1165 69 1191
rect 135 1165 165 1191
rect -345 812 -315 843
rect -249 812 -219 843
rect -153 817 -123 843
rect -57 817 -27 843
rect -153 812 -27 817
rect 39 812 69 843
rect 135 812 165 843
rect -363 796 -219 812
rect -363 762 -347 796
rect -313 762 -219 796
rect -363 746 -219 762
rect -172 796 -27 812
rect -172 762 -155 796
rect -121 762 -27 796
rect -172 746 -27 762
rect 21 796 165 812
rect 21 762 37 796
rect 71 762 165 796
rect 21 746 165 762
rect -356 602 -241 746
rect -172 713 -108 746
rect -174 707 -108 713
rect -356 568 -295 602
rect -258 568 -241 602
rect -356 550 -241 568
rect -198 705 -108 707
rect -198 671 -158 705
rect -121 671 -108 705
rect 21 699 97 746
rect -198 654 -108 671
rect -198 550 -145 654
rect -56 612 97 699
rect -102 596 97 612
rect -102 562 -56 596
rect -21 592 97 596
rect -21 562 48 592
rect -102 552 48 562
rect -294 524 -264 550
rect -198 524 -168 550
rect -102 546 24 552
rect -102 524 -72 546
rect -6 524 24 546
rect 90 524 120 550
rect 186 524 216 550
rect -294 202 -264 224
rect -312 186 -246 202
rect -198 198 -168 224
rect -102 198 -72 224
rect -6 198 24 224
rect 90 198 120 224
rect 186 198 216 224
rect -312 152 -296 186
rect -262 152 -246 186
rect -312 136 -246 152
rect 68 182 135 198
rect 68 148 84 182
rect 119 148 135 182
rect 68 132 135 148
rect 186 182 253 198
rect 186 148 202 182
rect 237 148 253 182
rect 186 132 253 148
<< polycont >>
rect -347 762 -313 796
rect -155 762 -121 796
rect 37 762 71 796
rect -295 568 -258 602
rect -158 671 -121 705
rect -56 562 -21 596
rect -296 152 -262 186
rect 84 148 119 182
rect 202 148 237 182
<< locali >>
rect -395 1159 -361 1169
rect -395 839 -361 855
rect -299 1153 -265 1169
rect -299 839 -265 849
rect -203 1159 -169 1169
rect -203 839 -169 855
rect -107 1153 -73 1169
rect -107 839 -73 849
rect -11 1159 23 1169
rect -11 839 23 855
rect 85 1153 119 1169
rect 85 839 119 849
rect 181 1159 215 1169
rect 181 839 215 855
rect -363 762 -347 796
rect -313 762 -297 796
rect -174 762 -155 796
rect -121 762 -105 796
rect 21 762 37 796
rect 71 762 87 796
rect -174 705 -105 762
rect -174 671 -158 705
rect -121 671 -105 705
rect -174 668 -105 671
rect -311 568 -295 602
rect -258 568 -242 602
rect -102 562 -56 596
rect -21 562 24 596
rect -344 512 -310 528
rect -344 220 -310 236
rect -56 512 -22 528
rect -56 220 -22 236
rect 232 512 266 528
rect 232 220 266 236
rect -312 152 -296 186
rect -262 152 -246 186
rect 68 148 84 182
rect 119 148 135 182
rect 186 148 202 182
rect 237 148 253 182
<< viali >>
rect -395 1153 -361 1159
rect -395 1027 -361 1153
rect -299 855 -265 981
rect -299 849 -265 855
rect -203 1153 -169 1159
rect -203 1027 -169 1153
rect -107 855 -73 981
rect -107 849 -73 855
rect -11 1153 23 1159
rect -11 1027 23 1153
rect 85 855 119 981
rect 85 849 119 855
rect 181 1153 215 1159
rect 181 1027 215 1153
rect 37 762 71 796
rect -158 671 -121 705
rect -295 568 -258 602
rect -56 562 -21 596
rect -344 236 -310 512
rect -56 236 -22 512
rect 232 236 266 512
rect -296 152 -262 186
rect 84 148 119 182
rect 202 148 237 182
<< metal1 >>
rect -407 1165 228 1227
rect -407 1159 227 1165
rect -407 1027 -395 1159
rect -361 1027 -203 1159
rect -169 1027 -11 1159
rect 23 1027 181 1159
rect 215 1027 227 1159
rect -407 1019 227 1027
rect -315 981 351 989
rect -315 849 -299 981
rect -265 849 -107 981
rect -73 849 85 981
rect 119 849 351 981
rect -315 843 351 849
rect -443 796 97 815
rect -443 762 37 796
rect 71 762 97 796
rect -443 746 97 762
rect -80 741 97 746
rect -443 705 -108 718
rect -443 671 -158 705
rect -121 671 -108 705
rect -443 649 -108 671
rect -442 602 -207 621
rect -442 568 -295 602
rect -258 568 -207 602
rect -442 552 -207 568
rect -442 512 -304 524
rect -442 236 -344 512
rect -310 236 -304 512
rect -442 223 -304 236
rect -442 220 -318 223
rect -442 16 -340 220
rect -276 192 -207 552
rect -312 186 -207 192
rect -312 152 -296 186
rect -262 152 -207 186
rect -312 104 -207 152
rect -179 387 -108 649
rect -80 596 24 741
rect -80 562 -56 596
rect -21 562 24 596
rect -80 552 24 562
rect 125 599 351 843
rect 125 524 198 599
rect -62 512 198 524
rect -179 195 -109 387
rect -62 236 -56 512
rect -22 236 198 512
rect -62 224 198 236
rect 226 512 351 524
rect 226 236 232 512
rect 266 332 351 512
rect 266 236 350 332
rect 226 224 350 236
rect 275 223 350 224
rect -179 182 135 195
rect -179 148 84 182
rect 119 148 135 182
rect -179 132 135 148
rect 186 182 253 195
rect 186 148 202 182
rect 237 148 253 182
rect 186 104 253 148
rect -312 45 253 104
rect 281 16 350 223
rect -442 -53 350 16
<< labels >>
rlabel metal1 -443 779 -443 779 7 A
port 1 w
rlabel metal1 -443 649 -410 718 7 B
port 2 w
rlabel metal1 -442 552 -409 568 7 C
port 3 w
rlabel metal1 -442 -53 350 16 5 VSS
port 4 s
rlabel metal1 -407 1166 228 1227 1 VDD
port 5 n
rlabel metal1 298 599 351 989 3 Y
port 6 e
<< end >>
