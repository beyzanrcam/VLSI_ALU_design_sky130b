* NGSPICE file created from NAND3.ext - technology: sky130B

.subckt efen3 a_n173_n300# a_81_n326# a_111_n300# a_n15_n326# a_n111_n326# VSUBS
X0 a_111_n300# a_81_n326# a_15_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X1 a_n81_n300# a_n111_n326# a_n173_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X2 a_15_n300# a_n15_n326# a_n81_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
.ends

.subckt efemosp a_111_n258# w_n353_n261# a_n273_n258# a_n317_n161# a_n81_n258# a_n225_n161#
X0 a_n317_n161# a_111_n258# a_n225_n161# w_n353_n261# sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1 a_n225_n161# a_111_n258# a_n317_n161# w_n353_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2 a_n225_n161# a_n273_n258# a_n317_n161# w_n353_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3 a_n317_n161# a_n81_n258# a_n225_n161# w_n353_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4 a_n317_n161# a_n273_n258# a_n225_n161# w_n353_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X5 a_n225_n161# a_n81_n258# a_n317_n161# w_n353_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
.ends

.subckt NAND3 A B C VSS VDD Y
Xefen3_0 VSS A Y B C VSS efen3
Xefemosp_0 A VDD C VDD B Y efemosp
.ends

