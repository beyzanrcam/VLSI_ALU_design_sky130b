magic
tech sky130B
magscale 1 2
timestamp 1733171354
<< nwell >>
rect 113 1369 1412 2357
rect 113 722 847 1369
rect 867 722 1412 1369
rect 113 573 1412 722
<< psubdiff >>
rect 387 -128 1151 -88
rect 387 -186 637 -128
rect 909 -186 1151 -128
rect 387 -262 1151 -186
<< nsubdiff >>
rect 175 2209 500 2284
rect 175 2146 259 2209
rect 401 2146 500 2209
rect 175 2072 500 2146
<< psubdiffcont >>
rect 637 -186 909 -128
<< nsubdiffcont >>
rect 259 2146 401 2209
<< locali >>
rect 175 2210 500 2218
rect 175 2145 258 2210
rect 402 2145 500 2210
rect 175 2137 500 2145
rect 266 645 568 679
rect 620 645 922 679
rect 974 645 1276 679
rect 518 306 552 645
rect 754 447 788 645
rect 787 413 788 447
rect 518 238 552 272
rect 754 238 788 413
rect 990 552 1024 645
rect 990 238 1024 518
rect 442 204 626 238
rect 678 204 862 238
rect 914 204 1098 238
rect 399 -105 433 -34
rect 635 -105 669 -37
rect 871 -105 905 -35
rect 1107 -105 1141 -36
rect 387 -128 1151 -105
rect 387 -186 637 -128
rect 909 -186 1151 -128
rect 387 -204 1151 -186
<< viali >>
rect 258 2209 402 2210
rect 258 2146 259 2209
rect 259 2146 401 2209
rect 401 2146 402 2209
rect 258 2145 402 2146
rect 753 413 787 447
rect 518 272 552 306
rect 990 518 1024 552
rect 637 -186 909 -128
<< metal1 >>
rect 246 2210 414 2216
rect 246 2145 258 2210
rect 402 2145 414 2210
rect 246 2010 414 2145
rect 217 1413 499 2010
rect 689 1413 1207 2010
rect 577 1362 853 1363
rect 335 1350 853 1362
rect 335 727 847 1350
rect 335 726 617 727
rect 1043 726 1325 1362
rect 247 552 1036 613
rect 247 518 990 552
rect 1024 518 1036 552
rect 247 515 1036 518
rect 983 511 1036 515
rect 247 447 807 487
rect 247 413 753 447
rect 787 413 807 447
rect 247 389 807 413
rect 246 306 570 353
rect 246 272 518 306
rect 552 272 570 306
rect 246 255 570 272
rect 1167 166 1325 726
rect 524 -34 1325 166
rect 625 -128 921 -120
rect 625 -186 637 -128
rect 909 -186 921 -128
rect 625 -193 921 -186
use sky130_fd_pr__nfet_01v8_WPN2C2  sky130_fd_pr__nfet_01v8_WPN2C2_0
timestamp 1733169655
transform 1 0 770 0 1 97
box -383 -157 383 157
use sky130_fd_pr__pfet_01v8_FMUCNY  sky130_fd_pr__pfet_01v8_FMUCNY_0
timestamp 1733168815
transform 1 0 771 0 1 1332
box -596 -706 596 740
<< labels >>
flabel metal1 1189 433 1305 551 1 FreeSerif 320 0 0 0 Y
port 1 n
flabel nwell 277 2145 382 2212 1 FreeSerif 320 0 0 0 VDD
port 2 n
flabel metal1 744 -181 804 -134 1 FreeSerif 320 0 0 0 VSS
port 3 n
flabel metal1 253 272 320 340 1 FreeSerif 320 0 0 0 A
port 4 n
flabel metal1 256 405 323 473 1 FreeSerif 320 0 0 0 B
port 5 n
flabel metal1 256 524 323 592 1 FreeSerif 320 0 0 0 C
port 6 n
<< end >>
