* NGSPICE file created from OR8.ext - technology: sky130B

.subckt sky130_fd_pr__nfet_01v8_6H9P4D a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt efepmos_W107-L15-F3 a_n129_n204# a_n173_n107# w_n209_n207# a_n81_n107#
X0 a_n81_n107# a_n129_n204# a_n173_n107# w_n209_n207# sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1 a_n81_n107# a_n129_n204# a_n173_n107# w_n209_n207# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2 a_n173_n107# a_n129_n204# a_n81_n107# w_n209_n207# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
.ends

.subckt inv A VSS VDD Y
Xsky130_fd_pr__nfet_01v8_6H9P4D_0 Y VSS A VSS sky130_fd_pr__nfet_01v8_6H9P4D
Xefepmos_W107-L15-F3_0 A VDD VDD Y efepmos_W107-L15-F3
.ends

.subckt NOT8 A7 A6 A5 A4 A3 A2 A1 A0 S0 S1 S2 S3 S4 S5 S6 S7 inv_7/VDD VSUBS
Xinv_0 A3 VSUBS inv_7/VDD S3 inv
Xinv_1 A7 VSUBS inv_7/VDD S7 inv
Xinv_2 A6 VSUBS inv_7/VDD S6 inv
Xinv_3 A5 VSUBS inv_7/VDD S5 inv
Xinv_4 A4 VSUBS inv_7/VDD S4 inv
Xinv_5 A2 VSUBS inv_7/VDD S2 inv
Xinv_6 A1 VSUBS inv_7/VDD S1 inv
Xinv_7 A0 VSUBS inv_7/VDD S0 inv
.ends

.subckt nmos_2shared_W200-L015-F1 a_63_n200# a_n63_n226# a_n33_n200# a_33_n226# a_n125_n200#
+ VSUBS
X0 a_n33_n200# a_n63_n226# a_n125_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1 a_63_n200# a_33_n226# a_n33_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
.ends

.subckt pmos_p2-w321-L015-f3 a_n317_n107# w_n353_n143# a_n225_n107# a_33_n138# a_n255_n138#
X0 a_n225_n107# a_33_n138# a_n317_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1 a_n225_n107# a_n255_n138# a_n317_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2 a_n317_n107# a_33_n138# a_n225_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3 a_n317_n107# a_n255_n138# a_n225_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4 a_n225_n107# a_n255_n138# a_n317_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X5 a_n317_n107# a_33_n138# a_n225_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
.ends

.subckt NAND2 A B VSS VDD Y
Xnmos_2shared_W200-L015-F1_0 VSS B a_994_146# A Y VSS nmos_2shared_W200-L015-F1
Xpmos_p2-w321-L015-f3_0 VDD VDD Y B A pmos_p2-w321-L015-f3
.ends

.subckt NAND8 A0 B0 A1 B1 A2 B2 A3 B3 A4 B4 A5 B5 A6 B6 A7 B7 P0 P1 P2 P3 P4 P5 P6
+ P7
XNAND2_7 B6 A6 VSUBS NAND2_9/VDD P6 NAND2
XNAND2_8 B1 A1 VSUBS NAND2_9/VDD P1 NAND2
XNAND2_9 B2 A2 VSUBS NAND2_9/VDD P2 NAND2
XNAND2_0 B7 A7 VSUBS NAND2_9/VDD P7 NAND2
XNAND2_1 B4 A4 VSUBS NAND2_9/VDD P4 NAND2
XNAND2_2 B3 A3 VSUBS NAND2_9/VDD P3 NAND2
XNAND2_4 B0 A0 VSUBS NAND2_9/VDD P0 NAND2
XNAND2_6 B5 A5 VSUBS NAND2_9/VDD P5 NAND2
.ends

.subckt OR8 B7 B6 B5 B4 B3 B2 B1 B0 A7 A6 A5 A4 A3 A2 A1 A0 S0 S1 S2 S3 S4 S5 S6 S7
XNOT8_0 A7 A6 A5 A4 A3 A2 A1 A0 NOT8_0/S0 NOT8_0/S1 NOT8_0/S2 NOT8_0/S3 NOT8_0/S4
+ NOT8_0/S5 NOT8_0/S6 NOT8_0/S7 NOT8_1/inv_7/VDD VSUBS NOT8
XNOT8_1 B7 B6 B5 B4 B3 B2 B1 B0 NOT8_1/S0 NOT8_1/S1 NOT8_1/S2 NOT8_1/S3 NOT8_1/S4
+ NOT8_1/S5 NOT8_1/S6 NOT8_1/S7 NOT8_1/inv_7/VDD VSUBS NOT8
XNAND8_0 NOT8_1/S7 NOT8_0/S7 NOT8_1/S6 NOT8_0/S6 NOT8_1/S5 NOT8_0/S5 NOT8_1/S4 NOT8_0/S4
+ NOT8_1/S3 NOT8_0/S3 NOT8_1/S2 NOT8_0/S2 NOT8_1/S1 NOT8_0/S1 NOT8_1/S0 NOT8_0/S0
+ S7 S6 S5 S4 S3 S2 S1 S0 NAND8
.ends

