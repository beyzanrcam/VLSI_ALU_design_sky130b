magic
tech sky130B
magscale 1 2
timestamp 1736094670
<< nmos >>
rect -159 -400 -129 400
rect -63 -400 -33 400
rect 33 -400 63 400
rect 129 -400 159 400
<< ndiff >>
rect -221 388 -159 400
rect -221 -388 -209 388
rect -175 -388 -159 388
rect -221 -400 -159 -388
rect -129 -400 -63 400
rect -33 -400 33 400
rect 63 -400 129 400
rect 159 388 221 400
rect 159 -388 175 388
rect 209 -388 221 388
rect 159 -400 221 -388
<< ndiffc >>
rect -209 -388 -175 388
rect 175 -388 209 388
<< poly >>
rect -159 400 -129 426
rect -63 400 -33 426
rect 33 400 63 426
rect 129 400 159 426
rect -159 -426 -129 -400
rect -63 -426 -33 -400
rect 33 -426 63 -400
rect 129 -426 159 -400
<< locali >>
rect -209 388 -175 404
rect -209 -404 -175 -388
rect 175 388 209 404
rect 175 -404 209 -388
<< viali >>
rect -209 -388 -175 388
rect 175 -388 209 388
<< metal1 >>
rect -215 388 -169 400
rect -215 -388 -209 388
rect -175 -388 -169 388
rect -215 -400 -169 -388
rect 169 388 215 400
rect 169 -388 175 388
rect 209 -388 215 388
rect 169 -400 215 -388
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 0.150 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
