magic
tech sky130B
magscale 1 2
timestamp 1736085364
<< nwell >>
rect 108 1772 218 2024
<< nsubdiff >>
rect 108 1901 218 2024
rect 108 1775 193 1901
rect 108 1772 218 1775
<< viali >>
rect 2164 1306 2364 1368
<< metal1 >>
rect 600 3429 740 3687
rect 998 3429 1045 3687
rect 72 3072 110 3130
rect 74 2978 112 3036
rect 72 2884 110 2946
rect 1379 2855 1445 3375
rect 74 2790 112 2852
rect 1379 2789 1713 2855
rect 72 1923 218 2757
rect 1396 2378 1713 2789
rect -7 1910 218 1923
rect -7 1766 6 1910
rect 150 1766 218 1910
rect 1647 1837 1713 2378
rect 1750 2403 1907 2416
rect 1750 2270 1761 2403
rect 1894 2276 1907 2403
rect 1894 2270 3122 2276
rect 1750 2259 3122 2270
rect 1760 2171 3122 2259
rect 1760 1985 1828 2171
rect 2908 2088 3122 2171
rect 1760 1980 1834 1985
rect 1647 1771 1983 1837
rect -7 1753 218 1766
rect 72 918 218 1753
rect 1631 1666 1960 1732
rect 1631 1296 1697 1666
rect 3146 1530 3206 1680
rect 2804 1433 2830 1434
rect 74 824 112 886
rect 1332 844 1697 1296
rect 2138 1382 2388 1384
rect 2138 1368 3108 1382
rect 2138 1306 2164 1368
rect 2364 1306 3108 1368
rect 2138 1297 3108 1306
rect 2138 1288 2388 1297
rect 2227 1224 2233 1288
rect 2297 1224 2303 1288
rect 1391 817 1697 844
rect 76 730 114 792
rect 76 636 114 698
rect 78 542 116 604
rect 602 -12 676 247
rect 935 -12 1045 247
<< via1 >>
rect 740 3429 998 3687
rect 6 1766 150 1910
rect 1761 2270 1894 2403
rect 2233 1224 2297 1288
rect 676 -12 935 247
<< metal2 >>
rect 705 3687 1043 3730
rect 705 3429 740 3687
rect 998 3429 1043 3687
rect 705 3396 1043 3429
rect 1750 2403 1907 2416
rect 1750 2270 1761 2403
rect 1894 2270 1907 2403
rect 1750 2259 1907 2270
rect -7 1910 163 1923
rect -7 1766 6 1910
rect 150 1766 163 1910
rect -7 1753 163 1766
rect 2102 1288 2429 1419
rect 2102 1224 2233 1288
rect 2297 1224 2429 1288
rect 2102 1091 2429 1224
rect 651 247 971 277
rect 651 -12 676 247
rect 935 -12 971 247
rect 651 -43 971 -12
<< via2 >>
rect 740 3429 998 3687
rect 1761 2270 1894 2403
rect 6 1766 150 1910
rect 2233 1224 2297 1288
rect 686 -12 935 247
<< metal3 >>
rect 705 3692 1043 3730
rect 705 3424 735 3692
rect 1003 3424 1043 3692
rect 705 3396 1043 3424
rect 1750 2408 1907 2416
rect 1750 2265 1756 2408
rect 1899 2265 1907 2408
rect 1750 2259 1907 2265
rect -7 1915 163 1923
rect -7 1761 1 1915
rect 155 1761 163 1915
rect -7 1753 163 1761
rect 2102 1293 2429 1419
rect 2102 1219 2228 1293
rect 2302 1219 2429 1293
rect 2102 1091 2429 1219
rect 651 252 971 277
rect 651 -17 681 252
rect 940 -17 971 252
rect 651 -43 971 -17
<< via3 >>
rect 735 3687 1003 3692
rect 735 3429 740 3687
rect 740 3429 998 3687
rect 998 3429 1003 3687
rect 735 3424 1003 3429
rect 1756 2403 1899 2408
rect 1756 2270 1761 2403
rect 1761 2270 1894 2403
rect 1894 2270 1899 2403
rect 1756 2265 1899 2270
rect 1 1910 155 1915
rect 1 1766 6 1910
rect 6 1766 150 1910
rect 150 1766 155 1910
rect 1 1761 155 1766
rect 2228 1288 2302 1293
rect 2228 1224 2233 1288
rect 2233 1224 2297 1288
rect 2297 1224 2302 1288
rect 2228 1219 2302 1224
rect 681 247 940 252
rect 681 -12 686 247
rect 686 -12 935 247
rect 935 -12 940 247
rect 681 -17 940 -12
<< metal4 >>
rect 1755 2408 1900 2409
rect 1755 2265 1756 2408
rect 1899 2265 1900 2408
rect 1755 2264 1900 2265
rect 0 1915 156 1916
rect 0 1761 1 1915
rect 155 1761 156 1915
rect 0 1760 156 1761
<< via4 >>
rect 733 3692 1005 3694
rect 733 3424 735 3692
rect 735 3424 1003 3692
rect 1003 3424 1005 3692
rect 733 3422 1005 3424
rect 2129 1293 2401 1392
rect 2129 1219 2228 1293
rect 2228 1219 2302 1293
rect 2302 1219 2401 1293
rect 2129 1120 2401 1219
rect 675 252 947 254
rect 675 -17 681 252
rect 681 -17 940 252
rect 940 -17 947 252
rect 675 -18 947 -17
<< metal5 >>
rect 674 3694 1202 3802
rect 674 3422 733 3694
rect 1005 3422 1202 3694
rect 674 3380 1202 3422
rect 2059 1392 2506 1471
rect 2059 1120 2129 1392
rect 2401 1120 2506 1392
rect 2059 1061 2506 1120
rect 589 254 1081 299
rect 589 -18 675 254
rect 947 -18 1081 254
rect 589 -74 1081 -18
use inv  inv_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/inv
timestamp 1735843251
transform 1 0 2808 0 1 1608
box 0 -311 412 486
use nor2  nor2_1 ~/Documents/vlsi/vlsi_sky130b/design/mag/NOR/NOR2
timestamp 1736020690
transform 1 0 1718 0 1 1768
box 0 -480 1090 580
use nor4  nor4_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NOR/NOR4
timestamp 1736019943
transform 1 0 674 0 -1 3804
box -602 118 790 1966
use nor4  nor4_1
timestamp 1736019943
transform 1 0 674 0 1 -128
box -602 118 790 1966
<< labels >>
flabel metal1 84 3082 96 3118 0 FreeSans 160 0 0 0 A0
port 0 nsew
flabel metal1 86 2990 98 3026 0 FreeSans 160 0 0 0 A1
port 1 nsew
flabel metal1 86 2896 98 2932 0 FreeSans 160 0 0 0 A2
port 2 nsew
flabel metal1 86 2800 98 2836 0 FreeSans 160 0 0 0 A3
port 3 nsew
flabel metal1 80 836 104 876 0 FreeSans 160 0 0 0 A4
port 4 nsew
flabel metal1 86 740 110 780 0 FreeSans 160 0 0 0 A5
port 5 nsew
flabel metal1 84 644 108 684 0 FreeSans 160 0 0 0 A6
port 6 nsew
flabel metal1 84 552 108 592 0 FreeSans 160 0 0 0 A7
port 8 nsew
flabel metal1 3156 1542 3196 1664 0 FreeSans 160 0 0 0 Z
port 10 nsew
flabel metal5 718 3426 996 3670 0 FreeSans 160 0 0 0 VSS
flabel metal5 682 -10 960 234 0 FreeSans 160 0 0 0 VSS
flabel metal5 2150 1116 2428 1360 0 FreeSans 160 0 0 0 VSS
flabel metal4 1810 2268 1854 2378 0 FreeSans 160 0 0 0 VDD
flabel metal4 94 1782 138 1892 0 FreeSans 160 0 0 0 VDD
<< end >>
