magic
tech sky130B
magscale 1 2
timestamp 1736181444
<< nwell >>
rect 356 372 1062 892
<< nmos >>
rect 626 212 1026 242
rect 626 116 1026 146
<< pmos >>
rect 454 434 484 648
rect 550 434 580 648
rect 646 434 676 648
rect 742 434 772 648
rect 838 434 868 648
rect 934 434 964 648
<< ndiff >>
rect 626 292 1026 304
rect 626 258 638 292
rect 1014 258 1026 292
rect 626 242 1026 258
rect 626 146 1026 212
rect 626 100 1026 116
rect 626 66 638 100
rect 1014 66 1026 100
rect 626 54 1026 66
<< pdiff >>
rect 392 636 454 648
rect 392 446 404 636
rect 438 446 454 636
rect 392 434 454 446
rect 484 636 550 648
rect 484 446 500 636
rect 534 446 550 636
rect 484 434 550 446
rect 580 636 646 648
rect 580 446 596 636
rect 630 446 646 636
rect 580 434 646 446
rect 676 636 742 648
rect 676 446 692 636
rect 726 446 742 636
rect 676 434 742 446
rect 772 636 838 648
rect 772 446 788 636
rect 822 446 838 636
rect 772 434 838 446
rect 868 636 934 648
rect 868 446 884 636
rect 918 446 934 636
rect 868 434 934 446
rect 964 636 1026 648
rect 964 446 980 636
rect 1014 446 1026 636
rect 964 434 1026 446
<< ndiffc >>
rect 638 258 1014 292
rect 638 66 1014 100
<< pdiffc >>
rect 404 446 438 636
rect 500 446 534 636
rect 596 446 630 636
rect 692 446 726 636
rect 788 446 822 636
rect 884 446 918 636
rect 980 446 1014 636
<< psubdiff >>
rect 626 30 1026 54
rect 626 -44 653 30
rect 988 -44 1026 30
rect 626 -63 1026 -44
<< nsubdiff >>
rect 396 791 1013 852
rect 396 744 606 791
rect 846 744 1013 791
rect 396 702 1013 744
<< psubdiffcont >>
rect 653 -44 988 30
<< nsubdiffcont >>
rect 606 744 846 791
<< poly >>
rect 454 648 484 679
rect 550 648 580 679
rect 646 648 676 679
rect 742 648 772 679
rect 838 648 868 679
rect 934 648 964 679
rect 454 408 484 434
rect 550 408 580 434
rect 646 408 676 434
rect 453 387 676 408
rect 453 352 470 387
rect 504 378 676 387
rect 742 408 772 434
rect 838 408 868 434
rect 934 408 964 434
rect 742 387 964 408
rect 504 352 520 378
rect 453 341 520 352
rect 742 352 759 387
rect 793 378 964 387
rect 793 352 809 378
rect 742 341 809 352
rect 453 146 496 341
rect 538 263 604 279
rect 538 228 554 263
rect 588 242 604 263
rect 588 228 626 242
rect 538 212 626 228
rect 1026 212 1052 242
rect 453 130 626 146
rect 453 95 554 130
rect 588 116 626 130
rect 1026 116 1052 146
rect 588 95 604 116
rect 453 79 604 95
<< polycont >>
rect 470 352 504 387
rect 759 352 793 387
rect 554 228 588 263
rect 554 95 588 130
<< locali >>
rect 532 744 606 791
rect 846 744 946 791
rect 404 642 438 652
rect 404 430 438 446
rect 500 636 534 652
rect 500 430 534 440
rect 596 642 630 652
rect 596 430 630 446
rect 692 636 726 652
rect 692 430 726 440
rect 788 642 822 652
rect 788 430 822 446
rect 884 636 918 652
rect 884 430 918 440
rect 980 642 1014 652
rect 980 430 1014 446
rect 453 352 470 387
rect 504 352 520 387
rect 742 381 759 387
rect 554 352 759 381
rect 793 352 809 387
rect 453 146 496 352
rect 554 347 809 352
rect 554 263 588 347
rect 622 258 638 292
rect 1014 258 1030 292
rect 554 212 588 228
rect 453 130 588 146
rect 453 95 554 130
rect 453 79 588 95
rect 622 66 638 100
rect 1014 66 1030 100
rect 626 -44 653 30
rect 988 -44 1026 30
<< viali >>
rect 606 744 846 791
rect 404 636 438 642
rect 404 562 438 636
rect 500 446 534 520
rect 500 440 534 446
rect 596 636 630 642
rect 596 562 630 636
rect 692 446 726 520
rect 692 440 726 446
rect 788 636 822 642
rect 788 562 822 636
rect 884 446 918 520
rect 884 440 918 446
rect 980 636 1014 642
rect 980 562 1014 636
rect 470 352 504 387
rect 759 352 793 387
rect 554 228 588 263
rect 638 258 1014 292
rect 638 66 1014 100
rect 653 -44 988 25
<< metal1 >>
rect 532 791 869 803
rect 532 744 606 791
rect 846 744 869 791
rect 532 684 869 744
rect 391 648 1025 684
rect 391 642 1026 648
rect 391 562 404 642
rect 438 562 596 642
rect 630 562 788 642
rect 822 562 980 642
rect 1014 562 1026 642
rect 391 556 1026 562
rect 391 555 1025 556
rect 484 520 1062 526
rect 484 440 500 520
rect 534 440 692 520
rect 726 440 884 520
rect 918 440 1062 520
rect 484 434 1062 440
rect 356 387 520 405
rect 356 352 470 387
rect 504 352 520 387
rect 356 270 520 352
rect 548 387 808 406
rect 548 352 759 387
rect 793 352 808 387
rect 548 332 808 352
rect 548 263 598 332
rect 884 304 1062 434
rect 548 241 554 263
rect 356 228 554 241
rect 588 228 598 263
rect 626 292 1062 304
rect 626 258 638 292
rect 1014 258 1062 292
rect 626 252 1062 258
rect 356 105 598 228
rect 626 100 1026 106
rect 626 66 638 100
rect 1014 66 1026 100
rect 626 25 1026 66
rect 626 -44 653 25
rect 988 -44 1026 25
rect 626 -63 1026 -44
<< end >>
