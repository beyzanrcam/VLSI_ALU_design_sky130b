magic
tech sky130B
magscale 1 2
timestamp 1736620191
<< nwell >>
rect 108 1772 218 2024
rect 1449 1873 1743 2305
rect 2418 1873 2863 2304
<< nsubdiff >>
rect 108 1901 218 2024
rect 108 1775 193 1901
rect 108 1772 218 1775
<< metal1 >>
rect 600 3429 740 3687
rect 998 3429 1045 3687
rect 72 3072 110 3130
rect 74 2978 112 3036
rect 72 2884 110 2946
rect 1379 2855 1445 3375
rect 74 2790 112 2852
rect 1379 2789 1713 2855
rect 72 1923 218 2757
rect 1396 2378 1713 2789
rect -7 1910 218 1923
rect -7 1766 6 1910
rect 150 1766 218 1910
rect 1647 1771 1713 2378
rect 1970 2403 2127 2416
rect 1970 2270 1981 2403
rect 2114 2276 2127 2403
rect 2114 2270 2832 2276
rect 1970 2259 2832 2270
rect 1980 2253 2832 2259
rect 1760 2177 2832 2253
rect 1760 2171 2382 2177
rect -7 1753 218 1766
rect 2419 1753 2517 2027
rect 2802 1759 2862 1909
rect 72 918 218 1753
rect 1647 1732 1713 1742
rect 1647 1666 1714 1732
rect 1647 1296 1713 1666
rect 2381 1484 2432 1555
rect 2503 1484 2661 1555
rect 74 824 112 886
rect 1332 844 1713 1296
rect 1391 817 1713 844
rect 76 730 114 792
rect 76 636 114 698
rect 78 542 116 604
rect 602 -12 676 247
rect 935 -12 1045 247
<< via1 >>
rect 740 3429 998 3687
rect 6 1766 150 1910
rect 1981 2270 2114 2403
rect 2432 1484 2503 1555
rect 676 -12 935 247
<< metal2 >>
rect 705 3687 1043 3730
rect 705 3429 740 3687
rect 998 3429 1043 3687
rect 705 3396 1043 3429
rect 1970 2403 2127 2416
rect 1970 2270 1981 2403
rect 2114 2270 2127 2403
rect 1970 2259 2127 2270
rect -7 1910 163 1923
rect -7 1766 6 1910
rect 150 1766 163 1910
rect -7 1753 163 1766
rect 2421 1555 2514 1566
rect 2421 1484 2432 1555
rect 2503 1484 2514 1555
rect 2421 1473 2514 1484
rect 651 247 971 277
rect 651 -12 676 247
rect 935 -12 971 247
rect 651 -43 971 -12
<< via2 >>
rect 740 3429 998 3687
rect 1981 2270 2114 2403
rect 6 1766 150 1910
rect 2432 1484 2503 1555
rect 686 -12 935 247
<< metal3 >>
rect 705 3692 1043 3730
rect 705 3424 735 3692
rect 1003 3424 1043 3692
rect 705 3396 1043 3424
rect 1970 2408 2127 2416
rect 1970 2265 1976 2408
rect 2119 2265 2127 2408
rect 1970 2259 2127 2265
rect -7 1915 163 1923
rect -7 1761 1 1915
rect 155 1761 163 1915
rect -7 1753 163 1761
rect 2406 1560 2532 1579
rect 2406 1479 2427 1560
rect 2508 1479 2532 1560
rect 2406 1459 2532 1479
rect 651 252 971 277
rect 651 -17 681 252
rect 940 -17 971 252
rect 651 -43 971 -17
<< via3 >>
rect 735 3687 1003 3692
rect 735 3429 740 3687
rect 740 3429 998 3687
rect 998 3429 1003 3687
rect 735 3424 1003 3429
rect 1976 2403 2119 2408
rect 1976 2270 1981 2403
rect 1981 2270 2114 2403
rect 2114 2270 2119 2403
rect 1976 2265 2119 2270
rect 1 1910 155 1915
rect 1 1766 6 1910
rect 6 1766 150 1910
rect 150 1766 155 1910
rect 1 1761 155 1766
rect 2427 1555 2508 1560
rect 2427 1484 2432 1555
rect 2432 1484 2503 1555
rect 2503 1484 2508 1555
rect 2427 1479 2508 1484
rect 681 247 940 252
rect 681 -12 686 247
rect 686 -12 935 247
rect 935 -12 940 247
rect 681 -17 940 -12
<< metal4 >>
rect 137 2408 2144 2426
rect 137 2265 1976 2408
rect 2119 2265 2144 2408
rect 137 2254 2144 2265
rect 1898 2251 2144 2254
rect -7 1915 168 1925
rect -7 1761 1 1915
rect 155 1761 168 1915
rect -7 1753 168 1761
<< via4 >>
rect 733 3692 1005 3694
rect 733 3424 735 3692
rect 735 3424 1003 3692
rect 1003 3424 1005 3692
rect 733 3422 1005 3424
rect 2332 1560 2604 1656
rect 2332 1479 2427 1560
rect 2427 1479 2508 1560
rect 2508 1479 2604 1560
rect 2332 1384 2604 1479
rect 675 252 947 254
rect 675 -17 681 252
rect 681 -17 940 252
rect 940 -17 947 252
rect 675 -18 947 -17
<< metal5 >>
rect 71 3694 2859 3814
rect 71 3422 733 3694
rect 1005 3422 2859 3694
rect 71 1656 2859 3422
rect 71 1384 2332 1656
rect 2604 1384 2859 1656
rect 71 254 2859 1384
rect 71 -18 675 254
rect 947 -18 2859 254
rect 71 -79 2859 -18
use inv  inv_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/inv
timestamp 1736620191
transform 1 0 2451 0 1 1795
box 0 -311 412 486
use NAND2  NAND2_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NAND/NAND2
timestamp 1736620191
transform 1 0 1357 0 1 1501
box 356 -17 1062 804
use nor4  nor4_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NOR/NOR4
timestamp 1736019943
transform 1 0 674 0 -1 3804
box -602 118 790 1966
use nor4  nor4_1
timestamp 1736019943
transform 1 0 674 0 1 -128
box -602 118 790 1966
<< labels >>
flabel metal1 84 3082 96 3118 0 FreeSans 160 0 0 0 A0
port 0 nsew
flabel metal1 86 2990 98 3026 0 FreeSans 160 0 0 0 A1
port 1 nsew
flabel metal1 86 2896 98 2932 0 FreeSans 160 0 0 0 A2
port 2 nsew
flabel metal1 86 2800 98 2836 0 FreeSans 160 0 0 0 A3
port 3 nsew
flabel metal1 80 836 104 876 0 FreeSans 160 0 0 0 A4
port 4 nsew
flabel metal1 86 740 110 780 0 FreeSans 160 0 0 0 A5
port 5 nsew
flabel metal1 84 644 108 684 0 FreeSans 160 0 0 0 A6
port 6 nsew
flabel metal1 84 552 108 592 0 FreeSans 160 0 0 0 A7
port 8 nsew
flabel metal4 94 1782 138 1892 0 FreeSans 160 0 0 0 VDD
port 12 nsew
flabel metal1 2812 1771 2852 1893 0 FreeSans 160 0 0 0 Z
port 10 nsew
rlabel metal5 1497 -44 1903 197 5 VSS
port 11 s
<< end >>
