* NGSPICE file created from MULT.ext - technology: sky130B

.subckt nmos_2shared_W200-L015-F1 a_63_n200# a_n63_n226# a_n33_n200# a_33_n226# a_n125_n200#
+ VSUBS
X0 a_n33_n200# a_n63_n226# a_n125_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=6.2e+11p ps=4.62e+06u w=2e+06u l=150000u
X1 a_63_n200# a_33_n226# a_n33_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=4.62e+06u as=0p ps=0u w=2e+06u l=150000u
.ends

.subckt pmos_p2-w321-L015-f3 a_n317_n107# w_n353_n143# a_n225_n107# a_33_n138# a_n255_n138#
X0 a_n225_n107# a_33_n138# a_n317_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=1.0593e+12p pd=8.4e+06u as=1.3696e+12p ps=1.112e+07u w=1.07e+06u l=150000u
X1 a_n225_n107# a_n255_n138# a_n317_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.07e+06u l=150000u
X2 a_n317_n107# a_33_n138# a_n225_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.07e+06u l=150000u
X3 a_n317_n107# a_n255_n138# a_n225_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.07e+06u l=150000u
X4 a_n225_n107# a_n255_n138# a_n317_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.07e+06u l=150000u
X5 a_n317_n107# a_33_n138# a_n225_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.07e+06u l=150000u
.ends

.subckt NAND2 A B VSS VDD Y
Xnmos_2shared_W200-L015-F1_0 VSS B a_994_146# A Y VSS nmos_2shared_W200-L015-F1
Xpmos_p2-w321-L015-f3_0 VDD VDD Y B A pmos_p2-w321-L015-f3
.ends

.subckt sky130_fd_pr__nfet_01v8_6H9P4D a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt efepmos_W107-L15-F3 a_n129_n204# a_n173_n107# w_n209_n207# a_n81_n107#
X0 a_n81_n107# a_n129_n204# a_n173_n107# w_n209_n207# sky130_fd_pr__pfet_01v8 ad=6.848e+11p pd=5.56e+06u as=6.848e+11p ps=5.56e+06u w=1.07e+06u l=150000u
X1 a_n81_n107# a_n129_n204# a_n173_n107# w_n209_n207# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.07e+06u l=150000u
X2 a_n173_n107# a_n129_n204# a_n81_n107# w_n209_n207# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.07e+06u l=150000u
.ends

.subckt inv A VSS Y VDD
Xsky130_fd_pr__nfet_01v8_6H9P4D_0 Y VSS A VSS sky130_fd_pr__nfet_01v8_6H9P4D
Xefepmos_W107-L15-F3_0 A VDD VDD Y efepmos_W107-L15-F3
.ends

.subckt XOR2 A B Y a_99_341# VDD VSS
X0 VDD A a_129_987# VDD sky130_fd_pr__pfet_01v8 ad=3.52e+12p pd=2.456e+07u as=5.445e+12p ps=3.696e+07u w=2.75e+06u l=150000u
X1 a_129_987# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.75e+06u l=150000u
X2 a_129_987# a_n51_367# Y VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.7225e+12p ps=1.848e+07u w=2.75e+06u l=150000u
X3 Y a_99_341# a_129_987# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.75e+06u l=150000u
X4 Y a_n51_367# a_129_987# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.75e+06u l=150000u
X5 Y a_n51_367# a_129_987# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.75e+06u l=150000u
X6 a_129_987# a_99_341# Y VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.75e+06u l=150000u
X7 a_129_987# a_99_341# Y VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.75e+06u l=150000u
X8 VDD B a_129_987# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.75e+06u l=150000u
X9 a_129_367# a_99_341# VSS VSS sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=5.88e+06u as=8.32e+11p ps=7.76e+06u w=650000u l=150000u
X10 a_99_341# B VSS VSS sky130_fd_pr__nfet_01v8 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=150000u
X11 a_129_987# B VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.75e+06u l=150000u
X12 VDD B a_129_987# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.75e+06u l=150000u
X13 VSS A a_n51_367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=150000u
X14 a_129_987# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.75e+06u l=150000u
X15 a_99_341# B VDD VDD sky130_fd_pr__pfet_01v8 ad=7.975e+11p pd=6.08e+06u as=0p ps=0u w=2.75e+06u l=150000u
X16 VDD A a_n51_367# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.975e+11p ps=6.08e+06u w=2.75e+06u l=150000u
X17 VSS a_99_341# a_129_367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_129_367# a_99_341# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_129_367# a_n51_367# Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=5.88e+06u w=650000u l=150000u
X20 Y A a_705_367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=5.88e+06u w=650000u l=150000u
X21 Y a_n51_367# a_129_367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y a_n51_367# a_129_367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_705_367# A Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_705_367# A Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VSS B a_705_367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_705_367# B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VSS B a_705_367# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt FULL_ADDER COUT CIN A B VDD VSS OUT
XNAND2_0 B A VSS VDD NAND2_2/B NAND2
XNAND2_1 XOR2_1/A CIN VSS VDD NAND2_2/A NAND2
XNAND2_2 NAND2_2/A NAND2_2/B VSS VDD COUT NAND2
XXOR2_0 B A XOR2_1/A li_1358_495# VDD VSS XOR2
XXOR2_1 XOR2_1/A CIN OUT XOR2_1/a_99_341# VDD VSS XOR2
.ends

.subckt x4bit_ADDER A2 A1 A0 B0 B1 B2 S0 S1 S2 S3 C Cout A3 B3 VDD VSS
XFULL_ADDER_0 Cout FULL_ADDER_0/CIN A3 B3 VDD VSS S3 FULL_ADDER
XFULL_ADDER_1 FULL_ADDER_0/CIN FULL_ADDER_1/CIN A2 B2 VDD VSS S2 FULL_ADDER
XFULL_ADDER_2 FULL_ADDER_1/CIN FULL_ADDER_2/CIN A1 B1 VDD VSS S1 FULL_ADDER
XFULL_ADDER_3 FULL_ADDER_2/CIN C A0 B0 VDD VSS S0 FULL_ADDER
.ends

.subckt MULT A0 B2 B0 B3 A2 A1 A3 SO S1 S2 S5 S4 S3 S7 S6 VSS VDD B1
XNAND2_13 B2 A3 VSS VDD inv_13/A NAND2
XNAND2_7 B2 A1 VSS VDD inv_7/A NAND2
XNAND2_8 A0 B3 VSS VDD inv_8/A NAND2
XNAND2_14 A2 B3 VSS VDD inv_14/A NAND2
XNAND2_15 B3 A3 VSS VDD inv_15/A NAND2
XNAND2_9 B3 A1 VSS VDD inv_9/A NAND2
Xinv_10 inv_10/A VSS inv_10/Y VDD inv
Xinv_11 inv_11/A VSS inv_11/Y VDD inv
Xinv_12 inv_12/A VSS inv_12/Y VDD inv
Xinv_13 inv_13/A VSS inv_13/Y VDD inv
Xinv_14 inv_14/A VSS inv_14/Y VDD inv
Xinv_15 inv_15/A VSS inv_15/Y VDD inv
Xinv_0 inv_0/A VSS inv_0/Y VDD inv
Xinv_1 inv_1/A VSS inv_1/Y VDD inv
X4bit_ADDER_0 inv_10/Y inv_4/Y inv_5/Y inv_2/Y inv_1/Y inv_0/Y S1 4bit_ADDER_1/B0
+ 4bit_ADDER_1/B1 4bit_ADDER_1/B2 VSS 4bit_ADDER_1/B3 inv_11/Y VSS VDD VSS x4bit_ADDER
Xinv_2 inv_2/A VSS inv_2/Y VDD inv
X4bit_ADDER_1 inv_12/Y inv_7/Y inv_6/Y 4bit_ADDER_1/B0 4bit_ADDER_1/B1 4bit_ADDER_1/B2
+ S2 4bit_ADDER_2/B0 4bit_ADDER_2/B1 4bit_ADDER_2/B2 VSS 4bit_ADDER_2/B3 inv_13/Y
+ 4bit_ADDER_1/B3 VDD VSS x4bit_ADDER
Xinv_3 inv_3/A VSS SO VDD inv
X4bit_ADDER_2 inv_14/Y inv_9/Y inv_8/Y 4bit_ADDER_2/B0 4bit_ADDER_2/B1 4bit_ADDER_2/B2
+ S3 S4 S5 S6 VSS S7 inv_15/Y 4bit_ADDER_2/B3 VDD VSS x4bit_ADDER
Xinv_4 inv_4/A VSS inv_4/Y VDD inv
Xinv_5 inv_5/A VSS inv_5/Y VDD inv
Xinv_7 inv_7/A VSS inv_7/Y VDD inv
Xinv_6 inv_6/A VSS inv_6/Y VDD inv
XNAND2_1 B0 A2 VSS VDD inv_1/A NAND2
XNAND2_0 B0 A3 VSS VDD inv_0/A NAND2
Xinv_8 inv_8/A VSS inv_8/Y VDD inv
XNAND2_2 B0 A1 VSS VDD inv_2/A NAND2
Xinv_9 inv_9/A VSS inv_9/Y VDD inv
XNAND2_3 B0 A0 VSS VDD inv_3/A NAND2
XNAND2_10 A2 B1 VSS VDD inv_10/A NAND2
XNAND2_4 A0 B1 VSS VDD inv_5/A NAND2
XNAND2_11 B1 A3 VSS VDD inv_11/A NAND2
XNAND2_5 B1 A1 VSS VDD inv_4/A NAND2
XNAND2_12 A2 B2 VSS VDD inv_12/A NAND2
XNAND2_6 A0 B2 VSS VDD inv_6/A NAND2
.ends

