magic
tech sky130B
magscale 1 2
timestamp 1732814151
<< nmos >>
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
<< ndiff >>
rect -221 88 -159 100
rect -221 -88 -209 88
rect -175 -88 -159 88
rect -221 -100 -159 -88
rect -129 -100 -63 100
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 -100 129 100
rect 159 88 221 100
rect 159 -88 175 88
rect 209 -88 221 88
rect 159 -100 221 -88
<< ndiffc >>
rect -209 -88 -175 88
rect -17 -88 17 88
rect 175 -88 209 88
<< poly >>
rect -159 100 -129 126
rect -63 100 -33 126
rect 33 100 63 126
rect 129 100 159 126
rect -159 -126 -129 -100
rect -63 -126 -33 -100
rect 33 -126 63 -100
rect 129 -126 159 -100
<< locali >>
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 175 88 209 104
rect 175 -104 209 -88
<< viali >>
rect -209 -88 -175 88
rect -17 -88 17 88
rect 175 -88 209 88
<< metal1 >>
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.150 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
