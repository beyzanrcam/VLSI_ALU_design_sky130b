magic
tech sky130B
magscale 1 2
timestamp 1733616374
<< error_p >>
rect -545 169 641 207
rect -641 32 641 169
rect -737 -136 641 32
rect -641 -169 641 -136
rect -641 -207 545 -169
<< nwell >>
rect -545 169 641 207
rect -641 -136 641 169
rect -641 -207 -569 -136
rect -543 -169 641 -136
rect -543 -207 545 -169
<< pmos >>
rect -543 -107 -513 107
rect -447 -107 -417 107
rect -351 -107 -321 107
rect -255 -107 -225 107
rect -159 -107 -129 107
rect -63 -107 -33 107
rect 33 -107 63 107
rect 129 -107 159 107
rect 225 -107 255 107
rect 321 -107 351 107
rect 417 -107 447 107
rect 513 -107 543 107
<< pdiff >>
rect -605 95 -543 107
rect -605 -95 -593 95
rect -559 -95 -543 95
rect -605 -107 -543 -95
rect -513 -107 -447 107
rect -417 95 -351 107
rect -417 -95 -401 95
rect -367 -95 -351 95
rect -417 -107 -351 -95
rect -321 -107 -255 107
rect -225 95 -159 107
rect -225 -95 -209 95
rect -175 -95 -159 95
rect -225 -107 -159 -95
rect -129 -107 -63 107
rect -33 95 33 107
rect -33 -95 -17 95
rect 17 -95 33 95
rect -33 -107 33 -95
rect 63 -107 129 107
rect 159 95 225 107
rect 159 -95 175 95
rect 209 -95 225 95
rect 159 -107 225 -95
rect 255 -107 321 107
rect 351 95 417 107
rect 351 -95 367 95
rect 401 -95 417 95
rect 351 -107 417 -95
rect 447 -107 513 107
rect 543 95 605 107
rect 543 -95 559 95
rect 593 -95 605 95
rect 543 -107 605 -95
<< pdiffc >>
rect -593 -95 -559 95
rect -401 -95 -367 95
rect -209 -95 -175 95
rect -17 -95 17 95
rect 175 -95 209 95
rect 367 -95 401 95
rect 559 -95 593 95
<< poly >>
rect -543 107 -513 133
rect -447 107 -417 133
rect -351 107 -321 133
rect -255 107 -225 133
rect -159 107 -129 133
rect -63 107 -33 133
rect 33 107 63 133
rect 129 107 159 133
rect 225 107 255 133
rect 321 107 351 133
rect 417 107 447 133
rect 513 107 543 133
rect -543 -138 -513 -107
rect -447 -138 -417 -107
rect -351 -138 -321 -107
rect -255 -138 -225 -107
rect -159 -138 -129 -107
rect -63 -138 -33 -107
rect -543 -154 -33 -138
rect -543 -188 -161 -154
rect -127 -188 -33 -154
rect -543 -204 -33 -188
rect 33 -138 63 -107
rect 129 -138 159 -107
rect 225 -138 255 -107
rect 321 -138 351 -107
rect 417 -138 447 -107
rect 513 -138 543 -107
rect 33 -204 543 -138
<< polycont >>
rect -161 -188 -127 -154
<< locali >>
rect -593 95 -559 111
rect -593 -111 -559 -95
rect -401 95 -367 111
rect -401 -111 -367 -95
rect -209 95 -175 111
rect -209 -111 -175 -95
rect -17 95 17 111
rect -17 -111 17 -95
rect 175 95 209 111
rect 175 -111 209 -95
rect 367 95 401 111
rect 367 -111 401 -95
rect 559 95 593 111
rect 559 -111 593 -95
rect -177 -188 -161 -154
rect -127 -188 -111 -154
<< viali >>
rect -593 -95 -559 95
rect -401 -95 -367 95
rect -209 -95 -175 95
rect -17 -95 17 95
rect 175 -95 209 95
rect 367 -95 401 95
rect 559 -95 593 95
<< metal1 >>
rect -599 95 -553 107
rect -599 -95 -593 95
rect -559 -95 -553 95
rect -599 -107 -553 -95
rect -407 95 -361 107
rect -407 -95 -401 95
rect -367 -95 -361 95
rect -407 -107 -361 -95
rect -215 95 -169 107
rect -215 -95 -209 95
rect -175 -95 -169 95
rect -215 -107 -169 -95
rect -23 95 23 107
rect -23 -95 -17 95
rect 17 -95 23 95
rect -23 -107 23 -95
rect 169 95 215 107
rect 169 -95 175 95
rect 209 -95 215 95
rect 169 -107 215 -95
rect 361 95 407 107
rect 361 -95 367 95
rect 401 -95 407 95
rect 361 -107 407 -95
rect 553 95 599 107
rect 553 -95 559 95
rect 593 -95 599 95
rect 553 -107 599 -95
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.07 l 0.15 m 1 nf 12 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
