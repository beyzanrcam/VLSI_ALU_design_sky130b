* NGSPICE file created from nor2_pex.ext - technology: sky130B

.subckt nor2 A B VSS VDD Y
X0 Y.t0 A.t0 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1 a_128_103.t4 A.t1 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2 VDD.t7 A.t2 a_128_103.t3 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3 VDD.t5 A.t3 a_128_103.t2 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X4 a_128_103.t1 A.t4 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X5 Y.t3 B.t0 a_128_103.t7 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X6 a_128_103.t8 B.t1 Y.t4 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X7 Y.t5 B.t2 a_128_103.t9 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X8 Y.t2 B.t3 a_128_103.t6 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X9 a_128_103.t5 B.t4 Y.t1 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X10 a_128_103.t0 A.t5 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X11 VSS.t3 B.t5 Y.t6 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
R0 A.n0 A.t0 379.173
R1 A.n1 A.t5 312.599
R2 A.n0 A.t4 247.428
R3 A.n3 A.t3 247.428
R4 A.n2 A.t1 247.428
R5 A.n1 A.t2 247.428
R6 A A.n4 161.994
R7 A.n3 A.n2 65.1723
R8 A.n2 A.n1 65.1723
R9 A.n4 A.n3 33.2653
R10 A.n4 A.n0 31.9075
R11 VSS.n0 VSS.t2 437.267
R12 VSS.n0 VSS.t0 437.267
R13 VSS.n1 VSS.n0 390
R14 VSS.n1 VSS.t3 156.332
R15 VSS.n1 VSS.t1 156.332
R16 VSS VSS.n1 3.12068
R17 Y.n3 Y.t2 256.425
R18 Y.n2 Y.n0 231.24
R19 Y.n2 Y.n1 231.03
R20 Y Y.n4 66.6553
R21 Y.n0 Y.t4 25.395
R22 Y.n0 Y.t3 25.395
R23 Y.n1 Y.t1 25.395
R24 Y.n1 Y.t5 25.395
R25 Y.n4 Y.t6 19.8005
R26 Y.n4 Y.t0 19.8005
R27 Y Y.n3 0.2365
R28 Y.n3 Y.n2 0.145237
R29 VDD.n7 VDD.t1 220.395
R30 VDD.n5 VDD.n4 195
R31 VDD.n3 VDD.n2 195
R32 VDD.t10 VDD.t11 158.06
R33 VDD.t14 VDD.t10 158.06
R34 VDD.t13 VDD.t14 158.06
R35 VDD.t12 VDD.t13 158.06
R36 VDD.t2 VDD.t12 158.06
R37 VDD.t4 VDD.t2 158.06
R38 VDD.t8 VDD.t4 158.06
R39 VDD.t6 VDD.t0 158.06
R40 VDD.n3 VDD.n0 102.978
R41 VDD.n8 VDD.n7 102.266
R42 VDD.n1 VDD.t8 87.2622
R43 VDD.n5 VDD.n0 75.6711
R44 VDD.n8 VDD.n1 74.0005
R45 VDD.n1 VDD.t6 70.7977
R46 VDD.n7 VDD.n6 36.2404
R47 VDD.n6 VDD.n3 36.2404
R48 VDD.n6 VDD.n5 36.0299
R49 VDD.n2 VDD.t3 25.395
R50 VDD.n2 VDD.t5 25.395
R51 VDD.n4 VDD.t9 25.395
R52 VDD.n4 VDD.t7 25.395
R53 VDD VDD.n8 1.87165
R54 VDD.n8 VDD.n0 0.711611
R55 a_128_103.n1 a_128_103.n5 231.24
R56 a_128_103.n0 a_128_103.n2 231.24
R57 a_128_103.n1 a_128_103.n4 231.03
R58 a_128_103.n0 a_128_103.n3 231.03
R59 a_128_103.n6 a_128_103.n1 231.03
R60 a_128_103.n5 a_128_103.t3 25.395
R61 a_128_103.n5 a_128_103.t0 25.395
R62 a_128_103.n4 a_128_103.t7 25.395
R63 a_128_103.n4 a_128_103.t1 25.395
R64 a_128_103.n3 a_128_103.t9 25.395
R65 a_128_103.n3 a_128_103.t8 25.395
R66 a_128_103.n2 a_128_103.t6 25.395
R67 a_128_103.n2 a_128_103.t5 25.395
R68 a_128_103.n6 a_128_103.t2 25.395
R69 a_128_103.t4 a_128_103.n6 25.395
R70 a_128_103.n1 a_128_103.n0 0.421553
R71 B.n0 B.t3 312.599
R72 B.n3 B.t0 247.428
R73 B.n0 B.t4 247.428
R74 B.n1 B.t2 247.428
R75 B.n2 B.t1 247.428
R76 B.n4 B.t5 229.754
R77 B B.n4 162.262
R78 B.n4 B.n3 91.5805
R79 B.n1 B.n0 65.1723
R80 B.n2 B.n1 65.1723
R81 B.n3 B.n2 65.1723
C0 A VDD 0.60147f
C1 B VDD 0.007635f
C2 A Y 0.013854f
C3 B Y 0.252442f
C4 B A 0.608892f
C5 Y VDD 0.069015f
C6 Y VSS 0.833364f
C7 B VSS 0.544323f
C8 A VSS 0.38021f
C9 VDD VSS 2.13317f
.ends

