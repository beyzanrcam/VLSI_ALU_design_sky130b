magic
tech sky130B
magscale 1 2
timestamp 1733082494
<< error_p >>
rect -773 -278 773 312
<< nwell >>
rect -773 -278 773 312
<< pmos >>
rect -679 -178 -619 250
rect -561 -178 -501 250
rect -443 -178 -383 250
rect -325 -178 -265 250
rect -207 -178 -147 250
rect -89 -178 -29 250
rect 29 -178 89 250
rect 147 -178 207 250
rect 265 -178 325 250
rect 383 -178 443 250
rect 501 -178 561 250
rect 619 -178 679 250
<< pdiff >>
rect -737 238 -679 250
rect -737 -166 -725 238
rect -691 -166 -679 238
rect -737 -178 -679 -166
rect -619 -178 -561 250
rect -501 238 -443 250
rect -501 -166 -489 238
rect -455 -166 -443 238
rect -501 -178 -443 -166
rect -383 -178 -325 250
rect -265 238 -207 250
rect -265 -166 -253 238
rect -219 -166 -207 238
rect -265 -178 -207 -166
rect -147 -178 -89 250
rect -29 238 29 250
rect -29 -166 -17 238
rect 17 -166 29 238
rect -29 -178 29 -166
rect 89 -178 147 250
rect 207 238 265 250
rect 207 -166 219 238
rect 253 -166 265 238
rect 207 -178 265 -166
rect 325 -178 383 250
rect 443 238 501 250
rect 443 -166 455 238
rect 489 -166 501 238
rect 443 -178 501 -166
rect 561 -178 619 250
rect 679 238 737 250
rect 679 -166 691 238
rect 725 -166 737 238
rect 679 -178 737 -166
<< pdiffc >>
rect -725 -166 -691 238
rect -489 -166 -455 238
rect -253 -166 -219 238
rect -17 -166 17 238
rect 219 -166 253 238
rect 455 -166 489 238
rect 691 -166 725 238
<< poly >>
rect -679 250 -619 276
rect -561 250 -501 276
rect -443 250 -383 276
rect -325 250 -265 276
rect -207 250 -147 276
rect -89 250 -29 276
rect 29 250 89 276
rect 147 250 207 276
rect 265 250 325 276
rect 383 250 443 276
rect 501 250 561 276
rect 619 250 679 276
rect -679 -209 -619 -178
rect -561 -209 -501 -178
rect -443 -209 -383 -178
rect -325 -209 -265 -178
rect -207 -209 -147 -178
rect -89 -209 -29 -178
rect 29 -209 89 -178
rect 147 -209 207 -178
rect 265 -209 325 -178
rect 383 -209 443 -178
rect 501 -209 561 -178
rect 619 -209 679 -178
rect -682 -225 -616 -209
rect -682 -259 -666 -225
rect -632 -259 -616 -225
rect -682 -275 -616 -259
rect -564 -225 -498 -209
rect -564 -259 -548 -225
rect -514 -259 -498 -225
rect -564 -275 -498 -259
rect -446 -225 -380 -209
rect -446 -259 -430 -225
rect -396 -259 -380 -225
rect -446 -275 -380 -259
rect -328 -225 -262 -209
rect -328 -259 -312 -225
rect -278 -259 -262 -225
rect -328 -275 -262 -259
rect -210 -225 -144 -209
rect -210 -259 -194 -225
rect -160 -259 -144 -225
rect -210 -275 -144 -259
rect -92 -225 -26 -209
rect -92 -259 -76 -225
rect -42 -259 -26 -225
rect -92 -275 -26 -259
rect 26 -225 92 -209
rect 26 -259 42 -225
rect 76 -259 92 -225
rect 26 -275 92 -259
rect 144 -225 210 -209
rect 144 -259 160 -225
rect 194 -259 210 -225
rect 144 -275 210 -259
rect 262 -225 328 -209
rect 262 -259 278 -225
rect 312 -259 328 -225
rect 262 -275 328 -259
rect 380 -225 446 -209
rect 380 -259 396 -225
rect 430 -259 446 -225
rect 380 -275 446 -259
rect 498 -225 564 -209
rect 498 -259 514 -225
rect 548 -259 564 -225
rect 498 -275 564 -259
rect 616 -225 682 -209
rect 616 -259 632 -225
rect 666 -259 682 -225
rect 616 -275 682 -259
<< polycont >>
rect -666 -259 -632 -225
rect -548 -259 -514 -225
rect -430 -259 -396 -225
rect -312 -259 -278 -225
rect -194 -259 -160 -225
rect -76 -259 -42 -225
rect 42 -259 76 -225
rect 160 -259 194 -225
rect 278 -259 312 -225
rect 396 -259 430 -225
rect 514 -259 548 -225
rect 632 -259 666 -225
<< locali >>
rect -725 238 -691 254
rect -725 -182 -691 -166
rect -489 238 -455 254
rect -489 -182 -455 -166
rect -253 238 -219 254
rect -253 -182 -219 -166
rect -17 238 17 254
rect -17 -182 17 -166
rect 219 238 253 254
rect 219 -182 253 -166
rect 455 238 489 254
rect 455 -182 489 -166
rect 691 238 725 254
rect 691 -182 725 -166
rect -682 -259 -666 -225
rect -632 -259 -616 -225
rect -564 -259 -548 -225
rect -514 -259 -498 -225
rect -446 -259 -430 -225
rect -396 -259 -380 -225
rect -328 -259 -312 -225
rect -278 -259 -262 -225
rect -210 -259 -194 -225
rect -160 -259 -144 -225
rect -92 -259 -76 -225
rect -42 -259 -26 -225
rect 26 -259 42 -225
rect 76 -259 92 -225
rect 144 -259 160 -225
rect 194 -259 210 -225
rect 262 -259 278 -225
rect 312 -259 328 -225
rect 380 -259 396 -225
rect 430 -259 446 -225
rect 498 -259 514 -225
rect 548 -259 564 -225
rect 616 -259 632 -225
rect 666 -259 682 -225
<< viali >>
rect -725 65 -691 238
rect -489 -166 -455 6
rect -253 65 -219 238
rect -17 -166 17 6
rect 219 65 253 238
rect 455 -166 489 6
rect 691 65 725 238
<< metal1 >>
rect -731 238 -685 250
rect -731 65 -725 238
rect -691 65 -685 238
rect -259 238 -213 250
rect -259 65 -253 238
rect -219 65 -213 238
rect 213 238 259 250
rect 213 65 219 238
rect 253 65 259 238
rect 685 238 731 250
rect 685 65 691 238
rect 725 65 731 238
rect -495 -166 -489 6
rect -455 -166 -449 6
rect -495 -178 -449 -166
rect -23 -166 -17 6
rect 17 -166 23 6
rect -23 -178 23 -166
rect 449 -166 455 6
rect 489 -166 495 6
rect 449 -178 495 -166
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.14 l 0.30 m 1 nf 12 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
