magic
tech sky130B
magscale 1 2
timestamp 1736620191
<< nwell >>
rect 6413 2450 6512 2634
rect 9708 2491 9799 2635
rect -3594 2381 -2393 2416
rect -3594 1895 -2415 2381
rect -1868 1895 -689 2416
rect -3594 603 -2415 1124
rect -1868 603 -689 1124
<< nmos >>
rect -1598 1735 -1198 1765
rect -965 1739 -765 1769
rect -1598 1639 -1198 1669
rect -3324 443 -2924 473
rect -2691 447 -2491 477
rect -1598 443 -1198 473
rect -965 447 -765 477
rect -3324 347 -2924 377
rect -1598 347 -1198 377
<< pmos >>
rect -1770 1957 -1740 2171
rect -1674 1957 -1644 2171
rect -1578 1957 -1548 2171
rect -1482 1957 -1452 2171
rect -1386 1957 -1356 2171
rect -1290 1957 -1260 2171
rect -965 2185 -751 2215
rect -965 2089 -751 2119
rect -965 1993 -751 2023
rect -3496 665 -3466 879
rect -3400 665 -3370 879
rect -3304 665 -3274 879
rect -3208 665 -3178 879
rect -3112 665 -3082 879
rect -3016 665 -2986 879
rect -2691 893 -2477 923
rect -2691 797 -2477 827
rect -2691 701 -2477 731
rect -1770 665 -1740 879
rect -1674 665 -1644 879
rect -1578 665 -1548 879
rect -1482 665 -1452 879
rect -1386 665 -1356 879
rect -1290 665 -1260 879
rect -965 893 -751 923
rect -965 797 -751 827
rect -965 701 -751 731
<< ndiff >>
rect -1598 1815 -1198 1827
rect -1598 1781 -1586 1815
rect -1210 1781 -1198 1815
rect -965 1815 -765 1827
rect -1598 1765 -1198 1781
rect -965 1781 -953 1815
rect -777 1781 -765 1815
rect -965 1769 -765 1781
rect -1598 1669 -1198 1735
rect -965 1727 -765 1739
rect -965 1693 -953 1727
rect -777 1693 -765 1727
rect -965 1681 -765 1693
rect -1598 1623 -1198 1639
rect -1598 1589 -1586 1623
rect -1210 1589 -1198 1623
rect -1598 1577 -1198 1589
rect -3324 523 -2924 535
rect -3324 489 -3312 523
rect -2936 489 -2924 523
rect -2691 523 -2491 535
rect -3324 473 -2924 489
rect -2691 489 -2679 523
rect -2503 489 -2491 523
rect -2691 477 -2491 489
rect -3324 377 -2924 443
rect -2691 435 -2491 447
rect -2691 401 -2679 435
rect -2503 401 -2491 435
rect -2691 389 -2491 401
rect -1598 523 -1198 535
rect -1598 489 -1586 523
rect -1210 489 -1198 523
rect -965 523 -765 535
rect -1598 473 -1198 489
rect -965 489 -953 523
rect -777 489 -765 523
rect -965 477 -765 489
rect -1598 377 -1198 443
rect -965 435 -765 447
rect -965 401 -953 435
rect -777 401 -765 435
rect -965 389 -765 401
rect -3324 331 -2924 347
rect -3324 297 -3312 331
rect -2936 297 -2924 331
rect -1598 331 -1198 347
rect -3324 285 -2924 297
rect -1598 297 -1586 331
rect -1210 297 -1198 331
rect -1598 285 -1198 297
<< pdiff >>
rect -965 2265 -751 2277
rect -1832 2159 -1770 2171
rect -1832 1969 -1820 2159
rect -1786 1969 -1770 2159
rect -1832 1957 -1770 1969
rect -1740 2159 -1674 2171
rect -1740 1969 -1724 2159
rect -1690 1969 -1674 2159
rect -1740 1957 -1674 1969
rect -1644 2159 -1578 2171
rect -1644 1969 -1628 2159
rect -1594 1969 -1578 2159
rect -1644 1957 -1578 1969
rect -1548 2159 -1482 2171
rect -1548 1969 -1532 2159
rect -1498 1969 -1482 2159
rect -1548 1957 -1482 1969
rect -1452 2159 -1386 2171
rect -1452 1969 -1436 2159
rect -1402 1969 -1386 2159
rect -1452 1957 -1386 1969
rect -1356 2159 -1290 2171
rect -1356 1969 -1340 2159
rect -1306 1969 -1290 2159
rect -1356 1957 -1290 1969
rect -1260 2159 -1198 2171
rect -1260 1969 -1244 2159
rect -1210 1969 -1198 2159
rect -965 2231 -953 2265
rect -763 2231 -751 2265
rect -965 2215 -751 2231
rect -965 2169 -751 2185
rect -965 2135 -953 2169
rect -759 2135 -751 2169
rect -965 2119 -751 2135
rect -965 2073 -751 2089
rect -965 2039 -953 2073
rect -763 2039 -751 2073
rect -965 2023 -751 2039
rect -965 1977 -751 1993
rect -1260 1957 -1198 1969
rect -965 1943 -953 1977
rect -759 1943 -751 1977
rect -965 1931 -751 1943
rect -2691 973 -2477 985
rect -3558 867 -3496 879
rect -3558 677 -3546 867
rect -3512 677 -3496 867
rect -3558 665 -3496 677
rect -3466 867 -3400 879
rect -3466 677 -3450 867
rect -3416 677 -3400 867
rect -3466 665 -3400 677
rect -3370 867 -3304 879
rect -3370 677 -3354 867
rect -3320 677 -3304 867
rect -3370 665 -3304 677
rect -3274 867 -3208 879
rect -3274 677 -3258 867
rect -3224 677 -3208 867
rect -3274 665 -3208 677
rect -3178 867 -3112 879
rect -3178 677 -3162 867
rect -3128 677 -3112 867
rect -3178 665 -3112 677
rect -3082 867 -3016 879
rect -3082 677 -3066 867
rect -3032 677 -3016 867
rect -3082 665 -3016 677
rect -2986 867 -2924 879
rect -2986 677 -2970 867
rect -2936 677 -2924 867
rect -2691 939 -2679 973
rect -2489 939 -2477 973
rect -2691 923 -2477 939
rect -965 973 -751 985
rect -2691 877 -2477 893
rect -2691 843 -2679 877
rect -2485 843 -2477 877
rect -2691 827 -2477 843
rect -1832 867 -1770 879
rect -2691 781 -2477 797
rect -2691 747 -2679 781
rect -2489 747 -2477 781
rect -2691 731 -2477 747
rect -2691 685 -2477 701
rect -2986 665 -2924 677
rect -2691 651 -2679 685
rect -2485 651 -2477 685
rect -1832 677 -1820 867
rect -1786 677 -1770 867
rect -1832 665 -1770 677
rect -1740 867 -1674 879
rect -1740 677 -1724 867
rect -1690 677 -1674 867
rect -1740 665 -1674 677
rect -1644 867 -1578 879
rect -1644 677 -1628 867
rect -1594 677 -1578 867
rect -1644 665 -1578 677
rect -1548 867 -1482 879
rect -1548 677 -1532 867
rect -1498 677 -1482 867
rect -1548 665 -1482 677
rect -1452 867 -1386 879
rect -1452 677 -1436 867
rect -1402 677 -1386 867
rect -1452 665 -1386 677
rect -1356 867 -1290 879
rect -1356 677 -1340 867
rect -1306 677 -1290 867
rect -1356 665 -1290 677
rect -1260 867 -1198 879
rect -1260 677 -1244 867
rect -1210 677 -1198 867
rect -965 939 -953 973
rect -763 939 -751 973
rect -965 923 -751 939
rect -965 877 -751 893
rect -965 843 -953 877
rect -759 843 -751 877
rect -965 827 -751 843
rect -965 781 -751 797
rect -965 747 -953 781
rect -763 747 -751 781
rect -965 731 -751 747
rect -965 685 -751 701
rect -1260 665 -1198 677
rect -2691 639 -2477 651
rect -965 651 -953 685
rect -759 651 -751 685
rect -965 639 -751 651
<< ndiffc >>
rect -1586 1781 -1210 1815
rect -953 1781 -777 1815
rect -953 1693 -777 1727
rect -1586 1589 -1210 1623
rect -3312 489 -2936 523
rect -2679 489 -2503 523
rect -2679 401 -2503 435
rect -1586 489 -1210 523
rect -953 489 -777 523
rect -953 401 -777 435
rect -3312 297 -2936 331
rect -1586 297 -1210 331
<< pdiffc >>
rect -1820 1969 -1786 2159
rect -1724 1969 -1690 2159
rect -1628 1969 -1594 2159
rect -1532 1969 -1498 2159
rect -1436 1969 -1402 2159
rect -1340 1969 -1306 2159
rect -1244 1969 -1210 2159
rect -953 2231 -763 2265
rect -953 2135 -759 2169
rect -953 2039 -763 2073
rect -953 1943 -759 1977
rect -3546 677 -3512 867
rect -3450 677 -3416 867
rect -3354 677 -3320 867
rect -3258 677 -3224 867
rect -3162 677 -3128 867
rect -3066 677 -3032 867
rect -2970 677 -2936 867
rect -2679 939 -2489 973
rect -2679 843 -2485 877
rect -2679 747 -2489 781
rect -2679 651 -2485 685
rect -1820 677 -1786 867
rect -1724 677 -1690 867
rect -1628 677 -1594 867
rect -1532 677 -1498 867
rect -1436 677 -1402 867
rect -1340 677 -1306 867
rect -1244 677 -1210 867
rect -953 939 -763 973
rect -953 843 -759 877
rect -953 747 -763 781
rect -953 651 -759 685
<< psubdiff >>
rect -1598 1553 -1198 1577
rect -1598 1479 -1571 1553
rect -1236 1479 -1198 1553
rect -1598 1460 -1198 1479
rect -3324 261 -2924 285
rect -3324 187 -3297 261
rect -2962 187 -2924 261
rect -3324 168 -2924 187
rect -1598 261 -1198 285
rect -1598 187 -1571 261
rect -1236 187 -1198 261
rect -1598 168 -1198 187
<< nsubdiff >>
rect -1828 2314 -1211 2375
rect -1828 2267 -1618 2314
rect -1378 2267 -1211 2314
rect -1828 2225 -1211 2267
rect -3554 1022 -2937 1083
rect -3554 975 -3344 1022
rect -3104 975 -2937 1022
rect -1828 1022 -1211 1083
rect -3554 933 -2937 975
rect -1828 975 -1618 1022
rect -1378 975 -1211 1022
rect -1828 933 -1211 975
<< psubdiffcont >>
rect -1571 1479 -1236 1553
rect -3297 187 -2962 261
rect -1571 187 -1236 261
<< nsubdiffcont >>
rect -1618 2267 -1378 2314
rect -3344 975 -3104 1022
rect -1618 975 -1378 1022
<< poly >>
rect -1062 2217 -996 2233
rect -1770 2171 -1740 2202
rect -1674 2171 -1644 2202
rect -1578 2171 -1548 2202
rect -1482 2171 -1452 2202
rect -1386 2171 -1356 2202
rect -1290 2171 -1260 2202
rect -1062 1991 -1046 2217
rect -1012 2215 -996 2217
rect -1012 2185 -965 2215
rect -751 2185 -725 2215
rect -1012 2119 -996 2185
rect -1012 2089 -965 2119
rect -751 2089 -725 2119
rect -1012 2023 -996 2089
rect -1012 1993 -965 2023
rect -751 1993 -725 2023
rect -1012 1991 -996 1993
rect -1062 1975 -996 1991
rect -1770 1931 -1740 1957
rect -1674 1931 -1644 1957
rect -1578 1931 -1548 1957
rect -1771 1910 -1548 1931
rect -1771 1875 -1754 1910
rect -1720 1901 -1548 1910
rect -1482 1931 -1452 1957
rect -1386 1931 -1356 1957
rect -1290 1931 -1260 1957
rect -1482 1910 -1260 1931
rect -1720 1875 -1704 1901
rect -1771 1864 -1704 1875
rect -1482 1875 -1465 1910
rect -1431 1901 -1260 1910
rect -1431 1875 -1415 1901
rect -1482 1864 -1415 1875
rect -1771 1669 -1728 1864
rect -1686 1786 -1620 1802
rect -1686 1751 -1670 1786
rect -1636 1765 -1620 1786
rect -1062 1771 -995 1787
rect -1636 1751 -1598 1765
rect -1686 1735 -1598 1751
rect -1198 1735 -1172 1765
rect -1062 1737 -1046 1771
rect -1012 1769 -995 1771
rect -1012 1739 -965 1769
rect -765 1739 -739 1769
rect -1012 1737 -995 1739
rect -1062 1721 -995 1737
rect -1771 1653 -1598 1669
rect -1771 1618 -1670 1653
rect -1636 1639 -1598 1653
rect -1198 1639 -1172 1669
rect -1636 1618 -1620 1639
rect -1771 1602 -1620 1618
rect -2788 925 -2722 941
rect -3496 879 -3466 910
rect -3400 879 -3370 910
rect -3304 879 -3274 910
rect -3208 879 -3178 910
rect -3112 879 -3082 910
rect -3016 879 -2986 910
rect -2788 699 -2772 925
rect -2738 923 -2722 925
rect -1062 925 -996 941
rect -2738 893 -2691 923
rect -2477 893 -2451 923
rect -2738 827 -2722 893
rect -1770 879 -1740 910
rect -1674 879 -1644 910
rect -1578 879 -1548 910
rect -1482 879 -1452 910
rect -1386 879 -1356 910
rect -1290 879 -1260 910
rect -2738 797 -2691 827
rect -2477 797 -2451 827
rect -2738 731 -2722 797
rect -2738 701 -2691 731
rect -2477 701 -2451 731
rect -2738 699 -2722 701
rect -2788 683 -2722 699
rect -3496 639 -3466 665
rect -3400 639 -3370 665
rect -3304 639 -3274 665
rect -3497 618 -3274 639
rect -3497 583 -3480 618
rect -3446 609 -3274 618
rect -3208 639 -3178 665
rect -3112 639 -3082 665
rect -3016 639 -2986 665
rect -1062 699 -1046 925
rect -1012 923 -996 925
rect -1012 893 -965 923
rect -751 893 -725 923
rect -1012 827 -996 893
rect -1012 797 -965 827
rect -751 797 -725 827
rect -1012 731 -996 797
rect -1012 701 -965 731
rect -751 701 -725 731
rect -1012 699 -996 701
rect -1062 683 -996 699
rect -1770 639 -1740 665
rect -1674 639 -1644 665
rect -1578 639 -1548 665
rect -3208 618 -2986 639
rect -3446 583 -3430 609
rect -3497 572 -3430 583
rect -3208 583 -3191 618
rect -3157 609 -2986 618
rect -1771 618 -1548 639
rect -3157 583 -3141 609
rect -3208 572 -3141 583
rect -1771 583 -1754 618
rect -1720 609 -1548 618
rect -1482 639 -1452 665
rect -1386 639 -1356 665
rect -1290 639 -1260 665
rect -1482 618 -1260 639
rect -1720 583 -1704 609
rect -1771 572 -1704 583
rect -1482 583 -1465 618
rect -1431 609 -1260 618
rect -1431 583 -1415 609
rect -1482 572 -1415 583
rect -3497 377 -3454 572
rect -3412 494 -3346 510
rect -3412 459 -3396 494
rect -3362 473 -3346 494
rect -2788 479 -2721 495
rect -3362 459 -3324 473
rect -3412 443 -3324 459
rect -2924 443 -2898 473
rect -2788 445 -2772 479
rect -2738 477 -2721 479
rect -2738 447 -2691 477
rect -2491 447 -2465 477
rect -2738 445 -2721 447
rect -2788 429 -2721 445
rect -1771 377 -1728 572
rect -1686 494 -1620 510
rect -1686 459 -1670 494
rect -1636 473 -1620 494
rect -1062 479 -995 495
rect -1636 459 -1598 473
rect -1686 443 -1598 459
rect -1198 443 -1172 473
rect -1062 445 -1046 479
rect -1012 477 -995 479
rect -1012 447 -965 477
rect -765 447 -739 477
rect -1012 445 -995 447
rect -1062 429 -995 445
rect -3497 361 -3324 377
rect -3497 326 -3396 361
rect -3362 347 -3324 361
rect -2924 347 -2898 377
rect -1771 361 -1598 377
rect -3362 326 -3346 347
rect -3497 310 -3346 326
rect -1771 326 -1670 361
rect -1636 347 -1598 361
rect -1198 347 -1172 377
rect -1636 326 -1620 347
rect -1771 310 -1620 326
<< polycont >>
rect -1046 1991 -1012 2217
rect -1754 1875 -1720 1910
rect -1465 1875 -1431 1910
rect -1670 1751 -1636 1786
rect -1046 1737 -1012 1771
rect -1670 1618 -1636 1653
rect -2772 699 -2738 925
rect -3480 583 -3446 618
rect -1046 699 -1012 925
rect -3191 583 -3157 618
rect -1754 583 -1720 618
rect -1465 583 -1431 618
rect -3396 459 -3362 494
rect -2772 445 -2738 479
rect -1670 459 -1636 494
rect -1046 445 -1012 479
rect -3396 326 -3362 361
rect -1670 326 -1636 361
<< locali >>
rect -1692 2267 -1618 2314
rect -1378 2267 -1278 2314
rect -1062 2217 -1012 2234
rect -969 2231 -959 2265
rect -763 2231 -747 2265
rect -1820 2165 -1786 2175
rect -1820 1953 -1786 1969
rect -1724 2159 -1690 2175
rect -1724 1953 -1690 1963
rect -1628 2165 -1594 2175
rect -1628 1953 -1594 1969
rect -1532 2159 -1498 2175
rect -1532 1953 -1498 1963
rect -1436 2165 -1402 2175
rect -1436 1953 -1402 1969
rect -1340 2159 -1306 2175
rect -1340 1953 -1306 1963
rect -1244 2165 -1210 2175
rect -1244 1953 -1210 1969
rect -1062 1991 -1046 2217
rect -969 2135 -953 2169
rect -759 2135 -741 2169
rect -969 2039 -959 2073
rect -763 2039 -747 2073
rect -1771 1875 -1754 1910
rect -1720 1875 -1704 1910
rect -1482 1904 -1465 1910
rect -1670 1875 -1465 1904
rect -1431 1875 -1415 1910
rect -1771 1669 -1728 1875
rect -1670 1870 -1415 1875
rect -1670 1786 -1636 1870
rect -1602 1781 -1586 1815
rect -1210 1781 -1194 1815
rect -1670 1735 -1636 1751
rect -1062 1771 -1012 1991
rect -969 1943 -953 1977
rect -759 1943 -741 1977
rect -969 1781 -953 1815
rect -777 1781 -761 1815
rect -1062 1737 -1046 1771
rect -1062 1721 -1012 1737
rect -969 1693 -953 1727
rect -777 1693 -761 1727
rect -1771 1653 -1636 1669
rect -1771 1618 -1670 1653
rect -1771 1602 -1636 1618
rect -1602 1589 -1586 1623
rect -1210 1589 -1194 1623
rect -1598 1479 -1571 1553
rect -1236 1479 -1198 1553
rect -3418 975 -3344 1022
rect -3104 975 -3004 1022
rect -1692 975 -1618 1022
rect -1378 975 -1278 1022
rect -2788 925 -2738 942
rect -2695 939 -2685 973
rect -2489 939 -2473 973
rect -3546 873 -3512 883
rect -3546 661 -3512 677
rect -3450 867 -3416 883
rect -3450 661 -3416 671
rect -3354 873 -3320 883
rect -3354 661 -3320 677
rect -3258 867 -3224 883
rect -3258 661 -3224 671
rect -3162 873 -3128 883
rect -3162 661 -3128 677
rect -3066 867 -3032 883
rect -3066 661 -3032 671
rect -2970 873 -2936 883
rect -2970 661 -2936 677
rect -2788 699 -2772 925
rect -1062 925 -1012 942
rect -969 939 -959 973
rect -763 939 -747 973
rect -2695 843 -2679 877
rect -2485 843 -2467 877
rect -1820 873 -1786 883
rect -2695 747 -2685 781
rect -2489 747 -2473 781
rect -3497 583 -3480 618
rect -3446 583 -3430 618
rect -3208 612 -3191 618
rect -3396 583 -3191 612
rect -3157 583 -3141 618
rect -3497 377 -3454 583
rect -3396 578 -3141 583
rect -3396 494 -3362 578
rect -3328 489 -3312 523
rect -2936 489 -2920 523
rect -3396 443 -3362 459
rect -2788 479 -2738 699
rect -2695 651 -2679 685
rect -2485 651 -2467 685
rect -1820 661 -1786 677
rect -1724 867 -1690 883
rect -1724 661 -1690 671
rect -1628 873 -1594 883
rect -1628 661 -1594 677
rect -1532 867 -1498 883
rect -1532 661 -1498 671
rect -1436 873 -1402 883
rect -1436 661 -1402 677
rect -1340 867 -1306 883
rect -1340 661 -1306 671
rect -1244 873 -1210 883
rect -1244 661 -1210 677
rect -1062 699 -1046 925
rect -969 843 -953 877
rect -759 843 -741 877
rect -969 747 -959 781
rect -763 747 -747 781
rect -1771 583 -1754 618
rect -1720 583 -1704 618
rect -1482 612 -1465 618
rect -1670 583 -1465 612
rect -1431 583 -1415 618
rect -2695 489 -2679 523
rect -2503 489 -2487 523
rect -2788 445 -2772 479
rect -2788 429 -2738 445
rect -2695 401 -2679 435
rect -2503 401 -2487 435
rect -1771 377 -1728 583
rect -1670 578 -1415 583
rect -1670 494 -1636 578
rect -1602 489 -1586 523
rect -1210 489 -1194 523
rect -1670 443 -1636 459
rect -1062 479 -1012 699
rect -969 651 -953 685
rect -759 651 -741 685
rect -969 489 -953 523
rect -777 489 -761 523
rect -1062 445 -1046 479
rect -1062 429 -1012 445
rect -969 401 -953 435
rect -777 401 -761 435
rect -3497 361 -3362 377
rect -3497 326 -3396 361
rect -1771 361 -1636 377
rect -3497 310 -3362 326
rect -3328 297 -3312 331
rect -2936 297 -2920 331
rect -1771 326 -1670 361
rect -1771 310 -1636 326
rect -1602 297 -1586 331
rect -1210 297 -1194 331
rect -3324 187 -3297 261
rect -2962 187 -2924 261
rect -1598 187 -1571 261
rect -1236 187 -1198 261
<< viali >>
rect -1618 2267 -1378 2314
rect -959 2231 -953 2265
rect -953 2231 -880 2265
rect -1820 2159 -1786 2165
rect -1820 2085 -1786 2159
rect -1724 1969 -1690 2043
rect -1724 1963 -1690 1969
rect -1628 2159 -1594 2165
rect -1628 2085 -1594 2159
rect -1532 1969 -1498 2043
rect -1532 1963 -1498 1969
rect -1436 2159 -1402 2165
rect -1436 2085 -1402 2159
rect -1340 1969 -1306 2043
rect -1340 1963 -1306 1969
rect -1244 2159 -1210 2165
rect -1244 2085 -1210 2159
rect -1046 1991 -1012 2217
rect -836 2135 -759 2169
rect -959 2039 -953 2073
rect -953 2039 -880 2073
rect -1754 1875 -1720 1910
rect -1465 1875 -1431 1910
rect -1670 1751 -1636 1786
rect -1586 1781 -1210 1815
rect -836 1943 -759 1977
rect -953 1781 -777 1815
rect -1046 1737 -1012 1771
rect -953 1693 -777 1727
rect -1586 1589 -1210 1623
rect -1571 1479 -1236 1548
rect -3344 975 -3104 1022
rect -1618 975 -1378 1022
rect -2685 939 -2679 973
rect -2679 939 -2606 973
rect -3546 867 -3512 873
rect -3546 793 -3512 867
rect -3450 677 -3416 751
rect -3450 671 -3416 677
rect -3354 867 -3320 873
rect -3354 793 -3320 867
rect -3258 677 -3224 751
rect -3258 671 -3224 677
rect -3162 867 -3128 873
rect -3162 793 -3128 867
rect -3066 677 -3032 751
rect -3066 671 -3032 677
rect -2970 867 -2936 873
rect -2970 793 -2936 867
rect -2772 699 -2738 925
rect -959 939 -953 973
rect -953 939 -880 973
rect -2562 843 -2485 877
rect -1820 867 -1786 873
rect -1820 793 -1786 867
rect -2685 747 -2679 781
rect -2679 747 -2606 781
rect -3480 583 -3446 618
rect -3191 583 -3157 618
rect -3396 459 -3362 494
rect -3312 489 -2936 523
rect -2562 651 -2485 685
rect -1724 677 -1690 751
rect -1724 671 -1690 677
rect -1628 867 -1594 873
rect -1628 793 -1594 867
rect -1532 677 -1498 751
rect -1532 671 -1498 677
rect -1436 867 -1402 873
rect -1436 793 -1402 867
rect -1340 677 -1306 751
rect -1340 671 -1306 677
rect -1244 867 -1210 873
rect -1244 793 -1210 867
rect -1046 699 -1012 925
rect -836 843 -759 877
rect -959 747 -953 781
rect -953 747 -880 781
rect -1754 583 -1720 618
rect -1465 583 -1431 618
rect -2679 489 -2503 523
rect -2772 445 -2738 479
rect -2679 401 -2503 435
rect -1670 459 -1636 494
rect -1586 489 -1210 523
rect -836 651 -759 685
rect -953 489 -777 523
rect -1046 445 -1012 479
rect -953 401 -777 435
rect -3312 297 -2936 331
rect -1586 297 -1210 331
rect -3297 187 -2962 256
rect -1571 187 -1236 256
<< metal1 >>
rect -2397 3005 9807 3089
rect -2397 2233 -2284 3005
rect -2496 2103 -2284 2233
rect -2215 2858 6517 2942
rect -3989 1793 -3594 1928
rect -2888 1775 -2805 2049
rect -3418 1022 -3081 1034
rect -3418 975 -3344 1022
rect -3104 975 -3081 1022
rect -3418 915 -3081 975
rect -2695 973 -2473 1021
rect -2695 969 -2685 973
rect -2805 925 -2722 941
rect -3559 879 -2925 915
rect -3559 873 -2924 879
rect -3559 793 -3546 873
rect -3512 793 -3354 873
rect -3320 793 -3162 873
rect -3128 793 -2970 873
rect -2936 793 -2924 873
rect -3559 787 -2924 793
rect -3559 786 -2925 787
rect -2805 757 -2772 925
rect -3466 751 -2772 757
rect -3466 671 -3450 751
rect -3416 671 -3258 751
rect -3224 671 -3066 751
rect -3032 699 -2772 751
rect -2738 699 -2722 925
rect -2691 939 -2685 969
rect -2606 969 -2473 973
rect -2606 939 -2600 969
rect -2691 781 -2600 939
rect -2691 747 -2685 781
rect -2606 747 -2600 781
rect -2691 731 -2600 747
rect -2568 877 -2415 941
rect -2568 843 -2562 877
rect -2485 843 -2415 877
rect -3032 671 -2722 699
rect -2568 685 -2415 843
rect -3466 665 -2722 671
rect -3594 618 -3430 636
rect -3594 616 -3480 618
rect -3594 506 -3569 616
rect -3446 583 -3430 618
rect -3474 506 -3430 583
rect -3594 501 -3430 506
rect -3402 618 -3142 637
rect -3402 583 -3191 618
rect -3157 583 -3142 618
rect -3402 563 -3142 583
rect -3402 494 -3352 563
rect -3066 535 -2722 665
rect -3402 472 -3396 494
rect -3764 459 -3396 472
rect -3362 459 -3352 494
rect -3324 523 -2722 535
rect -3324 489 -3312 523
rect -2936 489 -2722 523
rect -3324 483 -2722 489
rect -2691 651 -2562 685
rect -2485 651 -2415 685
rect -2691 616 -2415 651
rect -2215 616 -2078 2858
rect -386 2710 3226 2794
rect -1692 2314 -1355 2326
rect -1692 2267 -1618 2314
rect -1378 2267 -1355 2314
rect -1692 2207 -1355 2267
rect -969 2265 -747 2313
rect -969 2261 -959 2265
rect -1079 2217 -996 2233
rect -1833 2171 -1199 2207
rect -1833 2165 -1198 2171
rect -1833 2085 -1820 2165
rect -1786 2085 -1628 2165
rect -1594 2085 -1436 2165
rect -1402 2085 -1244 2165
rect -1210 2085 -1198 2165
rect -1833 2079 -1198 2085
rect -1833 2078 -1199 2079
rect -1079 2049 -1046 2217
rect -1740 2043 -1046 2049
rect -1740 1963 -1724 2043
rect -1690 1963 -1532 2043
rect -1498 1963 -1340 2043
rect -1306 1991 -1046 2043
rect -1012 1991 -996 2217
rect -965 2231 -959 2261
rect -880 2261 -747 2265
rect -880 2231 -874 2261
rect -965 2073 -874 2231
rect -965 2039 -959 2073
rect -880 2039 -874 2073
rect -965 2023 -874 2039
rect -842 2169 -689 2233
rect -842 2135 -836 2169
rect -759 2135 -689 2169
rect -1306 1963 -996 1991
rect -842 1977 -689 2135
rect -1740 1957 -996 1963
rect -1868 1910 -1704 1928
rect -1868 1900 -1754 1910
rect -1868 1823 -1847 1900
rect -1720 1875 -1704 1910
rect -1742 1823 -1704 1875
rect -1868 1793 -1704 1823
rect -1676 1910 -1416 1929
rect -1676 1875 -1465 1910
rect -1431 1875 -1416 1910
rect -1676 1855 -1416 1875
rect -1676 1786 -1626 1855
rect -1340 1827 -996 1957
rect -1676 1764 -1670 1786
rect -1868 1751 -1670 1764
rect -1636 1751 -1626 1786
rect -1598 1815 -996 1827
rect -1598 1781 -1586 1815
rect -1210 1781 -996 1815
rect -1598 1775 -996 1781
rect -965 1943 -836 1977
rect -759 1943 -689 1977
rect -965 1867 -689 1943
rect -386 1867 -255 2710
rect 3117 2633 3226 2710
rect 3117 2538 3129 2633
rect 3218 2538 3226 2633
rect 3117 2527 3226 2538
rect 6407 2634 6517 2858
rect 6407 2450 6413 2634
rect 6512 2450 6517 2634
rect 9699 2635 9807 3005
rect 9699 2491 9708 2635
rect 9799 2491 9807 2635
rect 9699 2480 9807 2491
rect 6407 2443 6517 2450
rect -965 1815 -255 1867
rect -965 1781 -953 1815
rect -777 1781 -255 1815
rect -965 1775 -765 1781
rect -1868 1749 -1626 1751
rect -1868 1645 -1852 1749
rect -1735 1645 -1626 1749
rect -1079 1771 -996 1775
rect -1079 1737 -1046 1771
rect -1012 1737 -996 1771
rect -1079 1720 -996 1737
rect -965 1727 -765 1734
rect -965 1693 -953 1727
rect -777 1693 -765 1727
rect -737 1720 -255 1781
rect -965 1692 -765 1693
rect -969 1645 -761 1692
rect -1868 1628 -1626 1645
rect -1598 1623 -1198 1629
rect -1598 1589 -1586 1623
rect -1210 1589 -1198 1623
rect -1598 1548 -1198 1589
rect -1598 1479 -1571 1548
rect -1236 1479 -1198 1548
rect -1598 1460 -1198 1479
rect -160 1063 49 1083
rect -1692 1022 -1355 1034
rect -1692 975 -1618 1022
rect -1378 975 -1355 1022
rect -1692 915 -1355 975
rect -969 973 -747 1021
rect -969 969 -959 973
rect -1079 925 -996 941
rect -1833 879 -1199 915
rect -1833 873 -1198 879
rect -1833 793 -1820 873
rect -1786 793 -1628 873
rect -1594 793 -1436 873
rect -1402 793 -1244 873
rect -1210 793 -1198 873
rect -1833 787 -1198 793
rect -1833 786 -1199 787
rect -1079 757 -1046 925
rect -1740 751 -1046 757
rect -1740 671 -1724 751
rect -1690 671 -1532 751
rect -1498 671 -1340 751
rect -1306 699 -1046 751
rect -1012 699 -996 925
rect -965 939 -959 969
rect -880 969 -747 973
rect -880 939 -874 969
rect -160 961 -130 1063
rect -12 961 49 1063
rect -965 781 -874 939
rect -965 747 -959 781
rect -880 747 -874 781
rect -965 731 -874 747
rect -842 877 -689 941
rect -160 931 49 961
rect 3113 953 3316 1044
rect 6404 953 6607 1044
rect 9695 953 9898 1044
rect -842 843 -836 877
rect -759 843 -689 877
rect -1306 671 -996 699
rect -842 693 -689 843
rect -842 691 -604 693
rect -842 685 -433 691
rect -1740 665 -996 671
rect -2691 523 -2078 616
rect -2691 489 -2679 523
rect -2503 489 -2078 523
rect -1868 618 -1704 636
rect -1868 516 -1853 618
rect -1777 583 -1754 618
rect -1720 583 -1704 618
rect -1777 516 -1704 583
rect -1868 501 -1704 516
rect -1676 618 -1416 637
rect -1676 583 -1465 618
rect -1431 583 -1416 618
rect -1676 563 -1416 583
rect -2691 483 -2491 489
rect -3764 347 -3352 459
rect -2805 479 -2722 483
rect -2805 445 -2772 479
rect -2738 445 -2722 479
rect -2805 428 -2722 445
rect -2691 435 -2491 442
rect -2691 401 -2679 435
rect -2503 401 -2491 435
rect -2463 430 -2078 489
rect -1676 494 -1626 563
rect -1340 535 -996 665
rect -1676 472 -1670 494
rect -1868 459 -1670 472
rect -1636 459 -1626 494
rect -1598 523 -996 535
rect -1598 489 -1586 523
rect -1210 489 -996 523
rect -1598 483 -996 489
rect -965 651 -836 685
rect -759 651 -433 685
rect -965 645 -433 651
rect -965 523 -692 645
rect -965 489 -953 523
rect -777 489 -692 523
rect -965 483 -765 489
rect -1868 451 -1626 459
rect -2463 428 -2139 430
rect -2691 400 -2491 401
rect -2695 353 -2487 400
rect -1868 362 -1851 451
rect -1724 362 -1626 451
rect -1079 479 -996 483
rect -1079 445 -1046 479
rect -1012 445 -996 479
rect -1079 428 -996 445
rect -737 463 -692 489
rect -482 463 -433 645
rect -965 435 -765 442
rect -965 401 -953 435
rect -777 401 -765 435
rect -737 428 -433 463
rect -965 400 -765 401
rect -3764 149 -3739 347
rect -3593 336 -3352 347
rect -3593 149 -3503 336
rect -3324 331 -2924 337
rect -1868 336 -1626 362
rect -969 353 -761 400
rect -3324 297 -3312 331
rect -2936 297 -2924 331
rect -3324 256 -2924 297
rect -3324 187 -3297 256
rect -2962 187 -2924 256
rect -3324 168 -2924 187
rect -1598 331 -1198 337
rect -1598 297 -1586 331
rect -1210 297 -1198 331
rect -1598 256 -1198 297
rect -1598 187 -1571 256
rect -1236 187 -1198 256
rect -1598 168 -1198 187
rect -3764 134 -3503 149
rect 12934 91 12983 1042
rect 12986 953 13189 1044
rect 12441 1 12992 91
rect 12934 -3 12983 1
<< via1 >>
rect -3563 1642 -3431 1743
rect -3569 583 -3480 616
rect -3480 583 -3474 616
rect -3569 506 -3474 583
rect -1847 1875 -1754 1900
rect -1754 1875 -1742 1900
rect -1847 1823 -1742 1875
rect 3129 2538 3218 2633
rect 6413 2450 6512 2634
rect 9708 2491 9799 2635
rect -1852 1645 -1735 1749
rect -130 961 -12 1063
rect -1853 516 -1777 618
rect -1851 362 -1724 451
rect -692 463 -482 645
rect -3739 149 -3593 347
<< metal2 >>
rect -2337 1900 -1704 1928
rect -2337 1823 -1847 1900
rect -1742 1823 -1704 1900
rect -2337 1793 -1704 1823
rect -3759 1743 -3396 1764
rect -3759 1642 -3563 1743
rect -3431 1642 -3396 1743
rect -3759 1628 -3396 1642
rect -2037 1749 -1718 1764
rect -2037 1645 -1852 1749
rect -1735 1645 -1718 1749
rect -2037 1628 -1718 1645
rect -483 1633 -96 1640
rect -3759 1369 -3583 1628
rect -2037 1369 -1861 1628
rect -3761 1234 -1861 1369
rect -3759 636 -3583 1234
rect -2037 636 -1861 1234
rect -522 1500 -96 1633
rect -689 691 -604 693
rect -522 691 -431 1500
rect -737 645 -431 691
rect -3759 616 -3452 636
rect -3759 506 -3569 616
rect -3474 506 -3452 616
rect -3759 501 -3452 506
rect -2037 618 -1764 636
rect -2037 516 -1853 618
rect -1777 516 -1764 618
rect -2037 501 -1764 516
rect -2038 465 -1699 471
rect -2039 451 -1699 465
rect -3764 347 -3566 376
rect -3764 149 -3739 347
rect -3593 149 -3566 347
rect -3764 134 -3566 149
rect -2039 362 -1851 451
rect -1724 362 -1699 451
rect -737 463 -692 645
rect -482 463 -431 645
rect -737 428 -431 463
rect -166 1063 19 1079
rect -166 961 -130 1063
rect -12 961 19 1063
rect -2039 336 -1699 362
rect -2039 57 -1863 336
rect -2039 -89 -1864 57
rect -166 -125 19 961
rect 12985 16 13185 127
<< via2 >>
rect -3739 149 -3593 347
<< metal3 >>
rect -3764 347 -3566 376
rect -3764 149 -3739 347
rect -3593 149 -3566 347
rect -3764 134 -3566 149
<< metal5 >>
rect -48 -307 12985 2650
use FULL_ADDER  FULL_ADDER_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/ADDER
timestamp 1736620191
transform 1 0 118 0 1 1114
box -292 -1421 3108 1536
use FULL_ADDER  FULL_ADDER_1
timestamp 1736620191
transform 1 0 3409 0 1 1114
box -292 -1421 3108 1536
use FULL_ADDER  FULL_ADDER_2
timestamp 1736620191
transform 1 0 6700 0 1 1114
box -292 -1421 3108 1536
use FULL_ADDER  FULL_ADDER_3
timestamp 1736620191
transform 1 0 9991 0 1 1114
box -292 -1421 3108 1536
use inv  inv_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/inv
timestamp 1736620191
transform 1 0 -2805 0 1 1895
box 0 -311 412 486
use NAND2  NAND2_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/NAND/NAND2
timestamp 1736620191
transform 1 0 -3950 0 1 1523
box 356 -17 1062 804
<< labels >>
rlabel metal1 -689 1864 -689 1864 3 Y
port 3 e
rlabel metal1 -1065 1864 -1065 1864 7 A
port 2 e
rlabel metal1 -921 2313 -921 2313 1 VDD
port 1 n
rlabel metal1 -864 1645 -864 1645 5 VSS
port 4 s
rlabel metal1 -1065 572 -1065 572 7 A
port 2 e
rlabel metal1 -921 1021 -921 1021 1 VDD
port 1 n
rlabel metal1 -864 353 -864 353 5 VSS
port 4 s
rlabel metal1 -2415 572 -2415 572 3 Y
port 3 e
rlabel metal1 -2791 572 -2791 572 7 A
port 2 e
rlabel metal1 -2647 1021 -2647 1021 1 VDD
port 1 n
rlabel metal1 -2590 353 -2590 353 5 VSS
port 4 s
rlabel via1 -689 572 -689 572 3 Y
port 3 e
<< end >>
