magic
tech sky130B
magscale 1 2
timestamp 1736620191
<< metal1 >>
rect -174 3784 -65 4393
rect 2287 4268 2437 4400
rect 2518 4202 2524 4388
rect 2710 4202 2716 4388
rect 3117 3827 3226 4385
rect 5578 4259 5728 4391
rect 5810 4389 5991 4395
rect 5810 4202 5991 4208
rect 6408 3834 6517 4396
rect 8872 4270 9022 4402
rect 9108 4214 9114 4392
rect 9292 4214 9298 4392
rect 9699 3842 9808 4407
rect 12159 4268 12309 4400
rect 12385 4223 12391 4398
rect 12566 4223 12572 4398
rect 3111 3823 3232 3827
rect -180 3675 -174 3784
rect -65 3675 -59 3784
rect 3111 3712 3117 3823
rect 3226 3712 3232 3823
rect 6408 3717 6517 3723
rect 9693 3838 9814 3842
rect 9693 3727 9699 3838
rect 9808 3727 9814 3838
rect 12990 3831 13099 4396
rect 15453 4267 15603 4399
rect 16280 3851 16389 4401
rect 18742 4270 18892 4402
rect 18956 4231 18962 4406
rect 19137 4231 19143 4406
rect 19571 3851 19680 4399
rect 22032 4283 22182 4415
rect 22249 4394 22437 4400
rect 22249 4219 22257 4394
rect 22432 4219 22437 4394
rect 22249 4212 22437 4219
rect 16274 3845 16395 3851
rect 9693 3721 9814 3727
rect 12984 3827 13105 3831
rect 3111 3706 3232 3712
rect 12984 3716 12990 3827
rect 13099 3716 13105 3827
rect 16274 3736 16280 3845
rect 16389 3736 16395 3845
rect 16274 3730 16395 3736
rect 19565 3845 19686 3851
rect 19565 3736 19571 3845
rect 19680 3736 19686 3845
rect 22862 3835 22971 4396
rect 25320 4266 25470 4398
rect 25536 4213 25542 4385
rect 25714 4213 25720 4385
rect 25542 4068 25714 4074
rect 25536 3896 25542 4068
rect 25714 3896 25720 4068
rect 25542 3890 25714 3896
rect 19565 3730 19686 3736
rect 22856 3830 22977 3835
rect 12984 3710 13105 3716
rect 22856 3719 22862 3830
rect 22971 3719 22977 3830
rect 22856 3713 22977 3719
rect 25486 3220 26456 3311
rect 26365 1044 26456 3220
rect 29 959 97 1037
rect 3113 953 3316 1044
rect 6404 953 6607 1044
rect 9695 953 9898 1044
rect 12986 953 13189 1044
rect 16277 953 16480 1044
rect 19567 953 19770 1044
rect 22858 953 23061 1044
rect 26149 953 26456 1044
<< via1 >>
rect 2524 4202 2710 4388
rect 5810 4208 5991 4389
rect 9114 4214 9292 4392
rect 12391 4223 12566 4398
rect -174 3675 -65 3784
rect 3117 3712 3226 3823
rect 6408 3723 6517 3834
rect 9699 3727 9808 3838
rect 15673 4088 15848 4265
rect 18962 4231 19137 4406
rect 22257 4219 22432 4394
rect 12990 3716 13099 3827
rect 16280 3736 16389 3845
rect 19571 3736 19680 3845
rect 25542 4213 25714 4385
rect 25542 3896 25714 4068
rect 22862 3719 22971 3830
<< metal2 >>
rect 18962 4406 19137 4412
rect 12391 4398 12566 4404
rect 2524 4388 2710 4394
rect 9114 4392 9292 4398
rect 5804 4208 5810 4389
rect 5991 4208 5997 4389
rect 2524 4073 2710 4202
rect 5810 4073 5991 4208
rect 2524 4071 6007 4073
rect 9114 4071 9292 4214
rect 2524 4069 9302 4071
rect 12391 4069 12566 4223
rect 15667 4265 15859 4272
rect 15667 4088 15673 4265
rect 15848 4088 15859 4265
rect 2524 4068 12567 4069
rect 15667 4068 15859 4088
rect 18962 4068 19137 4231
rect 22249 4394 22437 4400
rect 22249 4219 22257 4394
rect 22432 4219 22437 4394
rect 22249 4212 22437 4219
rect 25542 4385 25714 4391
rect 22257 4068 22432 4212
rect 25542 4068 25714 4213
rect 2524 3896 25542 4068
rect 25714 3896 25720 4068
rect 2524 3893 22432 3896
rect 2524 3891 12567 3893
rect 2524 3890 9302 3891
rect 25542 3890 25714 3896
rect 2524 3887 6007 3890
rect 16274 3845 16395 3851
rect -174 3784 -65 3790
rect 6402 3723 6408 3834
rect 6517 3723 6523 3834
rect 16274 3736 16280 3845
rect 16389 3736 16395 3845
rect 16274 3730 16395 3736
rect 19565 3845 19686 3851
rect 19565 3736 19571 3845
rect 19680 3736 19686 3845
rect 19565 3730 19686 3736
rect -174 3669 -65 3675
rect 3122 22 3216 135
rect 6421 24 6515 137
rect 9710 25 9804 138
rect 12996 23 13090 136
rect 16292 28 16386 141
rect 19577 28 19671 141
rect 22871 26 22965 139
rect 26164 31 26258 144
<< metal4 >>
rect 630 4203 25315 4515
<< metal5 >>
rect -83 -380 26191 4514
use FULL_ADDER_XORED  FULL_ADDER_XORED_0
timestamp 1736620191
transform 1 0 118 0 1 1114
box -292 -1421 3108 3355
use FULL_ADDER_XORED  FULL_ADDER_XORED_1
timestamp 1736620191
transform 1 0 3409 0 1 1114
box -292 -1421 3108 3355
use FULL_ADDER_XORED  FULL_ADDER_XORED_2
timestamp 1736620191
transform 1 0 6700 0 1 1114
box -292 -1421 3108 3355
use FULL_ADDER_XORED  FULL_ADDER_XORED_3
timestamp 1736620191
transform 1 0 9991 0 1 1114
box -292 -1421 3108 3355
use FULL_ADDER_XORED  FULL_ADDER_XORED_4
timestamp 1736620191
transform 1 0 13282 0 1 1114
box -292 -1421 3108 3355
use FULL_ADDER_XORED  FULL_ADDER_XORED_5
timestamp 1736620191
transform 1 0 16572 0 1 1114
box -292 -1421 3108 3355
use FULL_ADDER_XORED  FULL_ADDER_XORED_6
timestamp 1736620191
transform 1 0 19863 0 1 1114
box -292 -1421 3108 3355
use FULL_ADDER_XORED  FULL_ADDER_XORED_7
timestamp 1736620191
transform 1 0 23154 0 1 1114
box -292 -1421 3108 3355
<< labels >>
rlabel metal4 9690 4249 9989 4459 5 VDD
port 28 s
rlabel metal5 13013 4410 13092 4510 5 VSS
port 27 s
rlabel metal1 35 965 87 1026 5 C
port 26 s
flabel metal2 3135 36 3210 118 0 FreeSans 160 0 0 0 S7
port 25 nsew
flabel metal2 6430 39 6505 121 0 FreeSans 160 0 0 0 S6
port 24 nsew
flabel metal2 9718 42 9793 124 0 FreeSans 160 0 0 0 S5
port 23 nsew
flabel metal2 13005 43 13080 125 0 FreeSans 160 0 0 0 S4
port 22 nsew
flabel metal2 16307 40 16382 122 0 FreeSans 160 0 0 0 S3
port 21 nsew
flabel metal2 19585 39 19660 121 0 FreeSans 160 0 0 0 S2
port 20 nsew
flabel metal2 22884 49 22959 131 0 FreeSans 160 0 0 0 S1
port 19 nsew
flabel metal2 26174 43 26249 125 0 FreeSans 160 0 0 0 S0
port 18 nsew
flabel metal1 -167 4310 -72 4376 0 FreeSans 160 0 0 0 A7
port 17 nsew
flabel metal1 3124 4304 3219 4370 0 FreeSans 160 0 0 0 A6
port 16 nsew
flabel metal1 6414 4312 6509 4378 0 FreeSans 160 0 0 0 A5
port 15 nsew
flabel metal1 9707 4314 9802 4380 0 FreeSans 160 0 0 0 A4
port 14 nsew
flabel metal1 12997 4312 13092 4378 0 FreeSans 160 0 0 0 A3
port 13 nsew
flabel metal1 16289 4306 16384 4372 0 FreeSans 160 0 0 0 A2
port 12 nsew
flabel metal1 19580 4310 19675 4376 0 FreeSans 160 0 0 0 A1
port 11 nsew
flabel metal1 22869 4316 22964 4382 0 FreeSans 160 0 0 0 A0
port 10 nsew
flabel metal1 2314 4293 2409 4359 0 FreeSans 160 0 0 0 B7
port 9 nsew
flabel metal1 5600 4287 5695 4353 0 FreeSans 160 0 0 0 B6
port 8 nsew
flabel metal1 8899 4291 8994 4357 0 FreeSans 160 0 0 0 B5
port 7 nsew
flabel metal1 12185 4284 12280 4350 0 FreeSans 160 0 0 0 B4
port 6 nsew
flabel metal1 15490 4289 15585 4355 0 FreeSans 160 0 0 0 B3
port 5 nsew
flabel metal1 18766 4302 18861 4368 0 FreeSans 160 0 0 0 B2
port 4 nsew
flabel metal1 22065 4308 22160 4374 0 FreeSans 160 0 0 0 B1
port 3 nsew
flabel metal1 25337 4298 25432 4364 0 FreeSans 160 0 0 0 B0
port 2 nsew
rlabel metal2 25542 4215 25714 4386 5 K
port 1 s
<< end >>
