magic
tech sky130B
magscale 1 2
timestamp 1735933295
<< nwell >>
rect -3709 381 -3708 813
rect -2408 380 -2407 812
rect -1202 411 -1201 843
rect -14 413 -13 845
rect 1114 428 1115 860
rect 2319 433 2320 865
rect 3503 434 3504 866
<< metal1 >>
rect -5260 250 -5171 927
rect -5090 279 -5018 927
rect -4380 313 -4172 395
rect -5260 114 -4997 250
rect -4615 -367 -4514 26
rect -4250 -133 -4172 313
rect -3950 250 -3861 927
rect -3780 279 -3708 927
rect -3008 305 -2867 387
rect -3950 114 -3708 250
rect -4615 -474 -4514 -468
rect -3299 -407 -3198 42
rect -2945 -141 -2867 305
rect -2649 249 -2560 926
rect -2479 278 -2407 926
rect -1701 307 -1565 389
rect -2649 113 -2407 249
rect -3299 -514 -3198 -508
rect -2005 -410 -1904 69
rect -1643 -139 -1565 307
rect -1443 280 -1354 957
rect -1273 309 -1201 957
rect -512 323 -365 405
rect -1443 144 -1201 280
rect -807 -401 -706 77
rect -443 -123 -365 323
rect -255 282 -166 959
rect -85 311 -13 959
rect 691 376 824 458
rect -255 146 -13 282
rect 365 -378 466 87
rect 746 -70 824 376
rect 873 297 962 974
rect 1036 427 1106 974
rect 1114 427 1115 461
rect 1036 326 1115 427
rect 1802 360 1926 442
rect 873 161 1115 297
rect 1506 -370 1607 96
rect 1848 -86 1926 360
rect 2078 302 2167 979
rect 2248 331 2320 979
rect 3022 368 3131 450
rect 2078 166 2320 302
rect 2718 -361 2819 108
rect 3053 -78 3131 368
rect 3262 303 3351 980
rect 3432 332 3504 980
rect 4204 376 4324 458
rect 3262 167 3504 303
rect 3914 -318 4015 103
rect 4246 -70 4324 376
rect 3914 -425 4015 -419
rect 2718 -468 2819 -462
rect 1506 -477 1607 -471
rect 365 -485 466 -479
rect -807 -508 -706 -502
rect -2005 -517 -1904 -511
<< via1 >>
rect -4615 -468 -4514 -367
rect -3299 -508 -3198 -407
rect -2005 -511 -1904 -410
rect -807 -502 -706 -401
rect 365 -479 466 -378
rect 1506 -471 1607 -370
rect 2718 -462 2819 -361
rect 3914 -419 4015 -318
<< metal2 >>
rect 3899 -318 4027 -306
rect -4630 -367 -4502 -355
rect -4630 -468 -4615 -367
rect -4514 -468 -4502 -367
rect 350 -378 478 -366
rect -4630 -478 -4502 -468
rect -3314 -407 -3186 -395
rect -3314 -508 -3299 -407
rect -3198 -508 -3186 -407
rect -3314 -518 -3186 -508
rect -2020 -410 -1892 -398
rect -2020 -511 -2005 -410
rect -1904 -511 -1892 -410
rect -2020 -521 -1892 -511
rect -822 -401 -694 -389
rect -822 -502 -807 -401
rect -706 -502 -694 -401
rect 350 -479 365 -378
rect 466 -479 478 -378
rect 350 -489 478 -479
rect 1491 -370 1619 -358
rect 1491 -471 1506 -370
rect 1607 -471 1619 -370
rect 1491 -481 1619 -471
rect 2703 -361 2831 -349
rect 2703 -462 2718 -361
rect 2819 -462 2831 -361
rect 3899 -419 3914 -318
rect 4015 -419 4027 -318
rect 3899 -429 4027 -419
rect 2703 -472 2831 -462
rect -822 -512 -694 -502
<< via2 >>
rect -4615 -468 -4514 -367
rect -3299 -508 -3198 -407
rect -2005 -511 -1904 -410
rect -807 -502 -706 -401
rect 365 -479 466 -378
rect 1506 -471 1607 -370
rect 2718 -462 2819 -361
rect 3914 -419 4015 -318
<< metal3 >>
rect 3883 -313 4039 -289
rect -4646 -362 -4490 -338
rect -4646 -473 -4620 -362
rect -4509 -473 -4490 -362
rect -4646 -501 -4490 -473
rect -3330 -402 -3174 -378
rect -3330 -513 -3304 -402
rect -3193 -513 -3174 -402
rect -3330 -541 -3174 -513
rect -2036 -405 -1880 -381
rect -2036 -516 -2010 -405
rect -1899 -516 -1880 -405
rect -2036 -544 -1880 -516
rect -838 -396 -682 -372
rect -838 -507 -812 -396
rect -701 -507 -682 -396
rect -838 -535 -682 -507
rect 334 -373 490 -349
rect 334 -484 360 -373
rect 471 -484 490 -373
rect 334 -512 490 -484
rect 1475 -365 1631 -341
rect 1475 -476 1501 -365
rect 1612 -476 1631 -365
rect 1475 -504 1631 -476
rect 2687 -356 2843 -332
rect 2687 -467 2713 -356
rect 2824 -467 2843 -356
rect 3883 -424 3909 -313
rect 4020 -424 4039 -313
rect 3883 -452 4039 -424
rect 2687 -495 2843 -467
<< via3 >>
rect -4620 -367 -4509 -362
rect -4620 -468 -4615 -367
rect -4615 -468 -4514 -367
rect -4514 -468 -4509 -367
rect -4620 -473 -4509 -468
rect -3304 -407 -3193 -402
rect -3304 -508 -3299 -407
rect -3299 -508 -3198 -407
rect -3198 -508 -3193 -407
rect -3304 -513 -3193 -508
rect -2010 -410 -1899 -405
rect -2010 -511 -2005 -410
rect -2005 -511 -1904 -410
rect -1904 -511 -1899 -410
rect -2010 -516 -1899 -511
rect -812 -401 -701 -396
rect -812 -502 -807 -401
rect -807 -502 -706 -401
rect -706 -502 -701 -401
rect -812 -507 -701 -502
rect 360 -378 471 -373
rect 360 -479 365 -378
rect 365 -479 466 -378
rect 466 -479 471 -378
rect 360 -484 471 -479
rect 1501 -370 1612 -365
rect 1501 -471 1506 -370
rect 1506 -471 1607 -370
rect 1607 -471 1612 -370
rect 1501 -476 1612 -471
rect 2713 -361 2824 -356
rect 2713 -462 2718 -361
rect 2718 -462 2819 -361
rect 2819 -462 2824 -361
rect 2713 -467 2824 -462
rect 3909 -318 4020 -313
rect 3909 -419 3914 -318
rect 3914 -419 4015 -318
rect 4015 -419 4020 -318
rect 3909 -424 4020 -419
<< via4 >>
rect -4724 -362 -4404 -257
rect -4724 -473 -4620 -362
rect -4620 -473 -4509 -362
rect -4509 -473 -4404 -362
rect -4724 -577 -4404 -473
rect -3408 -402 -3088 -297
rect -3408 -513 -3304 -402
rect -3304 -513 -3193 -402
rect -3193 -513 -3088 -402
rect -3408 -617 -3088 -513
rect -2114 -405 -1794 -300
rect -2114 -516 -2010 -405
rect -2010 -516 -1899 -405
rect -1899 -516 -1794 -405
rect -2114 -620 -1794 -516
rect -916 -396 -596 -291
rect -916 -507 -812 -396
rect -812 -507 -701 -396
rect -701 -507 -596 -396
rect -916 -611 -596 -507
rect 256 -373 576 -268
rect 256 -484 360 -373
rect 360 -484 471 -373
rect 471 -484 576 -373
rect 256 -588 576 -484
rect 1397 -365 1717 -260
rect 1397 -476 1501 -365
rect 1501 -476 1612 -365
rect 1612 -476 1717 -365
rect 1397 -580 1717 -476
rect 2609 -356 2929 -251
rect 2609 -467 2713 -356
rect 2713 -467 2824 -356
rect 2824 -467 2929 -356
rect 2609 -571 2929 -467
rect 3805 -313 4125 -208
rect 3805 -424 3909 -313
rect 3909 -424 4020 -313
rect 4020 -424 4125 -313
rect 3805 -528 4125 -424
<< metal5 >>
rect -4789 -257 -4344 -192
rect -4789 -577 -4724 -257
rect -4404 -577 -4344 -257
rect -4789 -640 -4344 -577
rect -3473 -297 -3028 -232
rect -3473 -617 -3408 -297
rect -3088 -617 -3028 -297
rect -3473 -680 -3028 -617
rect -2179 -300 -1734 -235
rect -2179 -620 -2114 -300
rect -1794 -620 -1734 -300
rect -2179 -683 -1734 -620
rect -981 -291 -536 -226
rect -981 -611 -916 -291
rect -596 -611 -536 -291
rect -981 -674 -536 -611
rect 191 -268 636 -203
rect 191 -588 256 -268
rect 576 -588 636 -268
rect 191 -651 636 -588
rect 1332 -260 1777 -195
rect 1332 -580 1397 -260
rect 1717 -580 1777 -260
rect 1332 -643 1777 -580
rect 2544 -251 2989 -186
rect 2544 -571 2609 -251
rect 2929 -571 2989 -251
rect 2544 -634 2989 -571
rect 3740 -208 4185 -143
rect 3740 -528 3805 -208
rect 4125 -528 4185 -208
rect 3740 -591 4185 -528
use NAND2  NAND2_0 ~/Desktop/vlsi_sky130b/design/mag/NAND/NAND2
timestamp 1735933295
transform 1 0 3148 0 1 62
box 356 -17 1062 804
use NAND2  NAND2_1
timestamp 1735933295
transform 1 0 -369 0 1 41
box 356 -17 1062 804
use NAND2  NAND2_2
timestamp 1735933295
transform 1 0 -1563 0 1 39
box 356 -17 1062 804
use NAND2  NAND2_4
timestamp 1735933295
transform 1 0 -5375 0 1 9
box 356 -17 1062 804
use NAND2  NAND2_6
timestamp 1735933295
transform 1 0 750 0 1 56
box 356 -17 1062 804
use NAND2  NAND2_7
timestamp 1735933295
transform 1 0 1963 0 1 61
box 356 -17 1062 804
use NAND2  NAND2_8
timestamp 1735933295
transform 1 0 -4066 0 1 9
box 356 -17 1062 804
use NAND2  NAND2_9
timestamp 1735933295
transform 1 0 -2763 0 1 8
box 356 -17 1062 804
<< labels >>
rlabel metal1 -3709 350 -3709 350 7 A
port 1 w
rlabel metal1 -3709 182 -3709 182 7 B
port 2 w
rlabel metal1 -2408 181 -2408 181 7 B
port 2 w
rlabel metal1 -2408 349 -2408 349 7 A
port 1 w
rlabel metal1 -1202 380 -1202 380 7 A
port 1 w
rlabel metal1 -1202 212 -1202 212 7 B
port 2 w
rlabel metal1 -14 214 -14 214 7 B
port 2 w
rlabel metal1 -14 382 -14 382 7 A
port 1 w
rlabel metal1 1114 229 1114 229 7 B
port 2 w
rlabel metal1 1114 397 1114 397 7 A
port 1 w
rlabel metal1 2319 402 2319 402 7 A
port 1 w
rlabel metal1 2319 234 2319 234 7 B
port 2 w
rlabel metal1 3503 403 3503 403 7 A
port 1 w
rlabel metal1 3503 235 3503 235 7 B
port 2 w
<< end >>
