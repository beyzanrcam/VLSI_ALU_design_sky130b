* NGSPICE file created from nor8.ext - technology: sky130B

.subckt sky130_fd_pr__pfet_01v8_64A2S3 a_n33_n428# a_447_n428# a_n605_n428# a_321_n484#
+ a_n543_n484# a_543_n428# a_159_n428# a_33_n484# a_n255_n484# a_255_n428# w_n641_n484#
+ a_351_n428# a_n417_n428# a_n513_n428# a_n129_n428# a_63_n428# a_n225_n428# a_n321_n428#
X0 a_447_n428# a_321_n484# a_351_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X1 a_n513_n428# a_n543_n484# a_n605_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=1.3268 ps=9.18 w=4.28 l=0.15
X2 a_63_n428# a_33_n484# a_n33_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X3 a_n129_n428# a_n255_n484# a_n225_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X4 a_n417_n428# a_n543_n484# a_n513_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X5 a_n33_n428# a_n255_n484# a_n129_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X6 a_351_n428# a_321_n484# a_255_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X7 a_255_n428# a_33_n484# a_159_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X8 a_n321_n428# a_n543_n484# a_n417_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X9 a_543_n428# a_321_n484# a_447_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=1.3268 pd=9.18 as=0.7062 ps=4.61 w=4.28 l=0.15
X10 a_159_n428# a_33_n484# a_63_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X11 a_n225_n428# a_n255_n484# a_n321_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_S9NJ5Q a_159_n100# a_n159_n126# a_33_n126# a_n129_n100#
+ a_n221_n100# a_63_n100# a_n63_n126# a_n33_n100# a_129_n126# VSUBS
X0 a_n129_n100# a_n159_n126# a_n221_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1 a_63_n100# a_33_n126# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2 a_n33_n100# a_n63_n126# a_n129_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_159_n100# a_129_n126# a_63_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt nor4 A B C D VSS Y VDD
Xsky130_fd_pr__pfet_01v8_64A2S3_0 m1_n20_1047# m1_268_1523# VDD D A Y m1_n20_1047#
+ C B m1_268_1523# VDD Y VDD m1_n308_1523# m1_n308_1523# m1_268_1523# m1_n20_1047#
+ m1_n308_1523# sky130_fd_pr__pfet_01v8_64A2S3
Xsky130_fd_pr__nfet_01v8_S9NJ5Q_0 VSS A C Y VSS Y B VSS D VSS sky130_fd_pr__nfet_01v8_S9NJ5Q
.ends

.subckt sky130_fd_pr__pfet_01v8_UFBY79 a_n33_n128# a_n509_n128# a_447_n128# a_159_n128#
+ a_255_n128# a_351_n128# a_n417_n128# a_n447_n225# a_n129_n128# a_63_n128# a_n225_n128#
+ a_33_n225# w_n545_n228# a_n321_n128#
X0 a_63_n128# a_33_n225# a_n33_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1 a_n129_n128# a_n447_n225# a_n225_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2 a_n417_n128# a_n447_n225# a_n509_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X3 a_351_n128# a_33_n225# a_255_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X4 a_n33_n128# a_n447_n225# a_n129_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X5 a_255_n128# a_33_n225# a_159_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X6 a_n321_n128# a_n447_n225# a_n417_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X7 a_159_n128# a_33_n225# a_63_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X8 a_n225_n128# a_n447_n225# a_n321_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X9 a_447_n128# a_33_n225# a_351_n128# w_n545_n228# sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_LZEQWH a_33_n126# a_n125_n100# a_63_n100# a_n63_n126#
+ a_n33_n100# VSUBS
X0 a_63_n100# a_33_n126# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X1 a_n33_n100# a_n63_n126# a_n125_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
.ends

.subckt nor2 A B VSS VDD Y
Xsky130_fd_pr__pfet_01v8_UFBY79_0 m1_760_245# VDD Y m1_760_245# Y m1_760_245# m1_760_245#
+ A VDD Y m1_760_245# B VDD VDD sky130_fd_pr__pfet_01v8_UFBY79
Xsky130_fd_pr__nfet_01v8_LZEQWH_0 A VSS VSS B Y VSS sky130_fd_pr__nfet_01v8_LZEQWH
.ends

.subckt nor8 A0 A1 A2 A3 A4 A5 A6 A7 Y
Xnor4_0 A4 A5 A6 A7 VSS nor4_0/Y VDD nor4
Xnor4_1 A0 A1 A2 A3 VSS nor4_1/Y VDD nor4
Xnor2_0 nor4_1/Y nor4_0/Y VSS VDD Y nor2
.ends

