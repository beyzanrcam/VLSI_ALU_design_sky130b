* NGSPICE file created from alu_pex.ext - technology: sky130B

.subckt alu_pex B0 B1 B2 B3 B4 B5 B6 A0 A1 A2 A3 A4 A5 A6 A7 Y0 Y1 Y2 Y3 Y4 Y5 Y6
+ S Z C V VSS Y7 B7 SEL0 SEL1 SEL2 SEL3 VDD
X0 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t8 a_n13531_3164.t2 a_n13501_3190.t5 VSS.t1345 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VSS.t2026 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t12 a_n10081_1406.t0 VSS.t2025 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2 mux8_2.NAND4F_0.Y.t4 SEL0.t0 VDD.t3102 VDD.t3101 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3 a_n12416_n11683.t2 a_n12446_n11709.t2 VSS.t1939 VSS.t1938 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 VDD.t4298 mux8_5.NAND4F_8.Y.t9 a_11865_n20887.t9 VDD.t4297 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X5 a_11865_n2775.t9 mux8_1.NAND4F_8.Y.t9 VDD.t4315 VDD.t4314 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X6 a_n18305_n6187.t1 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t7 VSS.t1948 VSS.t352 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X7 a_n20083_3190.t2 a_n20839_3190.t2 VSS.t1923 VSS.t1922 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X8 VDD.t4274 MULT_0.inv_13.A.t7 MULT_0.4bit_ADDER_1.A3.t3 VDD.t4273 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X9 mux8_2.NAND4F_5.Y.t4 SEL1.t0 VDD.t4336 VDD.t4335 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X10 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t3 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t7 VDD.t4280 VDD.t4279 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X11 mux8_7.NAND4F_8.Y.t8 mux8_7.NAND4F_2.Y.t9 VDD.t4262 VDD.t4261 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X12 VDD.t3100 SEL0.t1 mux8_5.NAND4F_6.Y.t6 VDD.t3099 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X13 VSS.t1886 a_n4385_3190.t2 a_n3629_3190.t2 VSS.t1885 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X14 VDD.t3939 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t7 a_n13192_2026.t9 VDD.t3938 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X15 VDD.t4187 A1.t0 MULT_0.NAND2_9.Y.t3 VDD.t4186 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X16 mux8_3.inv_0.A.t0 mux8_3.NAND4F_8.Y.t9 VSS.t1779 VSS.t1778 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X17 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t4 a_n18222_1406.t2 a_n18042_2026.t5 VDD.t3897 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X18 a_n24624_1406.t3 a_n24654_1380.t2 VSS.t1755 VSS.t1754 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X19 a_n13975_n7799.t5 a_n14155_n8419.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t5 VDD.t3689 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X20 a_n11276_n15299.t5 a_n12347_n15041.t2 XOR8_0.S0.t11 VSS.t1689 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X21 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t7 a_n11723_n9452.t0 VSS.t1687 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X22 VDD.t3654 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t12 a_n18998_n11063.t7 VDD.t3653 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X23 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t6 a_n24130_3190.t2 a_n23950_3810.t5 VDD.t3697 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X24 VDD.t4025 MULT_0.4bit_ADDER_1.B2.t12 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t6 VDD.t4024 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X25 mux8_4.NAND4F_5.Y.t1 SEL2.t0 VDD.t3701 VDD.t3700 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X26 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t3 MULT_0.inv_9.Y.t4 VDD.t4007 VDD.t4006 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X27 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t3 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t8 a_n13381_373.t1 VSS.t163 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X28 a_n13975_n8419.t5 a_n14005_n8445.t2 VSS.t1659 VSS.t1658 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X29 mux8_5.NAND4F_3.Y.t1 mux8_5.NAND4F_0.C.t4 VDD.t3624 VDD.t3623 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X30 mux8_4.NAND4F_7.Y.t4 NOT8_0.S3.t4 VDD.t3572 VDD.t3571 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X31 VDD.t3580 B4.t0 a_n12345_n26161.t1 VDD.t3579 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X32 a_n10684_n11063.t6 MULT_0.inv_8.Y.t4 VDD.t3513 VDD.t3512 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X33 VSS.t1625 B6.t0 a_n23960_n22530.t0 VSS.t686 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X34 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t11 a_n14155_n5154.t2 a_n13975_n5154.t5 VSS.t1873 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X35 VDD.t4043 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t3 VDD.t4042 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X36 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t2 a_n4385_3190.t3 a_n4205_3810.t2 VDD.t4185 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X37 XOR8_0.S4.t5 B4.t1 a_n11274_n25843.t2 VSS.t1642 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X38 a_5197_5532.t6 a_5167_4886.t2 V_FLAG_0.XOR2_0.Y.t9 VDD.t55 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X39 mux8_7.NAND4F_7.Y.t4 NOT8_0.S5.t4 a_10459_n26405.t0 VSS.t19 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X40 a_n11274_n23651.t2 a_n12345_n23393.t2 XOR8_0.S3.t4 VSS.t1593 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X41 VDD.t4332 mux8_2.NAND4F_0.Y.t9 mux8_2.NAND4F_8.Y.t5 VDD.t4331 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X42 a_n16690_n8419.t5 MULT_0.4bit_ADDER_1.A2.t4 VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X43 VDD.t4051 MULT_0.4bit_ADDER_2.B3.t7 a_n20737_n11683.t1 VDD.t4050 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X44 VSS.t1032 VSS.t1030 a_n8549_n11683.t2 VSS.t1031 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X45 XOR8_0.S6.t2 B6.t1 a_n11274_n31085.t0 VSS.t1626 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X46 a_n23960_n23839.t0 A7.t0 AND8_0.NOT8_0.A7.t3 VSS.t1158 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X47 mux8_1.NAND4F_6.Y.t6 SEL1.t1 VDD.t4338 VDD.t4337 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X48 VSS.t110 MULT_0.4bit_ADDER_0.A2.t4 a_n16690_n5154.t2 VSS.t109 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X49 VDD.t258 A2.t0 AND8_0.NOT8_0.A2.t5 VDD.t257 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X50 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t2 a_n24804_1406.t2 a_n24624_2026.t2 VDD.t57 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X51 a_11865_1753.t4 mux8_0.NAND4F_8.Y.t9 VDD.t3503 VDD.t3502 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X52 VDD.t3497 V_FLAG_0.NAND2_0.Y.t7 V.t3 VDD.t3496 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X53 VSS.t26 a_n15737_n8445.t2 a_n15707_n8419.t5 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X54 mux8_2.NAND4F_1.Y.t3 XOR8_0.S1.t12 VDD.t63 VDD.t62 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X55 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t5 MULT_0.4bit_ADDER_1.B2.t13 VDD.t4027 VDD.t4026 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X56 VDD.t641 mux8_0.NAND4F_0.C.t4 mux8_0.NAND4F_3.Y.t3 VDD.t640 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X57 a_n18072_1380.t0 A5.t0 VSS.t176 VSS.t175 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X58 mux8_7.NAND4F_5.Y.t7 mux8_7.NAND4F_4.B.t4 VDD.t2049 VDD.t2048 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X59 AND8_0.NOT8_0.A1.t3 A1.t1 VDD.t4189 VDD.t4188 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X60 VDD.t881 OR8_0.S0.t4 mux8_1.NAND4F_2.Y.t2 VDD.t880 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X61 a_n15707_n5154.t5 a_n15737_n5180.t2 VSS.t1831 VSS.t1830 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X62 VDD.t4300 mux8_5.NAND4F_8.Y.t10 a_11865_n20887.t8 VDD.t4299 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X63 VDD.t3581 B4.t2 right_shifter_0.buffer_4.inv_1.A.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X64 AND8_0.NOT8_0.A3.t5 A3.t0 VDD.t4067 VDD.t4066 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X65 VDD.t3114 VDD.t3113 left_shifter_0.S0.t3 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X66 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t3 a_n5059_1406.t2 a_n4879_2026.t2 VDD.t797 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X67 mux8_5.NAND4F_5.Y.t1 SEL2.t1 VDD.t3703 VDD.t3702 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X68 VDD.t763 SEL3.t0 a_n7676_3190.t1 VDD.t762 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X69 VSS.t1029 VSS.t1027 a_n8549_n5154.t2 VSS.t1028 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X70 a_8592_n25478.t1 SEL0.t2 a_8496_n25478.t1 VSS.t1989 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X71 mux8_5.NAND4F_7.Y.t6 NOT8_0.S4.t4 VDD.t3955 VDD.t3954 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X72 mux8_4.NAND4F_9.Y.t4 mux8_4.NAND4F_6.Y.t9 VDD.t229 VDD.t228 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X73 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t3 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t7 a_n19187_n12716.t1 VSS.t465 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X74 VSS.t1866 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t7 a_n18422_n8419.t5 VSS.t1865 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X75 VDD.t2317 B1.t0 a_n12314_n18115.t2 VDD.t2316 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X76 mux8_1.NAND4F_1.Y.t8 mux8_1.NAND4F_4.B.t4 VDD.t1260 VDD.t1259 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X77 mux8_1.NAND4F_9.Y.t8 mux8_1.NAND4F_7.Y.t9 VDD.t1324 VDD.t1323 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X78 a_n18422_n5154.t4 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t7 VSS.t1276 VSS.t1275 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X79 VDD.t3098 SEL0.t3 mux8_8.NAND4F_6.Y.t8 VDD.t3097 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X80 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t5 a_n14931_1406.t2 a_n14751_1406.t5 VSS.t1548 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X81 VDD.t3096 SEL0.t4 mux8_1.NAND4F_7.Y.t8 VDD.t3095 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X82 VDD.t3094 SEL0.t5 mux8_4.NAND4F_4.B.t3 VDD.t3026 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X83 a_n14077_3810.t5 B4.t3 VDD.t3583 VDD.t3582 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X84 V_FLAG_0.NAND2_0.Y.t0 V_FLAG_0.XOR2_2.Y.t12 VDD.t2272 VDD.t2271 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X85 VDD.t3384 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t12 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t2 VDD.t3383 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X86 VSS.t1147 a_n3350_1380.t2 a_n3320_1406.t2 VSS.t1146 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X87 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t5 a_n1768_1406.t2 a_n1588_1406.t2 VSS.t1274 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X88 OR8_0.S5.t3 OR8_0.NOT8_0.A5.t7 VDD.t2277 VDD.t311 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X89 VDD.t584 B0.t0 MULT_0.NAND2_2.Y.t2 VDD.t583 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X90 a_n11274_n29052.t4 a_n12345_n28506.t2 VSS.t934 VSS.t933 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X91 a_9432_n20950.t0 mux8_5.NAND4F_0.C.t5 a_9336_n20950.t0 VSS.t1664 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X92 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t12 VDD.t2251 VDD.t2250 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X93 VDD.t151 MULT_0.4bit_ADDER_2.B2.t12 a_n17446_n11683.t1 VDD.t150 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X94 mux8_3.NAND4F_8.Y.t4 mux8_3.NAND4F_4.Y.t9 VDD.t2643 VDD.t2642 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X95 VSS.t645 left_shifter_0.buffer_2.inv_1.A.t4 left_shifter_0.S7.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X96 a_11865_n7203.t4 mux8_2.NAND4F_8.Y.t9 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X97 V_FLAG_0.XOR2_2.Y.t3 a_3463_4888.t2 a_3493_5534.t11 VDD.t487 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X98 mux8_6.NAND4F_7.Y.t4 NOT8_0.S7.t4 a_10459_n35461.t0 VSS.t199 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X99 VDD.t1983 VSS.t2033 a_n9125_n4534.t9 VDD.t1982 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X100 mux8_5.NAND4F_9.Y.t6 mux8_5.NAND4F_6.Y.t9 VDD.t4246 VDD.t4245 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X101 a_10459_n30006.t1 SEL0.t6 a_10363_n30006.t1 VSS.t1988 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X102 a_n14077_3190.t2 SEL3.t1 VSS.t372 VSS.t371 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X103 a_n12605_n12716.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t12 VSS.t1041 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X104 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t0 MULT_0.inv_9.Y.t5 a_n13714_n12716.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X105 C.t0 mux8_0.inv_0.A.t7 VSS.t1515 VSS.t1514 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X106 VDD.t222 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t3 VDD.t221 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X107 MULT_0.NAND2_14.Y.t2 A2.t1 VDD.t260 VDD.t259 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X108 VDD.t2319 B1.t1 a_n12345_n17857.t1 VDD.t2318 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X109 a_n4205_3190.t2 SEL3.t2 VSS.t374 VSS.t373 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X110 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t0 MULT_0.4bit_ADDER_0.B0.t4 VDD.t284 VDD.t283 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X111 mux8_6.NAND4F_5.Y.t8 mux8_6.NAND4F_4.B.t4 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X112 a_n11274_n18115.t5 a_n12345_n17857.t2 XOR8_0.S1.t0 VSS.t128 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X113 a_9336_n12822.t0 SEL2.t2 VSS.t1700 VSS.t1382 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X114 a_n914_3810.t2 SEL3.t3 VDD.t765 VDD.t764 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X115 VSS.t1218 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t7 a_n11840_n5154.t2 VSS.t1217 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X116 VDD.t4069 A3.t1 MULT_0.NAND2_11.Y.t6 VDD.t4068 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X117 mux8_8.NAND4F_5.Y.t1 SEL2.t3 VDD.t3705 VDD.t3704 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X118 VSS.t213 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t12 a_n15887_n5154.t0 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X119 a_n22426_n9284.t0 B2.t0 VSS.t1285 VSS.t1284 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X120 mux8_8.NAND4F_7.Y.t7 NOT8_0.S6.t4 VDD.t2281 VDD.t2280 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X121 VDD.t3527 B6.t2 right_shifter_0.buffer_2.inv_1.A.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X122 mux8_7.NAND4F_9.Y.t4 mux8_7.NAND4F_5.Y.t9 a_11386_n26406.t1 VSS.t243 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X123 VDD.t3495 MULT_0.4bit_ADDER_1.B1.t12 a_n14155_n8419.t1 VDD.t3494 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X124 a_n12314_n26419.t5 B4.t4 VDD.t3585 VDD.t3584 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X125 VDD.t802 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t7 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t6 VDD.t801 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X126 mux8_2.NAND4F_1.Y.t4 XOR8_0.S1.t13 a_9528_n8194.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X127 AND8_0.S0.t3 AND8_0.NOT8_0.A0.t7 VDD.t1353 VDD.t1352 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X128 8bit_ADDER_0.S0.t2 a_n209_1406.t2 a_n29_1406.t2 VSS.t1451 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X129 VDD.t3528 B6.t3 left_shifter_0.buffer_2.inv_1.A.t3 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X130 left_shifter_0.S1.t3 left_shifter_0.buffer_6.inv_1.A.t4 VDD.t1238 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X131 VDD.t1245 mux8_0.NAND4F_0.Y.t9 mux8_0.NAND4F_8.Y.t2 VDD.t1244 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X132 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t2 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t12 VDD.t749 VDD.t748 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X133 MULT_0.4bit_ADDER_0.A1.t3 MULT_0.NAND2_5.Y.t7 VDD.t3148 VDD.t3147 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X134 mux8_5.NAND4F_0.Y.t3 mux8_5.A1.t12 VDD.t1365 VDD.t1364 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X135 a_n14490_373.t0 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t12 VSS.t708 VSS.t707 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X136 VDD.t3412 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t6 VDD.t3411 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X137 a_n18042_1406.t2 a_n18072_1380.t2 VSS.t1065 VSS.t1064 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X138 VDD.t1249 left_shifter_0.S1.t4 mux8_2.NAND4F_5.Y.t0 VDD.t1248 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X139 VDD.t4340 SEL1.t2 mux8_0.NAND4F_2.Y.t4 VDD.t4339 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X140 a_n9325_1406.t2 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t7 VSS.t859 VSS.t858 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X141 a_16431_n18523.t5 Y1.t4 a_16143_n18523.t2 VDD.t3167 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X142 mux8_8.inv_0.A.t4 mux8_8.NAND4F_9.Y.t9 a_11865_n29943.t4 VDD.t1110 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X143 a_n17677_n21025.t4 B4.t5 VDD.t3587 VDD.t3586 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X144 VDD.t3468 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t12 a_n23245_1406.t1 VDD.t3467 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X145 mux8_2.NAND4F_5.Y.t1 left_shifter_0.S1.t5 a_7644_n8194.t0 VSS.t396 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X146 VSS.t178 A5.t1 OR8_0.NOT8_0.A5.t6 VSS.t177 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X147 a_n18998_n11063.t11 a_n19028_n11709.t2 mux8_8.A1.t9 VDD.t2728 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X148 VDD.t2713 MULT_0.4bit_ADDER_1.B3.t7 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t2 VDD.t2712 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X149 a_11865_n25415.t4 mux8_7.NAND4F_9.Y.t9 mux8_7.inv_0.A.t5 VDD.t3281 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X150 a_n15907_1406.t2 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t12 mux8_7.A0.t10 VSS.t1770 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X151 a_11290_n25478.t0 mux8_7.NAND4F_3.Y.t9 a_11194_n25478.t1 VSS.t1272 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X152 a_n20113_3164.t1 B6.t4 VDD.t3530 VDD.t3529 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X153 VDD.t3187 MULT_0.4bit_ADDER_1.A0.t4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t6 VDD.t3186 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X154 VDD.t2633 MULT_0.NAND2_14.Y.t7 MULT_0.inv_14.Y.t3 VDD.t2632 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X155 VDD.t2418 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t8 a_n12416_n4534.t3 VDD.t2417 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X156 VDD.t3352 mux8_3.NAND4F_7.Y.t9 mux8_3.NAND4F_9.Y.t6 VDD.t3351 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X157 VSS.t1519 mux8_6.A0.t12 a_5773_4912.t5 VSS.t1518 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X158 a_n6035_1406.t5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t12 8bit_ADDER_0.S2.t6 VSS.t1237 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X159 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t2 a_n17296_n8445.t2 a_n17266_n7799.t2 VDD.t3288 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X160 a_n6950_3164.t1 B2.t1 VDD.t2574 VDD.t2573 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X161 VDD.t713 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t6 VDD.t712 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X162 mux8_8.NAND4F_9.Y.t4 mux8_8.NAND4F_6.Y.t9 VDD.t354 VDD.t353 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X163 mux8_6.NAND4F_8.Y.t4 mux8_6.NAND4F_4.Y.t9 VDD.t911 VDD.t910 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X164 a_3463_4888.t0 V_FLAG_0.XOR2_2.B.t12 VSS.t489 VSS.t488 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X165 mux8_0.NAND4F_2.D.t0 SEL2.t4 VSS.t1702 VSS.t1701 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X166 mux8_2.NAND4F_8.Y.t1 mux8_2.NAND4F_4.Y.t9 VDD.t915 VDD.t914 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X167 a_n17677_n18225.t9 B2.t2 VDD.t2576 VDD.t2575 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X168 OR8_0.NOT8_0.A0.t4 A0.t0 a_n17677_n15425.t4 VDD.t1653 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X169 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t3 a_n17446_n8419.t2 a_n17266_n8419.t5 VSS.t356 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X170 VSS.t1834 A3.t2 OR8_0.NOT8_0.A3.t6 VSS.t810 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X171 VDD.t1061 right_shifter_0.S0.t4 mux8_1.NAND4F_6.Y.t2 VDD.t1060 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X172 mux8_6.NAND4F_4.B.t0 SEL0.t7 VSS.t1987 VSS.t1986 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X173 ZFLAG_0.nor4_0.Y.t4 Y3.t4 VSS.t1220 VSS.t1219 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X174 VDD.t888 B5.t0 NOT8_0.S5.t0 VDD.t887 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X175 a_7644_n16422.t0 mux8_4.NAND4F_4.B.t4 a_7548_n16422.t0 VSS.t1544 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X176 a_n10786_3190.t5 B3.t0 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t9 VSS.t1100 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X177 VDD.t180 mux8_7.NAND4F_0.C.t4 mux8_7.NAND4F_1.Y.t3 VDD.t179 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X178 a_n16690_n5154.t3 MULT_0.4bit_ADDER_0.B2.t4 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t9 VSS.t1445 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X179 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t2 a_n16822_3164.t2 a_n16792_3190.t2 VSS.t1434 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X180 a_n18998_n11063.t6 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t13 VDD.t3656 VDD.t3655 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X181 VSS.t137 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t12 a_n13372_1406.t0 VSS.t136 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X182 a_7548_n20950.t1 SEL1.t3 a_7452_n20950.t1 VSS.t1950 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X183 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t2 MULT_0.4bit_ADDER_2.B3.t8 VDD.t4053 VDD.t4052 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X184 mux8_0.NAND4F_4.Y.t3 mux8_0.NAND4F_2.D.t4 VDD.t2888 VDD.t2887 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X185 a_n14751_2026.t8 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t13 VDD.t1438 VDD.t1437 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X186 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t5 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t8 VDD.t804 VDD.t803 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X187 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t3 MULT_0.4bit_ADDER_0.A1.t4 VDD.t2303 VDD.t2302 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X188 VDD.t1349 mux8_2.NAND4F_7.Y.t9 mux8_2.NAND4F_9.Y.t1 VDD.t1348 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X189 a_n11274_n23651.t3 a_n12345_n23105.t2 VSS.t1360 VSS.t1359 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X190 VSS.t1791 a_n7676_3190.t2 a_n6920_3190.t2 VSS.t1790 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X191 VDD.t2749 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t7 a_n16483_2026.t5 VDD.t2748 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X192 a_n22489_1406.t4 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t13 mux8_6.A0.t1 VSS.t1600 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X193 VSS.t1053 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t7 a_n11840_n11683.t5 VSS.t1052 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X194 XOR8_0.S6.t3 a_n12345_n31403.t2 a_n11274_n31661.t2 VSS.t940 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X195 a_n20659_3810.t2 SEL3.t4 VDD.t767 VDD.t766 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X196 VDD.t2837 A6.t0 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t3 VDD.t2836 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X197 VDD.t751 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t13 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t1 VDD.t750 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X198 a_n18998_n7799.t8 a_n19028_n8445.t2 MULT_0.4bit_ADDER_2.B2.t9 VDD.t1344 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X199 mux8_6.NAND4F_9.Y.t2 mux8_6.NAND4F_5.Y.t9 a_11386_n35462.t1 VSS.t234 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X200 VDD.t2140 B3.t1 NOT8_0.S3.t2 VDD.t887 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X201 a_n8200_1380.t1 A2.t2 VDD.t262 VDD.t261 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X202 VDD.t831 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t7 a_n15707_n11063.t5 VDD.t830 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X203 a_n9125_n5154.t5 a_n9305_n5154.t2 MULT_0.S1.t6 VSS.t170 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X204 VDD.t635 MULT_0.4bit_ADDER_0.A3.t4 a_n20557_n4534.t2 VDD.t634 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X205 a_n18998_n8419.t2 a_n19178_n8419.t2 MULT_0.4bit_ADDER_2.B2.t0 VSS.t124 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X206 VDD.t4244 MULT_0.4bit_ADDER_1.A3.t4 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t6 VDD.t4243 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X207 a_11865_n7203.t5 mux8_2.NAND4F_9.Y.t9 mux8_2.inv_0.A.t5 VDD.t2113 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X208 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t1 a_n10864_n11683.t2 a_n10684_n11063.t1 VDD.t1536 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X209 VSS.t1809 MULT_0.inv_9.Y.t6 a_n13399_n11683.t2 VSS.t1808 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X210 AND8_0.NOT8_0.A1.t4 B1.t2 VDD.t2321 VDD.t2320 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X211 MULT_0.4bit_ADDER_1.B2.t2 a_n19178_n5154.t2 a_n18998_n5154.t2 VSS.t337 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X212 VSS.t330 AND8_0.NOT8_0.A4.t7 AND8_0.S4.t0 VSS.t329 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X213 a_n7909_373.t0 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t12 VSS.t430 VSS.t118 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X214 a_n19187_n9452.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t13 VSS.t1139 VSS.t1138 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X215 a_n16690_n11683.t2 MULT_0.4bit_ADDER_2.B2.t13 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t2 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X216 VDD.t4071 A3.t3 AND8_0.NOT8_0.A3.t4 VDD.t4070 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X217 VSS.t1695 a_n24130_3190.t3 a_n23374_3190.t3 VSS.t1694 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X218 VSS.t376 SEL3.t5 a_n20839_3190.t0 VSS.t375 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X219 MULT_0.NAND2_5.Y.t2 B1.t3 VDD.t2323 VDD.t2322 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X220 VDD.t2142 B3.t2 MULT_0.NAND2_15.Y.t6 VDD.t2141 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X221 AND8_0.NOT8_0.A5.t2 B5.t1 VDD.t890 VDD.t889 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X222 a_n11460_1406.t2 a_n11490_1380.t2 VSS.t475 VSS.t474 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X223 a_11865_n34471.t9 mux8_6.NAND4F_9.Y.t9 mux8_6.inv_0.A.t2 VDD.t694 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X224 right_shifter_0.buffer_4.inv_1.A.t2 B4.t6 VDD.t3588 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X225 a_n21333_2026.t3 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t12 VDD.t3233 VDD.t3232 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X226 mux8_5.A1.t6 a_n12596_n11683.t2 a_n12416_n11683.t3 VSS.t615 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X227 a_11865_n20887.t7 mux8_5.NAND4F_8.Y.t11 VDD.t4302 VDD.t4301 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X228 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t6 a_n1618_1380.t2 a_n1588_2026.t8 VDD.t1252 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X229 a_9336_n2838.t0 mux8_1.NAND4F_2.D.t4 VSS.t850 VSS.t849 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X230 a_n18998_n11063.t5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t14 VDD.t3658 VDD.t3657 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X231 mux8_4.NAND4F_4.B.t2 SEL0.t8 VDD.t3093 VDD.t3026 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X232 VDD.t4009 MULT_0.inv_9.Y.t7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t2 VDD.t4008 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X233 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t0 a_n8350_1406.t2 a_n8170_2026.t8 VDD.t227 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X234 VDD.t1329 MULT_0.NAND2_1.Y.t7 MULT_0.4bit_ADDER_0.B1.t3 VDD.t236 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X235 a_n10684_n4534.t2 a_n10714_n5180.t2 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t5 VDD.t305 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X236 a_n9125_n4534.t0 a_n9155_n5180.t2 MULT_0.S1.t0 VDD.t308 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X237 OR8_0.NOT8_0.A6.t4 A6.t1 a_n17677_n23825.t1 VDD.t2838 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X238 VDD.t324 mux8_6.NAND4F_0.C.t4 mux8_6.NAND4F_1.Y.t3 VDD.t323 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X239 VDD.t3092 SEL0.t9 mux8_4.NAND4F_7.Y.t6 VDD.t3091 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X240 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t2 MULT_0.4bit_ADDER_2.B2.t14 VDD.t153 VDD.t152 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X241 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t4 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t7 VDD.t2247 VDD.t2246 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X242 VDD.t3515 MULT_0.inv_8.Y.t5 a_n10684_n11063.t5 VDD.t3514 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X243 VDD.t922 mux8_3.NAND4F_5.Y.t9 mux8_3.NAND4F_9.Y.t0 VDD.t921 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X244 VDD.t3707 SEL2.t5 mux8_3.NAND4F_7.Y.t1 VDD.t3706 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X245 mux8_4.A0.t6 a_n10081_1406.t2 a_n9901_1406.t2 VSS.t2022 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X246 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t0 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t14 VDD.t753 VDD.t752 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X247 VSS.t416 AND8_0.NOT8_0.A1.t7 AND8_0.S1.t0 VSS.t415 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X248 mux8_7.NAND4F_6.Y.t2 right_shifter_0.S5.t4 a_8592_n26406.t0 VSS.t1050 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X249 VSS.t830 A0.t1 a_n1012_1406.t2 VSS.t829 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X250 VDD.t2840 A6.t2 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t2 VDD.t2839 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X251 a_n8549_n11683.t1 VSS.t1024 VSS.t1026 VSS.t1025 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X252 a_10459_n26405.t1 SEL0.t10 a_10363_n26405.t1 VSS.t1994 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X253 VDD.t2253 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t12 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t6 VDD.t2252 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X254 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t0 a_n10240_3164.t2 a_n10786_3810.t5 VDD.t683 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X255 a_n20587_n5180.t0 MULT_0.4bit_ADDER_0.A3.t5 VSS.t313 VSS.t312 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X256 VSS.t1259 right_shifter_0.buffer_5.inv_1.A.t4 right_shifter_0.S2.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X257 a_n17368_3810.t8 B5.t2 VDD.t892 VDD.t891 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X258 a_n12345_n28506.t1 A5.t2 VDD.t377 VDD.t376 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X259 VDD.t2305 MULT_0.4bit_ADDER_0.A1.t5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t2 VDD.t2304 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X260 VSS.t1680 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t7 a_n15131_n8419.t5 VSS.t1679 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X261 VSS.t435 a_n6641_1380.t2 a_n6611_1406.t3 VSS.t434 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X262 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t0 a_n5059_1406.t3 a_n4879_1406.t2 VSS.t399 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X263 VDD.t4342 SEL1.t4 mux8_0.NAND4F_6.Y.t3 VDD.t4341 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X264 V_FLAG_0.NAND2_0.Y.t1 V_FLAG_0.XOR2_2.Y.t13 a_7173_4939.t0 VSS.t1155 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X265 VDD.t4344 SEL1.t5 mux8_7.NAND4F_5.Y.t5 VDD.t4343 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X266 VDD.t4346 SEL1.t6 mux8_7.NAND4F_0.C.t3 VDD.t4345 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X267 OR8_0.NOT8_0.A5.t5 A5.t3 a_n17677_n22425.t9 VDD.t378 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X268 VDD.t2621 MULT_0.NAND2_11.Y.t7 MULT_0.4bit_ADDER_0.A3.t3 VDD.t2620 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X269 a_n20557_n7799.t2 a_n20587_n8445.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t9 VDD.t2868 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X270 right_shifter_0.buffer_4.inv_1.A.t1 B4.t7 VDD.t3589 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X271 mux8_1.NAND4F_3.Y.t6 mux8_1.NAND4F_2.D.t5 VDD.t1706 VDD.t1705 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X272 mux8_5.A1.t7 a_n12596_n11683.t3 a_n12416_n11683.t4 VSS.t616 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X273 a_11865_n20887.t6 mux8_5.NAND4F_8.Y.t12 VDD.t4304 VDD.t4303 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X274 XOR8_0.S1.t7 a_n12345_n17857.t3 a_n11274_n18115.t4 VSS.t1246 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X275 mux8_2.NAND4F_2.Y.t6 OR8_0.S1.t4 a_8592_n7266.t1 VSS.t304 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X276 a_11386_n7266.t1 mux8_2.NAND4F_2.Y.t9 a_11290_n7266.t0 VSS.t764 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X277 VSS.t378 SEL3.t6 a_3313_4914.t0 VSS.t377 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X278 MULT_0.NAND2_1.Y.t3 A2.t3 VDD.t264 VDD.t263 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X279 a_n20557_n8419.t5 a_n20737_n8419.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t3 VSS.t1416 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X280 a_n368_3164.t1 B0.t1 VDD.t586 VDD.t585 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X281 a_8496_n25478.t0 SEL1.t7 a_8400_n25478.t0 VSS.t1951 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X282 VDD.t3090 SEL0.t11 mux8_5.NAND4F_7.Y.t8 VDD.t3089 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X283 a_n338_3190.t5 a_n368_3164.t2 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t5 VSS.t1412 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X284 a_n9901_2026.t2 a_n9931_1380.t2 mux8_4.A0.t10 VDD.t2183 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X285 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t2 a_n20737_n5154.t2 a_n20557_n5154.t2 VSS.t361 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X286 MULT_0.4bit_ADDER_2.B3.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t7 VDD.t143 VDD.t142 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X287 XOR8_0.S3.t7 B3.t3 a_n11274_n23075.t5 VSS.t1101 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X288 AND8_0.S3.t3 AND8_0.NOT8_0.A3.t7 VDD.t2384 VDD.t678 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X289 a_n18042_2026.t0 A5.t4 VDD.t380 VDD.t379 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X290 a_n13222_1380.t0 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t9 VSS.t1783 VSS.t1782 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X291 mux8_1.NAND4F_4.Y.t4 mux8_1.NAND4F_2.D.t6 VDD.t1708 VDD.t1707 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X292 VDD.t3941 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t10 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t6 VDD.t3940 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X293 right_shifter_0.buffer_2.inv_1.A.t2 B6.t5 VDD.t3531 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X294 a_n7496_3190.t2 SEL3.t7 VSS.t869 VSS.t868 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X295 a_n16483_2026.t0 a_n16663_1406.t2 mux8_7.A0.t0 VDD.t139 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X296 OR8_0.NOT8_0.A3.t5 A3.t4 a_n17677_n19625.t4 VDD.t4072 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X297 VDD.t4135 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t12 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t2 VDD.t4134 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X298 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t0 A4.t0 a_n14490_373.t1 VSS.t707 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X299 a_n12416_n4534.t11 a_n12446_n5180.t2 MULT_0.4bit_ADDER_1.B0.t5 VDD.t3342 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X300 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t12 VDD.t661 VDD.t660 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X301 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t1 MULT_0.4bit_ADDER_2.B2.t15 VDD.t155 VDD.t154 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X302 a_11865_1753.t3 mux8_0.NAND4F_8.Y.t10 VDD.t3505 VDD.t3504 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X303 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t0 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t13 VDD.t298 VDD.t297 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X304 mux8_0.NAND4F_5.Y.t3 mux8_0.NAND4F_4.B.t4 VDD.t847 VDD.t846 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X305 a_n6611_2026.t10 a_n6641_1380.t3 8bit_ADDER_0.S2.t1 VDD.t884 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X306 a_9432_n16422.t0 mux8_4.NAND4F_0.C.t4 a_9336_n16422.t1 VSS.t1496 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X307 VDD.t3591 B4.t8 a_n17677_n21025.t3 VDD.t3590 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X308 mux8_5.NAND4F_2.Y.t8 SEL0.t12 VDD.t3088 VDD.t3087 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X309 VDD.t1385 B7.t0 a_1887_5534.t8 VDD.t1384 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X310 a_11865_n20887.t0 mux8_5.NAND4F_9.Y.t9 mux8_5.inv_0.A.t5 VDD.t686 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X311 VDD.t2278 OR8_0.NOT8_0.A5.t8 OR8_0.S5.t2 VDD.t313 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X312 a_9336_n20950.t1 mux8_5.NAND4F_2.D.t4 VSS.t676 VSS.t675 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X313 MULT_0.NAND2_2.Y.t3 A1.t2 a_n20446_n2915.t1 VSS.t502 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X314 XOR8_0.S7.t8 a_n12347_n34023.t2 a_n11276_n34281.t5 VSS.t485 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X315 AND8_0.NOT8_0.A5.t6 A5.t5 VDD.t382 VDD.t381 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X316 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t1 A6.t3 VDD.t2842 VDD.t2841 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X317 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t13 VDD.t2255 VDD.t2254 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X318 mux8_6.A1.t3 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t7 VDD.t2071 VDD.t2070 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X319 mux8_6.NAND4F_6.Y.t2 right_shifter_0.S7.t4 a_8592_n35462.t0 VSS.t127 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X320 VDD.t2512 right_shifter_0.C.t4 mux8_0.NAND4F_6.Y.t4 VDD.t2511 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X321 a_n20557_n7799.t8 MULT_0.4bit_ADDER_1.A3.t5 VDD.t3935 VDD.t3934 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X322 mux8_3.NAND4F_4.B.t0 SEL0.t13 VSS.t1993 VSS.t1992 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X323 a_8592_n30006.t0 SEL0.t14 a_8496_n30006.t1 VSS.t1991 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X324 a_10459_n35461.t1 SEL0.t15 a_10363_n35461.t1 VSS.t1990 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X325 AND8_0.NOT8_0.A4.t2 B4.t9 VDD.t3593 VDD.t3592 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X326 MULT_0.inv_6.A.t3 B2.t3 a_n24162_n7992.t0 VSS.t838 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X327 a_n10108_n5154.t5 MULT_0.4bit_ADDER_0.B0.t5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t8 VSS.t129 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X328 mux8_2.NAND4F_9.Y.t7 mux8_2.NAND4F_5.Y.t9 VDD.t4294 VDD.t4293 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X329 VDD.t3348 mux8_5.A0.t12 mux8_5.NAND4F_3.Y.t6 VDD.t3347 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X330 a_n19981_n8419.t2 MULT_0.4bit_ADDER_1.B3.t8 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t0 VSS.t1332 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X331 VDD.t2578 B2.t4 a_n17677_n18225.t8 VDD.t2577 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X332 a_n17677_n15425.t3 A0.t2 OR8_0.NOT8_0.A0.t3 VDD.t1654 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X333 a_7548_n2838.t0 SEL1.t8 a_7452_n2838.t1 VSS.t1952 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X334 VDD.t1045 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t14 a_n18998_n7799.t5 VDD.t1044 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X335 VDD.t2144 B3.t4 MULT_0.NAND2_14.Y.t3 VDD.t2143 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X336 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t0 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t12 a_n10884_1406.t5 VSS.t297 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X337 a_n8170_1406.t5 a_n8200_1380.t2 VSS.t154 VSS.t153 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X338 VDD.t4191 A1.t3 MULT_0.inv_7.A.t6 VDD.t4190 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X339 a_n12345_n31115.t1 A6.t4 VDD.t2844 VDD.t2843 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X340 mux8_5.A0.t5 a_n13372_1406.t2 a_n13192_1406.t2 VSS.t669 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X341 mux8_3.inv_0.A.t1 mux8_3.NAND4F_9.Y.t9 a_11865_n11831.t9 VDD.t2615 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X342 VDD.t4348 SEL1.t9 mux8_6.NAND4F_0.C.t3 VDD.t4347 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X343 VSS.t331 right_shifter_0.buffer_3.inv_1.A.t4 right_shifter_0.S4.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X344 VDD.t4350 SEL1.t10 mux8_6.NAND4F_5.Y.t6 VDD.t4349 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X345 a_n23095_1380.t0 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t7 VSS.t959 VSS.t958 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X346 a_n9125_n11683.t5 a_n9305_n11683.t2 mux8_4.A1.t11 VSS.t1054 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X347 a_n9125_n4534.t6 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t12 VDD.t1602 VDD.t1601 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X348 VDD.t3086 SEL0.t16 mux8_8.NAND4F_7.Y.t5 VDD.t3085 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X349 right_shifter_0.buffer_2.inv_1.A.t1 B6.t6 VDD.t3532 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X350 a_n17266_n7799.t7 MULT_0.4bit_ADDER_1.B2.t14 VDD.t4029 VDD.t4028 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X351 a_11386_n26406.t0 mux8_7.NAND4F_6.Y.t9 a_11290_n26406.t1 VSS.t1084 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X352 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t1 MULT_0.4bit_ADDER_0.B1.t4 a_n13399_n5154.t5 VSS.t653 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X353 VDD.t1317 mux8_5.inv_0.A.t7 Y4.t3 VDD.t1316 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X354 V_FLAG_0.XOR2_2.Y.t6 a_3313_4914.t2 a_3493_5534.t6 VDD.t1096 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X355 VDD.t3943 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t11 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t5 VDD.t3942 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X356 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t1 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t13 VDD.t4137 VDD.t4136 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X357 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t4 a_n20737_n8419.t3 a_n20557_n8419.t4 VSS.t1417 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X358 a_n14077_3190.t5 B4.t10 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t9 VSS.t1643 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X359 mux8_8.NAND4F_4.Y.t6 SEL1.t11 VDD.t4352 VDD.t4351 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X360 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t1 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t14 VDD.t300 VDD.t299 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X361 VDD.t3084 SEL0.t17 mux8_5.NAND4F_0.Y.t8 VDD.t3083 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X362 MULT_0.inv_7.A.t5 A1.t4 VDD.t4193 VDD.t4192 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X363 VSS.t1772 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t13 a_n16663_1406.t0 VSS.t1771 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X364 a_16143_n18523.t1 Y1.t5 a_16431_n18523.t4 VDD.t3168 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X365 a_n13192_2026.t3 a_n13222_1380.t2 mux8_5.A0.t11 VDD.t772 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X366 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t3 A2.t4 a_n7909_373.t1 VSS.t118 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X367 a_n12499_373.t0 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t7 VSS.t1666 VSS.t453 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X368 VDD.t1656 A0.t3 MULT_0.NAND2_4.Y.t6 VDD.t1655 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X369 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t11 a_n17548_3190.t2 a_n17368_3810.t11 VDD.t2854 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X370 a_8400_1690.t0 mux8_0.NAND4F_2.D.t5 VSS.t1436 VSS.t1435 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X371 VDD.t1710 mux8_1.NAND4F_2.D.t7 mux8_1.NAND4F_4.Y.t3 VDD.t1709 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X372 VDD.t1145 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t7 a_n19774_2026.t3 VDD.t1144 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X373 mux8_7.inv_0.A.t4 mux8_7.NAND4F_9.Y.t10 a_11865_n25415.t3 VDD.t3282 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X374 a_n23950_3810.t6 SEL3.t8 VDD.t1746 VDD.t1745 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X375 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t2 a_n7676_3190.t3 a_n7496_3810.t5 VDD.t3958 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X376 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t4 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t14 VDD.t2257 VDD.t2256 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X377 VDD.t286 MULT_0.4bit_ADDER_0.B0.t6 a_n10684_n4534.t8 VDD.t285 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X378 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t3 MULT_0.4bit_ADDER_1.A3.t6 a_n20296_n9452.t1 VSS.t1336 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X379 a_10459_n3765.t1 SEL0.t18 a_10363_n3765.t1 VSS.t1997 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X380 a_11194_n25478.t0 mux8_7.NAND4F_0.Y.t9 VSS.t480 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X381 a_n15737_n5180.t1 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t7 VDD.t3989 VDD.t3988 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X382 a_n15131_n5154.t2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t13 MULT_0.4bit_ADDER_1.B1.t2 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X383 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t6 VSS.t2034 VDD.t1981 VDD.t1980 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X384 a_n12314_n31661.t2 A6.t5 VDD.t2813 VDD.t2812 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X385 a_11290_762.t0 mux8_0.NAND4F_1.Y.t9 a_11194_762.t0 VSS.t174 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X386 VDD.t3709 SEL2.t6 mux8_7.NAND4F_2.D.t3 VDD.t3708 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X387 mux8_8.NAND4F_4.B.t0 SEL0.t19 VSS.t1996 VSS.t1995 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X388 mux8_0.NAND4F_9.Y.t4 mux8_0.NAND4F_1.Y.t10 VDD.t1069 VDD.t1068 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X389 mux8_2.NAND4F_0.C.t3 SEL1.t12 VDD.t4354 VDD.t4353 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X390 a_n20083_3190.t5 a_n20113_3164.t2 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t11 VSS.t1327 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X391 a_n9314_n12716.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t13 VSS.t1558 VSS.t428 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X392 VDD.t1626 A4.t1 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t3 VDD.t1625 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X393 mux8_1.NAND4F_1.Y.t1 SEL2.t7 VDD.t3711 VDD.t3710 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X394 a_7548_n16422.t1 SEL1.t13 a_7452_n16422.t1 VSS.t1953 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X395 Y0.t3 mux8_1.inv_0.A.t7 VDD.t1100 VDD.t1099 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X396 buffer_0.inv_1.A.t3 Y7.t4 VDD.t1091 VDD.t1090 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X397 mux8_7.NAND4F_1.Y.t2 mux8_7.NAND4F_0.C.t5 VDD.t182 VDD.t181 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X398 a_n14751_1406.t0 a_n14781_1380.t2 VSS.t266 VSS.t265 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X399 VDD.t3576 mux8_5.NAND4F_3.Y.t9 mux8_5.NAND4F_8.Y.t7 VDD.t3575 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X400 a_n24624_2026.t11 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t12 VDD.t3640 VDD.t3639 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X401 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t8 a_n15896_n6187.t1 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X402 mux8_0.inv_0.A.t1 mux8_0.NAND4F_9.Y.t9 a_11865_1753.t5 VDD.t3122 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X403 a_n12416_n4534.t8 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t12 VDD.t4172 VDD.t4171 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X404 mux8_2.NAND4F_4.B.t3 SEL0.t20 VDD.t3082 VDD.t2982 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X405 XOR8_0.S4.t11 a_n12345_n26161.t2 a_n11274_n26419.t5 VSS.t1876 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X406 mux8_0.NAND4F_3.Y.t4 8bit_ADDER_0.C.t7 VDD.t1579 VDD.t1578 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X407 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t4 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t12 VDD.t3945 VDD.t3944 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X408 a_1887_4914.t3 a_1857_4888.t2 VSS.t1366 VSS.t1365 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X409 VDD.t1262 mux8_1.NAND4F_4.B.t5 mux8_1.NAND4F_3.Y.t8 VDD.t1261 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X410 mux8_1.NAND4F_5.Y.t1 SEL2.t8 VDD.t3713 VDD.t3712 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X411 a_11386_n35462.t0 mux8_6.NAND4F_6.Y.t9 a_11290_n35462.t1 VSS.t123 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X412 VDD.t302 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t15 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t2 VDD.t301 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X413 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t0 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t14 VDD.t4139 VDD.t4138 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X414 VDD.t3293 mux8_0.inv_0.A.t8 C.t3 VDD.t3292 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X415 mux8_1.NAND4F_8.Y.t5 mux8_1.NAND4F_4.Y.t9 a_11386_n2838.t0 VSS.t785 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X416 a_11290_n30006.t0 mux8_8.NAND4F_3.Y.t9 a_11194_n30006.t1 VSS.t712 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X417 VDD.t2707 mux8_8.inv_0.A.t7 Y6.t3 VDD.t2706 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X418 mux8_5.NAND4F_0.C.t3 SEL1.t14 VDD.t4356 VDD.t4355 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X419 a_n12345_n17569.t1 A1.t5 VDD.t4195 VDD.t4194 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X420 VDD.t1658 A0.t4 a_n12316_n15299.t2 VDD.t1657 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X421 a_n10684_n11063.t9 a_n10714_n11709.t2 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t9 VDD.t2005 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X422 a_n13399_n11683.t1 MULT_0.inv_9.Y.t8 VSS.t1811 VSS.t1810 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X423 MULT_0.4bit_ADDER_2.B3.t3 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t7 a_n18305_n9452.t1 VSS.t67 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X424 a_n23065_1406.t2 a_n23095_1380.t2 VSS.t799 VSS.t798 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X425 MULT_0.4bit_ADDER_0.A0.t0 MULT_0.NAND2_4.Y.t7 VSS.t558 VSS.t557 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X426 a_n9931_1380.t1 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t8 VDD.t1728 VDD.t1727 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X427 VDD.t3311 MULT_0.inv_15.Y.t4 a_n20557_n11063.t11 VDD.t3310 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X428 MULT_0.NAND2_15.Y.t5 B3.t5 VDD.t2146 VDD.t2145 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X429 a_11194_762.t1 mux8_0.NAND4F_7.Y.t9 VSS.t737 VSS.t618 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X430 a_n5918_373.t1 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t7 VSS.t1535 VSS.t211 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X431 mux8_6.inv_0.A.t1 mux8_6.NAND4F_9.Y.t10 a_11865_n34471.t8 VDD.t695 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X432 VSS.t1102 B3.t6 right_shifter_0.buffer_5.inv_1.A.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X433 mux8_1.NAND4F_0.Y.t4 mux8_1.NAND4F_0.C.t4 VDD.t1420 VDD.t1419 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X434 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t5 a_n13531_3164.t3 a_n14077_3810.t11 VDD.t2731 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X435 VSS.t169 right_shifter_0.buffer_7.inv_1.A.t4 right_shifter_0.S0.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X436 mux8_0.NAND4F_9.Y.t0 mux8_0.NAND4F_5.Y.t9 a_11386_762.t0 VSS.t626 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X437 a_n20659_3810.t5 B6.t7 VDD.t3534 VDD.t3533 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X438 a_n1588_1406.t3 a_n1618_1380.t3 VSS.t621 VSS.t620 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X439 VSS.t173 OR8_0.NOT8_0.A4.t7 OR8_0.S4.t0 VSS.t172 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X440 VDD.t2325 B1.t4 a_n4205_3810.t9 VDD.t2324 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X441 a_n15707_n11063.t6 a_n15887_n11683.t2 mux8_7.A1.t5 VDD.t1109 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X442 VDD.t3715 SEL2.t9 mux8_6.NAND4F_2.D.t3 VDD.t3714 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X443 a_n11723_n12716.t1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t8 VSS.t1567 VSS.t428 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X444 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t1 a_n8350_1406.t3 a_n8170_1406.t2 VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X445 VDD.t4149 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t8 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t5 VDD.t4148 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X446 a_n12347_n33735.t1 A7.t1 VDD.t2289 VDD.t2288 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X447 VDD.t1628 A4.t2 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t2 VDD.t1627 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X448 mux8_8.A1.t10 a_n19178_n11683.t2 a_n18998_n11063.t8 VDD.t2484 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X449 a_3493_5534.t3 V_FLAG_0.XOR2_2.B.t13 VDD.t975 VDD.t974 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X450 VDD.t1979 VSS.t2035 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t5 VDD.t1978 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X451 a_7452_n21878.t0 SEL2.t10 VSS.t1703 VSS.t677 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X452 OR8_0.S1.t0 OR8_0.NOT8_0.A1.t7 VDD.t2479 VDD.t2478 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X453 a_9528_1690.t0 mux8_0.NAND4F_4.B.t5 a_9432_1690.t0 VSS.t425 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X454 mux8_4.NAND4F_7.Y.t5 SEL0.t21 VDD.t3081 VDD.t3080 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X455 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t6 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t14 VDD.t1436 VDD.t1435 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X456 VDD.t598 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t12 a_n9125_n7799.t5 VDD.t597 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X457 mux8_6.NAND4F_1.Y.t2 mux8_6.NAND4F_0.C.t5 VDD.t326 VDD.t325 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X458 VDD.t266 A2.t5 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t6 VDD.t265 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X459 VDD.t3079 SEL0.t22 mux8_2.NAND4F_0.Y.t3 VDD.t3078 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X460 mux8_1.inv_0.A.t5 mux8_1.NAND4F_9.Y.t9 a_11865_n2775.t0 VDD.t1318 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X461 a_n11276_n34281.t0 a_n12347_n33735.t2 VSS.t780 VSS.t779 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X462 VDD.t416 NOT8_0.S7.t5 mux8_6.NAND4F_7.Y.t6 VDD.t415 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X463 mux8_3.NAND4F_9.Y.t1 mux8_3.NAND4F_5.Y.t10 VDD.t924 VDD.t923 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X464 mux8_3.NAND4F_7.Y.t0 SEL2.t11 VDD.t3717 VDD.t3716 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X465 mux8_0.NAND4F_7.Y.t8 SEL0.t23 VDD.t3077 VDD.t3076 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X466 VDD.t304 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t16 a_n13192_2026.t0 VDD.t303 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X467 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t6 a_n11640_1406.t2 a_n11460_2026.t11 VDD.t1575 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X468 a_n16513_1380.t0 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t8 VSS.t1351 VSS.t1350 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X469 a_16143_n19505.t2 Y5.t4 a_15855_n19505.t2 VDD.t1528 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X470 a_n19774_2026.t8 a_n19954_1406.t2 mux8_8.A0.t9 VDD.t1544 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X471 8bit_ADDER_0.S1.t11 a_n3500_1406.t2 a_n3320_2026.t11 VDD.t1542 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X472 VSS.t1023 VSS.t1021 a_n8549_n11683.t0 VSS.t1022 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X473 VDD.t2684 MULT_0.NAND2_15.Y.t7 MULT_0.inv_15.Y.t3 VDD.t2683 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X474 mux8_2.NAND4F_7.Y.t1 SEL2.t12 VDD.t3719 VDD.t3718 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X475 a_n8170_2026.t5 A2.t6 VDD.t268 VDD.t267 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X476 mux8_8.NAND4F_0.C.t3 SEL1.t15 VDD.t4358 VDD.t4357 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X477 VDD.t1134 mux8_8.NAND4F_2.D.t4 mux8_8.NAND4F_3.Y.t0 VDD.t1133 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X478 a_n20557_n7799.t5 MULT_0.4bit_ADDER_1.B3.t9 VDD.t2715 VDD.t2714 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X479 VDD.t3721 SEL2.t13 mux8_1.NAND4F_5.Y.t0 VDD.t3720 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X480 a_n13975_n5154.t0 a_n14005_n5180.t2 VSS.t751 VSS.t750 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X481 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t4 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t7 VDD.t4045 VDD.t4044 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X482 a_547_1406.t5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t15 8bit_ADDER_0.S0.t10 VSS.t1140 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X483 a_10363_n11894.t0 mux8_3.NAND4F_0.C.t4 a_10267_n11894.t0 VSS.t1321 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X484 mux8_6.NAND4F_0.C.t2 SEL1.t16 VDD.t4359 VDD.t4347 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X485 a_8400_n17350.t0 SEL2.t14 VSS.t1704 VSS.t60 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X486 VSS.t1628 B6.t8 NOT8_0.S6.t0 VSS.t1627 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X487 mux8_0.NAND4F_8.Y.t4 mux8_0.NAND4F_2.Y.t9 VDD.t1742 VDD.t1741 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X488 VDD.t849 mux8_0.NAND4F_4.B.t6 mux8_0.NAND4F_1.Y.t3 VDD.t848 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X489 a_n11840_n11683.t2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t13 mux8_5.A1.t5 VSS.t1042 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X490 mux8_2.NAND4F_8.Y.t0 mux8_2.NAND4F_3.Y.t9 VDD.t81 VDD.t80 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X491 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t15 VDD.t3660 VDD.t3659 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X492 a_11386_762.t1 mux8_0.NAND4F_6.Y.t9 a_11290_762.t1 VSS.t867 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X493 VDD.t4361 SEL1.t17 mux8_2.NAND4F_2.Y.t1 VDD.t4360 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X494 VSS.t7 MULT_0.4bit_ADDER_1.A2.t5 a_n16690_n8419.t4 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X495 mux8_4.NAND4F_0.C.t0 SEL1.t18 VSS.t1955 VSS.t1954 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X496 a_n19198_1406.t5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t12 mux8_8.A0.t0 VSS.t411 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X497 a_n12316_n34281.t2 A7.t2 VDD.t2291 VDD.t2290 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X498 mux8_5.NAND4F_7.Y.t7 SEL0.t24 VDD.t3075 VDD.t3074 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X499 mux8_0.NAND4F_2.Y.t2 VSS.t2036 VDD.t1977 VDD.t1976 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X500 VDD.t3594 B4.t11 NOT8_0.S4.t3 VDD.t887 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X501 mux8_1.NAND4F_4.Y.t2 AND8_0.S0.t4 VDD.t578 VDD.t577 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X502 a_n16690_n5154.t1 MULT_0.4bit_ADDER_0.A2.t5 VSS.t112 VSS.t111 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X503 VDD.t564 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t2 VDD.t563 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X504 VDD.t4363 SEL1.t19 mux8_0.NAND4F_4.Y.t8 VDD.t4362 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X505 VSS.t1160 A7.t3 a_n24048_1406.t2 VSS.t1159 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X506 a_n10684_n11063.t7 MULT_0.4bit_ADDER_2.B0.t12 VDD.t1883 VDD.t1882 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X507 a_n13975_n11683.t2 a_n14155_n11683.t2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t6 VSS.t1047 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X508 VSS.t440 B5.t3 right_shifter_0.buffer_3.inv_1.A.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X509 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t1 A4.t3 VDD.t1630 VDD.t1629 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X510 mux8_4.NAND4F_1.Y.t4 XOR8_0.S3.t12 a_9528_n17350.t0 VSS.t16 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X511 V_FLAG_0.XOR2_2.B.t1 A7.t4 a_2463_4914.t2 VSS.t1161 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X512 VSS.t1833 a_n15737_n5180.t3 a_n15707_n5154.t4 VSS.t1832 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X513 VDD.t210 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t9 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t3 VDD.t209 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X514 VDD.t2438 MULT_0.inv_14.Y.t4 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t6 VDD.t2437 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X515 VSS.t1212 a_n12345_n20526.t2 a_n11274_n21072.t2 VSS.t1211 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X516 a_n3350_1380.t0 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t9 VSS.t402 VSS.t401 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X517 VDD.t1434 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t15 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t5 VDD.t1433 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X518 VDD.t3884 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t12 a_n12416_n7799.t2 VDD.t3883 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X519 a_9336_n16422.t0 mux8_4.NAND4F_2.D.t4 VSS.t55 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X520 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t0 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t7 a_n12499_373.t1 VSS.t453 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X521 MULT_0.4bit_ADDER_1.A1.t3 MULT_0.inv_7.A.t7 VDD.t2078 VDD.t2077 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X522 VDD.t4365 SEL1.t20 mux8_5.NAND4F_2.Y.t6 VDD.t4364 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X523 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t6 MULT_0.4bit_ADDER_0.B2.t5 VDD.t2910 VDD.t2909 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X524 VDD.t2002 Y4.t4 a_15855_n19505.t5 VDD.t2001 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X525 OR8_0.S3.t3 OR8_0.NOT8_0.A3.t7 VDD.t729 VDD.t315 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X526 mux8_5.inv_0.A.t4 mux8_5.NAND4F_9.Y.t10 a_11865_n20887.t1 VDD.t687 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X527 VSS.t1455 mux8_0.NAND4F_9.Y.t10 mux8_0.inv_0.A.t2 VSS.t1454 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X528 a_n12314_n29052.t5 A5.t6 VDD.t384 VDD.t383 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X529 VDD.t1264 mux8_1.NAND4F_4.B.t6 mux8_1.NAND4F_1.Y.t7 VDD.t1263 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X530 mux8_5.NAND4F_2.D.t3 SEL2.t15 VDD.t3723 VDD.t3722 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X531 VSS.t1278 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t8 a_n18422_n5154.t3 VSS.t1277 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X532 VDD.t2815 A6.t6 a_n12314_n31661.t1 VDD.t2814 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X533 VDD.t3073 SEL0.t25 mux8_0.NAND4F_0.Y.t8 VDD.t3072 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X534 a_n24213_n2915.t0 B0.t2 VSS.t281 VSS.t280 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X535 a_n15737_n11709.t1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t8 VDD.t833 VDD.t832 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X536 MULT_0.SO.t0 MULT_0.NAND2_3.Y.t7 VSS.t76 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X537 mux8_1.NAND4F_7.Y.t4 NOT8_0.S0.t4 VDD.t808 VDD.t807 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X538 a_8496_n30006.t0 SEL1.t21 a_8400_n30006.t1 VSS.t1956 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X539 VDD.t4366 SEL1.t22 mux8_2.NAND4F_0.C.t2 VDD.t4353 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X540 mux8_3.NAND4F_4.Y.t4 SEL1.t23 VDD.t4368 VDD.t4367 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X541 a_n14077_3810.t2 SEL3.t9 VDD.t1748 VDD.t1747 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X542 a_1887_5534.t3 A7.t5 VDD.t2293 VDD.t2292 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X543 a_n16483_2026.t6 a_n16513_1380.t2 mux8_7.A0.t6 VDD.t1483 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X544 mux8_6.A0.t11 a_n23245_1406.t2 a_n23065_1406.t5 VSS.t1256 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X545 VDD.t4151 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t9 a_n18998_n7799.t11 VDD.t4150 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X546 a_n4205_3810.t6 SEL3.t10 VDD.t1750 VDD.t1749 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X547 VDD.t1102 mux8_1.inv_0.A.t8 Y0.t2 VDD.t1101 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X548 VDD.t2652 mux8_8.NAND4F_0.C.t4 mux8_8.NAND4F_0.Y.t1 VDD.t2651 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X549 a_n6611_2026.t0 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t7 VDD.t87 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X550 a_n15896_n6187.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t14 VSS.t216 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X551 MULT_0.4bit_ADDER_1.B1.t5 a_n15887_n5154.t2 a_n15707_n4534.t5 VDD.t2268 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X552 a_9336_n7266.t0 mux8_2.NAND4F_2.D.t4 VSS.t1471 VSS.t1470 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X553 VDD.t3071 SEL0.t26 mux8_2.NAND4F_4.B.t2 VDD.t2982 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X554 VDD.t35 mux8_2.NAND4F_8.Y.t10 a_11865_n7203.t3 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X555 mux8_4.A1.t10 a_n9305_n11683.t3 a_n9125_n11683.t4 VSS.t1055 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X556 a_n11274_n26419.t0 a_n12345_n25873.t2 VSS.t306 VSS.t305 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X557 a_10363_n34534.t0 mux8_6.NAND4F_0.C.t6 a_10267_n34534.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X558 left_shifter_0.buffer_7.inv_1.A.t3 B1.t5 VDD.t2326 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X559 VSS.t229 a_3463_4888.t3 a_3493_4914.t2 VSS.t228 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X560 a_n9125_n4534.t8 VSS.t2037 VDD.t1975 VDD.t1974 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X561 mux8_8.NAND4F_7.Y.t4 SEL0.t27 VDD.t3070 VDD.t3069 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X562 mux8_7.NAND4F_0.C.t0 SEL1.t24 VSS.t1958 VSS.t1957 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X563 C.t2 mux8_0.inv_0.A.t9 VDD.t3295 VDD.t3294 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X564 a_n23374_3190.t0 a_n23404_3164.t2 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t0 VSS.t393 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X565 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t4 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t16 VDD.t1432 VDD.t1431 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X566 a_n12316_n15299.t1 A0.t5 VDD.t1660 VDD.t1659 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X567 VDD.t1504 mux8_8.NAND4F_2.D.t5 mux8_8.NAND4F_4.Y.t3 VDD.t1503 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X568 VSS.t1104 B3.t7 a_n23992_n18833.t1 VSS.t1103 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X569 OR8_0.NOT8_0.A0.t6 B0.t3 VSS.t283 VSS.t282 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X570 a_n23065_2026.t5 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t8 VDD.t1873 VDD.t1872 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X571 a_n18042_1406.t1 a_n18072_1380.t3 VSS.t1067 VSS.t1066 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X572 mux8_5.NAND4F_0.Y.t7 SEL0.t28 VDD.t3068 VDD.t3067 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X573 a_n12345_n23105.t1 A3.t5 VDD.t4074 VDD.t4073 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X574 MULT_0.NAND2_11.Y.t5 A3.t6 VDD.t4076 VDD.t4075 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X575 VDD.t120 mux8_4.NAND4F_2.D.t5 mux8_4.NAND4F_0.Y.t1 VDD.t119 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X576 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t7 a_n5918_373.t0 VSS.t211 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X577 a_11865_n25415.t9 mux8_7.NAND4F_8.Y.t9 VDD.t4252 VDD.t4251 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X578 mux8_8.NAND4F_2.D.t3 SEL2.t16 VDD.t3725 VDD.t3724 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X579 a_n14005_n11709.t0 MULT_0.inv_9.Y.t9 VSS.t1813 VSS.t1812 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X580 a_8400_n30934.t0 SEL2.t17 VSS.t1705 VSS.t742 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X581 V_FLAG_0.XOR2_0.Y.t6 A7.t6 a_5773_4912.t2 VSS.t1162 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X582 VDD.t1752 SEL3.t11 a_n29_2026.t2 VDD.t1751 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X583 mux8_6.NAND4F_2.D.t2 SEL2.t18 VDD.t3726 VDD.t3714 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X584 a_n17677_n19625.t9 B3.t8 VDD.t2148 VDD.t2147 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X585 a_n9901_1406.t3 a_n9931_1380.t3 VSS.t1114 VSS.t1113 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X586 mux8_7.NAND4F_5.Y.t2 left_shifter_0.S5.t4 a_7644_n26406.t0 VSS.t242 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X587 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t6 a_n18072_1380.t4 a_n18042_2026.t6 VDD.t2045 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X588 a_n24624_1406.t0 a_n24804_1406.t3 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t5 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X589 MULT_0.4bit_ADDER_2.B3.t4 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t8 VDD.t572 VDD.t571 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X590 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t3 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t7 VDD.t1694 VDD.t1693 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X591 a_n17677_n23825.t0 A6.t7 OR8_0.NOT8_0.A6.t3 VDD.t2816 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X592 mux8_4.NAND4F_2.D.t0 SEL2.t19 VSS.t1707 VSS.t1706 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X593 mux8_6.NAND4F_4.Y.t6 SEL1.t25 VDD.t4370 VDD.t4369 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X594 VDD.t1093 Y7.t5 buffer_0.inv_1.A.t2 VDD.t1092 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X595 a_n10786_3810.t6 a_n10966_3190.t2 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t6 VDD.t1446 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X596 mux8_8.NAND4F_1.Y.t2 XOR8_0.S6.t12 a_9528_n30934.t0 VSS.t736 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X597 VDD.t909 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t8 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t1 VDD.t908 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X598 mux8_5.NAND4F_8.Y.t8 mux8_5.NAND4F_3.Y.t10 VDD.t3578 VDD.t3577 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X599 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t5 a_n16822_3164.t3 a_n17368_3810.t5 VDD.t2886 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X600 a_10363_1690.t0 mux8_0.NAND4F_0.C.t5 a_10267_1690.t1 VSS.t316 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X601 a_n12416_n4534.t2 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t10 VDD.t212 VDD.t211 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X602 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t0 MULT_0.4bit_ADDER_1.B0.t12 VDD.t2498 VDD.t2497 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X603 VDD.t2709 mux8_8.inv_0.A.t8 Y6.t2 VDD.t2708 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X604 mux8_1.NAND4F_5.Y.t4 left_shifter_0.S0.t4 VDD.t2381 VDD.t2380 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X605 VSS.t1044 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t14 a_n12596_n11683.t0 VSS.t1043 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X606 a_n4879_1406.t4 a_n4909_1380.t2 VSS.t1226 VSS.t1225 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X607 VSS.t1506 mux8_7.NAND4F_9.Y.t11 mux8_7.inv_0.A.t0 VSS.t1505 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X608 VDD.t2580 B2.t5 a_n7496_3810.t11 VDD.t2579 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X609 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t8 VDD.t715 VDD.t714 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X610 a_n12314_n23651.t5 A3.t7 VDD.t4078 VDD.t4077 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X611 MULT_0.inv_15.Y.t2 MULT_0.NAND2_15.Y.t8 VDD.t2685 VDD.t2683 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X612 mux8_0.NAND4F_2.D.t3 SEL2.t20 VDD.t3728 VDD.t3727 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X613 VDD.t917 mux8_2.NAND4F_4.Y.t10 mux8_2.NAND4F_8.Y.t2 VDD.t916 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X614 a_n17266_n8419.t4 a_n17446_n8419.t3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t4 VSS.t357 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X615 a_5197_5532.t3 A7.t7 VDD.t2295 VDD.t2294 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X616 left_shifter_0.buffer_5.inv_1.A.t3 B3.t9 VDD.t2149 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X617 VDD.t1662 A0.t6 AND8_0.NOT8_0.A0.t3 VDD.t1661 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X618 a_11194_n30006.t0 mux8_8.NAND4F_0.Y.t9 VSS.t78 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X619 mux8_4.A0.t9 a_n10081_1406.t3 a_n9901_2026.t11 VDD.t1566 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X620 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t11 B0.t4 a_n914_3190.t5 VSS.t284 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X621 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t6 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t7 VDD.t1359 VDD.t1358 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X622 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t3 a_n17446_n5154.t2 a_n17266_n5154.t2 VSS.t1222 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X623 VDD.t574 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t9 MULT_0.4bit_ADDER_2.B3.t5 VDD.t573 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X624 OR8_0.NOT8_0.A6.t6 B6.t9 VSS.t1629 VSS.t177 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X625 NOT8_0.S2.t3 B2.t6 VDD.t2581 VDD.t1011 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X626 MULT_0.inv_7.A.t3 A1.t6 a_n24162_n9284.t1 VSS.t1292 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X627 a_7548_n7266.t0 SEL1.t26 a_7452_n7266.t1 VSS.t1959 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X628 VDD.t4372 SEL1.t27 mux8_2.NAND4F_6.Y.t6 VDD.t4371 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X629 mux8_2.NAND4F_9.Y.t4 mux8_2.NAND4F_1.Y.t9 VDD.t657 VDD.t656 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X630 VDD.t3128 mux8_7.NAND4F_2.D.t4 mux8_7.NAND4F_0.Y.t7 VDD.t3127 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X631 mux8_5.NAND4F_0.Y.t4 mux8_5.A1.t13 a_10459_n20950.t0 VSS.t674 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X632 VDD.t3901 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t14 a_n16483_2026.t11 VDD.t3900 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X633 a_n19804_1380.t0 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t8 VSS.t568 VSS.t567 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X634 VDD.t1387 B7.t1 a_n23950_3810.t0 VDD.t1386 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X635 VDD.t1754 SEL3.t12 a_n20839_3190.t1 VDD.t1753 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X636 a_n20557_n11063.t10 MULT_0.inv_15.Y.t5 VDD.t3313 VDD.t3312 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X637 VDD.t2297 A7.t8 a_n12316_n34281.t1 VDD.t2296 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X638 VDD.t4080 A3.t8 MULT_0.NAND2_15.Y.t3 VDD.t4079 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X639 a_n21333_2026.t0 a_n21513_1406.t2 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t0 VDD.t724 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X640 8bit_ADDER_0.S2.t7 a_n6791_1406.t2 a_n6611_2026.t6 VDD.t1230 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X641 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t6 a_n4909_1380.t3 a_n4879_2026.t3 VDD.t1182 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X642 a_11865_n34471.t4 mux8_6.NAND4F_8.Y.t9 VDD.t983 VDD.t982 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X643 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t6 VSS.t2038 VDD.t1973 VDD.t1972 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X644 VDD.t1233 AND8_0.S6.t4 mux8_8.NAND4F_4.Y.t0 VDD.t1232 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X645 mux8_7.A1.t4 a_n15887_n11683.t3 a_n15707_n11063.t10 VDD.t1615 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X646 VSS.t467 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t8 a_n18422_n11683.t5 VSS.t466 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X647 a_n18998_n5154.t1 a_n19178_n5154.t3 MULT_0.4bit_ADDER_1.B2.t3 VSS.t338 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X648 VDD.t2797 mux8_3.NAND4F_2.D.t4 mux8_3.NAND4F_3.Y.t4 VDD.t2796 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X649 mux8_5.NAND4F_8.Y.t5 mux8_5.NAND4F_0.Y.t9 VDD.t3414 VDD.t3413 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X650 mux8_6.NAND4F_5.Y.t2 left_shifter_0.S7.t4 a_7644_n35462.t0 VSS.t167 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X651 a_n12446_n8445.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t8 VSS.t1929 VSS.t1928 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X652 a_n20557_n11683.t2 a_n20587_n11709.t2 VSS.t392 VSS.t391 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X653 mux8_7.A0.t1 a_n16663_1406.t3 a_n16483_1406.t2 VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X654 VSS.t299 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t13 a_n11640_1406.t0 VSS.t298 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X655 a_664_373.t1 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t7 VSS.t1564 VSS.t939 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X656 VDD.t2079 MULT_0.inv_7.A.t8 MULT_0.4bit_ADDER_1.A1.t2 VDD.t2077 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X657 mux8_7.NAND4F_2.D.t0 SEL2.t21 VSS.t1709 VSS.t1708 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X658 VDD.t2481 OR8_0.NOT8_0.A1.t8 OR8_0.S1.t1 VDD.t2480 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X659 VDD.t3463 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t9 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t5 VDD.t3462 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X660 VDD.t1971 VSS.t2039 a_n9125_n7799.t11 VDD.t1970 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X661 mux8_7.NAND4F_6.Y.t8 SEL0.t29 VDD.t3066 VDD.t3065 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X662 a_n12314_n18115.t8 A1.t7 VDD.t4197 VDD.t4196 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X663 a_n20757_1406.t2 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t13 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t2 VSS.t1490 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X664 VDD.t386 A5.t7 a_n12314_n29052.t4 VDD.t385 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X665 VDD.t184 mux8_7.NAND4F_0.C.t6 mux8_7.NAND4F_7.Y.t2 VDD.t183 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X666 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t4 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t8 VDD.t3995 VDD.t3994 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X667 a_15855_n19505.t4 Y4.t5 VDD.t2004 VDD.t2003 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X668 MULT_0.4bit_ADDER_0.B0.t0 MULT_0.NAND2_2.Y.t7 VSS.t526 VSS.t525 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X669 VDD.t3360 mux8_4.NAND4F_4.B.t5 mux8_4.NAND4F_4.Y.t3 VDD.t3359 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X670 a_9432_n2838.t0 mux8_1.NAND4F_0.C.t5 a_9336_n2838.t1 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X671 a_10459_n8193.t1 SEL0.t30 a_10363_n8193.t1 VSS.t1998 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X672 VDD.t2500 MULT_0.4bit_ADDER_1.B0.t13 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t1 VDD.t2499 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X673 NOT8_0.S2.t2 B2.t7 VDD.t2582 VDD.t1013 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X674 a_n17677_n15425.t9 B0.t5 VDD.t588 VDD.t587 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X675 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t9 a_n10864_n5154.t2 a_n10684_n4534.t9 VDD.t2650 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X676 MULT_0.S1.t11 a_n9305_n5154.t3 a_n9125_n4534.t3 VDD.t367 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X677 VDD.t4082 A3.t9 MULT_0.inv_13.A.t3 VDD.t4081 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X678 VDD.t1202 XOR8_0.S5.t12 mux8_7.NAND4F_1.Y.t4 VDD.t1201 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X679 mux8_8.NAND4F_3.Y.t6 mux8_8.NAND4F_2.D.t6 VDD.t1506 VDD.t1505 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X680 a_n12314_n21072.t8 a_n12345_n20526.t3 XOR8_0.S2.t5 VDD.t2414 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X681 VDD.t4374 SEL1.t28 mux8_3.NAND4F_0.C.t3 VDD.t4373 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X682 a_10267_n11894.t1 mux8_3.NAND4F_2.D.t5 VSS.t1379 VSS.t1378 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X683 a_11290_1690.t0 mux8_0.NAND4F_3.Y.t9 a_11194_1690.t1 VSS.t174 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X684 VSS.t469 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t9 a_n18422_n11683.t4 VSS.t468 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X685 V_FLAG_0.NAND2_0.Y.t6 V_FLAG_0.XOR2_0.Y.t12 VDD.t4125 VDD.t4124 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X686 a_n914_3810.t9 a_n368_3164.t3 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t8 VDD.t1644 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X687 VDD.t4084 A3.t10 a_n11460_2026.t5 VDD.t4083 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X688 VDD.t3730 SEL2.t22 mux8_1.NAND4F_2.D.t3 VDD.t3729 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X689 VDD.t3064 SEL0.t31 mux8_3.NAND4F_4.B.t3 VDD.t3001 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X690 mux8_5.A0.t8 a_n13372_1406.t3 a_n13192_2026.t6 VDD.t1164 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X691 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t3 MULT_0.4bit_ADDER_0.A0.t4 a_n10423_n6187.t1 VSS.t130 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X692 VDD.t1885 MULT_0.4bit_ADDER_2.B0.t13 a_n10684_n11063.t8 VDD.t1884 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X693 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t7 a_n14155_n11683.t3 a_n13975_n11683.t1 VSS.t1048 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X694 a_n12416_n4534.t4 a_n12596_n5154.t2 MULT_0.4bit_ADDER_1.B0.t6 VDD.t1151 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X695 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t4 MULT_0.4bit_ADDER_0.B1.t5 VDD.t1331 VDD.t1330 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X696 a_n12316_n15299.t3 a_n12347_n14753.t2 XOR8_0.S0.t3 VDD.t1148 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X697 a_9528_n17350.t1 mux8_4.NAND4F_4.B.t6 a_9432_n17350.t1 VSS.t1545 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X698 a_n7496_3810.t2 SEL3.t13 VDD.t1756 VDD.t1755 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X699 a_n17266_n11683.t5 a_n17296_n11709.t2 VSS.t1316 VSS.t1315 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X700 a_n8432_n12716.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t7 VSS.t429 VSS.t428 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X701 VDD.t1712 mux8_1.NAND4F_2.D.t8 mux8_1.NAND4F_3.Y.t5 VDD.t1711 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X702 VDD.t2328 B1.t6 MULT_0.NAND2_10.Y.t6 VDD.t2327 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X703 VSS.t344 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t9 a_n15131_n5154.t5 VSS.t343 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X704 AND8_0.S2.t3 AND8_0.NOT8_0.A2.t7 VDD.t3481 VDD.t674 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X705 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t6 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t10 VDD.t3465 VDD.t3464 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X706 VDD.t2668 mux8_3.NAND4F_0.C.t5 mux8_3.NAND4F_0.Y.t6 VDD.t2667 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X707 mux8_2.NAND4F_8.Y.t3 mux8_2.NAND4F_4.Y.t11 a_11386_n7266.t0 VSS.t454 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X708 VDD.t4282 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t9 a_n12416_n7799.t8 VDD.t4281 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X709 VDD.t894 B5.t4 a_n12314_n29052.t2 VDD.t893 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X710 VDD.t420 mux8_6.NAND4F_2.D.t4 mux8_6.NAND4F_3.Y.t1 VDD.t419 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X711 VDD.t3997 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t9 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t3 VDD.t3996 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X712 a_8400_n2838.t0 mux8_1.NAND4F_2.D.t9 VSS.t852 VSS.t851 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X713 a_15855_n19505.t3 Y4.t6 VDD.t2732 VDD.t2421 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=1.3268 ps=9.18 w=4.28 l=0.15
X714 MULT_0.NAND2_0.Y.t6 A3.t11 VDD.t4086 VDD.t4085 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X715 mux8_6.NAND4F_6.Y.t8 SEL0.t32 VDD.t3063 VDD.t3062 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X716 VDD.t1476 ZFLAG_0.NAND2_0.Y.t7 Z.t3 VDD.t1475 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X717 mux8_0.NAND4F_8.Y.t3 mux8_0.NAND4F_0.Y.t10 VDD.t1247 VDD.t1246 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X718 a_n20557_n5154.t1 a_n20737_n5154.t3 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t1 VSS.t362 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X719 VDD.t1632 A4.t4 a_n12314_n26419.t9 VDD.t1631 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X720 VSS.t150 OR8_0.NOT8_0.A0.t7 OR8_0.S0.t0 VSS.t149 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X721 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t0 B6.t10 a_n20659_3190.t5 VSS.t1630 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X722 VDD.t444 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t8 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t1 VDD.t443 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X723 VSS.t1817 MULT_0.4bit_ADDER_1.B2.t15 a_n17446_n8419.t0 VSS.t1816 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X724 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t2 MULT_0.4bit_ADDER_2.B0.t14 VDD.t1887 VDD.t1886 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X725 a_n10714_n5180.t0 MULT_0.4bit_ADDER_0.A0.t5 VDD.t1290 VDD.t1289 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X726 MULT_0.4bit_ADDER_1.B0.t7 a_n12596_n5154.t3 a_n12416_n4534.t5 VDD.t1152 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X727 VDD.t663 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t13 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t1 VDD.t662 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X728 VDD.t2051 mux8_7.NAND4F_4.B.t5 mux8_7.NAND4F_4.Y.t8 VDD.t2050 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X729 VDD.t2799 mux8_3.NAND4F_2.D.t6 mux8_3.NAND4F_4.Y.t7 VDD.t2798 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X730 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t9 VDD.t835 VDD.t834 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X731 a_n17677_n23825.t9 B6.t11 VDD.t3536 VDD.t3535 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X732 VDD.t3266 XOR8_0.S7.t12 mux8_6.NAND4F_1.Y.t6 VDD.t3265 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X733 a_n17005_n12716.t0 MULT_0.4bit_ADDER_2.B2.t16 VSS.t71 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X734 mux8_8.NAND4F_0.Y.t0 mux8_8.NAND4F_0.C.t5 VDD.t2654 VDD.t2653 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X735 a_9528_n2838.t1 mux8_1.NAND4F_4.B.t7 a_9432_n2838.t1 VSS.t627 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X736 VDD.t2329 B1.t7 right_shifter_0.buffer_7.inv_1.A.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X737 VDD.t4088 A3.t12 MULT_0.NAND2_0.Y.t5 VDD.t4087 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X738 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t15 VDD.t450 VDD.t449 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X739 VDD.t104 MULT_0.4bit_ADDER_1.A1.t4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t0 VDD.t103 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X740 Y6.t1 mux8_8.inv_0.A.t9 VDD.t2711 VDD.t2710 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X741 VDD.t1634 A4.t5 AND8_0.NOT8_0.A4.t3 VDD.t1633 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X742 a_n10210_3190.t2 a_n10240_3164.t3 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t1 VSS.t332 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X743 VDD.t2865 mux8_7.NAND4F_1.Y.t9 mux8_7.NAND4F_9.Y.t7 VDD.t2864 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X744 VDD.t4313 MULT_0.4bit_ADDER_1.A3.t7 a_n20557_n7799.t7 VDD.t4312 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X745 a_n8549_n11683.t3 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t14 mux8_4.A1.t5 VSS.t1559 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X746 a_10267_n34534.t0 mux8_6.NAND4F_2.D.t5 VSS.t201 VSS.t200 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X747 VDD.t4090 A3.t13 a_n12314_n23651.t4 VDD.t4089 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X748 VDD.t2330 B1.t8 left_shifter_0.buffer_7.inv_1.A.t2 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X749 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t1 MULT_0.4bit_ADDER_1.B3.t10 a_n19981_n8419.t1 VSS.t1333 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X750 VDD.t4296 mux8_2.NAND4F_5.Y.t10 mux8_2.NAND4F_9.Y.t6 VDD.t4295 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X751 a_n14751_2026.t5 a_n14931_1406.t3 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t8 VDD.t3377 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X752 VSS.t607 a_n21363_1380.t2 a_n21333_1406.t2 VSS.t606 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X753 mux8_8.NAND4F_3.Y.t3 mux8_8.A0.t12 VDD.t1496 VDD.t1495 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X754 S.t3 buffer_0.inv_1.A.t4 VDD.t1135 VDD.t1090 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X755 a_7644_n2838.t1 mux8_1.NAND4F_4.B.t8 a_7548_n2838.t1 VSS.t628 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X756 MULT_0.NAND2_4.Y.t0 B1.t9 a_n24162_n4727.t0 VSS.t831 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X757 VDD.t726 MULT_0.NAND2_8.Y.t7 MULT_0.inv_8.Y.t0 VDD.t725 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X758 VDD.t4376 SEL1.t29 mux8_0.NAND4F_5.Y.t8 VDD.t4375 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X759 a_n19981_n5154.t5 VSS.t1019 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t11 VSS.t1020 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X760 MULT_0.inv_7.A.t2 B2.t8 VDD.t2584 VDD.t2583 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X761 a_n17677_n22425.t4 B5.t5 VDD.t896 VDD.t895 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X762 a_n14077_3810.t6 a_n14257_3190.t2 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t0 VDD.t1531 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X763 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t2 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t10 VDD.t3999 VDD.t3998 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X764 mux8_4.NAND4F_0.Y.t0 mux8_4.NAND4F_2.D.t6 VDD.t122 VDD.t121 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X765 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t2 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t9 VDD.t446 VDD.t445 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X766 VDD.t3915 mux8_3.inv_0.A.t7 Y2.t3 VDD.t3914 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X767 VDD.t3538 B6.t12 a_n12314_n31661.t5 VDD.t3537 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X768 XOR8_0.S7.t5 a_n12347_n34023.t3 a_n12316_n34281.t5 VDD.t971 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X769 VDD.t328 mux8_6.NAND4F_0.C.t7 mux8_6.NAND4F_0.Y.t3 VDD.t327 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X770 a_n14005_n5180.t1 MULT_0.4bit_ADDER_0.A1.t6 VDD.t2307 VDD.t2306 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X771 VDD.t3362 mux8_4.NAND4F_4.B.t7 mux8_4.NAND4F_5.Y.t7 VDD.t3361 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X772 mux8_0.NAND4F_6.Y.t5 right_shifter_0.C.t5 VDD.t2514 VDD.t2513 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X773 a_n18998_n4534.t2 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t12 VDD.t2736 VDD.t2735 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X774 a_n10684_n7799.t3 a_n10714_n8445.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t7 VDD.t1347 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X775 a_n9125_n7799.t6 a_n9155_n8445.t2 MULT_0.S2.t2 VDD.t1190 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X776 a_n20557_n8419.t2 a_n20587_n8445.t3 VSS.t1420 VSS.t1419 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X777 OR8_0.NOT8_0.A1.t5 A1.t8 a_n17677_n16825.t9 VDD.t4198 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X778 VSS.t871 SEL3.t14 a_n10966_3190.t0 VSS.t870 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X779 a_11865_n2775.t8 mux8_1.NAND4F_8.Y.t10 VDD.t4317 VDD.t4316 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X780 VSS.t1172 B1.t10 a_n24012_n16501.t0 VSS.t1171 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X781 VDD.t4092 A3.t14 MULT_0.NAND2_0.Y.t4 VDD.t4091 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X782 VDD.t1292 MULT_0.4bit_ADDER_0.A0.t6 a_n10684_n4534.t3 VDD.t1291 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X783 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t0 a_n20737_n5154.t4 a_n20557_n5154.t0 VSS.t363 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X784 a_n10684_n8419.t5 a_n10864_n8419.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t0 VSS.t342 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X785 MULT_0.NAND2_4.Y.t5 A0.t7 VDD.t1664 VDD.t1663 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X786 a_7644_n26406.t1 mux8_7.NAND4F_4.B.t6 a_7548_n26406.t1 VSS.t93 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X787 a_n20659_3810.t11 a_n20113_3164.t3 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t8 VDD.t2687 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X788 mux8_1.NAND4F_4.Y.t6 SEL1.t30 VDD.t4378 VDD.t4377 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X789 VDD.t1158 MULT_0.NAND2_0.Y.t7 MULT_0.4bit_ADDER_0.B2.t0 VDD.t1157 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X790 VDD.t2214 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t0 VDD.t2213 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X791 VDD.t1696 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t8 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t4 VDD.t1695 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X792 VDD.t823 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t13 a_n19774_2026.t0 VDD.t822 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X793 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t7 a_664_373.t0 VSS.t939 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X794 VSS.t442 B5.t6 a_n23959_n21227.t0 VSS.t441 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X795 a_n1588_2026.t5 a_n1768_1406.t3 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t0 VDD.t2554 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X796 VDD.t1388 B7.t2 right_shifter_0.buffer_1.inv_1.A.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X797 VSS.t1644 B4.t12 left_shifter_0.buffer_4.inv_1.A.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X798 a_n10684_n4534.t7 MULT_0.4bit_ADDER_0.B0.t7 VDD.t288 VDD.t287 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X799 mux8_6.A1.t6 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t7 VDD.t966 VDD.t965 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X800 a_9528_n30934.t1 mux8_8.NAND4F_4.B.t4 a_9432_n30934.t0 VSS.t1467 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X801 VDD.t422 mux8_6.NAND4F_2.D.t6 mux8_6.NAND4F_4.Y.t0 VDD.t421 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X802 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t2 a_n8200_1380.t3 a_n8170_2026.t11 VDD.t334 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X803 mux8_1.NAND4F_7.Y.t5 NOT8_0.S0.t5 a_10459_n3765.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X804 XOR8_0.S5.t11 a_n12345_n28794.t2 a_n12314_n29052.t11 VDD.t3291 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X805 VDD.t3416 mux8_5.NAND4F_0.Y.t10 mux8_5.NAND4F_8.Y.t6 VDD.t3415 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X806 a_n20557_n11063.t5 a_n20737_n11683.t2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t3 VDD.t3453 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X807 VDD.t2026 mux8_6.NAND4F_1.Y.t9 mux8_6.NAND4F_9.Y.t5 VDD.t2025 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X808 VDD.t1684 left_shifter_0.C.t4 mux8_0.NAND4F_5.Y.t4 VDD.t1683 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X809 mux8_7.inv_0.A.t6 mux8_7.NAND4F_8.Y.t10 VSS.t1918 VSS.t1917 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X810 VSS.t873 SEL3.t15 a_547_1406.t2 VSS.t872 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X811 VDD.t436 AND8_0.S2.t4 mux8_3.NAND4F_4.Y.t0 VDD.t435 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X812 mux8_4.A0.t3 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t13 a_n9325_1406.t5 VSS.t2027 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X813 VDD.t2206 mux8_0.NAND4F_4.Y.t9 mux8_0.NAND4F_8.Y.t6 VDD.t2205 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X814 VDD.t2586 B2.t9 MULT_0.inv_12.A.t6 VDD.t2585 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X815 MULT_0.4bit_ADDER_2.B0.t3 a_n12596_n8419.t2 a_n12416_n8419.t2 VSS.t948 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X816 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t6 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t10 a_n15896_n12716.t1 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X817 a_n13975_n4534.t5 a_n14005_n5180.t3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t3 VDD.t1525 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X818 VDD.t4379 SEL1.t31 mux8_8.NAND4F_0.C.t2 VDD.t4357 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X819 VDD.t3540 B6.t13 a_n12345_n31403.t1 VDD.t3539 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X820 VDD.t3061 SEL0.t33 mux8_5.NAND4F_4.B.t3 VDD.t2937 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X821 VDD.t2150 B3.t10 left_shifter_0.buffer_5.inv_1.A.t2 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X822 VDD.t590 B0.t6 a_n17677_n15425.t8 VDD.t589 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X823 VSS.t706 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t17 a_n14931_1406.t0 VSS.t705 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X824 VDD.t3732 SEL2.t23 mux8_1.NAND4F_1.Y.t0 VDD.t3731 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X825 VDD.t1985 mux8_5.NAND4F_4.B.t4 mux8_5.NAND4F_5.Y.t5 VDD.t1984 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X826 mux8_8.A0.t6 a_n19954_1406.t3 a_n19774_1406.t5 VSS.t227 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X827 VSS.t180 A5.t8 a_n17466_1406.t5 VSS.t179 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X828 a_7452_n25478.t0 mux8_7.NAND4F_2.D.t5 VSS.t1457 VSS.t1456 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X829 XOR8_0.S2.t4 a_n12345_n20526.t4 a_n12314_n21072.t7 VDD.t2415 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X830 a_n12345_n20526.t1 A2.t7 VDD.t270 VDD.t269 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X831 mux8_4.NAND4F_0.Y.t4 mux8_4.A1.t12 a_10459_n16422.t0 VSS.t3 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X832 left_shifter_0.buffer_0.inv_1.A.t3 B2.t10 VDD.t2587 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X833 mux8_3.NAND4F_0.C.t2 SEL1.t32 VDD.t4380 VDD.t4373 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X834 mux8_0.NAND4F_4.Y.t5 VSS.t2040 VDD.t1969 VDD.t1968 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X835 a_n24048_1406.t5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t13 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t11 VSS.t1667 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X836 VSS.t120 A2.t8 a_n7594_1406.t5 VSS.t119 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X837 VDD.t448 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t10 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t3 VDD.t447 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X838 mux8_7.NAND4F_0.Y.t8 mux8_7.NAND4F_2.D.t6 VDD.t3130 VDD.t3129 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X839 a_2463_4914.t5 B7.t3 VSS.t684 VSS.t683 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X840 mux8_1.NAND4F_3.Y.t4 8bit_ADDER_0.S0.t12 VDD.t3356 VDD.t3355 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X841 a_10459_n20950.t1 SEL0.t34 a_10363_n20950.t1 VSS.t2000 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X842 VDD.t1520 mux8_2.inv_0.A.t7 Y1.t0 VDD.t1519 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X843 a_8496_n3766.t0 SEL1.t33 a_8400_n3766.t1 VSS.t1960 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X844 a_11194_n3766.t1 mux8_1.NAND4F_7.Y.t10 VSS.t652 VSS.t651 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X845 a_n12416_n7799.t9 a_n12446_n8445.t2 MULT_0.4bit_ADDER_2.B0.t9 VDD.t2433 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X846 a_n10090_373.t1 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t14 VSS.t2029 VSS.t860 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X847 mux8_3.NAND4F_4.B.t2 SEL0.t35 VDD.t3060 VDD.t3001 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X848 a_n29_2026.t5 a_n209_1406.t3 8bit_ADDER_0.S0.t5 VDD.t3119 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X849 VDD.t1500 mux8_0.NAND4F_7.Y.t10 mux8_0.NAND4F_9.Y.t7 VDD.t1499 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X850 a_n10423_n6187.t0 MULT_0.4bit_ADDER_0.B0.t8 VSS.t131 VSS.t130 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X851 VDD.t1688 mux8_6.inv_0.A.t7 Y7.t3 VDD.t1687 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X852 MULT_0.4bit_ADDER_1.B1.t11 a_n15737_n5180.t4 a_n15707_n4534.t11 VDD.t927 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X853 VDD.t244 MULT_0.4bit_ADDER_0.A2.t6 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t2 VDD.t243 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X854 VDD.t4153 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t10 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t4 VDD.t4152 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X855 mux8_8.NAND4F_4.Y.t1 AND8_0.S6.t5 VDD.t1235 VDD.t1234 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X856 a_n10714_n11709.t0 MULT_0.inv_8.Y.t6 VSS.t1617 VSS.t1616 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X857 XOR8_0.S0.t8 a_n12347_n15041.t3 a_n12316_n15299.t8 VDD.t3690 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X858 a_n18422_n11683.t3 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t10 VSS.t471 VSS.t470 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X859 VSS.t1335 MULT_0.4bit_ADDER_1.B3.t11 a_n20737_n8419.t0 VSS.t1334 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X860 mux8_3.NAND4F_3.Y.t3 mux8_3.NAND4F_2.D.t7 VDD.t2801 VDD.t2800 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X861 OR8_0.NOT8_0.A7.t4 A7.t9 a_n17677_n25225.t4 VDD.t2298 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X862 VDD.t3734 SEL2.t24 mux8_2.NAND4F_2.D.t3 VDD.t3733 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X863 a_7644_n35462.t1 mux8_6.NAND4F_4.B.t5 a_7548_n35462.t1 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X864 a_8592_n12822.t1 SEL0.t36 a_8496_n12822.t1 VSS.t1999 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X865 MULT_0.NAND2_5.Y.t3 A1.t9 a_n24162_n6019.t1 VSS.t1173 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X866 AND8_0.S5.t3 AND8_0.NOT8_0.A5.t7 VDD.t2636 VDD.t674 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X867 a_10363_n12821.t0 mux8_3.NAND4F_0.C.t6 a_10267_n12821.t1 VSS.t1321 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X868 VDD.t67 mux8_1.NAND4F_0.C.t6 mux8_1.NAND4F_0.Y.t3 VDD.t66 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X869 VDD.t4382 SEL1.t34 mux8_7.NAND4F_6.Y.t6 VDD.t4381 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X870 VDD.t1636 A4.t6 a_n14751_2026.t9 VDD.t1635 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X871 mux8_7.NAND4F_7.Y.t3 mux8_7.NAND4F_0.C.t7 VDD.t186 VDD.t185 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X872 V_FLAG_0.XOR2_2.B.t5 a_1707_4914.t2 a_1887_5534.t4 VDD.t1474 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X873 a_n23065_1406.t1 a_n23095_1380.t3 VSS.t801 VSS.t800 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X874 XOR8_0.S6.t4 a_n12345_n31403.t3 a_n12314_n31661.t11 VDD.t1828 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X875 VSS.t1561 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t15 a_n9305_n11683.t0 VSS.t1560 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X876 mux8_0.NAND4F_0.C.t0 SEL1.t35 VSS.t1962 VSS.t1961 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X877 VDD.t4200 A1.t10 a_n4879_2026.t10 VDD.t4199 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X878 a_n15707_n4534.t10 a_n15737_n5180.t5 MULT_0.4bit_ADDER_1.B1.t10 VDD.t928 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X879 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t11 VDD.t4155 VDD.t4154 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X880 8bit_ADDER_0.S1.t10 a_n3500_1406.t3 a_n3320_2026.t10 VDD.t1543 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X881 mux8_4.NAND4F_4.Y.t2 mux8_4.NAND4F_4.B.t8 VDD.t3364 VDD.t3363 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X882 mux8_3.NAND4F_5.Y.t3 SEL1.t36 VDD.t4384 VDD.t4383 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X883 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t2 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t13 VDD.t1604 VDD.t1603 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X884 VDD.t3059 SEL0.t37 mux8_8.NAND4F_4.B.t3 VDD.t2988 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X885 VDD.t3152 mux8_8.NAND4F_4.B.t5 mux8_8.NAND4F_5.Y.t7 VDD.t3151 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X886 VDD.t507 AND8_0.S7.t4 mux8_6.NAND4F_4.Y.t2 VDD.t506 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X887 VDD.t3542 B6.t14 a_n17677_n23825.t8 VDD.t3541 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X888 a_3493_4914.t5 a_3313_4914.t3 V_FLAG_0.XOR2_2.Y.t7 VSS.t541 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X889 VDD.t1212 mux8_5.NAND4F_4.Y.t9 mux8_5.NAND4F_8.Y.t0 VDD.t1211 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X890 a_n9125_n7799.t4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t13 VDD.t600 VDD.t599 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X891 a_8400_n11894.t0 mux8_3.NAND4F_2.D.t8 VSS.t1381 VSS.t1380 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X892 mux8_2.NAND4F_0.Y.t0 MULT_0.S1.t12 VDD.t2030 VDD.t2029 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X893 a_11865_n2775.t1 mux8_1.NAND4F_9.Y.t10 mux8_1.inv_0.A.t4 VDD.t1319 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X894 VDD.t2067 mux8_0.NAND4F_6.Y.t10 mux8_0.NAND4F_9.Y.t6 VDD.t2066 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X895 mux8_5.A0.t0 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t17 a_n12616_1406.t2 VSS.t138 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X896 VDD.t2773 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t8 a_n12416_n11063.t11 VDD.t2772 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X897 left_shifter_0.buffer_4.inv_1.A.t3 B4.t13 VDD.t3595 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X898 mux8_6.A0.t3 a_n23095_1380.t4 a_n23065_2026.t8 VDD.t1617 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X899 VDD.t2818 A6.t8 a_n21333_2026.t6 VDD.t2817 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X900 VSS.t1646 B4.t14 a_n23990_n20027.t1 VSS.t1645 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X901 VSS.t595 left_shifter_0.buffer_0.inv_1.A.t4 left_shifter_0.S3.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X902 VDD.t3736 SEL2.t25 mux8_2.NAND4F_7.Y.t0 VDD.t3735 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X903 a_n15707_n11063.t2 a_n15737_n11709.t2 mux8_7.A1.t11 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X904 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t7 MULT_0.4bit_ADDER_2.B0.t15 a_n10108_n11683.t2 VSS.t963 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X905 right_shifter_0.buffer_7.inv_1.A.t2 B1.t11 VDD.t2331 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X906 VSS.t404 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t10 a_n2744_1406.t5 VSS.t403 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X907 VSS.t286 B0.t7 left_shifter_0.buffer_6.inv_1.A.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X908 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t4 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t8 VDD.t3402 VDD.t3401 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X909 a_n24162_n4727.t1 A0.t8 VSS.t832 VSS.t831 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X910 a_n13399_n11683.t3 MULT_0.4bit_ADDER_2.B1.t12 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t3 VSS.t956 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X911 mux8_3.NAND4F_3.Y.t0 8bit_ADDER_0.S2.t12 a_9528_n11894.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X912 a_n3509_373.t0 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t15 VSS.t365 VSS.t364 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X913 mux8_1.NAND4F_5.Y.t6 SEL1.t37 VDD.t4386 VDD.t4385 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X914 a_7644_1690.t0 mux8_0.NAND4F_4.B.t7 a_7548_1690.t0 VSS.t426 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X915 VDD.t1823 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t8 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t1 VDD.t1822 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X916 VDD.t2502 MULT_0.4bit_ADDER_1.B0.t14 a_n10684_n7799.t6 VDD.t2501 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X917 VSS.t1318 a_n17296_n11709.t3 a_n17266_n11683.t4 VSS.t1317 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X918 a_9432_n26406.t0 mux8_7.NAND4F_0.C.t8 a_9336_n26406.t1 VSS.t88 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X919 VDD.t2820 A6.t9 AND8_0.NOT8_0.A6.t3 VDD.t2819 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X920 VDD.t3482 AND8_0.NOT8_0.A2.t8 AND8_0.S2.t2 VDD.t676 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X921 left_shifter_0.S2.t3 left_shifter_0.buffer_7.inv_1.A.t4 VDD.t3262 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X922 a_n13501_3190.t4 a_n13531_3164.t4 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t7 VSS.t1344 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X923 mux8_2.NAND4F_2.Y.t3 SEL0.t38 VDD.t3058 VDD.t3057 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X924 VDD.t2398 mux8_2.NAND4F_3.Y.t10 mux8_2.NAND4F_8.Y.t8 VDD.t2397 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X925 a_n15737_n8445.t1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t8 VDD.t3668 VDD.t3667 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X926 mux8_3.NAND4F_0.Y.t5 mux8_3.NAND4F_0.C.t7 VDD.t2670 VDD.t2669 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X927 VSS.t1387 A6.t10 a_n11274_n31085.t3 VSS.t1386 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X928 mux8_6.NAND4F_3.Y.t0 mux8_6.NAND4F_2.D.t7 VDD.t424 VDD.t423 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X929 Y2.t2 mux8_3.inv_0.A.t8 VDD.t3917 VDD.t3916 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X930 VDD.t610 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t14 a_n11460_2026.t8 VDD.t609 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X931 VDD.t580 AND8_0.S0.t5 mux8_1.NAND4F_4.Y.t1 VDD.t579 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X932 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t3 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t8 VDD.t1083 VDD.t1082 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X933 VDD.t1967 VSS.t2041 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t6 VDD.t1966 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X934 a_n12316_n34281.t4 a_n12347_n34023.t4 XOR8_0.S7.t4 VDD.t972 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X935 VDD.t4388 SEL1.t38 mux8_6.NAND4F_6.Y.t6 VDD.t4387 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X936 a_n3629_3190.t1 a_n4385_3190.t4 VSS.t1890 VSS.t1889 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X937 VSS.t114 MULT_0.4bit_ADDER_0.A2.t7 a_n16690_n5154.t0 VSS.t113 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X938 VDD.t3737 SEL2.t26 mux8_8.NAND4F_2.D.t2 VDD.t3724 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X939 a_n18042_2026.t4 a_n18222_1406.t3 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t3 VDD.t3898 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X940 VSS.t1757 a_n24654_1380.t3 a_n24624_1406.t2 VSS.t1756 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X941 a_n15707_n11063.t7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t12 VDD.t1276 VDD.t1275 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X942 a_n18998_n11683.t5 a_n19178_n11683.t3 mux8_8.A1.t11 VSS.t1255 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X943 MULT_0.4bit_ADDER_0.A3.t0 MULT_0.NAND2_11.Y.t8 VSS.t1301 VSS.t1300 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X944 mux8_3.NAND4F_3.Y.t2 8bit_ADDER_0.S2.t13 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X945 OR8_0.S2.t3 OR8_0.NOT8_0.A2.t7 VDD.t1545 VDD.t311 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X946 VDD.t3517 MULT_0.inv_8.Y.t7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t6 VDD.t3516 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X947 a_n17677_n16825.t8 A1.t11 OR8_0.NOT8_0.A1.t4 VDD.t4201 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X948 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t6 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t13 VDD.t4174 VDD.t4173 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X949 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t6 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t9 a_n15896_n9452.t1 VSS.t321 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X950 a_n11199_373.t1 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t15 VSS.t301 VSS.t300 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X951 mux8_1.NAND4F_0.Y.t8 SEL0.t39 VDD.t3056 VDD.t3055 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X952 mux8_7.NAND4F_4.Y.t7 mux8_7.NAND4F_4.B.t7 VDD.t198 VDD.t197 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X953 a_n12416_n7799.t1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t13 VDD.t3886 VDD.t3885 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X954 VDD.t837 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t11 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t4 VDD.t836 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X955 mux8_8.NAND4F_2.Y.t3 SEL1.t39 VDD.t4390 VDD.t4389 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X956 mux8_0.NAND4F_1.Y.t2 mux8_0.NAND4F_4.B.t8 VDD.t851 VDD.t850 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X957 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t8 a_n14155_n5154.t3 a_n13975_n4534.t8 VDD.t4162 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X958 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t3 MULT_0.4bit_ADDER_0.A3.t6 VDD.t637 VDD.t636 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X959 V_FLAG_0.XOR2_0.Y.t4 a_5017_4912.t2 a_5197_5532.t2 VDD.t2106 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X960 a_n17296_n11709.t1 MULT_0.inv_14.Y.t5 VDD.t2440 VDD.t2439 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X961 XOR8_0.S1.t8 a_n12345_n17857.t4 a_n12314_n18115.t9 VDD.t2457 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X962 mux8_1.NAND4F_1.Y.t6 XOR8_0.S0.t12 VDD.t3694 VDD.t3693 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X963 right_shifter_0.buffer_7.inv_1.A.t1 B1.t12 VDD.t2332 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X964 a_11290_n12822.t1 mux8_3.NAND4F_1.Y.t9 a_11194_n12822.t1 VSS.t596 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X965 VDD.t3054 SEL0.t40 mux8_0.NAND4F_4.B.t3 VDD.t2943 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X966 a_n914_3190.t2 SEL3.t16 VSS.t875 VSS.t874 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X967 a_8400_n34534.t0 mux8_6.NAND4F_2.D.t8 VSS.t203 VSS.t202 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X968 mux8_7.NAND4F_9.Y.t8 mux8_7.NAND4F_1.Y.t10 VDD.t2867 VDD.t2866 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X969 a_n24624_2026.t8 a_n24654_1380.t4 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t8 VDD.t3880 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X970 right_shifter_0.buffer_1.inv_1.A.t2 B7.t4 VDD.t1389 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X971 VDD.t898 B5.t7 a_n12345_n28794.t1 VDD.t897 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X972 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t5 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t9 VDD.t3404 VDD.t3403 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X973 VDD.t246 MULT_0.4bit_ADDER_0.A2.t8 a_n17266_n4534.t2 VDD.t245 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X974 VDD.t3154 mux8_8.NAND4F_4.B.t6 mux8_8.NAND4F_3.Y.t2 VDD.t3153 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X975 VDD.t1136 buffer_0.inv_1.A.t5 S.t2 VDD.t1092 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X976 mux8_0.NAND4F_3.Y.t2 mux8_0.NAND4F_0.C.t6 VDD.t643 VDD.t642 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X977 a_n23950_3810.t9 a_n23404_3164.t3 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t7 VDD.t2411 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X978 a_n218_373.t1 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t16 VSS.t1141 VSS.t880 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X979 VDD.t3331 mux8_1.NAND4F_0.Y.t9 mux8_1.NAND4F_8.Y.t6 VDD.t3330 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X980 XOR8_0.S2.t8 a_n12345_n20814.t2 a_n12314_n21072.t11 VDD.t2871 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X981 VDD.t1825 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t9 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t2 VDD.t1824 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X982 a_n6611_2026.t5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t13 VDD.t2436 VDD.t2435 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X983 a_n4879_2026.t1 a_n5059_1406.t4 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t2 VDD.t798 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X984 VDD.t1965 VSS.t2042 mux8_0.NAND4F_7.Y.t6 VDD.t1964 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X985 VSS.t21 a_5167_4886.t3 a_5197_4912.t5 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X986 a_n15707_n4534.t2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t16 VDD.t452 VDD.t451 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X987 a_9432_n7266.t0 mux8_2.NAND4F_0.C.t4 a_9336_n7266.t1 VSS.t1486 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X988 mux8_6.NAND4F_3.Y.t6 mux8_6.A0.t13 a_9528_n34534.t1 VSS.t1499 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X989 mux8_4.NAND4F_7.Y.t2 NOT8_0.S3.t5 a_10459_n17349.t0 VSS.t3 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X990 a_9432_n35462.t0 mux8_6.NAND4F_0.C.t8 a_9336_n35462.t1 VSS.t152 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X991 VSS.t491 V_FLAG_0.XOR2_2.B.t14 a_4069_4914.t5 VSS.t490 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X992 a_n10240_3164.t0 B3.t11 VSS.t1106 VSS.t1105 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X993 VDD.t1963 VSS.t2043 a_n9125_n4534.t7 VDD.t1962 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X994 a_n13714_n9452.t1 MULT_0.4bit_ADDER_1.B1.t13 VSS.t1611 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X995 mux8_6.NAND4F_0.Y.t2 mux8_6.NAND4F_0.C.t9 VDD.t330 VDD.t329 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X996 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t0 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t9 a_n10090_373.t0 VSS.t860 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X997 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t4 MULT_0.4bit_ADDER_2.B1.t13 VDD.t1893 VDD.t1892 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X998 a_n16483_1406.t5 a_n16513_1380.t3 VSS.t731 VSS.t730 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X999 a_n14175_1406.t5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t18 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t11 VSS.t704 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1000 a_n18998_n4534.t8 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t9 VDD.t2556 VDD.t2555 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1001 Y7.t2 mux8_6.inv_0.A.t8 VDD.t1690 VDD.t1689 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1002 mux8_4.NAND4F_5.Y.t8 mux8_4.NAND4F_4.B.t9 VDD.t3366 VDD.t3365 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1003 left_shifter_0.S3.t3 left_shifter_0.buffer_0.inv_1.A.t5 VDD.t1184 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1004 MULT_0.4bit_ADDER_1.A2.t0 MULT_0.inv_12.A.t7 VSS.t408 VSS.t407 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1005 Z.t0 ZFLAG_0.NAND2_0.Y.t8 VSS.t725 VSS.t724 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1006 VDD.t3247 mux8_4.NAND4F_0.C.t5 mux8_4.NAND4F_3.Y.t3 VDD.t3246 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1007 VDD.t3739 SEL2.t27 mux8_3.NAND4F_1.Y.t1 VDD.t3738 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1008 VDD.t2274 V_FLAG_0.XOR2_2.Y.t14 V_FLAG_0.NAND2_0.Y.t2 VDD.t2273 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1009 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t4 a_n21513_1406.t3 a_n21333_1406.t5 VSS.t597 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1010 a_n4303_1406.t2 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t15 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t10 VSS.t1858 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1011 a_n17677_n25225.t3 A7.t10 OR8_0.NOT8_0.A7.t3 VDD.t2299 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1012 mux8_3.NAND4F_7.Y.t2 NOT8_0.S2.t4 VDD.t1724 VDD.t1723 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1013 a_n3320_1406.t1 a_n3350_1380.t3 VSS.t1149 VSS.t1148 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1014 mux8_6.NAND4F_3.Y.t8 mux8_6.A0.t14 VDD.t3299 VDD.t3298 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1015 a_n4618_373.t0 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t16 VSS.t1860 VSS.t1859 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1016 VDD.t735 mux8_8.NAND4F_8.Y.t9 a_11865_n29943.t5 VDD.t734 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1017 mux8_7.NAND4F_9.Y.t1 mux8_7.NAND4F_7.Y.t9 VDD.t48 VDD.t47 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1018 a_7548_n26406.t0 SEL1.t40 a_7452_n26406.t1 VSS.t1963 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1019 right_shifter_0.buffer_1.inv_1.A.t1 B7.t5 VDD.t1390 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1020 a_3493_5534.t10 a_3463_4888.t4 V_FLAG_0.XOR2_2.Y.t4 VDD.t488 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1021 VDD.t2152 B3.t12 a_n12314_n23651.t8 VDD.t2151 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1022 VDD.t2301 A7.t11 AND8_0.NOT8_0.A7.t2 VDD.t2300 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1023 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t4 a_n20737_n11683.t3 a_n20557_n11063.t4 VDD.t3454 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1024 a_n12314_n31661.t10 a_n12345_n31403.t4 XOR8_0.S6.t5 VDD.t1829 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1025 a_n19028_n11709.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t11 VSS.t473 VSS.t472 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1026 mux8_6.NAND4F_9.Y.t6 mux8_6.NAND4F_1.Y.t10 VDD.t2028 VDD.t2027 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1027 VDD.t3406 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t10 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t6 VDD.t3405 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1028 a_8400_n7266.t0 mux8_2.NAND4F_2.D.t5 VSS.t1473 VSS.t1472 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1029 MULT_0.4bit_ADDER_0.A2.t0 MULT_0.NAND2_10.Y.t7 VSS.t210 VSS.t209 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1030 mux8_3.NAND4F_4.Y.t1 AND8_0.S2.t5 VDD.t438 VDD.t437 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1031 a_n20659_3190.t2 SEL3.t17 VSS.t877 VSS.t876 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X1032 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t3 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t10 VDD.t1827 VDD.t1826 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1033 mux8_5.NAND4F_5.Y.t6 mux8_5.NAND4F_4.B.t5 VDD.t1987 VDD.t1986 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1034 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t0 a_n1094_3190.t2 a_n914_3810.t3 VDD.t918 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1035 a_n11460_2026.t2 a_n11490_1380.t3 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t3 VDD.t953 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1036 a_10459_n16422.t1 SEL0.t41 a_10363_n16422.t1 VSS.t2001 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1037 mux8_1.NAND4F_2.D.t0 SEL2.t28 VSS.t1711 VSS.t1710 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1038 VDD.t214 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t11 a_n12416_n4534.t1 VDD.t213 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1039 VSS.t1570 A7.t12 a_n11276_n33705.t2 VSS.t1569 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1040 mux8_1.NAND4F_4.B.t3 SEL0.t42 VDD.t3053 VDD.t2933 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1041 VDD.t2383 left_shifter_0.S0.t5 mux8_1.NAND4F_5.Y.t3 VDD.t2382 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1042 a_8592_n20950.t1 SEL0.t43 a_8496_n20950.t1 VSS.t2003 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1043 VDD.t454 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t17 a_n15887_n5154.t1 VDD.t453 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X1044 a_9528_n7266.t1 mux8_2.NAND4F_4.B.t4 a_9432_n7266.t1 VSS.t1488 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1045 ZFLAG_0.nor4_1.Y.t6 Y6.t4 VSS.t1469 VSS.t1468 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1046 a_n17266_n5154.t1 a_n17446_n5154.t3 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t4 VSS.t1223 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1047 VSS.t862 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t10 a_n9325_1406.t1 VSS.t861 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1048 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t3 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t11 a_n3509_373.t1 VSS.t364 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1049 VDD.t737 mux8_8.NAND4F_8.Y.t10 a_11865_n29943.t6 VDD.t736 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1050 VDD.t188 mux8_7.NAND4F_0.C.t9 mux8_7.NAND4F_3.Y.t0 VDD.t187 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1051 VDD.t2154 B3.t13 a_n12345_n23393.t1 VDD.t2153 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X1052 a_n23990_n20027.t0 A4.t7 AND8_0.NOT8_0.A4.t4 VSS.t805 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1053 left_shifter_0.S5.t0 left_shifter_0.buffer_4.inv_1.A.t4 VDD.t1197 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1054 a_n13531_3164.t0 B4.t15 VSS.t1648 VSS.t1647 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1055 a_n1618_1380.t0 A0.t9 VSS.t834 VSS.t833 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1056 Y5.t0 mux8_7.inv_0.A.t7 VSS.t1271 VSS.t1270 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1057 AND8_0.NOT8_0.A6.t6 B6.t15 VDD.t3544 VDD.t3543 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1058 a_1857_4888.t1 B7.t6 VDD.t1392 VDD.t1391 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1059 a_7644_n7266.t1 mux8_2.NAND4F_4.B.t5 a_7548_n7266.t1 VSS.t1489 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1060 VSS.t1945 MULT_0.4bit_ADDER_1.A3.t8 a_n19981_n8419.t5 VSS.t1944 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1061 mux8_2.NAND4F_6.Y.t8 SEL0.t44 VDD.t3052 VDD.t3051 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1062 VDD.t659 mux8_2.NAND4F_1.Y.t10 mux8_2.NAND4F_9.Y.t3 VDD.t658 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1063 mux8_4.NAND4F_9.Y.t0 mux8_4.NAND4F_5.Y.t9 a_11386_n17350.t0 VSS.t1377 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1064 a_7548_n35462.t0 SEL1.t41 a_7452_n35462.t1 VSS.t1964 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1065 VSS.t182 A5.t9 a_n11274_n28476.t5 VSS.t181 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1066 a_8496_n12822.t0 SEL1.t42 a_8400_n12822.t1 VSS.t1965 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1067 mux8_6.NAND4F_9.Y.t8 mux8_6.NAND4F_7.Y.t9 VDD.t2065 VDD.t2064 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1068 VDD.t2637 AND8_0.NOT8_0.A5.t8 AND8_0.S5.t2 VDD.t676 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1069 VDD.t719 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t7 MULT_0.4bit_ADDER_1.B3.t0 VDD.t718 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1070 a_7452_n30006.t0 mux8_8.NAND4F_2.D.t7 VSS.t739 VSS.t738 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1071 Y6.t0 mux8_8.inv_0.A.t10 VSS.t1331 VSS.t1330 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1072 a_10267_n12821.t0 SEL2.t29 VSS.t1712 VSS.t1378 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1073 VSS.t37 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t8 a_n6035_1406.t1 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1074 mux8_8.NAND4F_7.Y.t8 NOT8_0.S6.t5 a_10459_n30933.t1 VSS.t1157 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1075 a_n17677_n16825.t4 B1.t13 VDD.t2334 VDD.t2333 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1076 VDD.t701 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t10 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t6 VDD.t700 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1077 VSS.t122 A2.t9 OR8_0.NOT8_0.A2.t5 VSS.t121 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X1078 VDD.t1326 mux8_1.NAND4F_7.Y.t11 mux8_1.NAND4F_9.Y.t7 VDD.t1325 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1079 a_n11274_n20496.t2 A2.t10 VSS.t245 VSS.t244 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1080 VDD.t3741 SEL2.t30 mux8_3.NAND4F_5.Y.t1 VDD.t3740 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1081 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t10 B3.t14 a_n10786_3190.t4 VSS.t1107 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1082 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t0 A3.t15 a_n11199_373.t0 VSS.t300 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1083 MULT_0.4bit_ADDER_2.B1.t8 a_n15887_n8419.t2 a_n15707_n7799.t5 VDD.t2396 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1084 a_11865_n16359.t9 mux8_4.NAND4F_9.Y.t9 mux8_4.inv_0.A.t5 VDD.t960 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1085 VDD.t4392 SEL1.t43 mux8_4.NAND4F_4.Y.t5 VDD.t4391 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1086 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t3 MULT_0.4bit_ADDER_0.A2.t9 a_n17005_n6187.t0 VSS.t115 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1087 a_n16792_3190.t1 a_n16822_3164.t4 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t1 VSS.t1410 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1088 mux8_8.NAND4F_5.Y.t8 mux8_8.NAND4F_4.B.t7 VDD.t3156 VDD.t3155 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1089 a_n17266_n4534.t9 a_n17296_n5180.t2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t0 VDD.t1853 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1090 mux8_6.NAND4F_4.Y.t3 AND8_0.S7.t5 VDD.t509 VDD.t508 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1091 a_n12446_n5180.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t12 VSS.t95 VSS.t94 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1092 a_n9125_n7799.t10 VSS.t2044 VDD.t1961 VDD.t1960 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1093 mux8_5.NAND4F_8.Y.t1 mux8_5.NAND4F_4.Y.t10 VDD.t1214 VDD.t1213 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1094 VDD.t1430 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t19 a_n14751_2026.t7 VDD.t1429 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1095 a_n6920_3190.t1 a_n7676_3190.t4 VSS.t1793 VSS.t1792 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1096 mux8_1.NAND4F_8.Y.t0 mux8_1.NAND4F_4.Y.t10 VDD.t769 VDD.t768 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1097 a_n8549_n8419.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t14 MULT_0.S2.t11 VSS.t289 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1098 a_n59_1380.t0 SEL3.t18 VSS.t879 VSS.t878 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1099 a_n12416_n11063.t10 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t9 VDD.t2775 VDD.t2774 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1100 VDD.t2210 NOT8_0.S1.t4 mux8_2.NAND4F_7.Y.t2 VDD.t2209 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1101 XOR8_0.S3.t3 a_n12345_n23393.t3 a_n12314_n23651.t2 VDD.t3452 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1102 VDD.t3418 A7.t13 a_1887_5534.t2 VDD.t3417 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1103 VDD.t2742 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t3 VDD.t2741 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1104 a_n11276_n14723.t5 B0.t8 XOR8_0.S0.t0 VSS.t287 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1105 mux8_2.NAND4F_7.Y.t3 NOT8_0.S1.t5 a_10459_n8193.t0 VSS.t1051 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1106 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t2 MULT_0.4bit_ADDER_1.B0.t15 VDD.t2504 VDD.t2503 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1107 VDD.t3249 mux8_4.NAND4F_0.C.t6 mux8_4.NAND4F_1.Y.t3 VDD.t3248 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1108 a_n9125_n4534.t4 a_n9305_n5154.t4 MULT_0.S1.t10 VDD.t368 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1109 MULT_0.inv_13.A.t4 A3.t16 VDD.t4094 VDD.t4093 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1110 VDD.t1570 AND8_0.NOT8_0.A6.t7 AND8_0.S6.t0 VDD.t1569 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1111 a_9528_n11894.t1 mux8_3.NAND4F_4.B.t4 a_9432_n11894.t0 VSS.t1268 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1112 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t0 SEL3.t19 a_n218_373.t0 VSS.t880 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1113 a_n12314_n21072.t5 B2.t11 VDD.t2589 VDD.t2588 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1114 MULT_0.4bit_ADDER_1.B2.t4 a_n19178_n5154.t4 a_n18998_n4534.t5 VDD.t691 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1115 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t9 a_n17296_n11709.t4 a_n17266_n11063.t8 VDD.t2649 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1116 VSS.t1527 MULT_0.inv_15.Y.t6 a_n19981_n11683.t5 VSS.t1526 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1117 XOR8_0.S5.t4 a_n12345_n28794.t3 a_n11274_n29052.t1 VSS.t600 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1118 VDD.t1394 B7.t7 NOT8_0.S7.t2 VDD.t1393 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1119 a_n23374_3190.t2 a_n24130_3190.t4 VSS.t1697 VSS.t1696 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1120 VDD.t2890 mux8_0.NAND4F_2.D.t6 mux8_0.NAND4F_0.Y.t5 VDD.t2889 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1121 mux8_3.NAND4F_2.Y.t6 SEL1.t44 VDD.t4394 VDD.t4393 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1122 a_9336_n26406.t0 SEL2.t31 VSS.t1713 VSS.t1462 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1123 VDD.t3263 left_shifter_0.buffer_7.inv_1.A.t5 left_shifter_0.S2.t2 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1124 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t5 a_n21513_1406.t4 a_n21333_2026.t7 VDD.t1195 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1125 VSS.t807 A4.t8 a_n11274_n25843.t3 VSS.t806 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1126 VDD.t877 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t13 a_n8350_1406.t1 VDD.t876 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X1127 VDD.t2336 B1.t14 MULT_0.NAND2_4.Y.t3 VDD.t2335 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1128 a_11290_n20950.t0 mux8_5.NAND4F_3.Y.t11 a_11194_n20950.t0 VSS.t1329 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1129 VDD.t318 OR8_0.NOT8_0.A6.t7 OR8_0.S6.t3 VDD.t317 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1130 a_n12416_n11063.t8 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t15 VDD.t2009 VDD.t2008 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1131 a_n15131_n11683.t2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t13 mux8_7.A1.t8 VSS.t629 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1132 a_n1588_2026.t7 a_n1618_1380.t4 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t7 VDD.t1253 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1133 VDD.t1666 A0.t10 MULT_0.NAND2_3.Y.t3 VDD.t1665 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1134 mux8_2.NAND4F_2.D.t0 SEL2.t32 VSS.t1715 VSS.t1714 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1135 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t5 a_n20839_3190.t3 a_n20659_3810.t8 VDD.t4276 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1136 VDD.t2083 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t12 a_n1588_2026.t9 VDD.t2082 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1137 mux8_8.A1.t0 a_n19178_n11683.t4 a_n18998_n11683.t4 VSS.t769 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1138 a_n4909_1380.t0 A1.t12 VSS.t1896 VSS.t1895 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1139 VDD.t2522 mux8_3.NAND4F_4.B.t5 mux8_3.NAND4F_3.Y.t6 VDD.t2521 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1140 VDD.t1546 OR8_0.NOT8_0.A2.t8 OR8_0.S2.t2 VDD.t313 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1141 MULT_0.NAND2_10.Y.t2 A2.t11 VDD.t515 VDD.t514 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1142 VDD.t1668 A0.t11 MULT_0.inv_6.A.t6 VDD.t1667 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1143 a_5167_4886.t0 mux8_6.A0.t15 VDD.t3301 VDD.t3300 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1144 a_n8170_2026.t7 a_n8350_1406.t4 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t8 VDD.t1517 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1145 a_8496_n8194.t0 SEL1.t45 a_8400_n8194.t1 VSS.t1966 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1146 a_11194_n8194.t0 mux8_2.NAND4F_7.Y.t10 VSS.t668 VSS.t667 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1147 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t6 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t15 VDD.t1563 VDD.t1562 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1148 VDD.t4396 SEL1.t46 mux8_7.NAND4F_4.Y.t6 VDD.t4395 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1149 VDD.t806 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t12 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t4 VDD.t805 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1150 a_n12416_n7799.t7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t10 VDD.t4284 VDD.t4283 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1151 VDD.t3626 mux8_5.NAND4F_0.C.t6 mux8_5.NAND4F_1.Y.t3 VDD.t3625 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1152 a_n20296_n12716.t0 MULT_0.4bit_ADDER_2.B3.t9 VSS.t1824 VSS.t1534 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1153 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t3 A1.t13 a_n4618_373.t1 VSS.t1859 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1154 a_n9901_1406.t1 a_n10081_1406.t4 mux8_4.A0.t5 VSS.t2024 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1155 a_n11840_n8419.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t14 MULT_0.4bit_ADDER_2.B0.t2 VSS.t1760 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1156 VDD.t1508 mux8_8.NAND4F_2.D.t8 mux8_8.NAND4F_2.Y.t1 VDD.t1507 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1157 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t7 a_n11640_1406.t3 a_n11460_1406.t3 VSS.t773 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1158 VSS.t1836 A3.t17 a_n11274_n23075.t2 VSS.t1835 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1159 AND8_0.NOT8_0.A7.t1 A7.t14 VDD.t3420 VDD.t3419 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1160 a_11194_n12822.t0 mux8_3.NAND4F_7.Y.t10 VSS.t1542 VSS.t722 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1161 a_n19774_1406.t2 a_n19804_1380.t2 VSS.t716 VSS.t715 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1162 VDD.t3682 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t8 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t3 VDD.t3681 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1163 a_n10786_3810.t4 a_n10240_3164.t4 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t2 VDD.t684 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1164 a_n21363_1380.t0 A6.t11 VSS.t1389 VSS.t1388 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1165 VDD.t1959 VSS.t2045 a_n9125_n11063.t11 VDD.t1958 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1166 mux8_8.NAND4F_9.Y.t0 mux8_8.NAND4F_5.Y.t9 a_11386_n30934.t0 VSS.t727 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1167 VDD.t50 mux8_7.NAND4F_7.Y.t10 mux8_7.NAND4F_9.Y.t0 VDD.t49 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1168 VDD.t3398 left_shifter_0.S2.t4 mux8_3.NAND4F_5.Y.t6 VDD.t3397 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1169 VSS.t1447 MULT_0.4bit_ADDER_0.B2.t6 a_n17446_n5154.t0 VSS.t1446 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1170 a_n9314_n9452.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t15 VSS.t291 VSS.t290 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1171 OR8_0.NOT8_0.A3.t4 A3.t18 a_n17677_n19625.t3 VDD.t4095 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X1172 a_n7594_1406.t2 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t14 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t6 VSS.t431 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1173 a_n20587_n5180.t1 MULT_0.4bit_ADDER_0.A3.t7 VDD.t639 VDD.t638 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1174 AND8_0.S4.t3 AND8_0.NOT8_0.A4.t8 VDD.t675 VDD.t674 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1175 a_n6611_1406.t2 a_n6641_1380.t4 VSS.t437 VSS.t436 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1176 mux8_8.NAND4F_3.Y.t1 mux8_8.NAND4F_4.B.t8 VDD.t3158 VDD.t3157 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1177 mux8_1.NAND4F_3.Y.t2 8bit_ADDER_0.S0.t13 a_9528_n2838.t0 VSS.t1543 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1178 VDD.t3921 mux8_3.NAND4F_8.Y.t10 a_11865_n11831.t4 VDD.t3920 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1179 VSS.t594 right_shifter_0.buffer_1.inv_1.A.t4 right_shifter_0.S6.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1180 mux8_4.NAND4F_6.Y.t2 right_shifter_0.S3.t4 a_8592_n17350.t0 VSS.t196 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1181 8bit_ADDER_0.S0.t6 a_n59_1380.t2 a_n29_2026.t6 VDD.t1441 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1182 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t1 MULT_0.4bit_ADDER_1.A1.t5 VDD.t106 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1183 a_9528_n34534.t0 mux8_6.NAND4F_4.B.t6 a_9432_n34534.t1 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1184 a_10459_n17349.t1 SEL0.t45 a_10363_n17349.t1 VSS.t2001 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1185 VDD.t1730 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t11 a_n9901_2026.t5 VDD.t1729 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1186 a_9336_n35462.t0 SEL2.t33 VSS.t1716 VSS.t204 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1187 VDD.t3050 SEL0.t46 mux8_1.NAND4F_4.B.t2 VDD.t2933 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1188 a_n10684_n11683.t5 a_n10714_n11709.t3 VSS.t1036 VSS.t1035 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1189 left_shifter_0.buffer_1.inv_1.A.t3 B7.t8 VDD.t1395 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1190 mux8_6.NAND4F_2.Y.t6 SEL1.t47 VDD.t4398 VDD.t4397 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1191 mux8_8.A0.t1 a_n19804_1380.t3 a_n19774_2026.t4 VDD.t1448 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1192 VDD.t388 A5.t10 a_n18042_2026.t1 VDD.t387 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X1193 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t5 a_n20737_n5154.t5 a_n20557_n4534.t3 VDD.t744 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1194 a_n23950_3190.t2 SEL3.t20 VSS.t882 VSS.t881 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X1195 VSS.t824 a_n14005_n11709.t2 a_n13975_n11683.t3 VSS.t823 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1196 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t11 B2.t12 a_n7496_3190.t5 VSS.t1286 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1197 mux8_1.NAND4F_4.Y.t0 AND8_0.S0.t6 a_7644_n2838.t0 VSS.t275 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1198 OR8_0.NOT8_0.A2.t4 A2.t12 a_n17677_n18225.t4 VDD.t516 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1199 VDD.t1895 MULT_0.4bit_ADDER_2.B1.t14 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t5 VDD.t1894 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1200 a_n24624_2026.t5 A7.t15 VDD.t3422 VDD.t3421 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1201 VDD.t1561 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t16 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t5 VDD.t1560 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1202 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t2 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t13 VDD.t2085 VDD.t2084 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1203 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t10 VSS.t1017 a_n19981_n5154.t4 VSS.t1018 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1204 VDD.t4400 SEL1.t48 mux8_4.NAND4F_5.Y.t6 VDD.t4399 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1205 VDD.t592 B0.t9 a_n12316_n15299.t11 VDD.t591 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1206 a_8400_762.t0 SEL2.t34 VSS.t1717 VSS.t1435 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1207 mux8_3.NAND4F_1.Y.t0 SEL2.t35 VDD.t3743 VDD.t3742 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1208 a_1887_5534.t9 a_1857_4888.t3 V_FLAG_0.XOR2_2.B.t8 VDD.t2769 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1209 VDD.t1758 SEL3.t21 a_n10966_3190.t1 VDD.t1757 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X1210 mux8_4.NAND4F_3.Y.t2 mux8_4.NAND4F_0.C.t7 VDD.t3251 VDD.t3250 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1211 MULT_0.4bit_ADDER_1.A0.t0 MULT_0.inv_6.A.t7 VSS.t536 VSS.t535 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1212 VDD.t3049 SEL0.t47 mux8_3.NAND4F_7.Y.t8 VDD.t3048 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1213 a_10267_n2838.t1 mux8_1.NAND4F_2.D.t10 VSS.t854 VSS.t853 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1214 VDD.t2656 mux8_8.NAND4F_0.C.t6 mux8_8.NAND4F_1.Y.t8 VDD.t2655 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1215 VSS.t1898 A1.t14 a_n11274_n17539.t5 VSS.t1897 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1216 mux8_1.NAND4F_9.Y.t2 mux8_1.NAND4F_5.Y.t9 VDD.t1598 VDD.t1597 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1217 VDD.t7 mux8_6.NAND4F_4.B.t7 mux8_6.NAND4F_3.Y.t5 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1218 a_16431_n19505.t5 Y6.t5 a_16143_n19505.t5 VDD.t3167 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X1219 AND8_0.S1.t3 AND8_0.NOT8_0.A1.t8 VDD.t825 VDD.t824 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1220 a_n24162_n6019.t0 B1.t15 VSS.t1174 VSS.t1173 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1221 a_11865_n29943.t7 mux8_8.NAND4F_8.Y.t11 VDD.t739 VDD.t738 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1222 VDD.t2186 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t7 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t3 VDD.t2185 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1223 a_n2627_373.t1 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t8 VSS.t673 VSS.t672 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1224 a_n12314_n26419.t8 a_n12345_n26161.t3 XOR8_0.S4.t8 VDD.t4165 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1225 a_n12605_n9452.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t15 VSS.t1762 VSS.t1761 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1226 VDD.t2011 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t16 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t2 VDD.t2010 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1227 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t1 a_n10864_n8419.t3 a_n10684_n7799.t0 VDD.t699 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1228 MULT_0.S2.t3 a_n9305_n8419.t2 a_n9125_n7799.t0 VDD.t1041 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1229 VSS.t1422 a_n20587_n8445.t4 a_n20557_n8419.t1 VSS.t1421 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1230 VDD.t414 mux8_6.NAND4F_7.Y.t10 mux8_6.NAND4F_9.Y.t7 VDD.t413 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1231 MULT_0.NAND2_0.Y.t2 B0.t10 VDD.t594 VDD.t593 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1232 VDD.t4319 mux8_1.NAND4F_8.Y.t11 a_11865_n2775.t7 VDD.t4318 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1233 a_n10108_n11683.t1 MULT_0.4bit_ADDER_2.B0.t16 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t8 VSS.t964 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1234 VDD.t2338 B1.t16 a_n17677_n16825.t3 VDD.t2337 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1235 a_n10684_n4534.t1 a_n10714_n5180.t3 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t4 VDD.t306 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1236 a_n20557_n5154.t5 a_n20587_n5180.t2 VSS.t1057 VSS.t1056 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1237 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t8 a_n10864_n8419.t4 a_n10684_n8419.t4 VSS.t844 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1238 MULT_0.S2.t4 a_n9305_n8419.t3 a_n9125_n8419.t5 VSS.t517 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1239 VSS.t247 A2.t13 a_n11274_n20496.t1 VSS.t246 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1240 a_1887_4914.t4 a_1707_4914.t3 V_FLAG_0.XOR2_2.B.t6 VSS.t945 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1241 a_n14175_1406.t2 A4.t9 VSS.t809 VSS.t808 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1242 VDD.t3923 mux8_3.NAND4F_8.Y.t11 a_11865_n11831.t3 VDD.t3922 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1243 a_n13192_1406.t1 a_n13372_1406.t4 mux8_5.A0.t4 VSS.t580 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1244 a_n17005_n6187.t1 MULT_0.4bit_ADDER_0.B2.t7 VSS.t1448 VSS.t115 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1245 VDD.t3144 OR8_0.S6.t4 mux8_8.NAND4F_2.Y.t6 VDD.t3143 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1246 VDD.t163 MULT_0.NAND2_3.Y.t8 MULT_0.SO.t3 VDD.t162 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1247 a_n10684_n5154.t5 a_n10864_n5154.t3 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t1 VSS.t548 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1248 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t8 VDD.t2216 VDD.t2215 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1249 a_n23065_2026.t11 a_n23245_1406.t3 mux8_6.A0.t8 VDD.t2487 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1250 VDD.t4097 A3.t19 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t3 VDD.t4096 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1251 VDD.t4402 SEL1.t49 mux8_5.NAND4F_5.Y.t8 VDD.t4401 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1252 a_8592_n16422.t1 SEL0.t48 a_8496_n16422.t1 VSS.t2002 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1253 a_n2744_1406.t2 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t16 8bit_ADDER_0.S1.t0 VSS.t366 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1254 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t6 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t16 VDD.t612 VDD.t611 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1255 VDD.t2038 mux8_7.NAND4F_5.Y.t10 mux8_7.NAND4F_9.Y.t6 VDD.t2037 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1256 VDD.t596 B0.t11 a_n12347_n15041.t0 VDD.t595 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X1257 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t3 MULT_0.4bit_ADDER_1.A0.t5 a_n10423_n9452.t1 VSS.t1263 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1258 MULT_0.inv_8.Y.t1 MULT_0.NAND2_8.Y.t8 VSS.t354 VSS.t353 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1259 VDD.t3424 A7.t16 a_5017_4912.t1 VDD.t3423 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X1260 a_8496_n20950.t0 SEL1.t50 a_8400_n20950.t1 VSS.t1967 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1261 a_n12416_n7799.t3 a_n12596_n8419.t3 MULT_0.4bit_ADDER_2.B0.t4 VDD.t1837 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1262 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t4 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t17 VDD.t1559 VDD.t1558 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1263 VDD.t3047 SEL0.t49 mux8_0.NAND4F_6.Y.t8 VDD.t3046 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1264 a_3493_5534.t2 SEL3.t22 VDD.t1760 VDD.t1759 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1265 MULT_0.inv_12.A.t5 B2.t13 VDD.t2591 VDD.t2590 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1266 XOR8_0.S0.t1 B0.t12 a_n11276_n14723.t4 VSS.t288 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1267 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t4 a_n14005_n5180.t4 a_n13975_n4534.t4 VDD.t1526 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1268 a_n12416_n8419.t5 a_n12446_n8445.t3 VSS.t1232 VSS.t1231 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1269 VDD.t108 MULT_0.4bit_ADDER_1.A1.t6 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t2 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1270 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t10 B4.t16 a_n14077_3190.t4 VSS.t1649 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1271 mux8_2.NAND4F_3.Y.t1 mux8_2.NAND4F_0.C.t5 VDD.t3201 VDD.t3200 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1272 VSS.t757 Y5.t5 ZFLAG_0.nor4_1.Y.t4 VSS.t756 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1273 a_n338_3190.t0 a_n1094_3190.t3 VSS.t456 VSS.t455 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1274 a_8592_762.t1 SEL0.t50 a_8496_762.t1 VSS.t2007 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1275 MULT_0.4bit_ADDER_1.B0.t8 a_n12596_n5154.t4 a_n12416_n5154.t2 VSS.t575 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1276 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t3 a_n3659_3164.t2 a_n3629_3190.t3 VSS.t603 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1277 a_n22425_n7992.t0 A2.t14 VSS.t248 VSS.t220 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1278 a_11865_n29943.t8 mux8_8.NAND4F_8.Y.t12 VDD.t741 VDD.t740 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X1279 VDD.t3947 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t13 a_n13192_2026.t8 VDD.t3946 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1280 a_n11274_n29052.t3 a_n12345_n28506.t3 VSS.t936 VSS.t935 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1281 mux8_7.NAND4F_3.Y.t1 mux8_7.NAND4F_0.C.t10 VDD.t190 VDD.t189 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1282 VDD.t2873 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t12 a_n18042_2026.t9 VDD.t2872 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1283 VSS.t156 a_n8200_1380.t4 a_n8170_1406.t4 VSS.t155 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1284 VDD.t1762 SEL3.t23 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t3 VDD.t1761 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1285 VSS.t293 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t16 a_n9305_n8419.t0 VSS.t292 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1286 VSS.t811 A4.t10 OR8_0.NOT8_0.A4.t5 VSS.t810 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X1287 VDD.t2625 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t13 a_n3320_2026.t8 VDD.t2624 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X1288 a_n11274_n25843.t4 A4.t11 VSS.t813 VSS.t812 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1289 a_11386_n17350.t1 mux8_4.NAND4F_6.Y.t10 a_11290_n17350.t0 VSS.t103 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1290 VDD.t1855 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t7 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t0 VDD.t1854 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1291 a_n10714_n8445.t1 MULT_0.4bit_ADDER_1.A0.t6 VDD.t3189 VDD.t3188 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1292 a_8592_n3766.t1 SEL0.t51 a_8496_n3766.t1 VSS.t2006 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1293 a_11290_n3766.t1 mux8_1.NAND4F_1.Y.t9 a_11194_n3766.t0 VSS.t464 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1294 a_n12316_n34281.t8 B7.t9 VDD.t1397 VDD.t1396 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1295 VSS.t614 left_shifter_0.buffer_6.inv_1.A.t5 left_shifter_0.S1.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1296 MULT_0.4bit_ADDER_2.B0.t5 a_n12596_n8419.t4 a_n12416_n7799.t4 VDD.t1838 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1297 mux8_0.NAND4F_5.Y.t5 left_shifter_0.C.t5 VDD.t1686 VDD.t1685 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1298 left_shifter_0.S7.t3 left_shifter_0.buffer_2.inv_1.A.t5 VDD.t1310 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1299 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t1 MULT_0.4bit_ADDER_0.A2.t10 VDD.t248 VDD.t247 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1300 mux8_8.NAND4F_6.Y.t2 right_shifter_0.S6.t4 a_8592_n30934.t0 VSS.t527 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1301 VDD.t518 A2.t15 MULT_0.NAND2_1.Y.t2 VDD.t517 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1302 a_n15707_n4534.t9 a_n15737_n5180.t6 MULT_0.4bit_ADDER_1.B1.t9 VDD.t929 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1303 a_10459_n30933.t0 SEL0.t52 a_10363_n30933.t1 VSS.t1988 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1304 mux8_3.NAND4F_1.Y.t4 XOR8_0.S2.t12 VDD.t1208 VDD.t1207 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1305 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t9 VDD.t3408 VDD.t3407 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1306 a_5197_5532.t5 a_5167_4886.t4 V_FLAG_0.XOR2_0.Y.t8 VDD.t56 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1307 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t10 a_n20113_3164.t4 a_n20083_3190.t3 VSS.t1325 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1308 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t1 a_n18222_1406.t4 a_n18042_1406.t5 VSS.t1767 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1309 a_11865_n29943.t3 mux8_8.NAND4F_9.Y.t10 mux8_8.inv_0.A.t3 VDD.t1111 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1310 VDD.t614 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t17 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t5 VDD.t613 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1311 VSS.t1016 VSS.t1014 a_n20737_n5154.t0 VSS.t1015 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1312 mux8_4.inv_0.A.t4 mux8_4.NAND4F_9.Y.t10 a_11865_n16359.t8 VDD.t961 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1313 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t1 a_n24804_1406.t4 a_n24624_2026.t1 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1314 VDD.t4404 SEL1.t51 mux8_8.NAND4F_5.Y.t6 VDD.t4403 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1315 a_n18305_n12716.t1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t8 VSS.t484 VSS.t483 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1316 VDD.t4203 A1.t15 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t6 VDD.t4202 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1317 VDD.t853 mux8_0.NAND4F_4.B.t9 mux8_0.NAND4F_3.Y.t0 VDD.t852 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1318 VDD.t491 mux8_6.NAND4F_5.Y.t10 mux8_6.NAND4F_9.Y.t4 VDD.t490 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1319 VDD.t3745 SEL2.t36 mux8_6.NAND4F_7.Y.t1 VDD.t3744 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1320 mux8_5.NAND4F_4.B.t0 SEL0.t53 VSS.t2005 VSS.t2004 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1321 VDD.t4141 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t17 a_n4879_2026.t7 VDD.t4140 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1322 VDD.t2777 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t10 a_n12416_n11063.t9 VDD.t2776 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X1323 mux8_0.NAND4F_0.C.t3 SEL1.t52 VDD.t4406 VDD.t4405 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1324 a_5197_4912.t2 a_5017_4912.t3 V_FLAG_0.XOR2_0.Y.t5 VSS.t1085 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1325 a_8496_762.t0 SEL1.t53 a_8400_762.t1 VSS.t1968 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1326 a_n17677_n19625.t2 A3.t20 OR8_0.NOT8_0.A3.t3 VDD.t4098 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1327 mux8_4.NAND4F_1.Y.t2 mux8_4.NAND4F_0.C.t8 VDD.t3253 VDD.t3252 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1328 mux8_4.NAND4F_0.Y.t6 mux8_4.A1.t13 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1329 a_n17368_3190.t2 SEL3.t24 VSS.t884 VSS.t883 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X1330 AND8_0.S6.t1 AND8_0.NOT8_0.A6.t8 VDD.t1572 VDD.t1571 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1331 VSS.t1764 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t16 a_n12596_n8419.t0 VSS.t1763 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1332 VDD.t4011 MULT_0.inv_9.Y.t10 a_n13975_n11063.t5 VDD.t4010 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1333 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t1 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t8 VDD.t1857 VDD.t1856 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1334 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t13 VDD.t2738 VDD.t2737 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1335 mux8_7.inv_0.A.t3 mux8_7.NAND4F_9.Y.t12 a_11865_n25415.t2 VDD.t3283 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X1336 a_n14005_n8445.t0 MULT_0.4bit_ADDER_1.A1.t7 VDD.t110 VDD.t109 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1337 a_n17266_n11063.t7 a_n17296_n11709.t5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t10 VDD.t2857 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1338 VDD.t2803 mux8_3.NAND4F_2.D.t9 mux8_3.NAND4F_2.Y.t4 VDD.t2802 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1339 a_n11274_n31661.t3 a_n12345_n31115.t2 VSS.t1310 VSS.t1309 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1340 a_n11276_n33705.t5 B7.t10 XOR8_0.S7.t11 VSS.t685 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1341 VDD.t3457 mux8_4.inv_0.A.t7 Y3.t0 VDD.t3456 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1342 a_11290_n16422.t0 mux8_4.NAND4F_3.Y.t9 a_11194_n16422.t0 VSS.t967 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1343 a_n11490_1380.t1 A3.t21 VDD.t4100 VDD.t4099 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1344 a_n18998_n7799.t4 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t15 VDD.t1047 VDD.t1046 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1345 NOT8_0.S1.t3 B1.t17 VDD.t2340 VDD.t2339 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1346 a_n14077_3810.t10 a_n13531_3164.t5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t4 VDD.t2730 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1347 a_n24654_1380.t0 A7.t17 VSS.t1572 VSS.t1571 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1348 AND8_0.NOT8_0.A2.t6 B2.t14 VDD.t2593 VDD.t2592 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1349 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t4 a_n1768_1406.t4 a_n1588_1406.t1 VSS.t278 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1350 a_11194_n20950.t1 mux8_5.NAND4F_0.Y.t11 VSS.t1568 VSS.t104 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1351 VDD.t3191 MULT_0.4bit_ADDER_1.A0.t7 a_n10684_n7799.t11 VDD.t3190 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1352 mux8_5.A1.t8 a_n12596_n11683.t4 a_n12416_n11063.t2 VDD.t1241 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1353 mux8_7.A1.t7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t14 a_n15131_n11683.t1 VSS.t630 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1354 OR8_0.S6.t2 OR8_0.NOT8_0.A6.t8 VDD.t320 VDD.t319 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1355 a_n4205_3810.t10 B1.t18 VDD.t2342 VDD.t2341 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1356 VDD.t4408 SEL1.t54 mux8_2.NAND4F_4.Y.t4 VDD.t4407 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1357 a_n8432_n9452.t1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t9 VSS.t1124 VSS.t1123 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1358 MULT_0.inv_9.Y.t0 MULT_0.NAND2_9.Y.t7 VSS.t1781 VSS.t1780 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1359 a_n12316_n15299.t10 B0.t13 VDD.t988 VDD.t987 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1360 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t4 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t18 VDD.t616 VDD.t615 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1361 a_n10684_n7799.t5 MULT_0.4bit_ADDER_1.B0.t16 VDD.t2506 VDD.t2505 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1362 mux8_3.NAND4F_3.Y.t5 mux8_3.NAND4F_4.B.t6 VDD.t2524 VDD.t2523 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1363 a_n17677_n25225.t9 B7.t11 VDD.t1399 VDD.t1398 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1364 OR8_0.NOT8_0.A5.t4 A5.t11 a_n17677_n22425.t8 VDD.t389 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X1365 VDD.t977 V_FLAG_0.XOR2_2.B.t15 a_3493_5534.t4 VDD.t976 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1366 left_shifter_0.C.t0 left_shifter_0.buffer_1.inv_1.A.t4 VDD.t136 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1367 XOR8_0.S1.t5 B1.t19 a_n11274_n17539.t2 VSS.t1175 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1368 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t5 A1.t16 VDD.t4205 VDD.t4204 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1369 mux8_5.NAND4F_1.Y.t2 mux8_5.NAND4F_0.C.t7 VDD.t3628 VDD.t3627 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1370 mux8_1.NAND4F_7.Y.t1 SEL2.t37 VDD.t3747 VDD.t3746 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1371 a_n11274_n28476.t2 B5.t8 XOR8_0.S5.t3 VSS.t443 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1372 a_n14751_2026.t0 a_n14781_1380.t3 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t0 VDD.t557 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1373 a_n4205_3190.t1 SEL3.t25 VSS.t886 VSS.t885 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X1374 mux8_0.NAND4F_9.Y.t5 mux8_0.NAND4F_6.Y.t11 VDD.t2069 VDD.t2068 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1375 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t5 VSS.t2046 VDD.t1957 VDD.t1956 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1376 mux8_8.NAND4F_2.Y.t0 mux8_8.NAND4F_2.D.t9 VDD.t1510 VDD.t1509 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1377 a_n13192_2026.t1 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t18 VDD.t348 VDD.t347 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1378 buffer_0.inv_1.A.t0 Y7.t6 VSS.t538 VSS.t537 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1379 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t9 a_n21363_1380.t3 a_n21333_2026.t9 VDD.t1215 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1380 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t7 a_n2627_373.t0 VSS.t672 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1381 a_n13975_n7799.t9 a_n14005_n8445.t3 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t9 VDD.t3620 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1382 a_n914_3810.t1 SEL3.t26 VDD.t1764 VDD.t1763 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1383 mux8_0.NAND4F_6.Y.t6 right_shifter_0.C.t6 a_8592_762.t0 VSS.t983 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1384 VDD.t1126 MULT_0.NAND2_4.Y.t8 MULT_0.4bit_ADDER_0.A0.t3 VDD.t1125 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1385 a_n9125_n11063.t10 VSS.t2047 VDD.t1955 VDD.t1954 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1386 a_11386_n30934.t1 mux8_8.NAND4F_6.Y.t10 a_11290_n30934.t0 VSS.t166 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1387 mux8_3.NAND4F_5.Y.t7 left_shifter_0.S2.t5 VDD.t3400 VDD.t3399 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1388 VDD.t3045 SEL0.t54 mux8_1.NAND4F_0.Y.t7 VDD.t3044 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1389 VDD.t4176 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t14 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t5 VDD.t4175 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1390 a_n13399_n8419.t5 MULT_0.4bit_ADDER_1.B1.t14 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t6 VSS.t1500 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1391 XOR8_0.S2.t9 a_n12345_n20814.t3 a_n11274_n21072.t3 VSS.t1425 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1392 VDD.t677 AND8_0.NOT8_0.A4.t9 AND8_0.S4.t2 VDD.t676 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1393 VDD.t1057 MULT_0.NAND2_2.Y.t8 MULT_0.4bit_ADDER_0.B0.t3 VDD.t1056 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1394 mux8_7.NAND4F_0.Y.t2 mux8_7.A1.t12 VDD.t1106 VDD.t1105 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1395 OR8_0.NOT8_0.A4.t4 A4.t12 a_n17677_n21025.t5 VDD.t1637 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1396 NOT8_0.S1.t2 B1.t20 VDD.t2344 VDD.t2343 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1397 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t2 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t9 VDD.t1859 VDD.t1858 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1398 a_n13975_n4534.t11 MULT_0.4bit_ADDER_0.B1.t6 VDD.t1333 VDD.t1332 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1399 VDD.t1533 8bit_ADDER_0.S1.t12 mux8_2.NAND4F_3.Y.t6 VDD.t1532 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1400 a_9432_1690.t1 mux8_0.NAND4F_0.C.t7 a_9336_1690.t1 VSS.t317 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1401 VDD.t1294 MULT_0.4bit_ADDER_0.A0.t7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t4 VDD.t1293 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1402 a_11865_n11831.t2 mux8_3.NAND4F_8.Y.t12 VDD.t3925 VDD.t3924 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1403 mux8_6.inv_0.A.t5 mux8_6.NAND4F_9.Y.t11 a_11865_n34471.t7 VDD.t696 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X1404 mux8_5.A1.t9 a_n12596_n11683.t5 a_n12416_n11063.t1 VDD.t1242 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1405 VSS.t418 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t12 a_n15131_n11683.t5 VSS.t417 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1406 VDD.t3043 SEL0.t55 mux8_0.NAND4F_2.Y.t8 VDD.t3042 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1407 NOT8_0.S6.t3 B6.t16 VDD.t3546 VDD.t3545 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1408 MULT_0.4bit_ADDER_2.B1.t11 a_n15737_n8445.t3 a_n15707_n7799.t11 VDD.t59 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1409 VDD.t4410 SEL1.t55 mux8_1.NAND4F_0.C.t3 VDD.t4409 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1410 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t2 a_n10864_n11683.t3 a_n10684_n11683.t2 VSS.t760 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1411 OR8_0.S4.t3 OR8_0.NOT8_0.A4.t8 VDD.t369 VDD.t311 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1412 a_n10240_3164.t1 B3.t15 VDD.t2156 VDD.t2155 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1413 VDD.t426 mux8_6.NAND4F_2.D.t9 mux8_6.NAND4F_2.Y.t1 VDD.t425 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1414 a_n17266_n4534.t1 MULT_0.4bit_ADDER_0.A2.t11 VDD.t250 VDD.t249 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1415 MULT_0.4bit_ADDER_2.B1.t3 a_n15887_n8419.t3 a_n15707_n8419.t0 VSS.t709 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1416 mux8_2.NAND4F_1.Y.t5 mux8_2.NAND4F_0.C.t6 VDD.t3203 VDD.t3202 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1417 a_n11723_n9452.t1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t7 VSS.t1919 VSS.t1687 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1418 VDD.t4412 SEL1.t56 mux8_1.NAND4F_2.Y.t6 VDD.t4411 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1419 mux8_1.NAND4F_8.Y.t3 mux8_1.NAND4F_3.Y.t9 VDD.t931 VDD.t930 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1420 VDD.t2087 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t14 a_n1768_1406.t0 VDD.t2086 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X1421 a_n4303_1406.t5 A1.t17 VSS.t1900 VSS.t1899 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1422 VDD.t4207 A1.t18 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t4 VDD.t4206 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1423 VDD.t1491 OR8_0.S2.t4 mux8_3.NAND4F_2.Y.t2 VDD.t1490 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1424 VSS.t1521 mux8_6.A0.t16 a_5773_4912.t4 VSS.t1520 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1425 VDD.t456 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t18 a_n15707_n4534.t1 VDD.t455 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1426 mux8_3.NAND4F_7.Y.t7 SEL0.t56 VDD.t3041 VDD.t3040 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1427 VSS.t714 a_n10966_3190.t3 a_n10210_3190.t5 VSS.t713 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1428 mux8_0.inv_0.A.t0 mux8_0.NAND4F_8.Y.t11 VSS.t1615 VSS.t1614 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1429 mux8_8.NAND4F_1.Y.t7 mux8_8.NAND4F_0.C.t7 VDD.t2658 VDD.t2657 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1430 mux8_6.NAND4F_3.Y.t4 mux8_6.NAND4F_4.B.t8 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1431 a_n11274_n25843.t1 B4.t17 XOR8_0.S4.t4 VSS.t1650 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1432 XOR8_0.S3.t5 a_n12345_n23393.t4 a_n11274_n23651.t1 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1433 a_16143_n19505.t4 Y6.t6 a_16431_n19505.t4 VDD.t3168 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X1434 VDD.t827 AND8_0.NOT8_0.A1.t9 AND8_0.S1.t2 VDD.t826 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1435 VSS.t80 a_n15737_n11709.t3 a_n15707_n11683.t5 VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1436 a_n11274_n31085.t1 B6.t17 XOR8_0.S6.t1 VSS.t1631 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1437 a_n15707_n7799.t10 a_n15737_n8445.t4 MULT_0.4bit_ADDER_2.B1.t10 VDD.t60 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1438 a_n10786_3190.t2 SEL3.t27 VSS.t888 VSS.t887 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1439 mux8_0.NAND4F_0.Y.t7 SEL0.t57 VDD.t3039 VDD.t3038 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1440 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t8 B5.t9 a_n17368_3190.t5 VSS.t444 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1441 VDD.t2558 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t10 a_n18998_n4534.t7 VDD.t2557 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1442 AND8_0.NOT8_0.A2.t4 A2.t16 VDD.t520 VDD.t519 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1443 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t17 VDD.t2013 VDD.t2012 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1444 VDD.t2494 right_shifter_0.buffer_5.inv_1.A.t5 right_shifter_0.S2.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1445 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t8 a_n6950_3164.t2 a_n6920_3190.t5 VSS.t1805 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1446 VSS.t368 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t17 a_n3500_1406.t0 VSS.t367 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1447 VDD.t4209 A1.t19 AND8_0.NOT8_0.A1.t2 VDD.t4208 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1448 VDD.t2751 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t9 a_n16483_2026.t4 VDD.t2750 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1449 a_n22489_1406.t3 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t14 mux8_6.A0.t0 VSS.t1601 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1450 VDD.t1953 VSS.t2048 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t4 VDD.t1952 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1451 VSS.t1619 MULT_0.inv_8.Y.t8 a_n10108_n11683.t5 VSS.t1618 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1452 a_11865_n11831.t1 mux8_3.NAND4F_8.Y.t13 VDD.t3927 VDD.t3926 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X1453 a_n20659_3810.t1 SEL3.t28 VDD.t1766 VDD.t1765 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1454 VDD.t4211 A1.t20 MULT_0.NAND2_2.Y.t6 VDD.t4210 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1455 VDD.t89 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t9 a_n6611_2026.t1 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X1456 mux8_8.NAND4F_2.Y.t7 OR8_0.S6.t5 VDD.t3146 VDD.t3145 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1457 a_n20587_n11709.t0 MULT_0.inv_15.Y.t7 VSS.t1529 VSS.t1528 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1458 a_n19187_n12716.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t16 VSS.t1673 VSS.t465 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1459 a_n12314_n18115.t1 B1.t21 VDD.t2346 VDD.t2345 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1460 a_8496_n16422.t0 SEL1.t57 a_8400_n16422.t1 VSS.t1969 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1461 a_n17296_n8445.t0 MULT_0.4bit_ADDER_1.A2.t6 VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1462 a_n9125_n11063.t8 a_n9305_n11683.t4 mux8_4.A1.t8 VDD.t2033 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1463 mux8_7.NAND4F_9.Y.t5 mux8_7.NAND4F_5.Y.t11 VDD.t2040 VDD.t2039 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1464 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t8 a_n23404_3164.t4 a_n23374_3190.t4 VSS.t1209 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1465 a_n11460_1406.t1 a_n11490_1380.t4 VSS.t477 VSS.t476 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X1466 VDD.t1951 VSS.t2049 mux8_0.NAND4F_1.Y.t8 VDD.t1950 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1467 MULT_0.4bit_ADDER_0.B2.t1 MULT_0.NAND2_0.Y.t8 VSS.t579 VSS.t578 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1468 a_n21333_2026.t2 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t14 VDD.t3235 VDD.t3234 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1469 left_shifter_0.buffer_3.inv_1.A.t3 B5.t10 VDD.t899 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1470 VDD.t1875 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t9 a_n23065_2026.t4 VDD.t1874 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X1471 a_n12345_n25873.t0 A4.t13 VSS.t815 VSS.t814 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1472 ZFLAG_0.nor4_1.Y.t5 Y4.t7 VSS.t1347 VSS.t1346 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1473 VSS.t1675 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t17 a_n19178_n11683.t0 VSS.t1674 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1474 a_11865_n11831.t8 mux8_3.NAND4F_9.Y.t10 mux8_3.inv_0.A.t2 VDD.t2616 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1475 a_n13975_n8419.t4 a_n14005_n8445.t4 VSS.t1661 VSS.t1660 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X1476 mux8_3.NAND4F_8.Y.t5 mux8_3.NAND4F_4.Y.t10 a_11386_n11894.t0 VSS.t461 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1477 a_10363_n25478.t0 mux8_7.NAND4F_0.C.t11 a_10267_n25478.t0 VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1478 mux8_4.NAND4F_2.Y.t8 SEL0.t58 VDD.t3037 VDD.t3036 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1479 mux8_3.NAND4F_6.Y.t6 SEL1.t58 VDD.t4414 VDD.t4413 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1480 a_n13531_3164.t1 B4.t18 VDD.t3597 VDD.t3596 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1481 VDD.t1223 OR8_0.S7.t4 mux8_6.NAND4F_2.Y.t2 VDD.t1222 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1482 VDD.t4047 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t8 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t5 VDD.t4046 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1483 mux8_2.NAND4F_3.Y.t4 8bit_ADDER_0.S1.t13 a_9528_n7266.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1484 VSS.t671 AND8_0.NOT8_0.A0.t8 AND8_0.S0.t0 VSS.t670 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1485 VDD.t1311 left_shifter_0.buffer_2.inv_1.A.t6 left_shifter_0.S7.t2 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1486 a_n13714_n12716.t1 MULT_0.4bit_ADDER_2.B1.t15 VSS.t968 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1487 VDD.t4416 SEL1.t59 mux8_2.NAND4F_5.Y.t3 VDD.t4415 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1488 VDD.t4286 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t11 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t2 VDD.t4285 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1489 VDD.t2526 mux8_3.NAND4F_4.B.t7 mux8_3.NAND4F_1.Y.t6 VDD.t2525 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1490 VSS.t1116 a_n9931_1380.t4 a_n9901_1406.t4 VSS.t1115 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1491 VDD.t240 mux8_4.A0.t12 mux8_4.NAND4F_3.Y.t8 VDD.t239 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1492 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t4 a_n14155_n8419.t3 a_n13975_n7799.t4 VDD.t3688 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1493 VSS.t970 MULT_0.4bit_ADDER_2.B1.t16 a_n14155_n11683.t0 VSS.t969 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1494 VDD.t2491 mux8_8.A1.t12 mux8_8.NAND4F_0.Y.t6 VDD.t2490 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1495 VDD.t4001 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t3 VDD.t4000 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1496 VSS.t836 A0.t12 a_n1012_1406.t1 VSS.t835 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1497 VDD.t1401 B7.t12 a_n17677_n25225.t8 VDD.t1400 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1498 a_n17677_n22425.t7 A5.t12 OR8_0.NOT8_0.A5.t3 VDD.t390 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1499 a_16431_n18523.t3 Y1.t6 a_16143_n18523.t0 VDD.t3169 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X1500 VDD.t680 right_shifter_0.buffer_3.inv_1.A.t5 right_shifter_0.S4.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1501 VSS.t500 B0.t14 NOT8_0.S0.t0 VSS.t499 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1502 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t7 a_n10966_3190.t4 a_n10786_3810.t7 VDD.t1447 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1503 mux8_2.NAND4F_4.Y.t0 AND8_0.S1.t4 a_7644_n7266.t0 VSS.t396 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1504 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t4 MULT_0.4bit_ADDER_1.B2.t16 VDD.t4031 VDD.t4030 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1505 mux8_8.inv_0.A.t2 mux8_8.NAND4F_9.Y.t11 a_11865_n29943.t2 VDD.t1112 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1506 a_n11274_n17539.t1 B1.t22 XOR8_0.S1.t6 VSS.t1176 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1507 a_n14781_1380.t1 A4.t14 VDD.t1639 VDD.t1638 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1508 VSS.t1663 a_n14005_n8445.t5 a_n13975_n8419.t3 VSS.t1662 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1509 a_n19981_n11683.t2 MULT_0.4bit_ADDER_2.B3.t10 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t9 VSS.t1825 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1510 a_11865_n16359.t2 mux8_4.NAND4F_8.Y.t9 VDD.t1478 VDD.t1477 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1511 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t7 a_n15014_n6187.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1512 a_n17368_3810.t4 a_n16822_3164.t5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t4 VDD.t2855 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1513 a_10267_1690.t0 mux8_0.NAND4F_2.D.t7 VSS.t1438 VSS.t1437 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1514 VSS.t315 MULT_0.4bit_ADDER_0.A3.t8 a_n19981_n5154.t2 VSS.t314 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1515 MULT_0.4bit_ADDER_1.B3.t6 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t8 VDD.t4326 VDD.t4325 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1516 a_n19028_n8445.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t12 VSS.t1868 VSS.t1867 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1517 a_8400_n21878.t0 SEL2.t38 VSS.t1718 VSS.t681 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1518 AND8_0.NOT8_0.A7.t5 B7.t13 VDD.t1403 VDD.t1402 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1519 a_n7496_3810.t10 B2.t15 VDD.t2595 VDD.t2594 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1520 VDD.t19 MULT_0.4bit_ADDER_1.A2.t7 a_n17266_n7799.t11 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X1521 a_10267_n7266.t0 mux8_2.NAND4F_2.D.t6 VSS.t1475 VSS.t1474 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1522 mux8_6.NAND4F_9.Y.t3 mux8_6.NAND4F_5.Y.t11 VDD.t493 VDD.t492 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1523 mux8_6.NAND4F_7.Y.t0 SEL2.t39 VDD.t3749 VDD.t3748 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1524 VDD.t2538 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t8 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t3 VDD.t2537 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1525 VDD.t3149 MULT_0.NAND2_5.Y.t8 MULT_0.4bit_ADDER_0.A1.t2 VDD.t3147 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1526 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t11 VDD.t703 VDD.t702 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1527 mux8_5.NAND4F_4.Y.t8 SEL1.t60 VDD.t4418 VDD.t4417 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1528 MULT_0.4bit_ADDER_0.A0.t2 MULT_0.NAND2_4.Y.t9 VDD.t1127 VDD.t1125 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1529 VDD.t4420 SEL1.t61 mux8_1.NAND4F_6.Y.t5 VDD.t4419 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1530 mux8_1.NAND4F_9.Y.t6 mux8_1.NAND4F_1.Y.t10 VDD.t1307 VDD.t1306 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1531 mux8_4.NAND4F_5.Y.t2 left_shifter_0.S3.t4 a_7644_n17350.t0 VSS.t957 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1532 a_n29_2026.t1 SEL3.t29 VDD.t1768 VDD.t1767 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1533 a_n914_3190.t4 B0.t15 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t10 VSS.t501 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1534 a_n9901_2026.t1 a_n9931_1380.t5 mux8_4.A0.t11 VDD.t2184 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1535 a_n15707_n7799.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t14 VDD.t665 VDD.t664 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1536 a_n11274_n21072.t4 a_n12345_n20814.t4 XOR8_0.S2.t10 VSS.t1426 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1537 mux8_5.NAND4F_1.Y.t6 XOR8_0.S4.t12 a_9528_n21878.t1 VSS.t1541 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1538 a_n24013_n15316.t0 A0.t13 AND8_0.NOT8_0.A0.t4 VSS.t837 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1539 VDD.t3035 SEL0.t59 mux8_4.NAND4F_0.Y.t8 VDD.t3034 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1540 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t5 a_n17446_n5154.t4 a_n17266_n4534.t8 VDD.t2427 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1541 a_n15707_n8419.t4 a_n15737_n8445.t5 VSS.t28 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X1542 VDD.t65 XOR8_0.S1.t14 mux8_2.NAND4F_1.Y.t2 VDD.t64 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1543 a_n13975_n11063.t4 MULT_0.inv_9.Y.t11 VDD.t4013 VDD.t4012 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1544 a_n18042_2026.t7 a_n18072_1380.t5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t7 VDD.t2046 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1545 VDD.t1949 VSS.t2050 a_n9125_n7799.t9 VDD.t1948 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1546 a_n7496_3190.t1 SEL3.t30 VSS.t890 VSS.t889 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X1547 VDD.t1161 mux8_8.NAND4F_2.Y.t9 mux8_8.NAND4F_8.Y.t5 VDD.t1160 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1548 mux8_7.NAND4F_2.Y.t6 SEL0.t60 VDD.t3033 VDD.t3032 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1549 VSS.t1288 B2.t16 a_n12345_n20814.t0 VSS.t1287 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1550 VDD.t771 mux8_1.NAND4F_4.Y.t11 mux8_1.NAND4F_8.Y.t1 VDD.t770 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1551 a_n23950_3810.t1 B7.t14 VDD.t1405 VDD.t1404 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1552 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t7 a_n24654_1380.t5 a_n24624_2026.t7 VDD.t3881 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1553 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t4 MULT_0.4bit_ADDER_1.B0.t17 a_n10108_n8419.t2 VSS.t1260 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1554 MULT_0.S2.t10 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t17 a_n8549_n8419.t1 VSS.t294 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1555 VDD.t2634 MULT_0.NAND2_14.Y.t8 MULT_0.inv_14.Y.t2 VDD.t2632 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1556 mux8_3.NAND4F_2.Y.t3 mux8_3.NAND4F_2.D.t10 VDD.t2805 VDD.t2804 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1557 a_11194_n16422.t1 mux8_4.NAND4F_0.Y.t9 VSS.t398 VSS.t397 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1558 a_n18998_n7799.t10 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t13 VDD.t4157 VDD.t4156 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1559 VDD.t3470 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t15 a_n23065_2026.t2 VDD.t3469 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1560 a_n6611_2026.t11 a_n6791_1406.t3 8bit_ADDER_0.S2.t10 VDD.t3379 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1561 VDD.t1821 ZFLAG_0.nor4_0.Y.t7 ZFLAG_0.NAND2_0.Y.t2 VDD.t1820 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1562 VDD.t2348 B1.t23 NOT8_0.S1.t1 VDD.t2347 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1563 VDD.t1407 B7.t15 a_1887_5534.t7 VDD.t1406 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X1564 a_n8549_n5154.t3 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t14 MULT_0.S1.t3 VSS.t1068 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1565 mux8_6.NAND4F_8.Y.t2 mux8_6.NAND4F_4.Y.t10 a_11386_n34534.t0 VSS.t234 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1566 a_n18422_n8419.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t16 MULT_0.4bit_ADDER_2.B2.t8 VSS.t520 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1567 a_11865_n7203.t2 mux8_2.NAND4F_8.Y.t11 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1568 OR8_0.NOT8_0.A3.t0 B3.t16 VSS.t1108 VSS.t810 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1569 VDD.t606 mux8_7.A0.t12 mux8_7.NAND4F_3.Y.t4 VDD.t605 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1570 a_n18998_n4534.t4 a_n19178_n5154.t5 MULT_0.4bit_ADDER_1.B2.t5 VDD.t692 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1571 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t2 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t8 VDD.t867 VDD.t866 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1572 MULT_0.NAND2_8.Y.t3 B3.t17 a_n24162_n11256.t1 VSS.t1109 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1573 VSS.t413 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t14 a_n19954_1406.t0 VSS.t412 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1574 VDD.t1889 mux8_4.NAND4F_3.Y.t10 mux8_4.NAND4F_8.Y.t1 VDD.t1888 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1575 VSS.t1391 A6.t12 a_n20757_1406.t5 VSS.t1390 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1576 XOR8_0.S4.t10 a_n12345_n26161.t4 a_n11274_n26419.t4 VSS.t1877 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1577 a_n11274_n23651.t4 a_n12345_n23105.t3 VSS.t1362 VSS.t1361 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1578 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t2 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t9 VDD.t2540 VDD.t2539 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1579 MULT_0.NAND2_2.Y.t1 B0.t16 VDD.t990 VDD.t989 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1580 MULT_0.NAND2_3.Y.t6 B0.t17 VDD.t992 VDD.t991 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1581 VDD.t1361 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t9 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t5 VDD.t1360 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1582 VDD.t522 A2.t17 MULT_0.NAND2_10.Y.t1 VDD.t521 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1583 MULT_0.inv_6.A.t5 A0.t14 VDD.t1670 VDD.t1669 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1584 a_11290_n8194.t1 mux8_2.NAND4F_1.Y.t11 a_11194_n8194.t1 VSS.t318 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1585 VDD.t1947 VSS.t2051 a_n9125_n11063.t9 VDD.t1946 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X1586 a_8592_n8194.t1 SEL0.t61 a_8496_n8194.t1 VSS.t2008 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1587 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t2 SEL3.t31 VDD.t1770 VDD.t1769 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1588 VDD.t4288 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t12 a_n12416_n7799.t6 VDD.t4287 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1589 AND8_0.NOT8_0.A3.t1 B3.t18 VDD.t2158 VDD.t2157 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1590 mux8_4.NAND4F_6.Y.t8 SEL0.t62 VDD.t3031 VDD.t3030 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1591 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t2 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t8 VDD.t224 VDD.t223 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1592 VDD.t3029 SEL0.t63 mux8_7.NAND4F_0.Y.t6 VDD.t3028 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1593 VDD.t3255 mux8_4.NAND4F_0.C.t9 mux8_4.NAND4F_7.Y.t7 VDD.t3254 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1594 VDD.t667 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t15 a_n15887_n8419.t1 VDD.t666 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X1595 mux8_3.NAND4F_2.Y.t0 OR8_0.S2.t5 a_8592_n11894.t0 VSS.t562 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1596 right_shifter_0.S2.t2 right_shifter_0.buffer_5.inv_1.A.t6 VDD.t2495 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1597 V_FLAG_0.XOR2_2.Y.t8 a_3313_4914.t4 a_3493_5534.t7 VDD.t1097 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1598 MULT_0.4bit_ADDER_2.B0.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t17 a_n11840_n8419.t1 VSS.t1765 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1599 a_n14077_3190.t1 SEL3.t32 VSS.t892 VSS.t891 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1600 VDD.t2159 B3.t19 right_shifter_0.buffer_5.inv_1.A.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1601 a_11194_1690.t0 mux8_0.NAND4F_0.Y.t11 VSS.t619 VSS.t618 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1602 a_n11840_n5154.t5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t15 MULT_0.4bit_ADDER_1.B0.t11 VSS.t1878 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1603 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t9 VDD.t3684 VDD.t3683 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1604 a_n12416_n11063.t5 a_n12446_n11709.t3 mux8_5.A1.t2 VDD.t4307 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1605 a_n15131_n11683.t4 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t13 VSS.t420 VSS.t419 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1606 a_n4205_3190.t5 B1.t24 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t9 VSS.t1177 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1607 a_n13192_2026.t4 a_n13222_1380.t3 mux8_5.A0.t10 VDD.t773 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1608 a_n11460_2026.t4 A3.t22 VDD.t4102 VDD.t4101 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1609 VDD.t362 right_shifter_0.buffer_7.inv_1.A.t5 right_shifter_0.S0.t1 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1610 a_8592_1690.t1 SEL0.t64 a_8496_1690.t1 VSS.t2007 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1611 a_n10684_n11683.t1 a_n10864_n11683.t4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t3 VSS.t761 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1612 VDD.t370 OR8_0.NOT8_0.A4.t9 OR8_0.S4.t2 VDD.t313 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1613 VDD.t1147 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t9 a_n19774_2026.t2 VDD.t1146 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1614 VSS.t1249 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t14 a_n6791_1406.t0 VSS.t1248 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1615 mux8_6.NAND4F_2.Y.t0 mux8_6.NAND4F_2.D.t10 VDD.t428 VDD.t427 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1616 VDD.t44 XOR8_0.S3.t13 mux8_4.NAND4F_1.Y.t6 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1617 XOR8_0.S0.t9 a_n12347_n15041.t4 a_n11276_n15299.t4 VSS.t1692 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1618 a_n3320_2026.t5 a_n3350_1380.t4 8bit_ADDER_0.S1.t5 VDD.t2266 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1619 a_n13975_n11063.t2 a_n14155_n11683.t4 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t8 VDD.t2022 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1620 VDD.t3027 SEL0.t65 mux8_4.NAND4F_4.B.t1 VDD.t3026 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1621 a_n23950_3810.t7 SEL3.t33 VDD.t1772 VDD.t1771 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1622 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t1 a_n7676_3190.t5 a_n7496_3810.t4 VDD.t3959 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1623 a_7452_n12822.t0 SEL2.t40 VSS.t1719 VSS.t1384 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1624 MULT_0.4bit_ADDER_0.B1.t2 MULT_0.NAND2_1.Y.t8 VDD.t237 VDD.t236 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1625 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t10 MULT_0.4bit_ADDER_2.B3.t11 a_n19981_n11683.t1 VSS.t1826 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1626 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t5 a_n17446_n8419.t4 a_n17266_n8419.t3 VSS.t358 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1627 mux8_3.NAND4F_2.Y.t1 OR8_0.S2.t6 VDD.t1493 VDD.t1492 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1628 mux8_8.NAND4F_5.Y.t2 left_shifter_0.S6.t4 a_7644_n30934.t1 VSS.t613 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1629 VDD.t705 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t12 a_n15707_n4534.t8 VDD.t704 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X1630 VDD.t52 NOT8_0.S5.t5 mux8_7.NAND4F_7.Y.t6 VDD.t51 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1631 VDD.t1328 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t10 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t1 VDD.t1327 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1632 a_n20659_3190.t4 B6.t18 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t1 VSS.t1632 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1633 VDD.t1557 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t18 a_n10081_1406.t1 VDD.t1556 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X1634 VDD.t2548 mux8_7.NAND4F_3.Y.t10 mux8_7.NAND4F_8.Y.t5 VDD.t2547 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1635 mux8_5.NAND4F_6.Y.t5 SEL0.t66 VDD.t3025 VDD.t3024 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1636 a_n12616_1406.t5 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t14 VSS.t1785 VSS.t1784 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1637 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t4 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t10 VDD.t1363 VDD.t1362 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1638 a_7452_n3766.t0 SEL2.t41 VSS.t1720 VSS.t855 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1639 a_n15707_n11683.t4 a_n15737_n11709.t4 VSS.t82 VSS.t81 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1640 VDD.t3630 mux8_5.NAND4F_0.C.t8 mux8_5.NAND4F_7.Y.t3 VDD.t3629 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1641 a_n20557_n4534.t4 a_n20737_n5154.t6 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t4 VDD.t745 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1642 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t1 MULT_0.4bit_ADDER_1.B3.t12 VDD.t2717 VDD.t2716 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1643 VSS.t1194 AND8_0.NOT8_0.A3.t8 AND8_0.S3.t0 VSS.t329 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1644 VSS.t1550 a_n59_1380.t3 a_n29_1406.t5 VSS.t1549 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1645 a_n24624_2026.t10 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t14 VDD.t3642 VDD.t3641 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1646 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t0 MULT_0.4bit_ADDER_1.A2.t8 a_n17005_n9452.t1 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1647 VDD.t1369 mux8_5.NAND4F_2.D.t5 mux8_5.NAND4F_3.Y.t2 VDD.t1368 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1648 VDD.t2779 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t11 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t3 VDD.t2778 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1649 a_n17266_n7799.t1 a_n17296_n8445.t3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t1 VDD.t3289 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1650 right_shifter_0.S2.t1 right_shifter_0.buffer_5.inv_1.A.t7 VDD.t2496 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1651 mux8_7.NAND4F_0.C.t2 SEL1.t62 VDD.t4421 VDD.t4345 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1652 VDD.t4131 XOR8_0.S4.t13 mux8_5.NAND4F_1.Y.t8 VDD.t4130 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1653 a_10363_n2838.t0 mux8_1.NAND4F_0.C.t7 a_10267_n2838.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1654 VDD.t1600 mux8_1.NAND4F_5.Y.t10 mux8_1.NAND4F_9.Y.t3 VDD.t1599 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1655 a_n11274_n18115.t0 a_n12345_n17569.t2 VSS.t640 VSS.t639 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1656 VSS.t759 a_n14257_3190.t3 a_n13501_3190.t1 VSS.t758 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1657 a_n15014_n6187.t1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t9 VSS.t534 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1658 VDD.t3023 SEL0.t67 mux8_8.NAND4F_2.Y.t5 VDD.t3022 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1659 VSS.t687 B7.t16 a_n23960_n23839.t1 VSS.t686 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1660 MULT_0.NAND2_10.Y.t0 A2.t18 VDD.t524 VDD.t523 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1661 VSS.t1479 MULT_0.4bit_ADDER_1.A0.t8 a_n10108_n8419.t5 VSS.t1478 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1662 VSS.t1633 B6.t19 left_shifter_0.buffer_2.inv_1.A.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1663 a_n11274_n23075.t4 B3.t20 XOR8_0.S3.t8 VSS.t1110 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1664 right_shifter_0.S4.t2 right_shifter_0.buffer_3.inv_1.A.t6 VDD.t681 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1665 a_n9125_n7799.t1 a_n9305_n8419.t4 MULT_0.S2.t5 VDD.t1042 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1666 mux8_4.A1.t7 a_n9305_n11683.t5 a_n9125_n11063.t7 VDD.t2733 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1667 mux8_6.NAND4F_2.Y.t3 OR8_0.S7.t5 a_8592_n34534.t0 VSS.t127 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1668 a_n17677_n19625.t8 B3.t21 VDD.t2161 VDD.t2160 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1669 VDD.t900 B5.t11 right_shifter_0.buffer_3.inv_1.A.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1670 VSS.t1059 a_n20587_n5180.t3 a_n20557_n5154.t4 VSS.t1058 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1671 a_n10684_n8419.t2 a_n10714_n8445.t3 VSS.t666 VSS.t665 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1672 a_n9125_n8419.t2 a_n9155_n8445.t3 VSS.t602 VSS.t601 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1673 MULT_0.4bit_ADDER_2.B2.t1 a_n19178_n8419.t3 a_n18998_n7799.t0 VDD.t275 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1674 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t1 a_n14257_3190.t4 a_n14077_3810.t7 VDD.t1613 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1675 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t2 a_n10864_n5154.t4 a_n10684_n5154.t4 VSS.t549 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1676 MULT_0.S1.t7 a_n9305_n5154.t5 a_n9125_n5154.t4 VSS.t171 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1677 VDD.t1647 MULT_0.S2.t12 mux8_3.NAND4F_0.Y.t0 VDD.t1646 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1678 VDD.t901 B5.t12 left_shifter_0.buffer_3.inv_1.A.t2 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1679 left_shifter_0.S0.t2 VDD.t3111 VDD.t3112 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1680 a_n18072_1380.t1 A5.t13 VDD.t392 VDD.t391 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1681 a_n20557_n4534.t9 a_n20587_n5180.t4 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t8 VDD.t2034 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1682 MULT_0.4bit_ADDER_2.B2.t2 a_n19178_n8419.t4 a_n18998_n8419.t1 VSS.t125 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1683 a_n914_3810.t8 B0.t18 VDD.t994 VDD.t993 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1684 a_n1588_1406.t4 a_n1618_1380.t5 VSS.t623 VSS.t622 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X1685 mux8_2.inv_0.A.t4 mux8_2.NAND4F_9.Y.t10 a_11865_n7203.t6 VDD.t2114 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1686 mux8_3.inv_0.A.t3 mux8_3.NAND4F_9.Y.t11 a_11865_n11831.t7 VDD.t2617 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1687 VDD.t1869 mux8_4.NAND4F_1.Y.t9 mux8_4.NAND4F_9.Y.t7 VDD.t1868 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1688 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t4 a_n3659_3164.t3 a_n4205_3810.t3 VDD.t1198 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1689 a_n20446_n2915.t0 B0.t19 VSS.t503 VSS.t502 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1690 VDD.t4423 SEL1.t63 mux8_4.NAND4F_2.Y.t6 VDD.t4422 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1691 VDD.t3751 SEL2.t42 mux8_3.NAND4F_6.Y.t1 VDD.t3750 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1692 a_n13399_n8419.t2 MULT_0.4bit_ADDER_1.A1.t8 VSS.t45 VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1693 a_11386_n11894.t1 mux8_3.NAND4F_2.Y.t9 a_11290_n11894.t1 VSS.t612 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1694 a_10267_n25478.t1 mux8_7.NAND4F_2.D.t7 VSS.t1459 VSS.t1458 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1695 VDD.t394 A5.t14 AND8_0.NOT8_0.A5.t5 VDD.t393 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1696 OR8_0.S0.t1 OR8_0.NOT8_0.A0.t8 VDD.t312 VDD.t311 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1697 mux8_8.NAND4F_6.Y.t7 SEL0.t68 VDD.t3021 VDD.t3020 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1698 mux8_6.NAND4F_2.Y.t4 OR8_0.S7.t6 VDD.t1225 VDD.t1224 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1699 VDD.t2350 B1.t25 MULT_0.NAND2_5.Y.t1 VDD.t2349 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1700 VDD.t2660 mux8_8.NAND4F_0.C.t8 mux8_8.NAND4F_7.Y.t2 VDD.t2659 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1701 VDD.t3205 mux8_2.NAND4F_0.C.t7 mux8_2.NAND4F_3.Y.t0 VDD.t3204 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1702 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t4 MULT_0.4bit_ADDER_1.B1.t15 VDD.t3270 VDD.t3269 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1703 a_n14005_n11709.t1 MULT_0.inv_9.Y.t12 VDD.t4015 VDD.t4014 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1704 a_n17677_n18225.t7 B2.t17 VDD.t2597 VDD.t2596 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X1705 OR8_0.NOT8_0.A0.t2 A0.t15 a_n17677_n15425.t2 VDD.t1671 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1706 VSS.t1699 a_n24130_3190.t5 a_n23374_3190.t1 VSS.t1698 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1707 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t7 a_n14931_1406.t4 a_n14751_2026.t4 VDD.t3375 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1708 a_n19081_373.t0 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t7 VSS.t778 VSS.t777 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1709 a_n12416_n5154.t5 a_n12446_n5180.t3 VSS.t1538 VSS.t1537 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1710 mux8_8.NAND4F_4.Y.t4 mux8_8.NAND4F_2.D.t10 VDD.t1512 VDD.t1511 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1711 VDD.t3632 mux8_5.NAND4F_0.C.t9 mux8_5.NAND4F_0.Y.t1 VDD.t3631 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1712 mux8_3.NAND4F_1.Y.t5 mux8_3.NAND4F_4.B.t8 VDD.t2528 VDD.t2527 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1713 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t16 VDD.t3386 VDD.t3385 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1714 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t7 a_n20113_3164.t5 a_n20659_3810.t10 VDD.t2688 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1715 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t3 a_n20737_n5154.t7 a_n20557_n4534.t5 VDD.t746 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1716 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t2 a_n1768_1406.t5 a_n1588_2026.t4 VDD.t581 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1717 VDD.t3991 XOR8_0.S6.t13 mux8_8.NAND4F_1.Y.t4 VDD.t3990 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1718 a_16143_n18523.t3 Y2.t4 a_15855_n18523.t5 VDD.t1529 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X1719 right_shifter_0.S4.t1 right_shifter_0.buffer_3.inv_1.A.t7 VDD.t682 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1720 VDD.t755 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t18 a_n3320_2026.t2 VDD.t754 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1721 a_n6641_1380.t0 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t10 VSS.t39 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1722 VDD.t812 MULT_0.inv_12.A.t8 MULT_0.4bit_ADDER_1.A2.t1 VDD.t811 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1723 VDD.t3116 mux8_3.NAND4F_2.Y.t10 mux8_3.NAND4F_8.Y.t7 VDD.t3115 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1724 VSS.t1070 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t15 a_n9305_n5154.t0 VSS.t1069 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1725 VSS.t47 MULT_0.4bit_ADDER_1.A1.t9 a_n13399_n8419.t1 VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1726 VSS.t522 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t17 a_n19178_n8419.t0 VSS.t521 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1727 a_4069_4914.t2 SEL3.t34 V_FLAG_0.XOR2_2.Y.t2 VSS.t893 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1728 VDD.t2697 mux8_5.NAND4F_1.Y.t9 mux8_5.NAND4F_9.Y.t7 VDD.t2696 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1729 MULT_0.NAND2_1.Y.t6 B0.t20 VDD.t996 VDD.t995 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1730 a_n20587_n8445.t1 MULT_0.4bit_ADDER_1.A3.t9 VDD.t4311 VDD.t4310 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1731 a_n9155_n11709.t0 VSS.t1011 VSS.t1013 VSS.t1012 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1732 a_10363_n30006.t0 mux8_8.NAND4F_0.C.t9 a_10267_n30006.t0 VSS.t1319 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1733 a_547_1406.t4 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t17 8bit_ADDER_0.S0.t9 VSS.t1142 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1734 mux8_2.NAND4F_0.Y.t5 mux8_2.NAND4F_2.D.t7 VDD.t3171 VDD.t3170 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1735 VDD.t2015 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t18 a_n12596_n11683.t1 VDD.t2014 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X1736 mux8_0.NAND4F_8.Y.t7 mux8_0.NAND4F_4.Y.t10 VDD.t2208 VDD.t2207 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1737 VDD.t1371 mux8_5.NAND4F_2.D.t6 mux8_5.NAND4F_4.Y.t6 VDD.t1370 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1738 a_7644_n17350.t1 mux8_4.NAND4F_4.B.t10 a_7548_n17350.t0 VSS.t1544 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1739 a_n19198_1406.t4 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t15 mux8_8.A0.t4 VSS.t1206 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1740 VSS.t1262 MULT_0.4bit_ADDER_1.B0.t18 a_n10864_n8419.t0 VSS.t1261 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1741 VDD.t2163 B3.t22 AND8_0.NOT8_0.A3.t2 VDD.t2162 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1742 a_n17368_3810.t2 SEL3.t35 VDD.t1774 VDD.t1773 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1743 OR8_0.NOT8_0.A5.t0 B5.t13 VSS.t445 VSS.t177 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1744 a_9528_n21878.t0 mux8_5.NAND4F_4.B.t6 a_9432_n21878.t1 VSS.t1033 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1745 mux8_4.NAND4F_0.Y.t7 SEL0.t69 VDD.t3019 VDD.t3018 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1746 VSS.t1574 A7.t18 a_n24048_1406.t1 VSS.t1573 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1747 a_n15131_n8419.t4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t10 VSS.t1682 VSS.t1681 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1748 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t16 VDD.t669 VDD.t668 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1749 VDD.t1776 SEL3.t36 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t1 VDD.t1775 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1750 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t5 a_n20737_n8419.t4 a_n20557_n7799.t9 VDD.t2859 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1751 a_n20296_n9452.t0 MULT_0.4bit_ADDER_1.B3.t13 VSS.t1337 VSS.t1336 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1752 mux8_8.NAND4F_8.Y.t4 mux8_8.NAND4F_2.Y.t10 VDD.t1163 VDD.t1162 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1753 VDD.t3339 mux8_6.A1.t7 mux8_6.NAND4F_0.Y.t6 VDD.t3338 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1754 a_n12347_n14753.t1 A0.t16 VDD.t1673 VDD.t1672 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1755 VSS.t458 a_n1094_3190.t4 a_n338_3190.t1 VSS.t457 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1756 VDD.t4425 SEL1.t64 mux8_7.NAND4F_2.Y.t3 VDD.t4424 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1757 left_shifter_0.buffer_2.inv_1.A.t2 B6.t20 VDD.t3547 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1758 mux8_7.NAND4F_2.D.t2 SEL2.t43 VDD.t3752 VDD.t3708 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1759 8bit_ADDER_0.S0.t4 a_n209_1406.t4 a_n29_2026.t4 VDD.t3120 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1760 a_11386_n34534.t1 mux8_6.NAND4F_2.Y.t9 a_11290_n34534.t0 VSS.t123 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1761 ZFLAG_0.NAND2_0.Y.t1 ZFLAG_0.nor4_0.Y.t8 VDD.t2424 VDD.t2423 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1762 a_n11276_n15299.t0 a_n12347_n14753.t3 VSS.t570 VSS.t569 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1763 right_shifter_0.buffer_5.inv_1.A.t2 B3.t23 VDD.t2164 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1764 a_n18042_2026.t10 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t13 VDD.t2875 VDD.t2874 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1765 right_shifter_0.S0.t2 right_shifter_0.buffer_7.inv_1.A.t6 VDD.t364 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1766 VDD.t935 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t12 a_n18998_n11063.t0 VDD.t934 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1767 VDD.t1139 right_shifter_0.S2.t4 mux8_3.NAND4F_6.Y.t4 VDD.t1138 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1768 VDD.t1945 VSS.t2052 mux8_0.NAND4F_0.Y.t4 VDD.t1944 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1769 a_n9901_2026.t4 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t12 VDD.t1732 VDD.t1731 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1770 VDD.t2740 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t14 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t6 VDD.t2739 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1771 VSS.t1880 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t16 a_n12596_n5154.t0 VSS.t1879 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1772 MULT_0.NAND2_8.Y.t2 A0.t17 VDD.t1675 VDD.t1674 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1773 VDD.t2101 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t3 VDD.t2100 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1774 a_n20557_n11063.t2 MULT_0.4bit_ADDER_2.B3.t12 VDD.t4055 VDD.t4054 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1775 left_shifter_0.S4.t3 left_shifter_0.buffer_5.inv_1.A.t4 VDD.t2551 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1776 a_n16483_2026.t7 a_n16513_1380.t4 mux8_7.A0.t7 VDD.t1484 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1777 mux8_4.NAND4F_8.Y.t0 mux8_4.NAND4F_3.Y.t11 VDD.t1891 VDD.t1890 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1778 mux8_6.A0.t7 a_n23245_1406.t4 a_n23065_1406.t4 VSS.t1257 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1779 VDD.t2542 mux8_7.inv_0.A.t8 Y5.t3 VDD.t2541 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1780 a_n10684_n7799.t2 a_n10714_n8445.t4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t5 VDD.t1080 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1781 VSS.t966 MULT_0.4bit_ADDER_2.B0.t17 a_n10864_n11683.t1 VSS.t965 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1782 VDD.t1443 mux8_8.NAND4F_1.Y.t9 mux8_8.NAND4F_9.Y.t5 VDD.t1442 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1783 VDD.t2766 mux8_6.NAND4F_2.Y.t10 mux8_6.NAND4F_8.Y.t7 VDD.t2765 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1784 a_n4205_3810.t7 SEL3.t37 VDD.t1778 VDD.t1777 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1785 VSS.t336 mux8_5.NAND4F_9.Y.t11 mux8_5.inv_0.A.t6 VSS.t335 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X1786 VDD.t3303 mux8_6.A0.t17 a_5197_5532.t7 VDD.t3302 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1787 a_n6611_2026.t9 a_n6641_1380.t5 8bit_ADDER_0.S2.t2 VDD.t885 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1788 mux8_2.NAND4F_4.Y.t7 mux8_2.NAND4F_4.B.t6 VDD.t3217 VDD.t3216 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1789 VSS.t895 SEL3.t38 a_n24130_3190.t0 VSS.t894 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1790 a_3463_4888.t1 V_FLAG_0.XOR2_2.B.t16 VDD.t979 VDD.t978 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1791 VDD.t4426 SEL1.t65 mux8_7.NAND4F_0.C.t1 VDD.t4345 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1792 a_n18305_n9452.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t8 VSS.t68 VSS.t67 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1793 VDD.t3754 SEL2.t44 mux8_1.NAND4F_7.Y.t0 VDD.t3753 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1794 VDD.t4057 MULT_0.4bit_ADDER_2.B3.t13 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t1 VDD.t4056 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1795 a_7452_n20950.t0 mux8_5.NAND4F_2.D.t7 VSS.t678 VSS.t677 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1796 VSS.t1034 right_shifter_0.buffer_0.inv_1.A.t4 right_shifter_0.S1.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1797 mux8_7.NAND4F_0.Y.t5 SEL0.t70 VDD.t3017 VDD.t3016 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1798 VDD.t4428 SEL1.t66 mux8_4.NAND4F_6.Y.t6 VDD.t4427 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1799 VDD.t350 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t19 a_n13372_1406.t1 VDD.t349 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X1800 mux8_4.NAND4F_7.Y.t8 mux8_4.NAND4F_0.C.t10 VDD.t3257 VDD.t3256 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1801 a_n15907_1406.t3 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t10 VSS.t1353 VSS.t1352 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1802 a_n1327_373.t0 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t15 VSS.t1078 VSS.t840 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1803 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t10 a_n14005_n8445.t6 a_n13975_n7799.t10 VDD.t3621 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1804 AND8_0.S7.t3 AND8_0.NOT8_0.A7.t7 VDD.t3485 VDD.t3484 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1805 a_n23065_2026.t7 a_n23095_1380.t5 mux8_6.A0.t4 VDD.t1618 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1806 VDD.t873 AND8_0.S4.t4 mux8_5.NAND4F_4.Y.t2 VDD.t872 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1807 right_shifter_0.buffer_5.inv_1.A.t1 B3.t24 VDD.t2165 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1808 a_n2744_1406.t4 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t14 VSS.t1303 VSS.t1302 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1809 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t0 a_n14155_n8419.t4 a_n13975_n8419.t2 VSS.t1688 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1810 right_shifter_0.S0.t3 right_shifter_0.buffer_7.inv_1.A.t7 VDD.t366 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1811 mux8_1.NAND4F_0.Y.t0 MULT_0.SO.t4 VDD.t97 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1812 VDD.t937 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t13 a_n18998_n11063.t1 VDD.t936 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X1813 VDD.t2167 B3.t25 a_n17677_n19625.t7 VDD.t2166 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1814 a_n13399_n5154.t4 MULT_0.4bit_ADDER_0.B1.t7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t2 VSS.t654 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1815 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t9 a_n14155_n11683.t5 a_n13975_n11063.t1 VDD.t2023 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1816 VSS.t1239 MULT_0.inv_14.Y.t6 a_n16690_n11683.t5 VSS.t1238 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1817 a_7548_1690.t1 SEL1.t67 a_7452_1690.t1 VSS.t1970 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1818 VSS.t1517 a_n17548_3190.t3 a_n16792_3190.t5 VSS.t1516 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1819 right_shifter_0.buffer_3.inv_1.A.t2 B5.t14 VDD.t902 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1820 a_n17266_n11063.t2 MULT_0.4bit_ADDER_2.B2.t17 VDD.t157 VDD.t156 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1821 mux8_4.NAND4F_8.Y.t5 mux8_4.NAND4F_0.Y.t10 VDD.t796 VDD.t795 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1822 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t5 MULT_0.4bit_ADDER_0.A0.t8 VDD.t1296 VDD.t1295 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1823 VDD.t3015 SEL0.t71 mux8_3.NAND4F_2.Y.t8 VDD.t3014 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1824 a_n19981_n11683.t0 MULT_0.4bit_ADDER_2.B3.t14 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t11 VSS.t1827 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1825 a_7644_n30934.t0 mux8_8.NAND4F_4.B.t9 a_7548_n30934.t0 VSS.t1466 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1826 AND8_0.NOT8_0.A5.t1 B5.t15 VDD.t904 VDD.t903 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1827 a_n11460_2026.t7 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t19 VDD.t618 VDD.t617 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1828 a_n12416_n11683.t5 a_n12596_n11683.t6 mux8_5.A1.t10 VSS.t617 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1829 VSS.t782 a_n12347_n33735.t3 a_n11276_n34281.t1 VSS.t781 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1830 VSS.t1892 a_n4385_3190.t5 a_n3629_3190.t0 VSS.t1891 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1831 a_n15707_n7799.t9 a_n15737_n8445.t6 MULT_0.4bit_ADDER_2.B1.t9 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1832 VDD.t2169 B3.t26 a_n10786_3810.t10 VDD.t2168 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1833 mux8_7.NAND4F_8.Y.t6 mux8_7.NAND4F_3.Y.t11 VDD.t2550 VDD.t2549 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1834 VDD.t4430 SEL1.t68 mux8_5.NAND4F_6.Y.t4 VDD.t4429 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1835 VSS.t446 B5.t16 NOT8_0.S5.t1 VSS.t223 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1836 mux8_7.A1.t1 a_n15887_n11683.t4 a_n15707_n11683.t2 VSS.t795 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1837 mux8_5.NAND4F_7.Y.t2 mux8_5.NAND4F_0.C.t10 VDD.t3634 VDD.t3633 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1838 left_shifter_0.S6.t3 left_shifter_0.buffer_3.inv_1.A.t4 VDD.t815 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1839 VDD.t252 MULT_0.4bit_ADDER_0.A2.t12 a_n17266_n4534.t0 VDD.t251 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1840 a_n15707_n8419.t1 a_n15887_n8419.t4 MULT_0.4bit_ADDER_2.B1.t4 VSS.t710 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1841 VDD.t3207 mux8_2.NAND4F_0.C.t8 mux8_2.NAND4F_1.Y.t6 VDD.t3206 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1842 VDD.t21 MULT_0.4bit_ADDER_1.A2.t9 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t1 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1843 a_n10786_3810.t2 SEL3.t39 VDD.t1780 VDD.t1779 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1844 VSS.t547 mux8_8.NAND4F_9.Y.t12 mux8_8.inv_0.A.t5 VSS.t546 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X1845 a_n17677_n15425.t1 A0.t18 OR8_0.NOT8_0.A0.t1 VDD.t1676 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1846 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t9 a_n17548_3190.t4 a_n17368_3810.t9 VDD.t1142 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1847 mux8_1.NAND4F_2.Y.t8 SEL0.t72 VDD.t3013 VDD.t3012 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1848 VDD.t933 mux8_1.NAND4F_3.Y.t10 mux8_1.NAND4F_8.Y.t4 VDD.t932 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1849 MULT_0.4bit_ADDER_1.B1.t8 a_n15887_n5154.t3 a_n15707_n5154.t2 VSS.t1154 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1850 mux8_5.NAND4F_3.Y.t3 mux8_5.NAND4F_2.D.t8 VDD.t1373 VDD.t1372 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1851 mux8_0.NAND4F_0.Y.t2 VSS.t1010 a_10459_1690.t0 VSS.t1002 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1852 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t0 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t7 a_n19081_373.t1 VSS.t777 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1853 a_9432_n17350.t0 mux8_4.NAND4F_0.C.t11 a_9336_n17350.t1 VSS.t1496 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1854 a_n4879_1406.t3 a_n4909_1380.t4 VSS.t593 VSS.t592 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X1855 VDD.t159 MULT_0.4bit_ADDER_2.B2.t18 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t0 VDD.t158 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1856 VDD.t4431 SEL1.t69 mux8_6.NAND4F_0.C.t1 VDD.t4347 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1857 a_n17677_n22425.t3 B5.t17 VDD.t3962 VDD.t3961 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1858 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t5 a_n6950_3164.t3 a_n7496_3810.t8 VDD.t3985 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1859 VSS.t2031 VDD.t4515 right_shifter_0.S7.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1860 VSS.t1111 B3.t27 NOT8_0.S3.t3 VSS.t223 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1861 VSS.t355 OR8_0.NOT8_0.A3.t8 OR8_0.S3.t0 VSS.t172 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1862 a_8592_n26406.t1 SEL0.t73 a_8496_n26406.t1 VSS.t1989 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1863 a_10363_n26405.t0 mux8_7.NAND4F_0.C.t12 a_10267_n26405.t1 VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1864 VSS.t897 SEL3.t40 a_n914_3190.t1 VSS.t896 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1865 mux8_4.A0.t8 a_n10081_1406.t5 a_n9901_2026.t10 VDD.t1565 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1866 VSS.t195 right_shifter_0.buffer_4.inv_1.A.t4 right_shifter_0.S3.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1867 VDD.t1678 A0.t19 a_n1588_2026.t2 VDD.t1677 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X1868 a_n9125_n11063.t0 a_n9155_n11709.t2 mux8_4.A1.t0 VDD.t905 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1869 VSS.t689 B7.t17 a_n12347_n34023.t0 VSS.t688 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1870 right_shifter_0.buffer_3.inv_1.A.t1 B5.t18 VDD.t3963 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1871 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t18 VDD.t602 VDD.t601 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1872 a_n11274_n21072.t1 a_n12345_n20526.t5 VSS.t1214 VSS.t1213 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X1873 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t9 a_n23404_3164.t5 a_n23950_3810.t10 VDD.t2412 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1874 mux8_3.NAND4F_4.Y.t8 mux8_3.NAND4F_2.D.t11 VDD.t2807 VDD.t2806 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1875 mux8_7.NAND4F_5.Y.t4 SEL1.t70 VDD.t4433 VDD.t4432 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1876 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t1 a_n5059_1406.t5 a_n4879_2026.t0 VDD.t799 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1877 VDD.t1256 mux8_0.NAND4F_5.Y.t10 mux8_0.NAND4F_9.Y.t2 VDD.t1255 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X1878 MULT_0.NAND2_2.Y.t5 A1.t21 VDD.t4213 VDD.t4212 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1879 VDD.t2461 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t15 a_n6611_2026.t4 VDD.t2460 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1880 a_n17677_n21025.t2 B4.t19 VDD.t3599 VDD.t3598 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X1881 a_5197_4912.t4 a_5167_4886.t5 VSS.t1855 VSS.t1854 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X1882 VDD.t1734 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t13 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t3 VDD.t1733 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1883 VDD.t2622 MULT_0.NAND2_11.Y.t9 MULT_0.4bit_ADDER_0.A3.t2 VDD.t2620 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1884 mux8_7.NAND4F_8.Y.t3 mux8_7.NAND4F_0.Y.t10 VDD.t957 VDD.t956 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1885 a_8400_n25478.t1 mux8_7.NAND4F_2.D.t8 VSS.t1461 VSS.t1460 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1886 mux8_4.NAND4F_9.Y.t8 mux8_4.NAND4F_1.Y.t10 VDD.t1871 VDD.t1870 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1887 VDD.t1782 SEL3.t41 a_3313_4914.t1 VDD.t1781 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X1888 mux8_3.NAND4F_6.Y.t0 SEL2.t45 VDD.t3756 VDD.t3755 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1889 VDD.t314 OR8_0.NOT8_0.A0.t9 OR8_0.S0.t2 VDD.t313 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1890 a_n12314_n31661.t8 a_n12345_n31115.t3 XOR8_0.S6.t9 VDD.t2639 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1891 a_n17296_n5180.t0 MULT_0.4bit_ADDER_0.A2.t13 VSS.t117 VSS.t116 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1892 VDD.t4435 SEL1.t71 mux8_8.NAND4F_6.Y.t6 VDD.t4434 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1893 VDD.t3011 SEL0.t74 mux8_6.NAND4F_2.Y.t8 VDD.t3010 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1894 mux8_8.NAND4F_7.Y.t3 mux8_8.NAND4F_0.C.t10 VDD.t2662 VDD.t2661 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1895 VDD.t3757 SEL2.t46 mux8_7.NAND4F_2.D.t1 VDD.t3708 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1896 mux8_7.A0.t2 a_n16663_1406.t4 a_n16483_1406.t1 VSS.t65 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1897 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t10 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t20 a_n14175_1406.t4 VSS.t703 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1898 a_n24162_n7992.t1 A0.t20 VSS.t839 VSS.t838 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1899 a_n13222_1380.t1 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t15 VDD.t3949 VDD.t3948 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1900 a_n20757_1406.t1 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t15 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t1 VSS.t1491 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1901 8bit_ADDER_0.S2.t11 a_n6791_1406.t4 a_n6611_1406.t5 VSS.t1557 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1902 VSS.t1902 A1.t22 a_n4303_1406.t4 VSS.t1901 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1903 mux8_7.NAND4F_3.Y.t2 mux8_7.A0.t13 a_9528_n25478.t0 VSS.t296 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1904 VDD.t526 A2.t19 a_n12314_n21072.t2 VDD.t525 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X1905 VDD.t1943 VSS.t2053 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t6 VDD.t1942 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1906 OR8_0.S5.t1 OR8_0.NOT8_0.A5.t9 VDD.t2279 VDD.t315 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1907 mux8_5.NAND4F_0.Y.t0 mux8_5.NAND4F_0.C.t11 VDD.t3636 VDD.t3635 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1908 a_n12446_n11709.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t12 VSS.t1372 VSS.t1371 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1909 a_n13975_n5154.t1 a_n14005_n5180.t5 VSS.t753 VSS.t752 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X1910 VDD.t2599 B2.t18 MULT_0.inv_6.A.t2 VDD.t2598 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1911 VSS.t308 a_n12345_n25873.t3 a_n11274_n26419.t1 VSS.t307 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1912 a_15855_n18523.t4 Y2.t5 a_16143_n18523.t4 VDD.t1530 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X1913 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t6 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t9 VDD.t4049 VDD.t4048 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1914 mux8_3.NAND4F_8.Y.t8 mux8_3.NAND4F_2.Y.t11 VDD.t3118 VDD.t3117 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1915 a_8592_n35462.t1 SEL0.t75 a_8496_n35462.t1 VSS.t2009 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1916 a_n17368_3190.t4 B5.t19 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t7 VSS.t1796 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1917 VDD.t1087 MULT_0.inv_6.A.t8 MULT_0.4bit_ADDER_1.A0.t1 VDD.t1086 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1918 a_10363_n35461.t0 mux8_6.NAND4F_0.C.t10 a_10267_n35461.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1919 VSS.t1290 B2.t19 a_n24007_n17714.t1 VSS.t1289 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1920 mux8_5.NAND4F_9.Y.t8 mux8_5.NAND4F_1.Y.t10 VDD.t2699 VDD.t2698 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1921 mux8_5.NAND4F_3.Y.t7 mux8_5.A0.t13 VDD.t3350 VDD.t3349 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1922 mux8_2.NAND4F_5.Y.t5 mux8_2.NAND4F_4.B.t7 VDD.t3219 VDD.t3218 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1923 a_10267_n30006.t1 mux8_8.NAND4F_2.D.t11 VSS.t741 VSS.t740 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1924 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t2 B7.t18 a_n23950_3190.t5 VSS.t690 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1925 VDD.t3297 mux8_0.inv_0.A.t10 C.t1 VDD.t3296 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1926 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t18 VDD.t3888 VDD.t3887 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1927 mux8_3.NAND4F_4.Y.t2 AND8_0.S2.t6 a_7644_n11894.t0 VSS.t208 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1928 AND8_0.NOT8_0.A4.t1 B4.t20 VDD.t3601 VDD.t3600 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1929 MULT_0.NAND2_14.Y.t4 B3.t28 VDD.t2171 VDD.t2170 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1930 VDD.t1680 A0.t21 a_n12316_n15299.t0 VDD.t1679 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1931 a_n13975_n7799.t6 MULT_0.4bit_ADDER_1.B1.t16 VDD.t3272 VDD.t3271 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1932 a_7452_n8194.t0 SEL2.t47 VSS.t1721 VSS.t1476 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1933 a_7548_n17350.t1 SEL1.t72 a_7452_n17350.t1 VSS.t1953 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1934 mux8_0.NAND4F_8.Y.t8 mux8_0.NAND4F_4.Y.t11 a_11386_1690.t1 VSS.t626 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1935 mux8_6.NAND4F_5.Y.t5 SEL1.t73 VDD.t4437 VDD.t4436 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1936 mux8_4.NAND4F_9.Y.t6 mux8_4.NAND4F_7.Y.t9 VDD.t4168 VDD.t4167 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1937 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t5 MULT_0.4bit_ADDER_1.A3.t10 VDD.t4250 VDD.t4249 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1938 a_n914_3810.t4 a_n1094_3190.t5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t1 VDD.t919 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1939 mux8_5.A0.t7 a_n13372_1406.t5 a_n13192_2026.t11 VDD.t2747 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1940 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t4 a_n11490_1380.t5 a_n11460_2026.t1 VDD.t954 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1941 a_n8170_2026.t2 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t15 VDD.t879 VDD.t878 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1942 VDD.t1736 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t14 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t2 VDD.t1735 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1943 a_n12314_n29052.t6 a_n12345_n28794.t4 XOR8_0.S5.t5 VDD.t1459 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1944 VSS.t755 a_n14005_n5180.t6 a_n13975_n5154.t2 VSS.t754 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1945 VDD.t4328 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t9 MULT_0.4bit_ADDER_1.B3.t5 VDD.t4327 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1946 mux8_6.NAND4F_4.Y.t1 mux8_6.NAND4F_2.D.t11 VDD.t430 VDD.t429 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1947 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t3 A0.t22 a_n1327_373.t1 VSS.t840 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1948 a_9432_n30934.t1 mux8_8.NAND4F_0.C.t11 a_9336_n30934.t1 VSS.t1320 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1949 a_n23095_1380.t1 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t10 VDD.t1877 VDD.t1876 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1950 a_n17266_n7799.t10 MULT_0.4bit_ADDER_1.A2.t10 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1951 a_11290_n26406.t0 mux8_7.NAND4F_1.Y.t11 a_11194_n26406.t1 VSS.t1272 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1952 a_n7496_3810.t1 SEL3.t42 VDD.t1784 VDD.t1783 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1953 a_n19028_n5180.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t11 VSS.t1280 VSS.t1279 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X1954 a_10363_n7266.t0 mux8_2.NAND4F_0.C.t9 a_10267_n7266.t1 VSS.t1487 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1955 a_n16690_n8419.t2 MULT_0.4bit_ADDER_1.B2.t17 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t10 VSS.t1818 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1956 mux8_1.NAND4F_6.Y.t8 SEL0.t76 VDD.t3009 VDD.t3008 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1957 VDD.t1309 mux8_1.NAND4F_1.Y.t11 mux8_1.NAND4F_9.Y.t5 VDD.t1308 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1958 VDD.t3758 SEL2.t48 mux8_6.NAND4F_2.D.t1 VDD.t3714 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1959 VSS.t1074 left_shifter_0.buffer_4.inv_1.A.t5 left_shifter_0.S5.t1 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1960 VDD.t671 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t17 a_n15707_n7799.t1 VDD.t670 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1961 VSS.t1652 B4.t21 a_n12345_n26161.t0 VSS.t1651 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X1962 VSS.t1291 B2.t20 left_shifter_0.buffer_0.inv_1.A.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1963 VSS.t1838 A3.t23 a_n10884_1406.t2 VSS.t1837 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1964 a_n10714_n11709.t1 MULT_0.inv_8.Y.t9 VDD.t3519 VDD.t3518 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X1965 OR8_0.NOT8_0.A6.t2 A6.t13 a_n17677_n23825.t4 VDD.t2821 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1966 a_n17266_n4534.t7 a_n17446_n5154.t5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t6 VDD.t2428 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1967 VDD.t3903 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t15 a_n16663_1406.t1 VDD.t3902 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X1968 a_n18998_n11063.t2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t14 VDD.t939 VDD.t938 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1969 mux8_3.NAND4F_6.Y.t3 right_shifter_0.S2.t5 VDD.t1141 VDD.t1140 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1970 a_n19198_1406.t2 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t10 VSS.t551 VSS.t550 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1971 VDD.t440 MULT_0.NAND2_10.Y.t8 MULT_0.4bit_ADDER_0.A2.t1 VDD.t439 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1972 a_n15707_n5154.t3 a_n15737_n5180.t7 VSS.t463 VSS.t462 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X1973 VDD.t1682 A0.t23 MULT_0.NAND2_8.Y.t1 VDD.t1681 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1974 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t8 VDD.t2103 VDD.t2102 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1975 mux8_5.NAND4F_9.Y.t4 mux8_5.NAND4F_7.Y.t9 VDD.t233 VDD.t232 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X1976 VDD.t4159 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t14 a_n18998_n7799.t9 VDD.t4158 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X1977 VDD.t2552 left_shifter_0.buffer_5.inv_1.A.t5 left_shifter_0.S4.t2 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1978 VDD.t3760 SEL2.t49 mux8_0.NAND4F_7.Y.t1 VDD.t3759 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1979 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t7 MULT_0.4bit_ADDER_0.B0.t9 a_n10108_n5154.t4 VSS.t132 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1980 MULT_0.S1.t4 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t16 a_n8549_n5154.t4 VSS.t1071 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1981 VDD.t2486 mux8_4.NAND4F_0.Y.t11 mux8_4.NAND4F_8.Y.t4 VDD.t2485 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1982 MULT_0.4bit_ADDER_2.B2.t7 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t18 a_n18422_n8419.t1 VSS.t523 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1983 VDD.t3761 SEL2.t50 mux8_0.NAND4F_2.D.t2 VDD.t3727 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1984 VDD.t39 mux8_2.NAND4F_8.Y.t12 a_11865_n7203.t1 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X1985 VDD.t2686 MULT_0.NAND2_15.Y.t9 MULT_0.inv_15.Y.t1 VDD.t2683 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1986 mux8_8.NAND4F_9.Y.t6 mux8_8.NAND4F_1.Y.t10 VDD.t1445 VDD.t1444 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1987 a_n9208_373.t0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t10 VSS.t955 VSS.t954 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1988 mux8_6.NAND4F_8.Y.t8 mux8_6.NAND4F_2.Y.t11 VDD.t2768 VDD.t2767 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1989 mux8_5.inv_0.A.t0 mux8_5.NAND4F_8.Y.t13 VSS.t1937 VSS.t1936 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1990 AND8_0.NOT8_0.A0.t2 B0.t21 VDD.t998 VDD.t997 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1991 a_n18422_n5154.t5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t15 MULT_0.4bit_ADDER_1.B2.t8 VSS.t1349 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1992 VDD.t4438 SEL1.t74 mux8_5.NAND4F_0.C.t2 VDD.t4355 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X1993 VDD.t3388 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t17 a_n9305_n11683.t1 VDD.t3387 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X1994 VSS.t1925 a_n20839_3190.t4 a_n20083_3190.t1 VSS.t1924 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X1995 a_n10210_3190.t1 a_n10240_3164.t5 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t3 VSS.t333 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1996 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t1 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t15 VDD.t1738 VDD.t1737 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1997 a_n23254_373.t0 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t16 VSS.t1602 VSS.t960 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1998 Y3.t1 mux8_4.inv_0.A.t8 VSS.t1597 VSS.t1596 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1999 a_7452_n16422.t0 mux8_4.NAND4F_2.D.t7 VSS.t57 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2000 a_n9155_n8445.t0 VSS.t1007 VSS.t1009 VSS.t1008 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X2001 VDD.t3763 SEL2.t51 mux8_7.NAND4F_1.Y.t1 VDD.t3762 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2002 VDD.t810 NOT8_0.S0.t6 mux8_1.NAND4F_7.Y.t6 VDD.t809 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2003 mux8_6.NAND4F_4.Y.t4 AND8_0.S7.t6 a_7644_n34534.t0 VSS.t167 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2004 VDD.t3965 B5.t20 a_n17677_n22425.t2 VDD.t3964 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2005 a_n24162_n9284.t0 B2.t21 VSS.t1293 VSS.t1292 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2006 a_n14751_2026.t6 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t21 VDD.t1428 VDD.t1427 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2007 VSS.t642 a_n12345_n17569.t3 a_n11274_n18115.t1 VSS.t641 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2008 VSS.t1795 a_n7676_3190.t6 a_n6920_3190.t0 VSS.t1794 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X2009 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t0 MULT_0.4bit_ADDER_2.B3.t15 VDD.t4059 VDD.t4058 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2010 mux8_5.NAND4F_7.Y.t4 NOT8_0.S4.t5 a_10459_n21877.t0 VSS.t674 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2011 a_n12446_n5180.t1 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t13 VDD.t216 VDD.t215 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2012 a_n12316_n34281.t11 a_n12347_n33735.t4 XOR8_0.S7.t0 VDD.t1594 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2013 VDD.t1000 B0.t22 MULT_0.NAND2_3.Y.t5 VDD.t999 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2014 a_n14077_3810.t1 SEL3.t43 VDD.t1786 VDD.t1785 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2015 a_11290_n35462.t0 mux8_6.NAND4F_1.Y.t11 a_11194_n35462.t0 VSS.t721 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2016 a_1887_5534.t1 A7.t19 VDD.t3426 VDD.t3425 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2017 mux8_5.NAND4F_4.Y.t1 AND8_0.S4.t5 VDD.t875 VDD.t874 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2018 a_n4205_3810.t1 a_n4385_3190.t6 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t1 VDD.t3952 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2019 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t10 a_n10714_n11709.t4 a_n10684_n11063.t10 VDD.t2006 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2020 MULT_0.inv_14.Y.t0 MULT_0.NAND2_14.Y.t9 VSS.t1307 VSS.t1306 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2021 VDD.t226 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t9 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t1 VDD.t225 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2022 a_n13975_n11063.t11 a_n14005_n11709.t3 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t0 VDD.t1650 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2023 a_n16690_n11683.t4 MULT_0.inv_14.Y.t7 VSS.t1241 VSS.t1240 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2024 mux8_0.NAND4F_0.Y.t6 mux8_0.NAND4F_2.D.t8 VDD.t2892 VDD.t2891 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2025 OR8_0.S7.t3 OR8_0.NOT8_0.A7.t7 VDD.t786 VDD.t785 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2026 VDD.t3507 mux8_0.NAND4F_8.Y.t12 a_11865_1753.t2 VDD.t3506 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2027 VDD.t4215 A1.t23 a_n12314_n18115.t7 VDD.t4214 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2028 a_n23065_2026.t1 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t17 VDD.t3472 VDD.t3471 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2029 VDD.t161 MULT_0.4bit_ADDER_2.B2.t19 a_n17266_n11063.t1 VDD.t160 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2030 MULT_0.4bit_ADDER_1.B0.t10 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t17 a_n11840_n5154.t4 VSS.t1881 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2031 a_n12314_n29052.t9 a_n12345_n28506.t4 XOR8_0.S5.t8 VDD.t1817 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2032 a_7548_n30934.t1 SEL1.t75 a_7452_n30934.t1 VSS.t1971 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2033 mux8_8.NAND4F_9.Y.t8 mux8_8.NAND4F_7.Y.t9 VDD.t2570 VDD.t2569 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2034 VDD.t4104 A3.t24 MULT_0.NAND2_11.Y.t4 VDD.t4103 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2035 VDD.t2388 ZFLAG_0.nor4_1.Y.t7 ZFLAG_0.NAND2_0.Y.t3 VDD.t2387 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2036 VDD.t959 mux8_7.NAND4F_0.Y.t11 mux8_7.NAND4F_8.Y.t4 VDD.t958 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2037 a_n20659_3810.t7 a_n20839_3190.t5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t4 VDD.t4277 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2038 a_n1588_2026.t10 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t16 VDD.t2089 VDD.t2088 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2039 VDD.t816 left_shifter_0.buffer_3.inv_1.A.t5 left_shifter_0.S6.t2 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2040 VSS.t1179 B1.t26 a_n12345_n17857.t0 VSS.t1178 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2041 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t9 a_n8350_1406.t5 a_n8170_2026.t6 VDD.t1518 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2042 a_n18998_n11063.t3 a_n19178_n11683.t5 mux8_8.A1.t1 VDD.t1548 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2043 mux8_8.inv_0.A.t6 mux8_8.NAND4F_8.Y.t13 VSS.t360 VSS.t359 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X2044 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t8 a_n15014_n9452.t0 VSS.t1822 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2045 a_9336_n17350.t0 SEL2.t52 VSS.t1722 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2046 a_n17266_n8419.t2 a_n17296_n8445.t4 VSS.t1508 VSS.t1507 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2047 a_n17266_n11683.t3 a_n17296_n11709.t6 VSS.t1415 VSS.t1414 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2048 VDD.t3765 SEL2.t53 mux8_6.NAND4F_1.Y.t1 VDD.t3764 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2049 VDD.t3007 SEL0.t77 mux8_7.NAND4F_4.B.t3 VDD.t2951 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2050 mux8_6.NAND4F_7.Y.t5 NOT8_0.S7.t6 VDD.t418 VDD.t417 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2051 VDD.t1219 mux8_3.NAND4F_6.Y.t9 mux8_3.NAND4F_9.Y.t3 VDD.t1218 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2052 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t7 a_n17446_n5154.t6 a_n17266_n5154.t0 VSS.t1224 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2053 VDD.t2787 mux8_4.NAND4F_4.Y.t9 mux8_4.NAND4F_8.Y.t8 VDD.t2786 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2054 a_n13192_1406.t5 a_n13222_1380.t4 VSS.t380 VSS.t379 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2055 a_n11460_1406.t4 a_n11640_1406.t4 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t8 VSS.t774 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2056 VDD.t576 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t10 MULT_0.4bit_ADDER_2.B3.t6 VDD.t575 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2057 a_n11274_n26419.t2 a_n12345_n25873.t4 VSS.t310 VSS.t309 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2058 a_8496_n26406.t0 SEL1.t76 a_8400_n26406.t1 VSS.t1951 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2059 VDD.t3603 B4.t22 a_n14077_3810.t4 VDD.t3602 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2060 mux8_8.A0.t11 a_n19954_1406.t4 a_n19774_1406.t4 VSS.t559 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2061 mux8_1.NAND4F_2.D.t2 SEL2.t54 VDD.t3766 VDD.t3729 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2062 a_10267_n26405.t0 SEL2.t55 VSS.t1723 VSS.t1458 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2063 a_n16513_1380.t1 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t11 VDD.t2753 VDD.t2752 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2064 a_n1012_1406.t3 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t17 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t9 VSS.t1079 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2065 VDD.t3670 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t11 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t5 VDD.t3669 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2066 MULT_0.NAND2_9.Y.t5 B3.t29 VDD.t2173 VDD.t2172 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2067 VSS.t250 A2.t20 a_n7594_1406.t4 VSS.t249 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2068 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t6 a_n17446_n8419.t5 a_n17266_n7799.t3 VDD.t732 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2069 VDD.t2912 MULT_0.4bit_ADDER_0.B2.t8 a_n17446_n5154.t1 VDD.t2911 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X2070 VDD.t717 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t9 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t4 VDD.t716 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2071 a_n24007_n17714.t0 A2.t21 AND8_0.NOT8_0.A2.t2 VSS.t251 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2072 left_shifter_0.buffer_6.inv_1.A.t3 B0.t23 VDD.t1001 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2073 VDD.t3768 SEL2.t56 mux8_7.NAND4F_5.Y.t1 VDD.t3767 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2074 VSS.t899 SEL3.t44 a_n14077_3190.t0 VSS.t898 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2075 mux8_5.A1.t4 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t19 a_n11840_n11683.t1 VSS.t1045 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2076 a_n29_2026.t11 a_n59_1380.t4 8bit_ADDER_0.S0.t11 VDD.t3378 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2077 a_n24363_373.t1 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t15 VSS.t1668 VSS.t1575 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2078 VDD.t3662 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t18 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t1 VDD.t3661 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2079 a_n10108_n8419.t4 MULT_0.4bit_ADDER_1.A0.t9 VSS.t1481 VSS.t1480 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2080 mux8_5.NAND4F_9.Y.t0 mux8_5.NAND4F_5.Y.t9 a_11386_n21878.t0 VSS.t577 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2081 VDD.t3769 SEL2.t57 mux8_5.NAND4F_2.D.t2 VDD.t3722 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2082 Z.t2 ZFLAG_0.NAND2_0.Y.t9 VDD.t1461 VDD.t1460 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2083 VDD.t4170 mux8_4.NAND4F_7.Y.t10 mux8_4.NAND4F_9.Y.t5 VDD.t4169 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2084 a_n12314_n26419.t0 a_n12345_n25873.t5 XOR8_0.S4.t0 VDD.t627 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2085 VDD.t2220 A0.t24 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t6 VDD.t2219 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2086 VSS.t636 MULT_0.4bit_ADDER_0.A0.t9 a_n10108_n5154.t0 VSS.t635 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X2087 a_n19774_2026.t5 a_n19804_1380.t4 mux8_8.A0.t2 VDD.t1449 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2088 VSS.t1493 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t16 a_n21513_1406.t0 VSS.t1492 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2089 a_n18998_n7799.t1 a_n19178_n8419.t5 MULT_0.4bit_ADDER_2.B2.t3 VDD.t276 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2090 VDD.t3428 A7.t20 a_n24624_2026.t4 VDD.t3427 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2091 a_n17266_n11683.t2 a_n17446_n11683.t2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t7 VSS.t647 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2092 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t4 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t8 VDD.t1583 VDD.t1582 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2093 a_n10684_n5154.t2 a_n10714_n5180.t4 VSS.t140 VSS.t139 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2094 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t5 MULT_0.inv_14.Y.t8 VDD.t2442 VDD.t2441 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2095 a_n9125_n5154.t0 a_n9155_n5180.t3 VSS.t144 VSS.t143 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2096 V_FLAG_0.XOR2_2.B.t9 a_1857_4888.t4 a_1887_5534.t10 VDD.t2770 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2097 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t7 a_n20587_n5180.t5 a_n20557_n4534.t10 VDD.t2035 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2098 a_n18998_n8419.t5 a_n19028_n8445.t3 VSS.t660 VSS.t659 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2099 a_n17677_n23825.t3 A6.t14 OR8_0.NOT8_0.A6.t1 VDD.t2822 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2100 a_n29_1406.t3 a_n59_1380.t5 VSS.t1197 VSS.t1196 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2101 a_11865_n7203.t7 mux8_2.NAND4F_9.Y.t11 mux8_2.inv_0.A.t3 VDD.t2115 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2102 a_9528_n25478.t1 mux8_7.NAND4F_4.B.t8 a_9432_n25478.t1 VSS.t92 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2103 mux8_5.NAND4F_2.Y.t5 SEL1.t77 VDD.t4440 VDD.t4439 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2104 VDD.t1409 B7.t19 a_n23950_3810.t2 VDD.t1408 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2105 a_n3350_1380.t1 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t15 VDD.t2627 VDD.t2626 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2106 MULT_0.4bit_ADDER_1.A3.t0 MULT_0.inv_13.A.t8 VSS.t1921 VSS.t1920 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2107 a_11865_n20887.t2 mux8_5.NAND4F_9.Y.t12 mux8_5.inv_0.A.t3 VDD.t688 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2108 a_n23992_n18833.t0 A3.t25 AND8_0.NOT8_0.A3.t6 VSS.t1839 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2109 MULT_0.4bit_ADDER_1.B2.t6 a_n19178_n5154.t6 a_n18998_n5154.t0 VSS.t339 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2110 VSS.t49 MULT_0.4bit_ADDER_1.A1.t10 a_n13399_n8419.t0 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2111 VDD.t3006 SEL0.t78 mux8_6.NAND4F_4.B.t3 VDD.t2949 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2112 MULT_0.4bit_ADDER_0.A2.t2 MULT_0.NAND2_10.Y.t9 VDD.t441 VDD.t439 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2113 VDD.t511 mux8_7.NAND4F_4.Y.t9 mux8_7.NAND4F_8.Y.t0 VDD.t510 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2114 AND8_0.NOT8_0.A4.t5 A4.t15 VDD.t1641 VDD.t1640 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2115 mux8_0.NAND4F_2.Y.t3 SEL1.t78 VDD.t4442 VDD.t4441 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2116 a_n13399_n5154.t2 MULT_0.4bit_ADDER_0.A1.t7 VSS.t1164 VSS.t1163 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2117 MULT_0.NAND2_5.Y.t0 B1.t27 VDD.t2352 VDD.t2351 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2118 a_8496_n35462.t0 SEL1.t79 a_8400_n35462.t1 VSS.t1972 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2119 a_n12314_n23651.t11 a_n12345_n23105.t4 XOR8_0.S3.t10 VDD.t2763 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2120 VSS.t1510 a_n17296_n8445.t5 a_n17266_n8419.t1 VSS.t1509 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2121 a_8400_n30006.t0 mux8_8.NAND4F_2.D.t12 VSS.t743 VSS.t742 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2122 a_10267_n35461.t0 SEL2.t58 VSS.t1724 VSS.t200 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2123 VDD.t1989 mux8_5.NAND4F_4.B.t7 mux8_5.NAND4F_3.Y.t4 VDD.t1988 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2124 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t4 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t8 a_n9208_373.t1 VSS.t954 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2125 VDD.t235 mux8_5.NAND4F_7.Y.t10 mux8_5.NAND4F_9.Y.t3 VDD.t234 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2126 mux8_7.A0.t11 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t16 a_n15907_1406.t1 VSS.t1773 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2127 VSS.t817 A4.t16 a_n14175_1406.t1 VSS.t816 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X2128 MULT_0.inv_8.Y.t2 MULT_0.NAND2_8.Y.t9 VDD.t727 VDD.t725 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2129 a_n19028_n11709.t1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t15 VDD.t941 VDD.t940 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2130 a_7644_n11894.t1 mux8_3.NAND4F_4.B.t9 a_7548_n11894.t0 VSS.t1269 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2131 V_FLAG_0.XOR2_2.B.t11 a_1707_4914.t4 a_1887_4914.t5 VSS.t1413 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2132 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t3 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t11 a_n23254_373.t1 VSS.t960 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2133 a_n20557_n4534.t8 VSS.t2054 VDD.t1941 VDD.t1940 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2134 VDD.t2175 B3.t30 MULT_0.NAND2_14.Y.t5 VDD.t2174 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2135 mux8_6.A0.t10 a_n23245_1406.t5 a_n23065_2026.t10 VDD.t2488 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2136 VSS.t1653 B4.t23 NOT8_0.S4.t0 VSS.t223 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2137 8bit_ADDER_0.S1.t2 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t19 a_n2744_1406.t1 VSS.t369 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2138 a_n10684_n4534.t10 a_n10864_n5154.t5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t10 VDD.t2862 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2139 VDD.t3771 SEL2.t59 mux8_6.NAND4F_5.Y.t1 VDD.t3770 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2140 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t5 A0.t25 VDD.t2222 VDD.t2221 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2141 mux8_8.NAND4F_3.Y.t4 mux8_8.A0.t13 a_9528_n30006.t1 VSS.t736 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2142 a_n12314_n31661.t4 B6.t21 VDD.t3549 VDD.t3548 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2143 VSS.t1166 MULT_0.4bit_ADDER_0.A1.t8 a_n13399_n5154.t1 VSS.t1165 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X2144 a_9336_n30934.t0 SEL2.t60 VSS.t1725 VSS.t744 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2145 XOR8_0.S7.t1 a_n12347_n33735.t5 a_n12316_n34281.t10 VDD.t1595 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2146 VDD.t2091 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t18 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t1 VDD.t2090 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2147 VDD.t1003 B0.t24 MULT_0.NAND2_1.Y.t5 VDD.t1002 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2148 VSS.t236 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t16 a_n19178_n5154.t0 VSS.t235 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2149 VDD.t1005 B0.t25 a_n914_3810.t7 VDD.t1004 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2150 VDD.t3173 mux8_2.NAND4F_2.D.t8 mux8_2.NAND4F_0.Y.t6 VDD.t3172 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2151 a_11194_n26406.t0 mux8_7.NAND4F_7.Y.t11 VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2152 VDD.t1788 SEL3.t45 a_3493_5534.t1 VDD.t1787 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2153 VDD.t1568 left_shifter_0.S5.t5 mux8_7.NAND4F_5.Y.t3 VDD.t1567 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2154 VSS.t1294 B2.t22 right_shifter_0.buffer_0.inv_1.A.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2155 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t5 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t9 VDD.t1585 VDD.t1584 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2156 VSS.t962 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t12 a_n22489_1406.t5 VSS.t961 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2157 VDD.t3672 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t12 a_n15707_n7799.t8 VDD.t3671 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2158 a_n3629_3190.t4 a_n3659_3164.t4 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t5 VSS.t604 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2159 VSS.t848 right_shifter_0.buffer_6.inv_1.A.t4 right_shifter_0.C.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2160 a_n18042_2026.t11 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t14 VDD.t2877 VDD.t2876 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2161 VDD.t1335 MULT_0.4bit_ADDER_0.B1.t8 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t5 VDD.t1334 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2162 a_n8170_1406.t3 a_n8200_1380.t5 VSS.t158 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2163 VDD.t1159 MULT_0.NAND2_0.Y.t9 MULT_0.4bit_ADDER_0.B2.t2 VDD.t1157 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2164 MULT_0.4bit_ADDER_1.B0.t0 a_n12596_n5154.t5 a_n12416_n4534.t0 VDD.t986 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2165 VSS.t1684 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t13 a_n15131_n8419.t3 VSS.t1683 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2166 VDD.t4021 mux8_4.NAND4F_5.Y.t10 mux8_4.NAND4F_9.Y.t2 VDD.t4020 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2167 VSS.t134 MULT_0.4bit_ADDER_0.B0.t10 a_n10864_n5154.t0 VSS.t133 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2168 VDD.t3005 SEL0.t79 mux8_3.NAND4F_6.Y.t8 VDD.t3004 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2169 a_n20557_n7799.t10 a_n20737_n8419.t5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t6 VDD.t2860 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2170 a_n12314_n18115.t3 a_n12345_n17569.t4 XOR8_0.S1.t1 VDD.t1303 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2171 mux8_1.NAND4F_3.Y.t0 mux8_1.NAND4F_0.C.t8 VDD.t69 VDD.t68 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2172 a_n15131_n5154.t4 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t13 VSS.t346 VSS.t345 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2173 MULT_0.4bit_ADDER_0.A1.t0 MULT_0.NAND2_5.Y.t9 VSS.t1465 VSS.t1464 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2174 VDD.t4254 mux8_7.NAND4F_8.Y.t11 a_11865_n25415.t8 VDD.t4253 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2175 XOR8_0.S5.t7 a_n12345_n28506.t5 a_n12314_n29052.t8 VDD.t1818 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2176 a_11194_n2838.t0 mux8_1.NAND4F_0.Y.t10 VSS.t1536 VSS.t651 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2177 mux8_2.inv_0.A.t2 mux8_2.NAND4F_9.Y.t12 a_11865_n7203.t8 VDD.t2116 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X2178 a_8496_n2838.t0 SEL1.t80 a_8400_n2838.t1 VSS.t1960 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2179 a_n12345_n28506.t0 A5.t15 VSS.t184 VSS.t183 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X2180 a_n15896_n12716.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t15 VSS.t631 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2181 V_FLAG_0.XOR2_0.Y.t7 a_5167_4886.t6 a_5197_5532.t4 VDD.t4123 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2182 VDD.t2572 mux8_8.NAND4F_7.Y.t10 mux8_8.NAND4F_9.Y.t7 VDD.t2571 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2183 a_n17677_n15425.t7 B0.t26 VDD.t1007 VDD.t1006 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2184 mux8_5.NAND4F_4.B.t2 SEL0.t80 VDD.t3003 VDD.t2937 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2185 VSS.t1904 A1.t24 OR8_0.NOT8_0.A1.t6 VSS.t1903 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X2186 a_n17466_1406.t2 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t15 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t9 VSS.t1428 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2187 a_n12314_n21072.t6 a_n12345_n20526.t6 XOR8_0.S2.t3 VDD.t2416 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2188 VDD.t1790 SEL3.t46 a_n24130_3190.t1 VDD.t1789 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X2189 a_n9901_2026.t8 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t19 VDD.t1555 VDD.t1554 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2190 VDD.t2224 A0.t26 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t4 VDD.t2223 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2191 mux8_7.NAND4F_1.Y.t0 SEL2.t61 VDD.t3773 VDD.t3772 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2192 a_n24624_2026.t0 a_n24804_1406.t5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t0 VDD.t3466 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2193 VDD.t4443 SEL1.t81 mux8_3.NAND4F_0.C.t1 VDD.t4373 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2194 a_7644_n34534.t1 mux8_6.NAND4F_4.B.t9 a_7548_n34534.t1 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2195 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t0 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t19 VDD.t2093 VDD.t2092 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2196 VDD.t1939 VSS.t2055 a_n20737_n5154.t1 VDD.t1938 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X2197 mux8_0.NAND4F_3.Y.t1 mux8_0.NAND4F_4.B.t10 VDD.t855 VDD.t854 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2198 VDD.t3315 MULT_0.inv_15.Y.t8 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t3 VDD.t3314 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2199 mux8_5.NAND4F_6.Y.t0 right_shifter_0.S4.t4 a_8592_n21878.t0 VSS.t87 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2200 VDD.t1154 mux8_5.NAND4F_5.Y.t10 mux8_5.NAND4F_9.Y.t2 VDD.t1153 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2201 a_10459_n21877.t1 SEL0.t81 a_10363_n21877.t1 VSS.t2000 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2202 VDD.t4106 A3.t26 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t2 VDD.t4105 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2203 a_n4879_2026.t6 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t18 VDD.t4143 VDD.t4142 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2204 VDD.t3774 SEL2.t62 mux8_1.NAND4F_2.D.t1 VDD.t3729 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2205 MULT_0.NAND2_3.Y.t0 A0.t27 a_n18686_n2915.t0 VSS.t509 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2206 VDD.t3002 SEL0.t82 mux8_3.NAND4F_4.B.t1 VDD.t3001 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2207 VSS.t633 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t16 a_n15887_n11683.t0 VSS.t632 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2208 V_FLAG_0.XOR2_0.Y.t0 a_5017_4912.t4 a_5197_4912.t1 VSS.t973 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2209 VDD.t1587 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t10 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t6 VDD.t1586 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2210 VDD.t3221 mux8_2.NAND4F_4.B.t8 mux8_2.NAND4F_4.Y.t8 VDD.t3220 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2211 a_11194_n35462.t1 mux8_6.NAND4F_7.Y.t11 VSS.t198 VSS.t197 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2212 a_n20557_n7799.t1 a_n20587_n8445.t5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t10 VDD.t2869 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2213 MULT_0.NAND2_14.Y.t6 B3.t31 a_n22425_n11256.t1 VSS.t261 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2214 a_n12316_n15299.t7 a_n12347_n15041.t5 XOR8_0.S0.t7 VDD.t3692 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2215 VDD.t358 left_shifter_0.S7.t5 mux8_6.NAND4F_5.Y.t4 VDD.t357 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2216 VDD.t2226 A0.t28 AND8_0.NOT8_0.A0.t5 VDD.t2225 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2217 mux8_3.NAND4F_5.Y.t0 SEL2.t63 VDD.t3776 VDD.t3775 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2218 VDD.t2600 B2.t23 NOT8_0.S2.t1 VDD.t887 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2219 mux8_2.NAND4F_2.D.t2 SEL2.t64 VDD.t3777 VDD.t3733 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2220 MULT_0.NAND2_8.Y.t6 B3.t32 VDD.t2177 VDD.t2176 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2221 VDD.t4256 mux8_7.NAND4F_8.Y.t12 a_11865_n25415.t7 VDD.t4255 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2222 a_n16483_1406.t4 a_n16513_1380.t5 VSS.t733 VSS.t732 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2223 a_11865_n2775.t6 mux8_1.NAND4F_8.Y.t12 VDD.t4321 VDD.t4320 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2224 VSS.t1243 MULT_0.inv_14.Y.t9 a_n16690_n11683.t3 VSS.t1242 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X2225 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t0 A7.t21 a_n24363_373.t0 VSS.t1575 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2226 VDD.t2602 B2.t24 MULT_0.inv_7.A.t1 VDD.t2601 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2227 VDD.t3967 B5.t21 a_n17368_3810.t7 VDD.t3966 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2228 VDD.t3317 MULT_0.inv_15.Y.t9 a_n20557_n11063.t9 VDD.t3316 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2229 MULT_0.NAND2_15.Y.t2 A3.t27 VDD.t4108 VDD.t4107 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2230 VSS.t1608 AND8_0.NOT8_0.A7.t8 AND8_0.S7.t0 VSS.t1607 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2231 VDD.t985 mux8_6.NAND4F_8.Y.t10 a_11865_n34471.t3 VDD.t984 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2232 XOR8_0.S4.t1 a_n12345_n25873.t6 a_n12314_n26419.t1 VDD.t628 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2233 a_n19804_1380.t1 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t11 VDD.t1116 VDD.t1115 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2234 a_n4303_1406.t1 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t19 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t9 VSS.t1861 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2235 a_n12314_n23651.t1 a_n12345_n23393.t5 XOR8_0.S3.t2 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2236 a_n3320_1406.t0 a_n3350_1380.t5 VSS.t1151 VSS.t1150 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2237 XOR8_0.S6.t10 a_n12345_n31115.t4 a_n12314_n31661.t7 VDD.t2640 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2238 a_n13975_n8419.t1 a_n14155_n8419.t5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t1 VSS.t1690 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2239 VDD.t2354 B1.t28 a_n4205_3810.t11 VDD.t2353 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2240 a_n15707_n11063.t0 a_n15737_n11709.t5 mux8_7.A1.t9 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2241 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t10 a_n14155_n5154.t4 a_n13975_n5154.t4 VSS.t1874 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2242 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t7 a_n20737_n8419.t6 a_n20557_n7799.t11 VDD.t2861 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2243 ZFLAG_0.nor4_0.Y.t0 Y0.t4 a_16431_n18523.t0 VDD.t560 sky130_fd_pr__pfet_01v8 ad=1.3268 pd=9.18 as=0.7062 ps=4.61 w=4.28 l=0.15
X2244 a_9432_n11894.t1 mux8_3.NAND4F_0.C.t8 a_9336_n11894.t1 VSS.t1322 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2245 a_n12345_n31115.t0 A6.t15 VSS.t1393 VSS.t1392 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X2246 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t4 a_n368_3164.t4 a_n338_3190.t4 VSS.t820 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2247 mux8_8.A1.t2 a_n19178_n11683.t6 a_n18998_n11063.t4 VDD.t1549 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2248 mux8_8.NAND4F_4.B.t2 SEL0.t83 VDD.t3000 VDD.t2988 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2249 a_n17677_n23825.t7 B6.t22 VDD.t3551 VDD.t3550 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2250 mux8_4.inv_0.A.t3 mux8_4.NAND4F_9.Y.t11 a_11865_n16359.t7 VDD.t962 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X2251 VSS.t901 SEL3.t47 a_n17368_3190.t1 VSS.t900 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2252 VSS.t1228 a_n20587_n11709.t3 a_n20557_n11683.t1 VSS.t1227 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2253 VSS.t1576 A7.t22 OR8_0.NOT8_0.A7.t5 VSS.t177 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X2254 OR8_0.S1.t2 OR8_0.NOT8_0.A1.t9 VDD.t2483 VDD.t2482 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2255 mux8_2.NAND4F_2.Y.t4 mux8_2.NAND4F_2.D.t9 VDD.t3175 VDD.t3174 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2256 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t3 a_n17446_n11683.t3 a_n17266_n11683.t1 VSS.t648 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2257 VDD.t620 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t20 a_n11640_1406.t1 VDD.t619 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X2258 mux8_6.NAND4F_4.B.t2 SEL0.t84 VDD.t2999 VDD.t2949 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2259 mux8_6.NAND4F_1.Y.t0 SEL2.t65 VDD.t3779 VDD.t3778 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2260 mux8_7.A0.t3 a_n16663_1406.t5 a_n16483_2026.t1 VDD.t140 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2261 VSS.t903 SEL3.t48 a_n4205_3190.t0 VSS.t902 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2262 VDD.t4445 SEL1.t82 mux8_1.NAND4F_4.Y.t5 VDD.t4444 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2263 VDD.t2998 SEL0.t85 mux8_6.NAND4F_7.Y.t8 VDD.t2997 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2264 mux8_4.NAND4F_8.Y.t7 mux8_4.NAND4F_4.Y.t10 VDD.t2789 VDD.t2788 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2265 mux8_3.NAND4F_9.Y.t4 mux8_3.NAND4F_6.Y.t10 VDD.t1221 VDD.t1220 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2266 VSS.t1670 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t16 a_n24804_1406.t0 VSS.t1669 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2267 a_n21333_2026.t10 a_n21363_1380.t4 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t10 VDD.t1216 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2268 VDD.t2285 mux8_8.NAND4F_5.Y.t10 mux8_8.NAND4F_9.Y.t2 VDD.t2284 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2269 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t2 MULT_0.4bit_ADDER_1.A2.t11 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2270 mux8_4.NAND4F_4.B.t0 SEL0.t86 VSS.t2013 VSS.t2012 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2271 VDD.t1792 SEL3.t49 a_n914_3810.t0 VDD.t1791 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2272 VSS.t1578 A7.t23 a_1707_4914.t0 VSS.t1577 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2273 OR8_0.NOT8_0.A2.t3 A2.t22 a_n17677_n18225.t3 VDD.t527 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X2274 a_n15707_n5154.t1 a_n15887_n5154.t4 MULT_0.4bit_ADDER_1.B1.t7 VSS.t1153 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2275 VDD.t2179 B3.t33 MULT_0.NAND2_9.Y.t6 VDD.t2178 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2276 mux8_7.NAND4F_1.Y.t5 XOR8_0.S5.t13 VDD.t1204 VDD.t1203 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2277 mux8_0.NAND4F_5.Y.t1 SEL2.t66 VDD.t3781 VDD.t3780 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2278 VDD.t1008 B0.t27 left_shifter_0.buffer_6.inv_1.A.t2 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2279 VDD.t2904 mux8_6.NAND4F_8.Y.t11 a_11865_n34471.t2 VDD.t2903 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2280 a_9336_1690.t0 mux8_0.NAND4F_2.D.t9 VSS.t1440 VSS.t1439 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2281 mux8_1.NAND4F_1.Y.t2 mux8_1.NAND4F_0.C.t9 VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2282 a_n11840_n11683.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t20 mux8_5.A1.t3 VSS.t1046 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2283 a_n12314_n29052.t1 B5.t22 VDD.t3969 VDD.t3968 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2284 VDD.t3931 MULT_0.NAND2_9.Y.t8 MULT_0.inv_9.Y.t3 VDD.t3930 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2285 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t19 VDD.t3664 VDD.t3663 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2286 a_n11274_n31085.t4 A6.t16 VSS.t1395 VSS.t1394 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2287 VDD.t3919 mux8_3.inv_0.A.t9 Y2.t1 VDD.t3918 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2288 a_n10884_1406.t4 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t21 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t1 VSS.t302 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2289 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t5 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t9 VDD.t2188 VDD.t2187 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2290 a_n22372_373.t1 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t7 VSS.t1328 VSS.t951 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2291 a_11386_n21878.t1 mux8_5.NAND4F_6.Y.t10 a_11290_n21878.t1 VSS.t701 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2292 a_n10684_n11063.t0 MULT_0.4bit_ADDER_2.B0.t18 VDD.t1073 VDD.t1072 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2293 VDD.t3358 8bit_ADDER_0.S0.t14 mux8_1.NAND4F_3.Y.t3 VDD.t3357 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2294 OR8_0.NOT8_0.A1.t3 A1.t25 a_n17677_n16825.t7 VDD.t4216 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2295 a_n15896_n9452.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t18 VSS.t322 VSS.t321 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2296 VDD.t1897 MULT_0.4bit_ADDER_2.B1.t17 a_n13975_n11063.t8 VDD.t1896 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2297 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t8 a_n17446_n11683.t4 a_n17266_n11683.t0 VSS.t646 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2298 VDD.t2444 MULT_0.inv_14.Y.t10 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t4 VDD.t2443 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2299 a_5773_4912.t3 mux8_6.A0.t18 VSS.t1523 VSS.t1522 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2300 8bit_ADDER_0.S2.t5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t16 a_n6035_1406.t4 VSS.t1250 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2301 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t1 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t19 VDD.t1049 VDD.t1048 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2302 VDD.t1375 mux8_5.NAND4F_2.D.t9 mux8_5.NAND4F_2.Y.t0 VDD.t1374 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2303 a_n10210_3190.t4 a_n10966_3190.t5 VSS.t1554 VSS.t1553 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2304 a_n12314_n18115.t10 a_n12345_n17857.t5 XOR8_0.S1.t9 VDD.t2458 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2305 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t1 A3.t28 VDD.t4110 VDD.t4109 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2306 a_n12416_n11683.t1 a_n12446_n11709.t4 VSS.t1941 VSS.t1940 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2307 a_9432_n34534.t0 mux8_6.NAND4F_0.C.t11 a_9336_n34534.t1 VSS.t152 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2308 mux8_5.inv_0.A.t2 mux8_5.NAND4F_9.Y.t13 a_11865_n20887.t3 VDD.t689 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2309 VSS.t691 B7.t20 left_shifter_0.buffer_1.inv_1.A.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2310 mux8_7.NAND4F_8.Y.t1 mux8_7.NAND4F_4.Y.t10 VDD.t513 VDD.t512 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2311 VDD.t2996 SEL0.t87 mux8_0.NAND4F_4.B.t2 VDD.t2943 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2312 a_n20083_3190.t4 a_n20113_3164.t6 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t9 VSS.t1326 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2313 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t8 B3.t34 a_n10786_3190.t3 VSS.t1112 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2314 a_n12345_n17569.t0 A1.t26 VSS.t1906 VSS.t1905 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X2315 mux8_7.NAND4F_4.B.t0 SEL0.t88 VSS.t2011 VSS.t2010 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2316 VSS.t504 B0.t28 right_shifter_0.buffer_6.inv_1.A.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2317 a_n17368_3810.t10 a_n17548_3190.t5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t10 VDD.t1143 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2318 VSS.t1126 A0.t29 a_n11276_n14723.t2 VSS.t1125 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X2319 a_n6920_3190.t4 a_n6950_3164.t4 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t7 VSS.t1806 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2320 mux8_5.NAND4F_3.Y.t5 mux8_5.NAND4F_4.B.t8 VDD.t1991 VDD.t1990 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2321 VDD.t1010 B0.t29 a_n17677_n15425.t6 VDD.t1009 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2322 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t5 a_n24130_3190.t6 a_n23950_3810.t4 VDD.t3698 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2323 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t6 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t13 VDD.t1879 VDD.t1878 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2324 mux8_6.NAND4F_1.Y.t7 XOR8_0.S7.t13 VDD.t3268 VDD.t3267 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2325 mux8_0.NAND4F_9.Y.t1 mux8_0.NAND4F_5.Y.t11 VDD.t1258 VDD.t1257 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2326 a_n10684_n11063.t11 a_n10714_n11709.t5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t11 VDD.t2007 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2327 a_7548_n11894.t1 SEL1.t83 a_7452_n11894.t1 VSS.t1973 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2328 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t6 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t16 VDD.t943 VDD.t942 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2329 a_n24012_n16501.t1 A1.t27 AND8_0.NOT8_0.A1.t0 VSS.t1907 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2330 VDD.t1514 mux8_8.NAND4F_2.D.t13 mux8_8.NAND4F_0.Y.t3 VDD.t1513 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2331 VDD.t1187 right_shifter_0.buffer_1.inv_1.A.t5 right_shifter_0.S6.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2332 VDD.t2053 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t17 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t1 VDD.t2052 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2333 VDD.t2190 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t10 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t6 VDD.t2189 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2334 mux8_4.A1.t4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t18 a_n8549_n11683.t4 VSS.t1562 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2335 a_9528_n30006.t0 mux8_8.NAND4F_4.B.t10 a_9432_n30006.t0 VSS.t1467 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2336 VDD.t2032 MULT_0.S1.t13 mux8_2.NAND4F_0.Y.t1 VDD.t2031 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2337 VSS.t1502 MULT_0.4bit_ADDER_1.B1.t17 a_n14155_n8419.t0 VSS.t1501 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2338 left_shifter_0.buffer_7.inv_1.A.t1 B1.t29 VDD.t2355 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2339 mux8_1.inv_0.A.t3 mux8_1.NAND4F_9.Y.t11 a_11865_n2775.t2 VDD.t1320 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2340 VDD.t3223 mux8_2.NAND4F_4.B.t9 mux8_2.NAND4F_5.Y.t6 VDD.t3222 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2341 NOT8_0.S0.t3 B0.t30 VDD.t1012 VDD.t1011 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2342 VDD.t645 mux8_0.NAND4F_0.C.t8 mux8_0.NAND4F_0.Y.t1 VDD.t644 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2343 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t4 a_n14931_1406.t5 a_n14751_1406.t4 VSS.t1546 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2344 MULT_0.NAND2_1.Y.t0 A2.t23 a_n22176_n2915.t0 VSS.t252 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2345 VDD.t3890 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t19 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t5 VDD.t3889 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2346 VDD.t1692 mux8_6.inv_0.A.t9 Y7.t1 VDD.t1691 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2347 a_11865_1753.t6 mux8_0.NAND4F_9.Y.t11 mux8_0.inv_0.A.t3 VDD.t3123 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2348 a_n12347_n33735.t0 A7.t24 VSS.t1580 VSS.t1579 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X2349 VDD.t3237 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t17 a_n21333_2026.t1 VDD.t3236 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2350 mux8_7.NAND4F_5.Y.t8 left_shifter_0.S5.t6 VDD.t2791 VDD.t2790 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2351 mux8_2.NAND4F_7.Y.t7 mux8_2.NAND4F_0.C.t10 VDD.t3209 VDD.t3208 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2352 OR8_0.NOT8_0.A7.t2 A7.t25 a_n17677_n25225.t2 VDD.t3429 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2353 VDD.t3782 SEL2.t67 mux8_2.NAND4F_2.D.t1 VDD.t3733 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2354 VDD.t3193 MULT_0.4bit_ADDER_1.A0.t10 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t5 VDD.t3192 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2355 mux8_4.NAND4F_9.Y.t1 mux8_4.NAND4F_5.Y.t11 VDD.t4023 VDD.t4022 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2356 VDD.t4447 SEL1.t84 mux8_1.NAND4F_5.Y.t5 VDD.t4446 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2357 VDD.t27 MULT_0.4bit_ADDER_1.A2.t12 a_n17266_n7799.t9 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2358 a_11865_n25415.t6 mux8_7.NAND4F_8.Y.t13 VDD.t4258 VDD.t4257 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2359 a_n12314_n23651.t7 B3.t35 VDD.t2181 VDD.t2180 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2360 XOR8_0.S6.t6 a_n12345_n31403.t5 a_n12314_n31661.t9 VDD.t1830 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2361 VDD.t2995 SEL0.t89 mux8_2.NAND4F_2.Y.t2 VDD.t2994 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2362 mux8_2.NAND4F_8.Y.t6 mux8_2.NAND4F_2.Y.t10 VDD.t2108 VDD.t2107 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2363 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t9 MULT_0.4bit_ADDER_1.B2.t18 a_n16690_n8419.t1 VSS.t1819 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2364 VSS.t1430 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t16 a_n18222_1406.t0 VSS.t1429 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2365 a_n16690_n5154.t4 MULT_0.4bit_ADDER_0.B2.t9 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t10 VSS.t1449 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2366 a_n9901_1406.t5 a_n9931_1380.t6 VSS.t1118 VSS.t1117 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2367 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t2 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t18 VDD.t3474 VDD.t3473 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2368 VDD.t2042 OR8_0.S4.t4 mux8_5.NAND4F_2.Y.t2 VDD.t2041 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2369 V.t0 V_FLAG_0.NAND2_0.Y.t8 VSS.t1613 VSS.t1612 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2370 a_n1012_1406.t0 A0.t30 VSS.t1128 VSS.t1127 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2371 VDD.t3553 B6.t23 a_n17677_n23825.t6 VDD.t3552 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2372 a_n19774_1406.t1 a_n19804_1380.t5 VSS.t718 VSS.t717 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2373 a_n10786_3810.t3 a_n10240_3164.t6 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t4 VDD.t685 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2374 mux8_2.NAND4F_6.Y.t1 SEL2.t68 VDD.t3784 VDD.t3783 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2375 VDD.t3555 B6.t24 a_n20659_3810.t4 VDD.t3554 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2376 VDD.t968 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t9 mux8_6.A1.t5 VDD.t967 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2377 a_n11276_n33705.t1 A7.t26 VSS.t1582 VSS.t1581 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2378 a_n7594_1406.t1 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t16 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t7 VSS.t432 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2379 a_7548_n34534.t0 SEL1.t85 a_7452_n34534.t1 VSS.t1964 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2380 NOT8_0.S0.t2 B0.t31 VDD.t1014 VDD.t1013 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2381 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t12 a_n19187_n6187.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2382 VDD.t1606 MULT_0.4bit_ADDER_0.A3.t9 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t2 VDD.t1605 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2383 a_n18422_n8419.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t20 MULT_0.4bit_ADDER_2.B2.t6 VSS.t524 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2384 VDD.t2604 B2.t25 a_n7496_3810.t9 VDD.t2603 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2385 VDD.t1608 MULT_0.4bit_ADDER_0.A3.t10 a_n20557_n4534.t1 VDD.t1607 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2386 VDD.t3696 XOR8_0.S0.t13 mux8_1.NAND4F_1.Y.t5 VDD.t3695 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2387 mux8_5.NAND4F_9.Y.t1 mux8_5.NAND4F_5.Y.t11 VDD.t1156 VDD.t1155 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2388 a_n19963_373.t1 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t16 VSS.t1207 VSS.t552 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2389 MULT_0.4bit_ADDER_1.B2.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t17 a_n18422_n5154.t0 VSS.t237 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2390 a_n17677_n18225.t2 A2.t24 OR8_0.NOT8_0.A2.t2 VDD.t528 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2391 VDD.t4449 SEL1.t86 mux8_4.NAND4F_0.C.t3 VDD.t4448 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2392 VDD.t1794 SEL3.t50 a_n29_2026.t0 VDD.t1793 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2393 VSS.t1144 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t18 a_n209_1406.t0 VSS.t1143 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2394 left_shifter_0.buffer_5.inv_1.A.t1 B3.t36 VDD.t2182 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2395 mux8_4.A0.t0 a_n9931_1380.t7 a_n9901_2026.t0 VDD.t333 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2396 mux8_6.NAND4F_5.Y.t3 left_shifter_0.S7.t6 VDD.t360 VDD.t359 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2397 VDD.t1426 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t22 a_n14931_1406.t1 VDD.t1425 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X2398 VSS.t1863 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t20 a_n5059_1406.t0 VSS.t1862 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2399 mux8_8.A0.t8 a_n19954_1406.t5 a_n19774_2026.t11 VDD.t2648 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2400 VDD.t396 A5.t16 a_n18042_2026.t2 VDD.t395 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2401 a_n9155_n5180.t0 VSS.t1004 VSS.t1006 VSS.t1005 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X2402 a_11865_n25415.t5 mux8_7.NAND4F_8.Y.t14 VDD.t4260 VDD.t4259 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X2403 VDD.t3557 B6.t25 AND8_0.NOT8_0.A6.t5 VDD.t3556 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2404 VSS.t905 SEL3.t51 a_n7496_3190.t0 VSS.t904 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2405 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t3 A7.t27 VDD.t3431 VDD.t3430 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2406 a_n11274_n28476.t4 A5.t17 VSS.t186 VSS.t185 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2407 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t9 a_n15014_n12716.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2408 a_10363_n20950.t0 mux8_5.NAND4F_0.C.t12 a_10267_n20950.t0 VSS.t1665 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2409 a_n24624_2026.t6 a_n24654_1380.t6 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t6 VDD.t3882 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2410 VDD.t530 A2.t25 a_n8170_2026.t4 VDD.t529 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2411 MULT_0.inv_9.Y.t2 MULT_0.NAND2_9.Y.t9 VDD.t3932 VDD.t3930 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2412 VSS.t1397 A6.t17 a_n11274_n31085.t5 VSS.t1396 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2413 mux8_0.NAND4F_7.Y.t0 SEL2.t69 VDD.t3786 VDD.t3785 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2414 mux8_0.NAND4F_9.Y.t8 mux8_0.NAND4F_7.Y.t11 VDD.t1502 VDD.t1501 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2415 VDD.t4112 A3.t29 MULT_0.NAND2_15.Y.t1 VDD.t4111 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2416 AND8_0.S0.t2 AND8_0.NOT8_0.A0.t9 VDD.t1355 VDD.t1354 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2417 a_1887_5534.t6 B7.t21 VDD.t1411 VDD.t1410 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2418 8bit_ADDER_0.C.t0 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t7 a_n22372_373.t0 VSS.t951 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2419 a_11865_n34471.t1 mux8_6.NAND4F_8.Y.t12 VDD.t2906 VDD.t2905 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2420 left_shifter_0.S1.t2 left_shifter_0.buffer_6.inv_1.A.t6 VDD.t1239 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2421 8bit_ADDER_0.S0.t1 a_n209_1406.t5 a_n29_1406.t1 VSS.t1452 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2422 VDD.t1881 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t14 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t5 VDD.t1880 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2423 VDD.t3160 mux8_8.NAND4F_4.B.t11 mux8_8.NAND4F_4.Y.t7 VDD.t3159 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2424 VDD.t373 mux8_0.NAND4F_3.Y.t10 mux8_0.NAND4F_8.Y.t0 VDD.t372 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2425 a_n9125_n4534.t1 a_n9155_n5180.t4 MULT_0.S1.t1 VDD.t309 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2426 mux8_7.A1.t10 a_n15737_n11709.t6 a_n15707_n11063.t1 VDD.t101 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2427 OR8_0.NOT8_0.A2.t6 B2.t26 VSS.t1295 VSS.t810 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X2428 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t1 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t19 VDD.t3476 VDD.t3475 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2429 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t8 VDD.t2249 VDD.t2248 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2430 a_16431_n18523.t1 Y0.t5 ZFLAG_0.nor4_0.Y.t1 VDD.t561 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X2431 VDD.t4218 A1.t28 MULT_0.NAND2_5.Y.t6 VDD.t4217 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2432 a_9336_n11894.t0 mux8_3.NAND4F_2.D.t12 VSS.t1383 VSS.t1382 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2433 VSS.t395 OR8_0.NOT8_0.A7.t8 OR8_0.S7.t0 VSS.t394 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2434 OR8_0.NOT8_0.A4.t3 A4.t17 a_n17677_n21025.t6 VDD.t1642 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X2435 a_n20557_n11683.t0 a_n20587_n11709.t4 VSS.t1230 VSS.t1229 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2436 mux8_0.NAND4F_4.Y.t7 SEL1.t87 VDD.t4451 VDD.t4450 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2437 a_11865_n25415.t1 mux8_7.NAND4F_9.Y.t13 mux8_7.inv_0.A.t2 VDD.t3284 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2438 XOR8_0.S1.t10 a_n12345_n17857.t6 a_n12314_n18115.t11 VDD.t2459 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2439 mux8_7.NAND4F_6.Y.t5 SEL1.t88 VDD.t4453 VDD.t4452 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2440 mux8_7.NAND4F_8.Y.t2 mux8_7.NAND4F_4.Y.t11 a_11386_n25478.t0 VSS.t243 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2441 a_2463_4914.t1 A7.t28 V_FLAG_0.XOR2_2.B.t2 VSS.t1583 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2442 MULT_0.NAND2_11.Y.t2 B1.t30 VDD.t2357 VDD.t2356 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2443 VDD.t3788 SEL2.t70 mux8_7.NAND4F_7.Y.t1 VDD.t3787 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2444 mux8_6.NAND4F_7.Y.t7 SEL0.t90 VDD.t2993 VDD.t2992 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2445 a_n23065_2026.t0 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t20 VDD.t3478 VDD.t3477 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2446 XOR8_0.S3.t11 a_n12345_n23105.t5 a_n12314_n23651.t10 VDD.t2764 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2447 mux8_8.NAND4F_9.Y.t1 mux8_8.NAND4F_5.Y.t11 VDD.t2287 VDD.t2286 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2448 a_n11276_n14723.t1 A0.t31 VSS.t1130 VSS.t1129 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2449 a_n3320_1406.t3 a_n3500_1406.t4 8bit_ADDER_0.S1.t8 VSS.t765 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2450 VDD.t200 mux8_7.NAND4F_4.B.t9 mux8_7.NAND4F_1.Y.t8 VDD.t199 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2451 a_n12345_n23105.t0 A3.t30 VSS.t1841 VSS.t1840 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X2452 VSS.t63 left_shifter_0.buffer_1.inv_1.A.t5 left_shifter_0.C.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2453 VDD.t3433 A7.t29 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t2 VDD.t3432 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2454 a_8496_n7266.t0 SEL1.t89 a_8400_n7266.t1 VSS.t1966 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2455 a_11194_n7266.t0 mux8_2.NAND4F_0.Y.t10 VSS.t1949 VSS.t667 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2456 a_n19981_n8419.t0 MULT_0.4bit_ADDER_1.B3.t14 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t2 VSS.t1338 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2457 Y1.t1 mux8_2.inv_0.A.t8 VSS.t749 VSS.t748 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2458 a_3493_5534.t8 a_3313_4914.t5 V_FLAG_0.XOR2_2.Y.t9 VDD.t1098 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2459 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t6 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t17 VDD.t3644 VDD.t3643 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2460 a_n17266_n5154.t3 a_n17296_n5180.t3 VSS.t1201 VSS.t1200 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2461 MULT_0.4bit_ADDER_2.B3.t1 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t9 VDD.t145 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2462 a_11865_n34471.t0 mux8_6.NAND4F_8.Y.t13 VDD.t2908 VDD.t2907 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X2463 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t11 B4.t24 a_n14077_3190.t3 VSS.t1654 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2464 VDD.t1796 SEL3.t52 a_n14077_3810.t0 VDD.t1795 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2465 a_n29_1406.t4 a_n59_1380.t6 VSS.t1199 VSS.t1198 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2466 XOR8_0.S7.t3 a_n12347_n34023.t5 a_n12316_n34281.t3 VDD.t973 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2467 a_n20757_1406.t4 A6.t18 VSS.t1399 VSS.t1398 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2468 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t10 B1.t31 a_n4205_3190.t4 VSS.t1180 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2469 mux8_5.A0.t9 a_n13222_1380.t5 a_n13192_2026.t5 VDD.t774 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2470 VDD.t839 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t14 a_n15707_n11063.t4 VDD.t838 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2471 a_8496_1690.t0 SEL1.t90 a_8400_1690.t1 VSS.t1968 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2472 a_n12416_n4534.t9 a_n12446_n5180.t4 MULT_0.4bit_ADDER_1.B0.t4 VDD.t3286 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2473 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t14 VDD.t3674 VDD.t3673 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2474 right_shifter_0.S6.t2 right_shifter_0.buffer_1.inv_1.A.t6 VDD.t1188 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2475 VDD.t3480 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t21 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t0 VDD.t3479 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2476 mux8_6.NAND4F_0.C.t0 SEL1.t91 VSS.t1975 VSS.t1974 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2477 VDD.t2629 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t16 a_n3320_2026.t7 VDD.t2628 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2478 a_n17266_n7799.t4 a_n17446_n8419.t6 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t7 VDD.t733 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2479 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t4 a_n10864_n11683.t5 a_n10684_n11063.t2 VDD.t1537 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2480 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t4 MULT_0.4bit_ADDER_2.B1.t18 a_n13399_n11683.t4 VSS.t971 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2481 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t7 VDD.t2516 VDD.t2515 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2482 a_3493_4914.t1 a_3463_4888.t5 VSS.t231 VSS.t230 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2483 a_n16690_n11683.t1 MULT_0.4bit_ADDER_2.B2.t20 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t1 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2484 AND8_0.S2.t1 AND8_0.NOT8_0.A2.t9 VDD.t3483 VDD.t678 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2485 VDD.t2809 mux8_3.NAND4F_2.D.t13 mux8_3.NAND4F_0.Y.t4 VDD.t2808 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2486 a_11865_n34471.t6 mux8_6.NAND4F_9.Y.t12 mux8_6.inv_0.A.t4 VDD.t697 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2487 mux8_5.NAND4F_2.Y.t1 mux8_5.NAND4F_2.D.t10 VDD.t1377 VDD.t1376 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2488 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t2 B6.t26 a_n20659_3190.t3 VSS.t1634 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2489 VSS.t1787 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t16 a_n12616_1406.t4 VSS.t1786 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X2490 VDD.t3790 SEL2.t71 mux8_3.NAND4F_2.D.t3 VDD.t3789 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2491 VSS.t1943 a_n12446_n11709.t5 a_n12416_n11683.t0 VSS.t1942 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2492 mux8_6.NAND4F_6.Y.t5 SEL1.t92 VDD.t4455 VDD.t4454 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2493 a_9336_n34534.t0 mux8_6.NAND4F_2.D.t12 VSS.t205 VSS.t204 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2494 a_11865_n20887.t5 mux8_5.NAND4F_8.Y.t14 VDD.t4306 VDD.t4305 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2495 VDD.t3792 SEL2.t72 mux8_4.NAND4F_2.D.t3 VDD.t3791 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2496 a_n10108_n5154.t1 MULT_0.4bit_ADDER_0.A0.t10 VSS.t638 VSS.t637 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2497 a_n11274_n23075.t1 A3.t31 VSS.t1843 VSS.t1842 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2498 VDD.t3435 A7.t30 AND8_0.NOT8_0.A7.t0 VDD.t3434 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2499 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t0 a_n18222_1406.t5 a_n18042_1406.t4 VSS.t1768 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2500 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t2 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t17 VDD.t338 VDD.t337 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2501 a_n19981_n8419.t4 MULT_0.4bit_ADDER_1.A3.t11 VSS.t1894 VSS.t1893 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2502 VDD.t2991 SEL0.t91 mux8_2.NAND4F_6.Y.t7 VDD.t2990 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2503 mux8_2.NAND4F_9.Y.t8 mux8_2.NAND4F_6.Y.t9 VDD.t2849 VDD.t2848 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2504 VDD.t1278 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t17 a_n15707_n11063.t8 VDD.t1277 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2505 MULT_0.NAND2_9.Y.t2 A1.t29 VDD.t4220 VDD.t4219 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2506 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t5 MULT_0.inv_8.Y.t10 VDD.t3521 VDD.t3520 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2507 VDD.t3646 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t18 a_n24624_2026.t9 VDD.t3645 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2508 VSS.t662 a_n19028_n8445.t4 a_n18998_n8419.t4 VSS.t661 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2509 VDD.t1581 8bit_ADDER_0.C.t8 mux8_0.NAND4F_3.Y.t5 VDD.t1580 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2510 mux8_5.NAND4F_5.Y.t2 left_shifter_0.S4.t4 a_7644_n21878.t1 VSS.t328 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2511 VDD.t3574 NOT8_0.S3.t6 mux8_4.NAND4F_7.Y.t3 VDD.t3573 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2512 VDD.t3437 A7.t31 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t1 VDD.t3436 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2513 a_n18998_n5154.t3 a_n19028_n5180.t2 VSS.t1405 VSS.t1404 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2514 VDD.t11 mux8_6.NAND4F_4.B.t10 mux8_6.NAND4F_1.Y.t5 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2515 a_n23960_n22530.t1 A6.t19 AND8_0.NOT8_0.A6.t0 VSS.t1158 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2516 a_n12446_n8445.t1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t13 VDD.t4290 VDD.t4289 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2517 VDD.t3523 MULT_0.inv_8.Y.t11 a_n10684_n11063.t4 VDD.t3522 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2518 VDD.t945 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t17 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t5 VDD.t944 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2519 a_5773_4912.t1 A7.t32 V_FLAG_0.XOR2_0.Y.t10 VSS.t1584 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2520 mux8_8.NAND4F_0.Y.t2 mux8_8.NAND4F_2.D.t14 VDD.t1516 VDD.t1515 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2521 VDD.t2672 mux8_3.NAND4F_0.C.t9 mux8_3.NAND4F_7.Y.t5 VDD.t2671 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2522 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t19 VDD.t3648 VDD.t3647 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2523 VSS.t1586 A7.t33 a_n11276_n33705.t0 VSS.t1585 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2524 VSS.t1168 MULT_0.4bit_ADDER_0.A1.t9 a_n13399_n5154.t0 VSS.t1167 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2525 a_16431_n19505.t3 Y6.t7 a_16143_n19505.t3 VDD.t3169 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X2526 right_shifter_0.S6.t1 right_shifter_0.buffer_1.inv_1.A.t7 VDD.t1189 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2527 a_n19187_n6187.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t18 VSS.t239 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2528 a_n20587_n11709.t1 MULT_0.inv_15.Y.t10 VDD.t3319 VDD.t3318 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2529 a_n17266_n8419.t0 a_n17296_n8445.t6 VSS.t1512 VSS.t1511 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2530 a_n8549_n11683.t5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t19 mux8_4.A1.t3 VSS.t1563 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2531 VDD.t532 A2.t26 AND8_0.NOT8_0.A2.t3 VDD.t531 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2532 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t4 a_n24804_1406.t6 a_n24624_1406.t4 VSS.t1598 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2533 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t0 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t12 a_n19963_373.t0 VSS.t552 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2534 VSS.t1203 a_n17296_n5180.t4 a_n17266_n5154.t4 VSS.t1202 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2535 a_n17677_n18225.t6 B2.t27 VDD.t2606 VDD.t2605 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2536 mux8_4.NAND4F_0.C.t2 SEL1.t93 VDD.t4456 VDD.t4448 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2537 VDD.t2359 B1.t32 MULT_0.NAND2_4.Y.t2 VDD.t2358 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2538 VDD.t1937 VSS.t2056 a_n20557_n4534.t7 VDD.t1936 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2539 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t5 a_n5059_1406.t6 a_n4879_1406.t1 VSS.t400 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2540 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t8 VDD.t2744 VDD.t2743 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2541 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t11 a_n10864_n5154.t6 a_n10684_n4534.t11 VDD.t2863 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2542 MULT_0.S1.t9 a_n9305_n5154.t6 a_n9125_n4534.t5 VDD.t1539 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2543 a_n4205_3810.t4 a_n3659_3164.t5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t6 VDD.t1199 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2544 a_10267_n3765.t0 SEL2.t73 VSS.t1726 VSS.t853 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2545 VDD.t4114 A3.t32 MULT_0.inv_13.A.t5 VDD.t4113 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2546 a_n11274_n17539.t4 A1.t30 VSS.t1909 VSS.t1908 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2547 VDD.t3439 A7.t34 a_5197_5532.t10 VDD.t3438 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2548 VDD.t3666 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t20 a_n19178_n11683.t1 VDD.t3665 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X2549 VSS.t188 A5.t18 a_n11274_n28476.t3 VSS.t187 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2550 VDD.t2518 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t8 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t1 VDD.t2517 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2551 mux8_7.NAND4F_2.Y.t1 OR8_0.S5.t4 a_8592_n25478.t0 VSS.t1050 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2552 VDD.t3957 NOT8_0.S4.t6 mux8_5.NAND4F_7.Y.t5 VDD.t3956 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2553 VDD.t432 mux8_6.NAND4F_2.D.t13 mux8_6.NAND4F_0.Y.t1 VDD.t431 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2554 XOR8_0.S4.t7 a_n12345_n26161.t5 a_n12314_n26419.t7 VDD.t3526 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2555 AND8_0.S3.t2 AND8_0.NOT8_0.A3.t9 VDD.t2385 VDD.t674 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2556 VDD.t981 V_FLAG_0.XOR2_2.B.t17 a_3493_5534.t5 VDD.t980 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2557 a_n9125_n11683.t0 a_n9155_n11709.t3 VSS.t448 VSS.t447 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2558 a_n16483_2026.t10 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t17 VDD.t3905 VDD.t3904 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2559 a_n14751_2026.t1 a_n14781_1380.t4 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t1 VDD.t558 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2560 MULT_0.NAND2_4.Y.t1 B1.t33 VDD.t2361 VDD.t2360 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2561 a_n17677_n16825.t2 B1.t34 VDD.t2363 VDD.t2362 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X2562 a_n11274_n20496.t5 B2.t28 XOR8_0.S2.t0 VSS.t1296 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2563 MULT_0.SO.t2 MULT_0.NAND2_3.Y.t9 VDD.t164 VDD.t162 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2564 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t6 MULT_0.4bit_ADDER_0.B1.t9 VDD.t1337 VDD.t1336 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2565 VDD.t2989 SEL0.t92 mux8_8.NAND4F_4.B.t1 VDD.t2988 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2566 mux8_5.NAND4F_2.Y.t3 OR8_0.S4.t5 VDD.t2044 VDD.t2043 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2567 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t6 a_n21513_1406.t5 a_n21333_2026.t8 VDD.t1196 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2568 a_n4879_2026.t4 a_n4909_1380.t5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t7 VDD.t1183 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2569 VDD.t3650 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t20 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t4 VDD.t3649 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2570 a_n12416_n4534.t7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t18 VDD.t4178 VDD.t4177 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2571 a_7452_n26406.t0 SEL2.t74 VSS.t1727 VSS.t1456 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2572 a_n17677_n21025.t7 A4.t18 OR8_0.NOT8_0.A4.t2 VDD.t1643 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2573 a_n3320_2026.t1 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t20 VDD.t757 VDD.t756 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2574 VDD.t1899 MULT_0.4bit_ADDER_2.B1.t19 a_n14155_n11683.t1 VDD.t1898 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X2575 VDD.t73 mux8_1.NAND4F_0.C.t10 mux8_1.NAND4F_3.Y.t1 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2576 VSS.t348 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t14 a_n15131_n5154.t3 VSS.t347 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2577 mux8_6.A1.t4 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t10 VDD.t970 VDD.t969 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2578 mux8_6.NAND4F_2.D.t0 SEL2.t75 VSS.t1729 VSS.t1728 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2579 V_FLAG_0.XOR2_2.Y.t1 SEL3.t53 a_4069_4914.t1 VSS.t906 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2580 a_n10423_n9452.t0 MULT_0.4bit_ADDER_1.B0.t19 VSS.t1264 VSS.t1263 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2581 a_n20557_n11063.t6 a_n20587_n11709.t5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t0 VDD.t2430 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2582 a_8592_n2838.t1 SEL0.t93 a_8496_n2838.t1 VSS.t2006 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2583 a_11290_n2838.t1 mux8_1.NAND4F_3.Y.t11 a_11194_n2838.t1 VSS.t464 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2584 VDD.t2055 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t18 a_n9305_n5154.t1 VDD.t2054 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X2585 VDD.t4275 MULT_0.inv_13.A.t9 MULT_0.4bit_ADDER_1.A3.t2 VDD.t4273 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2586 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t3 MULT_0.inv_8.Y.t12 a_n10423_n12716.t1 VSS.t428 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2587 VDD.t4033 MULT_0.4bit_ADDER_1.B2.t19 a_n17446_n8419.t1 VDD.t4032 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X2588 VDD.t2530 mux8_3.NAND4F_4.B.t10 mux8_3.NAND4F_4.Y.t5 VDD.t2529 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2589 a_n11276_n14723.t3 B0.t32 XOR8_0.S0.t2 VSS.t505 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2590 a_n16822_3164.t0 B5.t23 VSS.t1798 VSS.t1797 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X2591 VDD.t3794 SEL2.t76 mux8_0.NAND4F_1.Y.t1 VDD.t3793 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2592 VSS.t938 a_n12345_n28506.t6 a_n11274_n29052.t2 VSS.t937 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2593 OR8_0.NOT8_0.A4.t6 B4.t25 VSS.t1655 VSS.t810 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X2594 a_10363_n16422.t0 mux8_4.NAND4F_0.C.t12 a_10267_n16422.t1 VSS.t1497 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2595 mux8_1.NAND4F_0.Y.t6 mux8_1.NAND4F_2.D.t11 VDD.t1714 VDD.t1713 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2596 a_n9125_n11683.t1 a_n9155_n11709.t4 VSS.t450 VSS.t449 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2597 VSS.t819 A4.t19 a_n11274_n25843.t5 VSS.t818 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2598 VDD.t2283 NOT8_0.S6.t6 mux8_8.NAND4F_7.Y.t6 VDD.t2282 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2599 mux8_3.NAND4F_0.C.t0 SEL1.t94 VSS.t1977 VSS.t1976 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2600 a_n12316_n34281.t7 B7.t22 VDD.t1413 VDD.t1412 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2601 a_10267_n20950.t1 mux8_5.NAND4F_2.D.t11 VSS.t680 VSS.t679 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2602 VDD.t1357 AND8_0.NOT8_0.A0.t10 AND8_0.S0.t1 VDD.t1356 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2603 VDD.t1240 left_shifter_0.buffer_6.inv_1.A.t7 left_shifter_0.S1.t1 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2604 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t11 a_n20587_n8445.t6 a_n20557_n7799.t0 VDD.t2870 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2605 VDD.t3499 V_FLAG_0.NAND2_0.Y.t9 V.t2 VDD.t3498 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2606 VDD.t118 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t8 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t1 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2607 mux8_8.NAND4F_4.Y.t8 mux8_8.NAND4F_4.B.t12 VDD.t3162 VDD.t3161 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2608 VDD.t1367 mux8_5.A1.t14 mux8_5.NAND4F_0.Y.t2 VDD.t1366 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2609 a_n10786_3190.t1 SEL3.t54 VSS.t908 VSS.t907 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2610 VSS.t1604 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t22 a_n23245_1406.t0 VSS.t1603 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2611 VDD.t1740 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t16 a_n9901_2026.t3 VDD.t1739 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2612 ZFLAG_0.nor4_0.Y.t2 Y0.t6 a_16431_n18523.t2 VDD.t562 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X2613 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t7 a_n368_3164.t5 a_n914_3810.t10 VDD.t1645 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2614 VDD.t4323 mux8_1.NAND4F_8.Y.t13 a_11865_n2775.t5 VDD.t4322 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2615 VSS.t847 a_n9155_n8445.t4 a_n9125_n8419.t1 VSS.t846 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2616 mux8_0.inv_0.A.t4 mux8_0.NAND4F_9.Y.t12 a_11865_1753.t7 VDD.t3124 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X2617 MULT_0.inv_7.A.t0 B2.t29 VDD.t2608 VDD.t2607 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2618 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t5 a_n20737_n11683.t4 a_n20557_n11683.t5 VSS.t1594 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2619 a_7452_n35462.t0 SEL2.t77 VSS.t1730 VSS.t206 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2620 a_8400_n12822.t0 SEL2.t78 VSS.t1731 VSS.t1380 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2621 VDD.t1798 SEL3.t55 a_n17368_3810.t1 VDD.t1797 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2622 a_n1618_1380.t1 A0.t32 VDD.t2228 VDD.t2227 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2623 mux8_7.inv_0.A.t1 mux8_7.NAND4F_9.Y.t14 a_11865_n25415.t0 VDD.t3285 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2624 AND8_0.S5.t1 AND8_0.NOT8_0.A5.t9 VDD.t2638 VDD.t678 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2625 VDD.t4180 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t19 a_n12596_n5154.t1 VDD.t4179 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X2626 mux8_3.NAND4F_2.D.t2 SEL2.t79 VDD.t3795 VDD.t3789 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2627 VDD.t3797 SEL2.t80 mux8_7.NAND4F_6.Y.t1 VDD.t3796 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2628 mux8_4.NAND4F_2.D.t2 SEL2.t81 VDD.t3798 VDD.t3791 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2629 mux8_7.NAND4F_7.Y.t0 SEL2.t82 VDD.t3800 VDD.t3799 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2630 a_11386_n25478.t1 mux8_7.NAND4F_2.Y.t10 a_11290_n25478.t1 VSS.t1084 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2631 VSS.t1845 A3.t33 a_n11274_n23075.t0 VSS.t1844 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2632 AND8_0.NOT8_0.A7.t6 B7.t23 VDD.t1415 VDD.t1414 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2633 VDD.t1800 SEL3.t56 a_n4205_3810.t8 VDD.t1799 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2634 VDD.t91 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t11 a_n6611_2026.t2 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2635 VDD.t4457 SEL1.t95 mux8_0.NAND4F_0.C.t2 VDD.t4405 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2636 a_n20557_n7799.t4 MULT_0.4bit_ADDER_1.B3.t15 VDD.t2719 VDD.t2718 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2637 OR8_0.NOT8_0.A3.t2 A3.t34 a_n17677_n19625.t1 VDD.t4115 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2638 mux8_0.NAND4F_1.Y.t6 VSS.t1003 a_9528_762.t1 VSS.t776 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2639 a_n13975_n5154.t3 a_n14155_n5154.t5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t9 VSS.t1875 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2640 mux8_4.NAND4F_4.Y.t4 SEL1.t96 VDD.t4459 VDD.t4458 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2641 a_n10684_n7799.t7 a_n10864_n8419.t5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t9 VDD.t1699 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2642 mux8_3.NAND4F_1.Y.t2 XOR8_0.S2.t13 a_9528_n12822.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2643 a_n20557_n8419.t0 a_n20587_n8445.t7 VSS.t1424 VSS.t1423 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2644 VDD.t13 mux8_6.NAND4F_4.B.t11 mux8_6.NAND4F_4.Y.t8 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2645 VDD.t2610 B2.t30 a_n12314_n21072.t4 VDD.t2609 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2646 NOT8_0.S5.t2 B5.t24 VDD.t3970 VDD.t1011 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2647 VDD.t1016 B0.t33 MULT_0.NAND2_0.Y.t1 VDD.t1015 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2648 VDD.t3177 mux8_2.NAND4F_2.D.t10 mux8_2.NAND4F_2.Y.t5 VDD.t3176 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2649 mux8_7.NAND4F_1.Y.t7 mux8_7.NAND4F_4.B.t10 VDD.t202 VDD.t201 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2650 VDD.t1422 mux8_5.NAND4F_2.Y.t9 mux8_5.NAND4F_8.Y.t3 VDD.t1421 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2651 a_n14751_1406.t1 a_n14781_1380.t5 VSS.t268 VSS.t267 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2652 VSS.t1355 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t12 a_n15907_1406.t4 VSS.t1354 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X2653 VDD.t3459 mux8_4.inv_0.A.t9 Y3.t2 VDD.t3458 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2654 VDD.t1841 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t8 8bit_ADDER_0.C.t1 VDD.t1840 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2655 mux8_1.NAND4F_4.Y.t8 mux8_1.NAND4F_4.B.t9 VDD.t1266 VDD.t1265 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2656 VSS.t1312 a_n12345_n31115.t5 a_n11274_n31661.t4 VSS.t1311 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2657 XOR8_0.S7.t7 a_n12347_n34023.t6 a_n11276_n34281.t4 VSS.t486 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2658 a_n8200_1380.t0 A2.t27 VSS.t254 VSS.t253 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X2659 8bit_ADDER_0.C.t4 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t8 VDD.t2691 VDD.t2690 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2660 mux8_8.NAND4F_0.C.t0 SEL1.t97 VSS.t1979 VSS.t1978 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2661 VSS.t1884 right_shifter_0.buffer_2.inv_1.A.t4 right_shifter_0.S5.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2662 a_n59_1380.t1 SEL3.t57 VDD.t1802 VDD.t1801 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2663 VDD.t218 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t14 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t2 VDD.t217 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2664 a_n15707_n11063.t3 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t15 VDD.t841 VDD.t840 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2665 NOT8_0.S3.t0 B3.t37 VDD.t2118 VDD.t1011 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2666 mux8_8.NAND4F_8.Y.t6 mux8_8.NAND4F_4.Y.t9 a_11386_n30006.t1 VSS.t727 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2667 VDD.t2612 B2.t31 a_n17677_n18225.t5 VDD.t2611 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2668 MULT_0.4bit_ADDER_2.B0.t6 a_n12596_n8419.t5 a_n12416_n7799.t5 VDD.t1839 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2669 a_n10684_n11063.t3 a_n10864_n11683.t6 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t5 VDD.t1538 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2670 a_n13399_n11683.t5 MULT_0.4bit_ADDER_2.B1.t20 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t5 VSS.t972 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2671 VDD.t2614 B2.t32 MULT_0.inv_12.A.t4 VDD.t2613 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2672 S.t0 buffer_0.inv_1.A.t6 VSS.t561 VSS.t560 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2673 a_n13975_n4534.t3 a_n14005_n5180.t7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t5 VDD.t1527 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2674 VSS.t1234 a_n12446_n8445.t4 a_n12416_n8419.t4 VSS.t1233 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2675 VDD.t75 mux8_1.NAND4F_0.C.t11 mux8_1.NAND4F_1.Y.t3 VDD.t74 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2676 left_shifter_0.S2.t1 left_shifter_0.buffer_7.inv_1.A.t6 VDD.t3264 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2677 mux8_3.NAND4F_0.Y.t3 mux8_3.NAND4F_2.D.t14 VDD.t2811 VDD.t2810 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2678 XOR8_0.S5.t10 a_n12345_n28794.t5 a_n11274_n29052.t5 VSS.t944 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2679 a_n21333_1406.t1 a_n21363_1380.t5 VSS.t609 VSS.t608 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2680 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t1 a_n20587_n11709.t6 a_n20557_n11063.t7 VDD.t2431 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2681 mux8_6.inv_0.A.t3 mux8_6.NAND4F_9.Y.t13 a_11865_n34471.t5 VDD.t698 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2682 a_n10786_3810.t9 B3.t38 VDD.t2120 VDD.t2119 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2683 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t10 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t20 a_n1012_1406.t4 VSS.t1080 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2684 VDD.t3802 SEL2.t83 mux8_6.NAND4F_6.Y.t1 VDD.t3801 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2685 a_n12314_n26419.t4 B4.t26 VDD.t3605 VDD.t3604 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2686 NOT8_0.S6.t2 B6.t27 VDD.t3559 VDD.t3558 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2687 a_9528_762.t0 mux8_0.NAND4F_4.B.t11 a_9432_762.t0 VSS.t425 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2688 VDD.t3344 mux8_5.inv_0.A.t8 Y4.t2 VDD.t3343 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2689 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t11 a_n10966_3190.t6 a_n10786_3810.t11 VDD.t3381 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2690 a_n15707_n11063.t9 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t18 VDD.t1280 VDD.t1279 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2691 a_n18422_n11683.t2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t21 mux8_8.A1.t4 VSS.t1676 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2692 VSS.t272 Y0.t7 ZFLAG_0.nor4_0.Y.t3 VSS.t271 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X2693 a_n20659_3810.t9 a_n20113_3164.t7 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t6 VDD.t2689 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2694 mux8_1.NAND4F_6.Y.t3 right_shifter_0.S0.t5 a_8592_n3766.t0 VSS.t433 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2695 a_11386_n3766.t0 mux8_1.NAND4F_6.Y.t9 a_11290_n3766.t0 VSS.t311 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2696 VSS.t1636 B6.t28 a_n12345_n31403.t0 VSS.t1635 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2697 OR8_0.S2.t1 OR8_0.NOT8_0.A2.t9 VDD.t1547 VDD.t315 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2698 NOT8_0.S5.t3 B5.t25 VDD.t3971 VDD.t1013 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2699 VDD.t3525 MULT_0.inv_8.Y.t13 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t4 VDD.t3524 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2700 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t10 a_n8350_1406.t6 a_n8170_1406.t1 VSS.t746 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2701 MULT_0.4bit_ADDER_1.A1.t0 MULT_0.inv_7.A.t9 VSS.t1077 VSS.t1076 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2702 a_n4909_1380.t1 A1.t31 VDD.t4222 VDD.t4221 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2703 a_10459_1690.t1 SEL0.t94 a_10363_1690.t1 VSS.t2014 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2704 a_n13975_n11683.t4 a_n14005_n11709.t4 VSS.t826 VSS.t825 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2705 XOR8_0.S2.t1 B2.t33 a_n11274_n20496.t4 VSS.t1297 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2706 MULT_0.4bit_ADDER_0.B0.t2 MULT_0.NAND2_2.Y.t9 VDD.t1058 VDD.t1056 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2707 MULT_0.4bit_ADDER_1.B1.t4 a_n15887_n5154.t5 a_n15707_n4534.t4 VDD.t2270 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2708 VDD.t254 MULT_0.4bit_ADDER_0.A2.t14 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t0 VDD.t253 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2709 VDD.t1051 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t21 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t0 VDD.t1050 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2710 mux8_7.NAND4F_4.Y.t5 SEL1.t98 VDD.t4461 VDD.t4460 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2711 a_n12345_n20526.t0 A2.t28 VSS.t256 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X2712 a_n7496_3810.t7 a_n6950_3164.t5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t4 VDD.t3986 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2713 VDD.t2721 MULT_0.4bit_ADDER_1.B3.t16 a_n20737_n8419.t1 VDD.t2720 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X2714 VSS.t1870 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t15 a_n18422_n8419.t4 VSS.t1869 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X2715 mux8_3.NAND4F_2.D.t0 SEL2.t84 VSS.t1733 VSS.t1732 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2716 a_7644_n21878.t0 mux8_5.NAND4F_4.B.t9 a_7548_n21878.t0 VSS.t857 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2717 a_n17677_n21025.t1 B4.t27 VDD.t3607 VDD.t3606 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2718 mux8_6.NAND4F_1.Y.t4 mux8_6.NAND4F_4.B.t12 VDD.t2452 VDD.t2451 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2719 VDD.t2112 right_shifter_0.S5.t5 mux8_7.NAND4F_6.Y.t4 VDD.t2111 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2720 VSS.t482 mux8_4.NAND4F_9.Y.t12 mux8_4.inv_0.A.t6 VSS.t481 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X2721 VDD.t1843 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t9 8bit_ADDER_0.C.t2 VDD.t1842 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2722 NOT8_0.S3.t1 B3.t39 VDD.t2121 VDD.t1013 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2723 mux8_3.NAND4F_7.Y.t6 mux8_3.NAND4F_0.C.t10 VDD.t2674 VDD.t2673 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2724 a_n9901_2026.t9 a_n10081_1406.t6 mux8_4.A0.t7 VDD.t1564 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2725 a_16143_n19505.t1 Y5.t6 a_15855_n19505.t1 VDD.t1529 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X2726 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t9 a_n11640_1406.t5 a_n11460_2026.t10 VDD.t1576 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2727 8bit_ADDER_0.C.t5 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t9 VDD.t2693 VDD.t2692 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2728 mux8_1.NAND4F_0.C.t2 SEL1.t99 VDD.t4462 VDD.t4409 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2729 a_n19774_2026.t9 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t17 VDD.t2400 VDD.t2399 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2730 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t3 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t13 VDD.t1118 VDD.t1117 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2731 VSS.t693 B7.t24 NOT8_0.S7.t3 VSS.t692 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2732 XOR8_0.S0.t10 a_n12347_n15041.t6 a_n11276_n15299.t3 VSS.t1693 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2733 a_n21363_1380.t1 A6.t20 VDD.t2824 VDD.t2823 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2734 VDD.t2664 mux8_8.NAND4F_0.C.t12 mux8_8.NAND4F_3.Y.t7 VDD.t2663 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2735 a_n8170_2026.t10 a_n8200_1380.t6 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t3 VDD.t335 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2736 a_n6611_2026.t3 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t17 VDD.t2463 VDD.t2462 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2737 mux8_3.NAND4F_0.Y.t1 MULT_0.S2.t13 a_10459_n11894.t0 VSS.t822 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2738 a_8592_n17350.t1 SEL0.t95 a_8496_n17350.t1 VSS.t2002 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2739 a_10363_763.t0 mux8_0.NAND4F_0.C.t9 a_10267_763.t1 VSS.t316 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2740 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t19 VDD.t2057 VDD.t2056 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2741 a_10363_n17349.t0 mux8_4.NAND4F_0.C.t13 a_10267_n17349.t1 VSS.t1497 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2742 a_n9325_1406.t4 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t20 mux8_4.A0.t2 VSS.t2028 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2743 XOR8_0.S6.t7 a_n12345_n31403.t6 a_n11274_n31661.t1 VSS.t941 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2744 a_11865_n2775.t3 mux8_1.NAND4F_9.Y.t12 mux8_1.inv_0.A.t2 VDD.t1321 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2745 a_n17466_1406.t4 A5.t19 VSS.t190 VSS.t189 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2746 VDD.t2386 AND8_0.NOT8_0.A3.t10 AND8_0.S3.t1 VDD.t676 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2747 a_n16483_1406.t0 a_n16663_1406.t6 mux8_7.A0.t4 VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2748 VSS.t656 MULT_0.4bit_ADDER_0.B1.t10 a_n14155_n5154.t0 VSS.t655 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2749 a_n13975_n11683.t5 a_n14005_n11709.t5 VSS.t828 VSS.t827 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2750 VSS.t452 a_n9155_n11709.t5 a_n9125_n11683.t2 VSS.t451 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2751 mux8_6.NAND4F_0.Y.t0 mux8_6.NAND4F_2.D.t14 VDD.t434 VDD.t433 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2752 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t6 MULT_0.4bit_ADDER_2.B1.t21 VDD.t1901 VDD.t1900 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2753 VDD.t857 mux8_0.NAND4F_4.B.t12 mux8_0.NAND4F_4.Y.t0 VDD.t856 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2754 a_n17296_n5180.t1 MULT_0.4bit_ADDER_0.A2.t15 VDD.t256 VDD.t255 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2755 mux8_4.NAND4F_5.Y.t5 SEL1.t100 VDD.t4464 VDD.t4463 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2756 VSS.t2032 VDD.t4516 left_shifter_0.S0.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2757 a_n6035_1406.t3 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t18 8bit_ADDER_0.S2.t4 VSS.t1251 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2758 VDD.t3211 mux8_2.NAND4F_0.C.t11 mux8_2.NAND4F_7.Y.t8 VDD.t3210 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2759 AND8_0.NOT8_0.A1.t5 B1.t35 VDD.t2365 VDD.t2364 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2760 VDD.t124 mux8_4.NAND4F_2.D.t8 mux8_4.NAND4F_3.Y.t1 VDD.t123 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2761 VSS.t695 B7.t25 a_2463_4914.t4 VSS.t694 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2762 a_7173_4939.t1 V_FLAG_0.XOR2_0.Y.t13 VSS.t1857 VSS.t1856 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2763 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t4 MULT_0.4bit_ADDER_1.A0.t11 VDD.t3195 VDD.t3194 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2764 VDD.t2987 SEL0.t96 mux8_5.NAND4F_2.Y.t7 VDD.t2986 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2765 VDD.t4117 A3.t35 AND8_0.NOT8_0.A3.t3 VDD.t4116 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2766 8bit_ADDER_0.C.t3 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t10 VDD.t1845 VDD.t1844 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2767 mux8_1.NAND4F_5.Y.t8 mux8_1.NAND4F_4.B.t10 VDD.t1268 VDD.t1267 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2768 mux8_8.NAND4F_2.D.t0 SEL2.t85 VSS.t1735 VSS.t1734 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2769 OR8_0.S3.t2 OR8_0.NOT8_0.A3.t9 VDD.t730 VDD.t311 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2770 VDD.t280 right_shifter_0.S7.t5 mux8_6.NAND4F_6.Y.t4 VDD.t279 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2771 VDD.t2695 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t10 8bit_ADDER_0.C.t6 VDD.t2694 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2772 VDD.t1120 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t14 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t2 VDD.t1119 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2773 VDD.t2073 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t8 mux8_6.A1.t2 VDD.t2072 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2774 a_n13975_n4534.t10 MULT_0.4bit_ADDER_0.B1.t11 VDD.t1339 VDD.t1338 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2775 mux8_2.NAND4F_2.Y.t8 OR8_0.S1.t5 VDD.t949 VDD.t948 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2776 VDD.t2110 mux8_2.NAND4F_2.Y.t11 mux8_2.NAND4F_8.Y.t7 VDD.t2109 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2777 a_n23950_3190.t4 B7.t26 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t3 VSS.t696 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2778 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t6 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t18 VDD.t2402 VDD.t2401 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2779 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t11 MULT_0.4bit_ADDER_0.B2.t10 a_n16690_n5154.t5 VSS.t1450 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2780 VDD.t1282 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t19 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t2 VDD.t1281 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2781 mux8_8.NAND4F_2.Y.t8 OR8_0.S6.t6 a_8592_n30006.t1 VSS.t527 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2782 a_n9155_n11709.t1 VSS.t2057 VDD.t1935 VDD.t1934 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2783 mux8_3.NAND4F_4.Y.t6 mux8_3.NAND4F_4.B.t11 VDD.t2532 VDD.t2531 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2784 a_1887_5534.t5 a_1707_4914.t5 V_FLAG_0.XOR2_2.B.t7 VDD.t1846 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2785 a_n14751_2026.t10 A4.t20 VDD.t2192 VDD.t2191 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2786 a_11386_1690.t0 mux8_0.NAND4F_2.Y.t10 a_11290_1690.t1 VSS.t867 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2787 a_10267_763.t0 SEL2.t86 VSS.t1736 VSS.t1437 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2788 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t4 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t20 VDD.t4182 VDD.t4181 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2789 VDD.t3804 SEL2.t87 mux8_2.NAND4F_6.Y.t0 VDD.t3803 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2790 mux8_5.NAND4F_5.Y.t7 SEL1.t101 VDD.t4466 VDD.t4465 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2791 a_n13192_2026.t10 a_n13372_1406.t6 mux8_5.A0.t6 VDD.t2076 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2792 mux8_0.NAND4F_7.Y.t4 VSS.t1001 a_10459_763.t0 VSS.t1002 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2793 a_10267_n16422.t0 mux8_4.NAND4F_2.D.t9 VSS.t59 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2794 a_n11276_n34281.t3 a_n12347_n34023.t7 XOR8_0.S7.t6 VSS.t487 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2795 VDD.t398 A5.t20 AND8_0.NOT8_0.A5.t4 VDD.t397 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2796 a_n3320_2026.t4 a_n3350_1380.t6 8bit_ADDER_0.S1.t4 VDD.t2267 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2797 mux8_4.A1.t9 a_n9305_n11683.t6 a_n9125_n11683.t3 VSS.t1348 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2798 a_8400_n20950.t0 mux8_5.NAND4F_2.D.t12 VSS.t682 VSS.t681 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2799 VDD.t1804 SEL3.t58 a_n7496_3810.t0 VDD.t1803 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2800 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t5 VSS.t2058 VDD.t1933 VDD.t1932 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2801 mux8_6.NAND4F_0.Y.t4 mux8_6.A1.t8 a_10459_n34534.t0 VSS.t199 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2802 VDD.t1341 MULT_0.4bit_ADDER_0.B1.t12 a_n13975_n4534.t9 VDD.t1340 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2803 V_FLAG_0.XOR2_2.Y.t10 a_3313_4914.t6 a_3493_4914.t4 VSS.t542 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2804 a_n19028_n5180.t1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t13 VDD.t2560 VDD.t2559 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2805 a_n18422_n5154.t1 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t19 MULT_0.4bit_ADDER_1.B2.t1 VSS.t240 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2806 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t13 a_n12605_n12716.t1 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2807 mux8_5.NAND4F_4.Y.t5 mux8_5.NAND4F_2.D.t13 VDD.t1379 VDD.t1378 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2808 VDD.t4468 SEL1.t102 mux8_8.NAND4F_4.Y.t5 VDD.t4467 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2809 a_n12616_1406.t1 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t20 mux8_5.A0.t2 VSS.t162 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2810 mux8_1.inv_0.A.t1 mux8_1.NAND4F_9.Y.t13 a_11865_n2775.t4 VDD.t1322 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X2811 a_n17677_n25225.t7 B7.t27 VDD.t1417 VDD.t1416 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X2812 VDD.t3132 mux8_7.NAND4F_2.D.t9 mux8_7.NAND4F_3.Y.t7 VDD.t3131 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2813 OR8_0.NOT8_0.A5.t2 A5.t21 a_n17677_n22425.t6 VDD.t399 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2814 mux8_5.NAND4F_3.Y.t8 mux8_5.A0.t14 a_9528_n20950.t1 VSS.t1541 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2815 VSS.t554 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t15 a_n19198_1406.t1 VSS.t553 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X2816 a_9432_n21878.t0 mux8_5.NAND4F_0.C.t13 a_9336_n21878.t1 VSS.t1664 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2817 VDD.t2075 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t9 mux8_6.A1.t1 VDD.t2074 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2818 XOR8_0.S1.t11 a_n12345_n17857.t7 a_n11274_n18115.t3 VSS.t1247 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2819 VDD.t3259 mux8_4.NAND4F_0.C.t14 mux8_4.NAND4F_0.Y.t3 VDD.t3258 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2820 a_11290_n17350.t1 mux8_4.NAND4F_1.Y.t11 a_11194_n17350.t1 VSS.t967 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2821 VDD.t340 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t18 a_n8170_2026.t1 VDD.t339 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2822 VSS.t1000 VSS.t998 a_n8549_n8419.t5 VSS.t999 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X2823 MULT_0.inv_13.A.t6 A3.t36 a_n22426_n9284.t1 VSS.t1284 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2824 a_n21072_373.t0 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t18 VSS.t1494 VSS.t1400 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2825 a_n15707_n4534.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t19 VDD.t458 VDD.t457 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2826 mux8_2.NAND4F_7.Y.t6 SEL0.t97 VDD.t2985 VDD.t2984 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2827 VDD.t1122 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t16 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t1 VDD.t1121 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2828 a_8592_n30934.t1 SEL0.t98 a_8496_n30934.t1 VSS.t1991 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2829 mux8_7.NAND4F_6.Y.t0 SEL2.t88 VDD.t3806 VDD.t3805 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2830 MULT_0.NAND2_9.Y.t0 A1.t32 a_n24162_n12548.t0 VSS.t1910 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2831 a_10363_n30933.t0 mux8_8.NAND4F_0.C.t13 a_10267_n30933.t1 VSS.t1319 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2832 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t3 a_n10714_n5180.t5 a_n10684_n4534.t0 VDD.t307 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2833 MULT_0.S1.t2 a_n9155_n5180.t5 a_n9125_n4534.t2 VDD.t310 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2834 a_10267_n8193.t0 SEL2.t89 VSS.t1737 VSS.t1474 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2835 VSS.t1800 B5.t26 a_n12345_n28794.t0 VSS.t1799 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2836 VDD.t1128 MULT_0.NAND2_4.Y.t10 MULT_0.4bit_ADDER_0.A0.t1 VDD.t1125 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2837 MULT_0.NAND2_14.Y.t1 A2.t29 VDD.t534 VDD.t533 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2838 VSS.t794 a_n14257_3190.t5 a_n13501_3190.t2 VSS.t793 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2839 VDD.t1075 MULT_0.4bit_ADDER_2.B0.t19 a_n10864_n11683.t0 VDD.t1074 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X2840 XOR8_0.S2.t11 a_n12345_n20814.t5 a_n11274_n21072.t5 VSS.t1427 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2841 a_n18998_n4534.t9 a_n19028_n5180.t3 MULT_0.4bit_ADDER_1.B2.t9 VDD.t2845 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2842 VDD.t126 mux8_4.NAND4F_2.D.t10 mux8_4.NAND4F_4.Y.t1 VDD.t125 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2843 a_9528_n12822.t1 mux8_3.NAND4F_4.B.t12 a_9432_n12822.t0 VSS.t1268 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2844 a_10459_763.t1 SEL0.t99 a_10363_763.t1 VSS.t2014 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2845 VDD.t3609 B4.t28 a_n17677_n21025.t0 VDD.t3608 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2846 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t2 a_n18222_1406.t6 a_n18042_2026.t3 VDD.t3899 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2847 a_n24624_1406.t1 a_n24654_1380.t7 VSS.t1759 VSS.t1758 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2848 mux8_8.NAND4F_5.Y.t5 SEL1.t103 VDD.t4470 VDD.t4469 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2849 mux8_6.NAND4F_4.Y.t7 mux8_6.NAND4F_4.B.t13 VDD.t2454 VDD.t2453 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2850 VDD.t1095 Y7.t7 buffer_0.inv_1.A.t1 VDD.t1094 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2851 VDD.t2367 B1.t36 MULT_0.NAND2_11.Y.t1 VDD.t2366 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2852 mux8_5.NAND4F_8.Y.t4 mux8_5.NAND4F_2.Y.t10 VDD.t1424 VDD.t1423 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2853 MULT_0.inv_14.Y.t1 MULT_0.NAND2_14.Y.t10 VDD.t2635 VDD.t2632 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2854 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t4 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t8 VDD.t3325 VDD.t3324 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2855 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t2 a_n14257_3190.t6 a_n14077_3810.t8 VDD.t1614 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2856 VDD.t4471 SEL1.t104 mux8_1.NAND4F_0.C.t1 VDD.t4409 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2857 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t0 a_n4385_3190.t7 a_n4205_3810.t0 VDD.t3953 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2858 VDD.t2369 B1.t37 MULT_0.NAND2_10.Y.t5 VDD.t2368 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2859 a_5197_5532.t0 a_5017_4912.t5 V_FLAG_0.XOR2_0.Y.t1 VDD.t1906 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2860 a_11386_n30006.t0 mux8_8.NAND4F_2.Y.t11 a_11290_n30006.t1 VSS.t166 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2861 VDD.t3808 SEL2.t90 mux8_4.NAND4F_1.Y.t1 VDD.t3807 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2862 a_11290_n7266.t1 mux8_2.NAND4F_3.Y.t11 a_11194_n7266.t1 VSS.t318 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2863 mux8_7.NAND4F_4.Y.t0 AND8_0.S5.t4 a_7644_n25478.t0 VSS.t242 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2864 a_8592_n7266.t0 SEL0.t100 a_8496_n7266.t1 VSS.t2008 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2865 a_n24162_n11256.t0 A0.t33 VSS.t1131 VSS.t1109 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2866 a_n9931_1380.t0 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t17 VSS.t864 VSS.t863 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X2867 a_n19981_n5154.t3 VSS.t996 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t9 VSS.t997 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2868 VSS.t1931 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t14 a_n11840_n8419.t5 VSS.t1930 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X2869 VDD.t147 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t10 MULT_0.4bit_ADDER_2.B3.t2 VDD.t146 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2870 VDD.t2446 MULT_0.inv_14.Y.t11 a_n17266_n11063.t11 VDD.t2445 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2871 a_11865_1753.t1 mux8_0.NAND4F_8.Y.t13 VDD.t3509 VDD.t3508 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2872 VDD.t192 mux8_7.NAND4F_0.C.t13 mux8_7.NAND4F_0.Y.t1 VDD.t191 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2873 mux8_0.NAND4F_6.Y.t2 SEL1.t105 VDD.t4473 VDD.t4472 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2874 VSS.t1364 a_n12345_n23105.t6 a_n11274_n23651.t5 VSS.t1363 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2875 VDD.t2894 mux8_0.NAND4F_2.D.t10 mux8_0.NAND4F_3.Y.t7 VDD.t2893 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2876 a_n20557_n11063.t8 a_n20587_n11709.t7 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t2 VDD.t2432 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2877 a_n11274_n31661.t0 a_n12345_n31403.t7 XOR8_0.S6.t8 VSS.t942 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2878 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t3 a_n20839_3190.t6 a_n20659_3810.t6 VDD.t4278 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2879 MULT_0.4bit_ADDER_1.B0.t3 a_n12446_n5180.t5 a_n12416_n4534.t10 VDD.t3287 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2880 a_n12416_n11063.t0 a_n12596_n11683.t7 mux8_5.A1.t11 VDD.t1243 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2881 mux8_6.NAND4F_6.Y.t0 SEL2.t91 VDD.t3810 VDD.t3809 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2882 a_n24654_1380.t1 A7.t35 VDD.t3441 VDD.t3440 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2883 VDD.t3561 B6.t29 NOT8_0.S6.t1 VDD.t3560 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2884 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t1 a_n1768_1406.t6 a_n1588_2026.t3 VDD.t582 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2885 mux8_7.A1.t3 a_n15887_n11683.t5 a_n15707_n11063.t11 VDD.t1616 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2886 mux8_8.A1.t6 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t22 a_n18422_n11683.t1 VSS.t1677 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2887 VDD.t2676 mux8_3.NAND4F_0.C.t11 mux8_3.NAND4F_3.Y.t8 VDD.t2675 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2888 VDD.t2371 B1.t38 AND8_0.NOT8_0.A1.t6 VDD.t2370 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2889 a_4069_4914.t4 V_FLAG_0.XOR2_2.B.t18 VSS.t493 VSS.t492 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2890 VDD.t3134 mux8_7.NAND4F_2.D.t10 mux8_7.NAND4F_4.Y.t4 VDD.t3133 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2891 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t6 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t16 a_n19187_n9452.t1 VSS.t1138 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2892 VDD.t3812 SEL2.t92 mux8_5.NAND4F_1.Y.t1 VDD.t3811 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2893 a_7548_n21878.t1 SEL1.t106 a_7452_n21878.t1 VSS.t1950 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2894 VDD.t647 mux8_0.NAND4F_0.C.t10 mux8_0.NAND4F_7.Y.t3 VDD.t646 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2895 VDD.t1998 right_shifter_0.buffer_0.inv_1.A.t5 right_shifter_0.S1.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2896 VDD.t4272 MULT_0.4bit_ADDER_1.A3.t12 a_n20557_n7799.t6 VDD.t4271 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2897 mux8_7.NAND4F_6.Y.t3 right_shifter_0.S5.t6 VDD.t845 VDD.t844 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2898 VSS.t382 a_n13222_1380.t6 a_n13192_1406.t4 VSS.t381 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2899 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t10 a_n11640_1406.t6 a_n11460_1406.t5 VSS.t775 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2900 mux8_4.inv_0.A.t0 mux8_4.NAND4F_8.Y.t10 VSS.t729 VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X2901 VDD.t1541 mux8_2.NAND4F_6.Y.t10 mux8_2.NAND4F_9.Y.t2 VDD.t1540 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2902 V_FLAG_0.NAND2_0.Y.t5 V_FLAG_0.XOR2_0.Y.t14 VDD.t4127 VDD.t4126 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2903 a_n19774_1406.t3 a_n19954_1406.t6 mux8_8.A0.t10 VSS.t804 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2904 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t8 a_n17446_n5154.t7 a_n17266_n4534.t6 VDD.t2429 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2905 VSS.t1888 MULT_0.4bit_ADDER_1.A3.t13 a_n19981_n8419.t3 VSS.t1887 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2906 mux8_2.NAND4F_6.Y.t2 right_shifter_0.S1.t4 VDD.t624 VDD.t623 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2907 a_7452_n2838.t0 mux8_1.NAND4F_2.D.t12 VSS.t856 VSS.t855 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2908 a_15855_n19505.t0 Y5.t7 a_16143_n19505.t0 VDD.t1530 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X2909 8bit_ADDER_0.S1.t7 a_n3500_1406.t5 a_n3320_1406.t4 VSS.t766 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2910 a_11290_n30934.t1 mux8_8.NAND4F_1.Y.t11 a_11194_n30934.t0 VSS.t712 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2911 a_n19981_n5154.t1 MULT_0.4bit_ADDER_0.A3.t11 VSS.t787 VSS.t786 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2912 VSS.t1815 MULT_0.inv_9.Y.t13 a_n13399_n11683.t0 VSS.t1814 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X2913 VDD.t2793 AND8_0.S3.t4 mux8_4.NAND4F_4.Y.t7 VDD.t2792 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2914 VDD.t2534 mux8_3.NAND4F_4.B.t13 mux8_3.NAND4F_5.Y.t4 VDD.t2533 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2915 a_n7594_1406.t3 A2.t30 VSS.t258 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2916 MULT_0.NAND2_11.Y.t0 B1.t39 VDD.t2373 VDD.t2372 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2917 VSS.t1093 B3.t40 a_n12345_n23393.t0 VSS.t1092 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2918 AND8_0.S4.t1 AND8_0.NOT8_0.A4.t10 VDD.t679 VDD.t678 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2919 VDD.t238 MULT_0.NAND2_1.Y.t9 MULT_0.4bit_ADDER_0.B1.t1 VDD.t236 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2920 mux8_8.NAND4F_3.Y.t8 mux8_8.NAND4F_0.C.t14 VDD.t2666 VDD.t2665 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2921 VSS.t1407 a_n19028_n5180.t4 a_n18998_n5154.t4 VSS.t1406 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2922 VDD.t707 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t15 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t4 VDD.t706 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2923 a_10459_n11894.t1 SEL0.t101 a_10363_n11894.t1 VSS.t2015 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2924 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t20 VDD.t1284 VDD.t1283 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2925 a_8496_n17350.t0 SEL1.t107 a_8400_n17350.t1 VSS.t1969 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2926 a_10267_n17349.t0 SEL2.t93 VSS.t1738 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2927 VSS.t910 SEL3.t59 a_n20659_3190.t1 VSS.t909 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2928 a_n9125_n7799.t7 a_n9155_n8445.t5 MULT_0.S2.t1 VDD.t1701 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2929 a_n17266_n5154.t5 a_n17296_n5180.t5 VSS.t1205 VSS.t1204 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X2930 a_n10108_n8419.t1 MULT_0.4bit_ADDER_1.B0.t20 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t3 VSS.t1265 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2931 NOT8_0.S4.t2 B4.t29 VDD.t3610 VDD.t1011 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2932 VDD.t1298 MULT_0.4bit_ADDER_0.A0.t11 a_n10684_n4534.t4 VDD.t1297 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2933 a_n8549_n8419.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t19 MULT_0.S2.t9 VSS.t295 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2934 VDD.t4224 A1.t33 MULT_0.inv_7.A.t4 VDD.t4223 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2935 a_n17005_n9452.t0 MULT_0.4bit_ADDER_1.B2.t20 VSS.t1820 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2936 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t10 a_n14155_n11683.t6 a_n13975_n11683.t0 VSS.t1049 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2937 a_9336_n3766.t0 SEL2.t94 VSS.t1739 VSS.t849 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2938 MULT_0.NAND2_4.Y.t4 A0.t34 VDD.t2230 VDD.t2229 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2939 VDD.t4017 MULT_0.inv_9.Y.t14 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t1 VDD.t4016 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2940 VDD.t3814 SEL2.t95 mux8_4.NAND4F_5.Y.t0 VDD.t3813 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2941 MULT_0.NAND2_10.Y.t3 B1.t40 a_n22426_n4727.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2942 VDD.t2746 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t9 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t5 VDD.t2745 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2943 a_n17677_n22425.t5 A5.t22 OR8_0.NOT8_0.A5.t1 VDD.t400 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2944 VSS.t1656 B4.t30 right_shifter_0.buffer_4.inv_1.A.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2945 a_n10684_n4534.t6 MULT_0.4bit_ADDER_0.B0.t11 VDD.t290 VDD.t289 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2946 a_n9125_n4534.t10 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t20 VDD.t2059 VDD.t2058 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2947 mux8_4.NAND4F_3.Y.t0 mux8_4.NAND4F_2.D.t11 VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2948 a_10363_n3765.t0 mux8_1.NAND4F_0.C.t12 a_10267_n3765.t1 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2949 MULT_0.4bit_ADDER_0.A3.t1 MULT_0.NAND2_11.Y.t10 VDD.t2623 VDD.t2620 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2950 MULT_0.inv_13.A.t0 B2.t34 VDD.t464 VDD.t463 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2951 VDD.t3110 VDD.t3109 right_shifter_0.S7.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2952 VDD.t3305 mux8_6.A0.t19 a_5197_5532.t8 VDD.t3304 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2953 a_n4879_2026.t9 A1.t34 VDD.t4226 VDD.t4225 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2954 VDD.t3816 SEL2.t96 mux8_8.NAND4F_1.Y.t1 VDD.t3815 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2955 VDD.t332 mux8_6.NAND4F_0.C.t12 mux8_6.NAND4F_3.Y.t3 VDD.t331 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2956 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t2 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t9 VDD.t2520 VDD.t2519 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2957 VDD.t731 OR8_0.NOT8_0.A3.t10 OR8_0.S3.t1 VDD.t313 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2958 AND8_0.S1.t1 AND8_0.NOT8_0.A1.t10 VDD.t829 VDD.t828 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2959 MULT_0.4bit_ADDER_1.B2.t7 a_n19178_n5154.t7 a_n18998_n4534.t3 VDD.t693 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2960 mux8_6.NAND4F_6.Y.t3 right_shifter_0.S7.t6 VDD.t282 VDD.t281 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2961 VDD.t2896 mux8_0.NAND4F_2.D.t11 mux8_0.NAND4F_2.Y.t5 VDD.t2895 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2962 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t0 A6.t21 a_n21072_373.t1 VSS.t1400 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2963 a_n12446_n11709.t1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t14 VDD.t2781 VDD.t2780 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2964 XOR8_0.S3.t0 a_n12345_n23393.t6 a_n11274_n23651.t0 VSS.t1610 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2965 VDD.t800 right_shifter_0.buffer_4.inv_1.A.t5 right_shifter_0.S3.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2966 VSS.t1340 a_n19028_n11709.t3 a_n18998_n11683.t2 VSS.t1339 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2967 a_n13975_n4534.t2 MULT_0.4bit_ADDER_0.A1.t10 VDD.t2309 VDD.t2308 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2968 a_n24162_n12548.t1 B3.t41 VSS.t1095 VSS.t1094 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2969 a_n17677_n19625.t0 A3.t37 OR8_0.NOT8_0.A3.t1 VDD.t4118 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X2970 a_1887_4914.t2 a_1857_4888.t5 VSS.t1368 VSS.t1367 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2971 a_n15907_1406.t0 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t18 mux8_7.A0.t9 VSS.t1774 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2972 a_n10108_n11683.t4 MULT_0.inv_8.Y.t14 VSS.t1621 VSS.t1620 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2973 VDD.t503 AND8_0.S5.t5 mux8_7.NAND4F_4.Y.t1 VDD.t502 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X2974 VDD.t4475 SEL1.t108 mux8_3.NAND4F_4.Y.t3 VDD.t4474 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2975 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t21 VDD.t1286 VDD.t1285 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2976 a_n11274_n21072.t0 a_n12345_n20526.t7 VSS.t1216 VSS.t1215 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2977 a_n16822_3164.t1 B5.t27 VDD.t3973 VDD.t3972 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2978 a_n23065_2026.t6 a_n23095_1380.t6 mux8_6.A0.t5 VDD.t1619 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2979 VDD.t759 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t21 a_n3500_1406.t1 VDD.t758 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X2980 a_n6035_1406.t2 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t12 VSS.t41 VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2981 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t5 VSS.t2059 VDD.t1931 VDD.t1930 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2982 mux8_2.NAND4F_6.Y.t3 right_shifter_0.S1.t5 a_8592_n8194.t0 VSS.t304 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2983 a_11386_n8194.t0 mux8_2.NAND4F_6.Y.t11 a_11290_n8194.t0 VSS.t764 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2984 VDD.t3818 SEL2.t97 mux8_5.NAND4F_5.Y.t0 VDD.t3817 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2985 a_8400_n16422.t0 mux8_4.NAND4F_2.D.t12 VSS.t61 VSS.t60 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2986 VSS.t1829 MULT_0.4bit_ADDER_2.B3.t16 a_n20737_n11683.t0 VSS.t1828 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X2987 a_n12416_n7799.t10 a_n12446_n8445.t5 MULT_0.4bit_ADDER_2.B0.t10 VDD.t2434 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X2988 VDD.t2097 mux8_7.NAND4F_6.Y.t10 mux8_7.NAND4F_9.Y.t2 VDD.t2096 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X2989 NOT8_0.S4.t1 B4.t31 VDD.t3611 VDD.t1013 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X2990 a_10459_n34534.t1 SEL0.t102 a_10363_n34534.t1 VSS.t1990 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2991 VDD.t2311 MULT_0.4bit_ADDER_0.A1.t11 a_n13975_n4534.t1 VDD.t2310 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X2992 a_n11840_n8419.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t20 MULT_0.4bit_ADDER_2.B0.t1 VSS.t1766 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2993 VSS.t564 a_n17548_3190.t6 a_n16792_3190.t3 VSS.t563 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2994 VDD.t495 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t20 a_n19178_n5154.t1 VDD.t494 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X2995 VDD.t3686 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t10 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t1 VDD.t3685 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X2996 mux8_4.NAND4F_3.Y.t6 mux8_4.A0.t13 a_9528_n16422.t1 VSS.t16 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2997 a_n11460_2026.t6 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t22 VDD.t622 VDD.t621 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X2998 a_n22489_1406.t0 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t15 VSS.t84 VSS.t83 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2999 mux8_7.NAND4F_3.Y.t8 mux8_7.NAND4F_2.D.t11 VDD.t3136 VDD.t3135 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3000 VDD.t1716 mux8_1.NAND4F_2.D.t13 mux8_1.NAND4F_0.Y.t5 VDD.t1715 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3001 MULT_0.4bit_ADDER_1.A2.t2 MULT_0.inv_12.A.t9 VDD.t813 VDD.t811 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3002 a_9336_n21878.t0 SEL2.t98 VSS.t1740 VSS.t675 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3003 a_9528_n20950.t0 mux8_5.NAND4F_4.B.t10 a_9432_n20950.t1 VSS.t1033 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3004 a_n10786_3810.t1 SEL3.t60 VDD.t1806 VDD.t1805 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3005 VSS.t1637 B6.t30 right_shifter_0.buffer_2.inv_1.A.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3006 mux8_4.NAND4F_0.Y.t2 mux8_4.NAND4F_0.C.t15 VDD.t3261 VDD.t3260 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3007 VDD.t292 MULT_0.4bit_ADDER_0.B0.t12 a_n10864_n5154.t1 VDD.t291 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3008 a_11194_n17350.t0 mux8_4.NAND4F_7.Y.t11 VSS.t1641 VSS.t397 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3009 a_n15707_n4534.t7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t16 VDD.t709 VDD.t708 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3010 left_shifter_0.S7.t1 left_shifter_0.buffer_2.inv_1.A.t7 VDD.t1312 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3011 VSS.t912 SEL3.t61 a_547_1406.t1 VSS.t911 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3012 a_8496_n30934.t0 SEL1.t109 a_8400_n30934.t1 VSS.t1956 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3013 VDD.t1865 left_shifter_0.S3.t5 mux8_4.NAND4F_5.Y.t3 VDD.t1864 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3014 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t9 VDD.t1130 VDD.t1129 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3015 a_10267_n30933.t0 SEL2.t99 VSS.t1741 VSS.t740 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3016 mux8_4.NAND4F_3.Y.t7 mux8_4.A0.t14 VDD.t242 VDD.t241 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3017 a_7548_n3766.t0 SEL1.t110 a_7452_n3766.t1 VSS.t1952 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3018 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t8 VDD.t4003 VDD.t4002 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3019 mux8_0.NAND4F_1.Y.t0 SEL2.t100 VDD.t3820 VDD.t3819 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3020 mux8_8.NAND4F_0.Y.t5 mux8_8.A1.t13 VDD.t2493 VDD.t2492 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3021 VSS.t1133 A0.t35 OR8_0.NOT8_0.A0.t5 VSS.t1132 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X3022 VDD.t1553 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t21 a_n9901_2026.t7 VDD.t1552 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3023 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t10 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t17 a_n17466_1406.t1 VSS.t1431 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3024 VDD.t2232 A0.t36 a_n1588_2026.t1 VDD.t2231 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3025 a_n9125_n8419.t0 a_n9155_n8445.t6 VSS.t947 VSS.t946 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3026 VSS.t74 MULT_0.4bit_ADDER_2.B2.t21 a_n17446_n11683.t0 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X3027 a_11865_n29943.t1 mux8_8.NAND4F_9.Y.t13 mux8_8.inv_0.A.t1 VDD.t1113 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3028 VDD.t1480 mux8_4.NAND4F_8.Y.t11 a_11865_n16359.t3 VDD.t1479 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3029 VDD.t3822 SEL2.t101 mux8_8.NAND4F_5.Y.t0 VDD.t3821 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3030 VSS.t146 a_n9155_n5180.t6 a_n9125_n5154.t1 VSS.t145 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3031 VDD.t4477 SEL1.t111 mux8_6.NAND4F_4.Y.t5 VDD.t4476 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3032 a_10459_n2838.t1 SEL0.t103 a_10363_n2838.t1 VSS.t1997 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3033 MULT_0.NAND2_11.Y.t3 A3.t38 a_n22426_n6019.t1 VSS.t1183 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3034 VDD.t272 mux8_6.NAND4F_6.Y.t10 mux8_6.NAND4F_9.Y.t0 VDD.t271 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3035 VDD.t2826 A6.t22 a_n12314_n31661.t0 VDD.t2825 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X3036 right_shifter_0.S1.t2 right_shifter_0.buffer_0.inv_1.A.t6 VDD.t1999 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3037 a_5197_4912.t3 a_5167_4886.t7 VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3038 VDD.t2723 MULT_0.4bit_ADDER_1.B3.t17 a_n20557_n7799.t3 VDD.t2722 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3039 VSS.t572 a_n12347_n14753.t4 a_n11276_n15299.t1 VSS.t571 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3040 mux8_4.A0.t4 a_n10081_1406.t7 a_n9901_1406.t0 VSS.t2023 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3041 VDD.t4478 SEL1.t112 mux8_2.NAND4F_0.C.t1 VDD.t4353 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3042 VDD.t3150 MULT_0.NAND2_5.Y.t10 MULT_0.4bit_ADDER_0.A1.t1 VDD.t3147 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3043 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t10 a_n10864_n8419.t6 a_n10684_n7799.t8 VDD.t1700 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3044 MULT_0.S2.t6 a_n9305_n8419.t5 a_n9125_n7799.t2 VDD.t1043 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3045 VDD.t1487 left_shifter_0.S4.t5 mux8_5.NAND4F_5.Y.t3 VDD.t1486 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3046 mux8_4.NAND4F_1.Y.t0 SEL2.t102 VDD.t3824 VDD.t3823 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3047 a_7644_n25478.t1 mux8_7.NAND4F_4.B.t11 a_7548_n25478.t1 VSS.t93 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3048 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t3 VSS.t995 a_n9314_n12716.t1 VSS.t428 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3049 VDD.t2473 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t8 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t3 VDD.t2472 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3050 MULT_0.NAND2_0.Y.t0 B0.t34 VDD.t1018 VDD.t1017 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3051 a_n20557_n5154.t3 a_n20587_n5180.t6 VSS.t1061 VSS.t1060 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3052 mux8_2.NAND4F_2.Y.t0 SEL1.t113 VDD.t4480 VDD.t4479 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3053 VSS.t531 a_n10714_n8445.t5 a_n10684_n8419.t1 VSS.t530 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3054 left_shifter_0.buffer_0.inv_1.A.t2 B2.t35 VDD.t465 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3055 VDD.t1104 mux8_1.inv_0.A.t9 Y0.t1 VDD.t1103 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3056 VSS.t735 a_n16513_1380.t6 a_n16483_1406.t3 VSS.t734 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3057 VDD.t1270 mux8_1.NAND4F_4.B.t11 mux8_1.NAND4F_4.Y.t7 VDD.t1269 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3058 VDD.t2983 SEL0.t104 mux8_2.NAND4F_4.B.t1 VDD.t2982 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3059 a_n15737_n8445.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t15 VSS.t1686 VSS.t1685 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3060 a_n17266_n11063.t10 MULT_0.inv_14.Y.t12 VDD.t2448 VDD.t2447 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3061 mux8_7.NAND4F_0.Y.t0 mux8_7.NAND4F_0.C.t14 VDD.t194 VDD.t193 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3062 a_n21333_1406.t4 a_n21513_1406.t6 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t7 VSS.t598 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3063 8bit_ADDER_0.S2.t9 a_n6791_1406.t5 a_n6611_1406.t4 VSS.t1513 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3064 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t8 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t21 a_n4303_1406.t0 VSS.t1864 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3065 a_n11274_n26419.t3 a_n12345_n26161.t6 XOR8_0.S4.t9 VSS.t1624 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3066 Y5.t2 mux8_7.inv_0.A.t9 VDD.t2544 VDD.t2543 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3067 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t1 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t15 VDD.t220 VDD.t219 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3068 a_n12416_n7799.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t21 VDD.t3892 VDD.t3891 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3069 VDD.t4481 SEL1.t114 mux8_5.NAND4F_0.C.t1 VDD.t4355 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3070 VDD.t1482 mux8_4.NAND4F_8.Y.t12 a_11865_n16359.t4 VDD.t1481 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3071 a_n338_3190.t3 a_n368_3164.t6 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t3 VSS.t821 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3072 mux8_7.NAND4F_3.Y.t3 mux8_7.A0.t14 VDD.t608 VDD.t607 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3073 a_n22426_n4727.t0 A2.t31 VSS.t260 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3074 VDD.t2914 MULT_0.4bit_ADDER_0.B2.t11 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t5 VDD.t2913 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3075 MULT_0.inv_12.A.t2 A2.t32 VDD.t536 VDD.t535 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3076 mux8_3.NAND4F_3.Y.t7 mux8_3.NAND4F_0.C.t12 VDD.t2678 VDD.t2677 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3077 a_n18422_n11683.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t23 mux8_8.A1.t5 VSS.t1678 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3078 a_n17368_3190.t0 SEL3.t62 VSS.t914 VSS.t913 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3079 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t7 a_n14155_n5154.t6 a_n13975_n4534.t7 VDD.t4163 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3080 mux8_2.NAND4F_3.Y.t8 mux8_2.NAND4F_4.B.t10 VDD.t3225 VDD.t3224 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3081 mux8_2.NAND4F_8.Y.t4 mux8_2.NAND4F_0.Y.t11 VDD.t4334 VDD.t4333 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3082 a_n12416_n8419.t3 a_n12446_n8445.t6 VSS.t1236 VSS.t1235 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3083 VDD.t3274 MULT_0.4bit_ADDER_1.B1.t18 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t5 VDD.t3273 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3084 Y2.t0 mux8_3.inv_0.A.t10 VSS.t1777 VSS.t1776 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3085 VDD.t604 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t20 a_n9305_n8419.t1 VDD.t603 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3086 VSS.t916 SEL3.t63 a_n23950_3190.t1 VSS.t915 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3087 a_n7496_3190.t4 B2.t36 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t10 VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3088 a_n6800_373.t0 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t19 VSS.t1252 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3089 VSS.t1087 a_n12446_n5180.t6 a_n12416_n5154.t4 VSS.t1086 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3090 VDD.t1132 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t10 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t6 VDD.t1131 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3091 mux8_5.NAND4F_1.Y.t0 SEL2.t103 VDD.t3826 VDD.t3825 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3092 VSS.t507 B0.t35 a_n12347_n15041.t1 VSS.t506 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X3093 a_n17266_n11063.t0 MULT_0.4bit_ADDER_2.B2.t22 VDD.t1816 VDD.t1815 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3094 mux8_8.NAND4F_4.Y.t2 AND8_0.S6.t6 a_7644_n30006.t0 VSS.t613 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3095 right_shifter_0.S1.t1 right_shifter_0.buffer_0.inv_1.A.t7 VDD.t2000 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3096 mux8_3.NAND4F_7.Y.t3 NOT8_0.S2.t5 a_10459_n12821.t0 VSS.t822 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3097 VDD.t2404 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t19 a_n19954_1406.t1 VDD.t2403 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3098 VDD.t2981 SEL0.t105 mux8_7.NAND4F_6.Y.t7 VDD.t2980 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3099 VDD.t2828 A6.t23 a_n21333_2026.t5 VDD.t2827 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3100 right_shifter_0.S7.t2 VDD.t3107 VDD.t3108 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3101 mux8_1.NAND4F_9.Y.t4 mux8_1.NAND4F_5.Y.t11 a_11386_n3766.t1 VSS.t785 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3102 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t9 a_n11723_n12716.t0 VSS.t428 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3103 mux8_1.NAND4F_2.Y.t3 mux8_1.NAND4F_2.D.t14 VDD.t1718 VDD.t1717 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3104 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t0 MULT_0.4bit_ADDER_0.A1.t12 a_n13714_n6187.t0 VSS.t657 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3105 a_11194_n30934.t1 mux8_8.NAND4F_7.Y.t11 VSS.t1283 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3106 a_n17677_n19625.t6 B3.t42 VDD.t2123 VDD.t2122 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3107 VSS.t1801 B5.t28 left_shifter_0.buffer_3.inv_1.A.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3108 OR8_0.NOT8_0.A1.t2 A1.t35 a_n17677_n16825.t6 VDD.t4227 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X3109 mux8_3.NAND4F_5.Y.t5 mux8_3.NAND4F_4.B.t14 VDD.t2536 VDD.t2535 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3110 mux8_4.NAND4F_4.Y.t6 AND8_0.S3.t5 VDD.t2795 VDD.t2794 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3111 a_n15707_n4534.t3 a_n15887_n5154.t6 MULT_0.4bit_ADDER_1.B1.t3 VDD.t2269 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3112 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t4 MULT_0.4bit_ADDER_0.B2.t12 VDD.t2916 VDD.t2915 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3113 a_n18998_n11683.t1 a_n19028_n11709.t4 VSS.t1342 VSS.t1341 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3114 right_shifter_0.S3.t2 right_shifter_0.buffer_4.inv_1.A.t6 VDD.t952 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3115 VDD.t1861 left_shifter_0.S6.t5 mux8_8.NAND4F_5.Y.t3 VDD.t1860 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3116 VDD.t2475 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t9 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t2 VDD.t2474 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3117 VSS.t1182 B1.t41 NOT8_0.S1.t0 VSS.t1181 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3118 a_8592_n11894.t1 SEL0.t106 a_8496_n11894.t1 VSS.t1999 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3119 VSS.t1282 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t14 a_n18422_n5154.t2 VSS.t1281 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3120 MULT_0.NAND2_15.Y.t4 B3.t43 VDD.t2125 VDD.t2124 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3121 a_n11276_n34281.t2 a_n12347_n33735.t6 VSS.t784 VSS.t783 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3122 VDD.t3975 B5.t29 AND8_0.NOT8_0.A5.t0 VDD.t3974 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3123 mux8_5.A1.t1 a_n12446_n11709.t6 a_n12416_n11063.t4 VDD.t4308 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3124 VSS.t422 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t16 a_n15131_n11683.t3 VSS.t421 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3125 left_shifter_0.buffer_4.inv_1.A.t2 B4.t32 VDD.t3612 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3126 mux8_5.A0.t3 a_n13372_1406.t7 a_n13192_1406.t0 VSS.t1075 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3127 VSS.t1847 A3.t39 a_n10884_1406.t1 VSS.t1846 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3128 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t6 a_n10864_n11683.t7 a_n10684_n11683.t0 VSS.t762 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3129 OR8_0.S4.t1 OR8_0.NOT8_0.A4.t10 VDD.t371 VDD.t315 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3130 mux8_4.NAND4F_1.Y.t5 XOR8_0.S3.t14 VDD.t46 VDD.t45 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3131 a_n16672_373.t1 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t19 VSS.t1775 VSS.t1356 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3132 VDD.t4482 SEL1.t115 mux8_8.NAND4F_0.C.t1 VDD.t4357 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3133 OR8_0.NOT8_0.A0.t0 A0.t37 a_n17677_n15425.t0 VDD.t2233 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3134 VDD.t2465 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t20 a_n6791_1406.t1 VDD.t2464 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3135 a_n17266_n11063.t5 a_n17446_n11683.t5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t6 VDD.t1314 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3136 VDD.t3894 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t22 a_n12596_n8419.t1 VDD.t3893 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3137 mux8_7.NAND4F_5.Y.t0 SEL2.t104 VDD.t3828 VDD.t3827 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3138 mux8_7.NAND4F_7.Y.t5 NOT8_0.S5.t6 VDD.t54 VDD.t53 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3139 Y4.t0 mux8_5.inv_0.A.t9 VSS.t1540 VSS.t1539 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3140 VSS.t1556 a_n10966_3190.t7 a_n10210_3190.t3 VSS.t1555 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3141 VDD.t814 MULT_0.inv_12.A.t10 MULT_0.4bit_ADDER_1.A2.t3 VDD.t811 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3142 mux8_8.NAND4F_1.Y.t0 SEL2.t105 VDD.t3830 VDD.t3829 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3143 right_shifter_0.S7.t1 VDD.t3105 VDD.t3106 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3144 a_n13501_3190.t3 a_n13531_3164.t6 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t6 VSS.t1343 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3145 mux8_6.NAND4F_3.Y.t2 mux8_6.NAND4F_0.C.t13 VDD.t566 VDD.t565 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3146 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t21 VDD.t497 VDD.t496 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3147 VDD.t3443 A7.t36 a_n12316_n34281.t0 VDD.t3442 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X3148 VDD.t2979 SEL0.t107 mux8_6.NAND4F_6.Y.t7 VDD.t2978 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3149 VSS.t1927 a_n20839_3190.t7 a_n20083_3190.t0 VSS.t1926 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3150 a_n13192_2026.t7 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t17 VDD.t3951 VDD.t3950 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3151 a_n18998_n11683.t0 a_n19028_n11709.t5 VSS.t1193 VSS.t1192 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3152 right_shifter_0.S3.t1 right_shifter_0.buffer_4.inv_1.A.t7 VDD.t747 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3153 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t15 VDD.t2783 VDD.t2782 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3154 VDD.t2259 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t19 a_n29_2026.t10 VDD.t2258 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3155 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t1 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t10 VDD.t2477 VDD.t2476 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3156 a_n23950_3810.t3 a_n24130_3190.t7 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t4 VDD.t3699 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3157 mux8_7.NAND4F_4.Y.t2 AND8_0.S5.t6 VDD.t505 VDD.t504 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3158 VSS.t1623 MULT_0.inv_8.Y.t15 a_n10108_n11683.t3 VSS.t1622 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3159 VDD.t843 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t17 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t3 VDD.t842 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3160 mux8_5.NAND4F_1.Y.t7 XOR8_0.S4.t14 VDD.t4133 VDD.t4132 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3161 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t20 VDD.t2406 VDD.t2405 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3162 a_9432_n25478.t0 mux8_7.NAND4F_0.C.t15 a_9336_n25478.t0 VSS.t88 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3163 VDD.t1272 mux8_1.NAND4F_4.B.t12 mux8_1.NAND4F_5.Y.t7 VDD.t1271 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3164 VDD.t2080 MULT_0.inv_7.A.t10 MULT_0.4bit_ADDER_1.A1.t1 VDD.t2077 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3165 mux8_8.NAND4F_2.Y.t4 SEL0.t108 VDD.t2977 VDD.t2976 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3166 VSS.t1156 OR8_0.NOT8_0.A5.t10 OR8_0.S5.t0 VSS.t172 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3167 VDD.t1929 VSS.t2060 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t4 VDD.t1928 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3168 mux8_3.NAND4F_9.Y.t2 mux8_3.NAND4F_5.Y.t11 a_11386_n12822.t1 VSS.t461 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3169 VDD.t402 A5.t23 a_n12314_n29052.t3 VDD.t401 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X3170 VDD.t3831 SEL2.t106 mux8_5.NAND4F_2.D.t1 VDD.t3722 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3171 mux8_1.NAND4F_7.Y.t2 mux8_1.NAND4F_0.C.t13 VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3172 VDD.t951 OR8_0.S1.t6 mux8_2.NAND4F_2.Y.t7 VDD.t950 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3173 a_8592_n34534.t1 SEL0.t109 a_8496_n34534.t1 VSS.t2009 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3174 mux8_7.NAND4F_9.Y.t3 mux8_7.NAND4F_6.Y.t11 VDD.t2099 VDD.t2098 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3175 mux8_0.NAND4F_4.B.t0 SEL0.t110 VSS.t2017 VSS.t2016 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3176 a_n14751_1406.t3 a_n14931_1406.t6 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t3 VSS.t1547 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3177 mux8_0.NAND4F_0.Y.t0 mux8_0.NAND4F_0.C.t11 VDD.t649 VDD.t648 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3178 MULT_0.NAND2_0.Y.t3 A3.t40 a_n24213_n2915.t1 VSS.t1848 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3179 a_n11276_n15299.t2 a_n12347_n14753.t5 VSS.t574 VSS.t573 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3180 mux8_0.inv_0.A.t5 mux8_0.NAND4F_9.Y.t13 a_11865_1753.t8 VDD.t3125 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3181 a_n13975_n7799.t11 a_n14005_n8445.t7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t11 VDD.t3622 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3182 VDD.t1498 mux8_8.A0.t14 mux8_8.NAND4F_3.Y.t5 VDD.t1497 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3183 VDD.t1137 buffer_0.inv_1.A.t7 S.t1 VDD.t1094 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3184 mux8_3.NAND4F_0.Y.t2 MULT_0.S2.t14 VDD.t1649 VDD.t1648 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3185 a_7452_n7266.t0 mux8_2.NAND4F_2.D.t11 VSS.t1477 VSS.t1476 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3186 left_shifter_0.buffer_3.inv_1.A.t1 B5.t30 VDD.t3976 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3187 a_9528_n16422.t0 mux8_4.NAND4F_4.B.t11 a_9432_n16422.t1 VSS.t1545 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3188 mux8_2.NAND4F_6.Y.t5 SEL1.t116 VDD.t4484 VDD.t4483 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3189 a_n12314_n21072.t1 A2.t33 VDD.t538 VDD.t537 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3190 VDD.t99 MULT_0.SO.t5 mux8_1.NAND4F_0.Y.t1 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3191 a_11865_n11831.t6 mux8_3.NAND4F_9.Y.t12 mux8_3.inv_0.A.t4 VDD.t2618 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3192 mux8_6.NAND4F_5.Y.t0 SEL2.t107 VDD.t3833 VDD.t3832 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3193 mux8_5.inv_0.A.t1 mux8_5.NAND4F_9.Y.t14 a_11865_n20887.t4 VDD.t690 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X3194 a_11290_n11894.t0 mux8_3.NAND4F_3.Y.t9 a_11194_n11894.t1 VSS.t596 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3195 mux8_4.NAND4F_2.Y.t5 SEL1.t117 VDD.t4486 VDD.t4485 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3196 a_n1588_2026.t11 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t21 VDD.t2095 VDD.t2094 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3197 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t4 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t19 VDD.t3239 VDD.t3238 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3198 VDD.t1927 VSS.t2061 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t4 VDD.t1926 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3199 MULT_0.4bit_ADDER_1.A0.t2 MULT_0.inv_6.A.t9 VDD.t1088 VDD.t1086 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3200 VDD.t2546 mux8_7.inv_0.A.t10 Y5.t1 VDD.t2545 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3201 VDD.t1300 MULT_0.4bit_ADDER_0.A0.t12 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t6 VDD.t1299 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3202 mux8_1.NAND4F_6.Y.t1 SEL2.t108 VDD.t3835 VDD.t3834 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3203 MULT_0.4bit_ADDER_2.B1.t5 a_n15887_n8419.t5 a_n15707_n7799.t4 VDD.t1439 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3204 VDD.t3614 B4.t33 AND8_0.NOT8_0.A4.t0 VDD.t3613 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3205 mux8_4.NAND4F_5.Y.t4 left_shifter_0.S3.t6 VDD.t1867 VDD.t1866 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3206 left_shifter_0.S3.t2 left_shifter_0.buffer_0.inv_1.A.t6 VDD.t1185 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3207 VDD.t2408 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t21 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t4 VDD.t2407 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3208 a_n12316_n15299.t4 a_n12347_n14753.t6 XOR8_0.S0.t4 VDD.t1149 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3209 VDD.t2680 mux8_3.NAND4F_0.C.t13 mux8_3.NAND4F_1.Y.t8 VDD.t2679 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3210 VDD.t3368 mux8_4.NAND4F_4.B.t12 mux8_4.NAND4F_3.Y.t5 VDD.t3367 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3211 VDD.t3616 B4.t34 a_n14077_3810.t3 VDD.t3615 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3212 mux8_1.NAND4F_0.C.t0 SEL1.t118 VSS.t1981 VSS.t1980 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3213 a_n17266_n4534.t10 a_n17296_n5180.t6 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t1 VDD.t2394 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3214 MULT_0.4bit_ADDER_2.B1.t6 a_n15887_n8419.t6 a_n15707_n8419.t2 VSS.t711 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3215 mux8_2.NAND4F_1.Y.t7 mux8_2.NAND4F_4.B.t11 VDD.t3227 VDD.t3226 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3216 mux8_2.NAND4F_9.Y.t0 mux8_2.NAND4F_7.Y.t11 VDD.t1351 VDD.t1350 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3217 VDD.t2975 SEL0.t111 mux8_8.NAND4F_0.Y.t8 VDD.t2974 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3218 VDD.t4005 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t10 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t1 VDD.t4004 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3219 VDD.t2276 V_FLAG_0.XOR2_2.Y.t15 V_FLAG_0.NAND2_0.Y.t3 VDD.t2275 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3220 VSS.t720 a_n19804_1380.t6 a_n19774_1406.t0 VSS.t719 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3221 mux8_8.NAND4F_1.Y.t3 XOR8_0.S6.t14 VDD.t3993 VDD.t3992 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3222 a_n1588_1406.t0 a_n1768_1406.t7 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t3 VSS.t279 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3223 a_n17781_373.t0 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t18 VSS.t1432 VSS.t192 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3224 ZFLAG_0.nor4_1.Y.t0 Y7.t8 a_16431_n19505.t2 VDD.t560 sky130_fd_pr__pfet_01v8 ad=1.3268 pd=9.18 as=0.7062 ps=4.61 w=4.28 l=0.15
X3225 AND8_0.NOT8_0.A3.t0 B3.t44 VDD.t2127 VDD.t2126 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3226 VDD.t2973 SEL0.t112 mux8_1.NAND4F_2.Y.t7 VDD.t2972 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3227 mux8_1.NAND4F_8.Y.t2 mux8_1.NAND4F_2.Y.t9 VDD.t926 VDD.t925 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3228 a_9336_n8194.t0 SEL2.t109 VSS.t1742 VSS.t1470 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3229 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t7 VDD.t1465 VDD.t1464 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3230 mux8_8.inv_0.A.t0 mux8_8.NAND4F_9.Y.t14 a_11865_n29943.t0 VDD.t1114 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3231 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t19 a_n7594_1406.t0 VSS.t159 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3232 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t2 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t13 a_n6800_373.t1 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3233 a_n8549_n8419.t4 VSS.t992 VSS.t994 VSS.t993 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3234 XOR8_0.S5.t9 a_n12345_n28794.t6 a_n12314_n29052.t10 VDD.t1835 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3235 a_n23959_n21227.t1 A5.t24 AND8_0.NOT8_0.A5.t3 VSS.t191 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3236 a_11865_n16359.t0 mux8_4.NAND4F_8.Y.t13 VDD.t1227 VDD.t1226 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3237 VDD.t2971 SEL0.t113 mux8_2.NAND4F_7.Y.t5 VDD.t2970 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3238 a_n6641_1380.t1 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t14 VDD.t93 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3239 mux8_1.NAND4F_4.B.t0 SEL0.t114 VSS.t2021 VSS.t2020 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3240 VSS.t991 VSS.t989 a_n8549_n5154.t1 VSS.t990 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3241 VDD.t3836 SEL2.t110 mux8_8.NAND4F_2.D.t1 VDD.t3724 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3242 VDD.t2194 A4.t21 a_n12314_n26419.t10 VDD.t2193 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X3243 a_10363_n8193.t0 mux8_2.NAND4F_0.C.t12 a_10267_n8193.t1 VSS.t1487 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3244 VSS.t1096 B3.t45 left_shifter_0.buffer_5.inv_1.A.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3245 a_3493_5534.t9 a_3463_4888.t6 V_FLAG_0.XOR2_2.Y.t5 VDD.t489 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3246 mux8_6.NAND4F_9.Y.t1 mux8_6.NAND4F_6.Y.t11 VDD.t274 VDD.t273 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3247 a_n29_2026.t7 a_n59_1380.t7 8bit_ADDER_0.S0.t7 VDD.t2393 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3248 VDD.t2129 B3.t46 a_n17677_n19625.t5 VDD.t2128 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3249 VSS.t460 a_n1094_3190.t6 a_n338_3190.t2 VSS.t459 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3250 a_n13714_n6187.t1 MULT_0.4bit_ADDER_0.B1.t13 VSS.t658 VSS.t657 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3251 VDD.t1288 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t22 a_n15887_n11683.t1 VDD.t1287 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3252 MULT_0.4bit_ADDER_1.B2.t10 a_n19028_n5180.t5 a_n18998_n4534.t10 VDD.t2846 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3253 VDD.t1610 MULT_0.4bit_ADDER_0.A3.t12 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t1 VDD.t1609 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3254 VDD.t466 B2.t37 right_shifter_0.buffer_0.inv_1.A.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3255 mux8_5.NAND4F_5.Y.t4 left_shifter_0.S4.t6 VDD.t1489 VDD.t1488 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3256 VDD.t1702 right_shifter_0.buffer_6.inv_1.A.t5 right_shifter_0.C.t1 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3257 a_n19774_2026.t6 a_n19804_1380.t7 mux8_8.A0.t3 VDD.t1450 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3258 VDD.t1589 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t21 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t1 VDD.t1588 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3259 a_7548_n25478.t0 SEL1.t119 a_7452_n25478.t1 VSS.t1963 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3260 VDD.t468 B2.t38 left_shifter_0.buffer_0.inv_1.A.t1 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3261 mux8_6.NAND4F_0.Y.t5 mux8_6.A1.t9 VDD.t3341 VDD.t3340 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3262 VDD.t3445 A7.t37 a_n24624_2026.t3 VDD.t3444 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3263 VDD.t3335 mux8_8.NAND4F_3.Y.t10 mux8_8.NAND4F_8.Y.t1 VDD.t3334 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3264 mux8_7.NAND4F_2.Y.t2 SEL1.t120 VDD.t4488 VDD.t4487 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3265 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t20 VDD.t3241 VDD.t3240 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3266 VDD.t4229 A1.t36 MULT_0.NAND2_2.Y.t4 VDD.t4228 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3267 a_n9155_n5180.t1 VSS.t2062 VDD.t1925 VDD.t1924 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3268 VDD.t2235 A0.t38 MULT_0.NAND2_3.Y.t2 VDD.t2234 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3269 VDD.t2450 MULT_0.inv_14.Y.t13 a_n17266_n11063.t9 VDD.t2449 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X3270 a_n17296_n8445.t1 MULT_0.4bit_ADDER_1.A2.t13 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3271 VDD.t4120 A3.t41 a_n12314_n23651.t3 VDD.t4119 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X3272 a_n29_1406.t0 a_n209_1406.t6 8bit_ADDER_0.S0.t0 VSS.t1453 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3273 a_11290_n34534.t1 mux8_6.NAND4F_3.Y.t9 a_11194_n34534.t0 VSS.t721 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3274 VDD.t3837 SEL2.t111 mux8_0.NAND4F_2.D.t1 VDD.t3727 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3275 MULT_0.NAND2_10.Y.t4 B1.t42 VDD.t2375 VDD.t2374 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3276 VDD.t470 B2.t39 MULT_0.inv_6.A.t1 VDD.t469 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3277 mux8_0.NAND4F_8.Y.t1 mux8_0.NAND4F_3.Y.t11 VDD.t375 VDD.t374 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3278 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t0 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t13 a_n16672_373.t0 VSS.t1356 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3279 VDD.t1020 B0.t36 AND8_0.NOT8_0.A0.t1 VDD.t1019 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3280 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t8 VDD.t1467 VDD.t1466 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3281 mux8_0.NAND4F_2.Y.t7 SEL0.t115 VDD.t2969 VDD.t2968 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3282 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t3 VSS.t987 a_n9314_n6187.t1 VSS.t988 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3283 VDD.t204 mux8_7.NAND4F_4.B.t12 mux8_7.NAND4F_3.Y.t6 VDD.t203 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3284 left_shifter_0.S5.t2 left_shifter_0.buffer_4.inv_1.A.t6 VDD.t2062 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3285 a_11865_n16359.t1 mux8_4.NAND4F_8.Y.t14 VDD.t1229 VDD.t1228 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X3286 a_n17677_n22425.t1 B5.t31 VDD.t3978 VDD.t3977 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3287 a_n11840_n8419.t4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t15 VSS.t1933 VSS.t1932 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3288 VSS.t1401 A6.t24 OR8_0.NOT8_0.A6.t5 VSS.t177 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X3289 VDD.t2898 mux8_0.NAND4F_2.D.t12 mux8_0.NAND4F_4.Y.t2 VDD.t2897 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3290 VDD.t4061 MULT_0.4bit_ADDER_2.B3.t17 a_n20557_n11063.t1 VDD.t4060 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3291 a_n11274_n18115.t2 a_n12345_n17569.t5 VSS.t644 VSS.t643 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3292 a_n13975_n7799.t7 MULT_0.4bit_ADDER_1.B1.t19 VDD.t3276 VDD.t3275 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3293 VSS.t97 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t16 a_n11840_n5154.t1 VSS.t96 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3294 mux8_3.NAND4F_6.Y.t2 right_shifter_0.S2.t6 a_8592_n12822.t0 VSS.t562 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3295 V_FLAG_0.XOR2_2.B.t4 a_1707_4914.t6 a_1887_4914.t0 VSS.t410 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3296 VSS.t1120 A4.t22 a_n14175_1406.t0 VSS.t1119 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3297 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t5 a_n17446_n11683.t6 a_n17266_n11063.t4 VDD.t1315 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3298 a_7644_n30006.t1 mux8_8.NAND4F_4.B.t13 a_7548_n30006.t0 VSS.t1466 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3299 a_10459_n12821.t1 SEL0.t116 a_10363_n12821.t1 VSS.t2015 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3300 mux8_6.A0.t9 a_n23245_1406.t6 a_n23065_2026.t9 VDD.t2489 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3301 VSS.t1912 A1.t37 a_n4303_1406.t3 VSS.t1911 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3302 MULT_0.inv_6.A.t0 B2.t40 VDD.t472 VDD.t471 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3303 8bit_ADDER_0.S1.t6 a_n3500_1406.t6 a_n3320_1406.t5 VSS.t767 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3304 VSS.t918 SEL3.t64 a_n14257_3190.t0 VSS.t917 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X3305 a_11865_n16359.t6 mux8_4.NAND4F_9.Y.t13 mux8_4.inv_0.A.t2 VDD.t963 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3306 VDD.t4490 SEL1.t121 mux8_3.NAND4F_5.Y.t2 VDD.t4489 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3307 mux8_8.NAND4F_5.Y.t4 left_shifter_0.S6.t6 VDD.t1863 VDD.t1862 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3308 mux8_4.NAND4F_6.Y.t5 SEL1.t122 VDD.t4492 VDD.t4491 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3309 VDD.t3839 SEL2.t112 mux8_4.NAND4F_7.Y.t1 VDD.t3838 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3310 a_n16792_3190.t0 a_n16822_3164.t6 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t0 VSS.t1411 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3311 VDD.t3243 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t21 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t6 VDD.t3242 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3312 VDD.t3278 MULT_0.4bit_ADDER_1.B1.t20 a_n13975_n7799.t8 VDD.t3277 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3313 a_7548_n8194.t0 SEL1.t123 a_7452_n8194.t1 VSS.t1959 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3314 a_8496_n11894.t0 SEL1.t124 a_8400_n11894.t1 VSS.t1965 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3315 VDD.t3841 SEL2.t113 mux8_0.NAND4F_6.Y.t1 VDD.t3840 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3316 VDD.t4231 A1.t38 a_n12314_n18115.t6 VDD.t4230 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X3317 a_n17266_n4534.t5 MULT_0.4bit_ADDER_0.B2.t13 VDD.t2918 VDD.t2917 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3318 mux8_2.NAND4F_0.C.t0 SEL1.t125 VSS.t1983 VSS.t1982 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3319 a_n19028_n8445.t1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t17 VDD.t4161 VDD.t4160 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3320 VDD.t626 right_shifter_0.S1.t6 mux8_2.NAND4F_6.Y.t4 VDD.t625 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3321 VDD.t3487 AND8_0.NOT8_0.A7.t9 AND8_0.S7.t2 VDD.t3486 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3322 a_n16483_2026.t3 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t14 VDD.t2755 VDD.t2754 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3323 VSS.t1403 A6.t25 a_n20757_1406.t3 VSS.t1402 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3324 VDD.t95 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t15 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t3 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3325 VDD.t3937 MULT_0.4bit_ADDER_1.A3.t14 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t4 VDD.t3936 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3326 mux8_6.A0.t2 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t23 a_n22489_1406.t2 VSS.t1605 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3327 a_n12416_n11063.t3 a_n12446_n11709.t7 mux8_5.A1.t0 VDD.t4309 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3328 VDD.t3617 B4.t35 left_shifter_0.buffer_4.inv_1.A.t1 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3329 a_n3629_3190.t5 a_n3659_3164.t6 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t7 VSS.t605 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3330 VDD.t1808 SEL3.t65 a_n20659_3810.t0 VDD.t1807 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3331 VSS.t789 MULT_0.4bit_ADDER_0.A3.t13 a_n19981_n5154.t0 VSS.t788 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3332 MULT_0.4bit_ADDER_1.B3.t4 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t10 VDD.t4330 VDD.t4329 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3333 a_n10108_n11683.t0 MULT_0.4bit_ADDER_2.B0.t20 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t0 VSS.t528 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3334 a_n3320_2026.t6 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t17 VDD.t2631 VDD.t2630 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3335 mux8_2.NAND4F_4.B.t0 SEL0.t117 VSS.t2019 VSS.t2018 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3336 a_10459_n7266.t0 SEL0.t118 a_10363_n7266.t1 VSS.t1998 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3337 VDD.t3370 mux8_4.NAND4F_4.B.t13 mux8_4.NAND4F_1.Y.t8 VDD.t3369 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3338 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t17 a_n12605_n6187.t0 VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3339 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t20 VDD.t460 VDD.t459 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3340 a_n15014_n9452.t1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t10 VSS.t1823 VSS.t1822 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3341 VDD.t2967 SEL0.t119 mux8_1.NAND4F_6.Y.t7 VDD.t2966 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3342 mux8_1.NAND4F_9.Y.t1 mux8_1.NAND4F_6.Y.t10 VDD.t631 VDD.t630 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3343 VDD.t540 A2.t34 a_n12314_n21072.t0 VDD.t539 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3344 VDD.t171 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t16 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t4 VDD.t170 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3345 a_n15707_n7799.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t19 VDD.t673 VDD.t672 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3346 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t4 a_n17446_n11683.t7 a_n17266_n11063.t3 VDD.t1313 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3347 VSS.t1531 MULT_0.inv_15.Y.t11 a_n19981_n11683.t4 VSS.t1530 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3348 mux8_7.NAND4F_4.B.t2 SEL0.t120 VDD.t2965 VDD.t2951 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3349 mux8_0.NAND4F_7.Y.t2 mux8_0.NAND4F_0.C.t12 VDD.t651 VDD.t650 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3350 mux8_3.NAND4F_2.Y.t7 SEL0.t121 VDD.t2964 VDD.t2963 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3351 a_n23374_3190.t5 a_n23404_3164.t6 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t10 VSS.t1210 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3352 mux8_0.NAND4F_5.Y.t7 SEL1.t126 VDD.t4494 VDD.t4493 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3353 VDD.t2962 SEL0.t122 mux8_7.NAND4F_7.Y.t8 VDD.t2961 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3354 VSS.t479 a_n11490_1380.t6 a_n11460_1406.t0 VSS.t478 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3355 VSS.t920 SEL3.t66 a_n1094_3190.t0 VSS.t919 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X3356 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t6 a_n10714_n8445.t6 a_n10684_n7799.t1 VDD.t1081 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3357 MULT_0.S2.t0 a_n9155_n8445.t7 a_n9125_n7799.t8 VDD.t1836 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3358 mux8_5.NAND4F_6.Y.t3 SEL1.t127 VDD.t4496 VDD.t4495 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3359 a_n18042_1406.t3 a_n18222_1406.t7 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t5 VSS.t1769 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3360 VDD.t1089 MULT_0.inv_6.A.t10 MULT_0.4bit_ADDER_1.A0.t3 VDD.t1086 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3361 mux8_5.NAND4F_8.Y.t2 mux8_5.NAND4F_4.Y.t11 a_11386_n20950.t0 VSS.t577 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3362 VDD.t1522 mux8_2.inv_0.A.t9 Y1.t2 VDD.t1521 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3363 a_n12416_n11063.t7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t21 VDD.t2017 VDD.t2016 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3364 a_n15707_n11683.t1 a_n15887_n11683.t6 mux8_7.A1.t2 VSS.t796 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3365 VDD.t3843 SEL2.t114 mux8_5.NAND4F_7.Y.t1 VDD.t3842 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3366 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t11 a_n10864_n8419.t7 a_n10684_n8419.t3 VSS.t845 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3367 MULT_0.S2.t7 a_n9305_n8419.t6 a_n9125_n8419.t4 VSS.t518 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3368 a_n10684_n4534.t5 MULT_0.4bit_ADDER_0.A0.t13 VDD.t1302 VDD.t1301 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3369 a_n18998_n7799.t7 a_n19028_n8445.t5 MULT_0.4bit_ADDER_2.B2.t10 VDD.t1345 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3370 a_9432_n3766.t0 mux8_1.NAND4F_0.C.t14 a_9336_n3766.t1 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3371 a_n10108_n5154.t3 MULT_0.4bit_ADDER_0.B0.t13 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t6 VSS.t135 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3372 VDD.t3 8bit_ADDER_0.S2.t14 mux8_3.NAND4F_3.Y.t1 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3373 mux8_8.A1.t3 a_n19178_n11683.t7 a_n18998_n11683.t3 VSS.t770 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3374 XOR8_0.S0.t5 a_n12347_n14753.t7 a_n12316_n15299.t5 VDD.t1150 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3375 a_n8549_n5154.t5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t21 MULT_0.S1.t5 VSS.t1072 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3376 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t10 VDD.t2218 VDD.t2217 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3377 VDD.t2785 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t16 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t6 VDD.t2784 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3378 OR8_0.NOT8_0.A7.t1 A7.t38 a_n17677_n25225.t1 VDD.t3446 sky130_fd_pr__pfet_01v8 ad=0.3968 pd=3.18 as=0.2112 ps=1.61 w=1.28 l=0.15
X3379 a_11865_n7203.t0 mux8_2.NAND4F_8.Y.t13 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3380 VDD.t474 B2.t41 MULT_0.inv_13.A.t1 VDD.t473 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3381 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t9 a_n8432_n12716.t1 VSS.t428 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3382 VDD.t1993 mux8_5.NAND4F_4.B.t11 mux8_5.NAND4F_1.Y.t5 VDD.t1992 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3383 a_n4879_2026.t5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t22 VDD.t4145 VDD.t4144 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3384 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t3 A5.t25 a_n17781_373.t1 VSS.t192 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3385 V_FLAG_0.XOR2_0.Y.t2 a_5017_4912.t6 a_5197_4912.t0 VSS.t974 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3386 a_9336_n25478.t1 mux8_7.NAND4F_2.D.t12 VSS.t1463 VSS.t1462 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3387 a_n18998_n4534.t1 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t22 VDD.t499 VDD.t498 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3388 a_n12314_n29052.t0 B5.t32 VDD.t3980 VDD.t3979 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3389 VDD.t4498 SEL1.t128 mux8_8.NAND4F_2.Y.t2 VDD.t4497 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3390 VDD.t1463 ZFLAG_0.NAND2_0.Y.t10 Z.t1 VDD.t1462 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3391 VDD.t83 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t16 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t0 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3392 a_11386_n12822.t0 mux8_3.NAND4F_6.Y.t11 a_11290_n12822.t0 VSS.t612 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3393 a_n22426_n6019.t0 B1.t43 VSS.t1184 VSS.t1183 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3394 a_n12314_n26419.t11 A4.t23 VDD.t2196 VDD.t2195 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3395 a_n24048_1406.t4 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t21 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t10 VSS.t1671 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3396 VDD.t2313 MULT_0.4bit_ADDER_0.A1.t13 a_n13975_n4534.t0 VDD.t2312 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3397 mux8_2.NAND4F_3.Y.t2 mux8_2.NAND4F_2.D.t12 VDD.t3179 VDD.t3178 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3398 a_n12416_n8419.t1 a_n12596_n8419.t6 MULT_0.4bit_ADDER_2.B0.t7 VSS.t949 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3399 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t6 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t21 VDD.t2467 VDD.t2466 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3400 mux8_4.A1.t1 a_n9155_n11709.t6 a_n9125_n11063.t1 VDD.t906 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3401 a_8496_n34534.t0 SEL1.t129 a_8400_n34534.t1 VSS.t1972 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3402 VDD.t3982 B5.t33 a_n17368_3810.t6 VDD.t3981 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3403 MULT_0.NAND2_3.Y.t4 B0.t37 VDD.t1022 VDD.t1021 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3404 VDD.t2920 MULT_0.4bit_ADDER_0.B2.t14 a_n17266_n4534.t4 VDD.t2919 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3405 a_n6611_1406.t1 a_n6641_1380.t6 VSS.t439 VSS.t438 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3406 a_n4879_1406.t0 a_n5059_1406.t7 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t4 VSS.t576 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3407 VDD.t2960 SEL0.t123 mux8_3.NAND4F_0.Y.t8 VDD.t2959 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3408 OR8_0.NOT8_0.A6.t0 A6.t26 a_n17677_n23825.t2 VDD.t2829 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3409 mux8_2.NAND4F_4.Y.t5 mux8_2.NAND4F_2.D.t13 VDD.t3181 VDD.t3180 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3410 mux8_2.NAND4F_9.Y.t5 mux8_2.NAND4F_5.Y.t11 a_11386_n8194.t1 VSS.t454 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3411 mux8_3.inv_0.A.t5 mux8_3.NAND4F_9.Y.t13 a_11865_n11831.t5 VDD.t2619 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3412 VSS.t1273 left_shifter_0.buffer_5.inv_1.A.t6 left_shifter_0.S4.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3413 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t3 MULT_0.inv_14.Y.t14 a_n17005_n12716.t1 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3414 a_5197_5532.t11 A7.t39 VDD.t3448 VDD.t3447 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3415 a_8400_n3766.t0 SEL2.t115 VSS.t1743 VSS.t851 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3416 VDD.t442 MULT_0.NAND2_10.Y.t10 MULT_0.4bit_ADDER_0.A2.t3 VDD.t439 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3417 right_shifter_0.buffer_0.inv_1.A.t2 B2.t42 VDD.t475 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3418 MULT_0.4bit_ADDER_2.B0.t11 a_n12446_n8445.t7 a_n12416_n7799.t11 VDD.t3382 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3419 VDD.t2198 A4.t24 AND8_0.NOT8_0.A4.t6 VDD.t2197 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3420 VSS.t1185 B1.t44 left_shifter_0.buffer_7.inv_1.A.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3421 VDD.t130 mux8_4.NAND4F_2.D.t13 mux8_4.NAND4F_2.Y.t1 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3422 a_n10714_n8445.t0 MULT_0.4bit_ADDER_1.A0.t12 VSS.t1483 VSS.t1482 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3423 a_11194_n11894.t0 mux8_3.NAND4F_0.Y.t9 VSS.t723 VSS.t722 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3424 OR8_0.S0.t3 OR8_0.NOT8_0.A0.t10 VDD.t316 VDD.t315 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3425 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t9 B0.t38 a_n914_3190.t3 VSS.t508 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3426 a_n10684_n11683.t4 a_n10714_n11709.t6 VSS.t1038 VSS.t1037 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3427 a_9432_n30006.t1 mux8_8.NAND4F_0.C.t15 a_9336_n30006.t0 VSS.t1320 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3428 left_shifter_0.buffer_1.inv_1.A.t2 B7.t28 VDD.t1418 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3429 right_shifter_0.C.t2 right_shifter_0.buffer_6.inv_1.A.t6 VDD.t1703 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3430 MULT_0.4bit_ADDER_2.B0.t8 a_n12596_n8419.t7 a_n12416_n8419.t0 VSS.t950 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3431 mux8_8.NAND4F_6.Y.t5 SEL1.t130 VDD.t4500 VDD.t4499 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3432 mux8_6.NAND4F_2.Y.t7 SEL0.t124 VDD.t2958 VDD.t2957 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3433 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t1 MULT_0.4bit_ADDER_2.B0.t21 VDD.t1077 VDD.t1076 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3434 VDD.t3845 SEL2.t116 mux8_8.NAND4F_7.Y.t1 VDD.t3844 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3435 VDD.t1023 B0.t39 right_shifter_0.buffer_6.inv_1.A.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3436 a_n11840_n5154.t3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t21 MULT_0.4bit_ADDER_1.B0.t9 VSS.t1882 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3437 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t6 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t8 VDD.t4266 VDD.t4265 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3438 mux8_7.A0.t5 a_n16663_1406.t7 a_n16483_2026.t2 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3439 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t2 a_n14781_1380.t6 a_n14751_2026.t2 VDD.t559 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3440 VDD.t728 MULT_0.NAND2_8.Y.t10 MULT_0.inv_8.Y.t3 VDD.t725 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3441 VDD.t1186 left_shifter_0.buffer_0.inv_1.A.t7 left_shifter_0.S3.t1 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3442 AND8_0.NOT8_0.A0.t0 B0.t40 VDD.t1025 VDD.t1024 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3443 VDD.t3511 mux8_0.NAND4F_8.Y.t14 a_11865_1753.t0 VDD.t3510 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3444 a_n21333_2026.t11 a_n21363_1380.t6 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t11 VDD.t1217 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3445 VDD.t4233 A1.t39 a_n4879_2026.t8 VDD.t4232 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3446 a_n9314_n6187.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t22 VSS.t1073 VSS.t988 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3447 VDD.t1381 mux8_5.NAND4F_2.D.t14 mux8_5.NAND4F_0.Y.t5 VDD.t1380 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3448 mux8_4.NAND4F_3.Y.t4 mux8_4.NAND4F_4.B.t14 VDD.t3372 VDD.t3371 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3449 mux8_3.NAND4F_1.Y.t7 mux8_3.NAND4F_0.C.t14 VDD.t2682 VDD.t2681 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3450 8bit_ADDER_0.S2.t8 a_n6791_1406.t6 a_n6611_2026.t7 VDD.t1231 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3451 mux8_8.NAND4F_0.Y.t7 SEL0.t125 VDD.t2956 VDD.t2955 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3452 VDD.t3984 B5.t34 a_n17677_n22425.t0 VDD.t3983 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3453 VDD.t3164 mux8_8.NAND4F_4.B.t14 mux8_8.NAND4F_1.Y.t6 VDD.t3163 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3454 VDD.t2831 A6.t27 AND8_0.NOT8_0.A6.t2 VDD.t2830 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3455 VDD.t1726 NOT8_0.S2.t6 mux8_3.NAND4F_7.Y.t4 VDD.t1725 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3456 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t1 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t17 VDD.t85 VDD.t84 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3457 a_9528_n3766.t1 mux8_1.NAND4F_4.B.t13 a_9432_n3766.t1 VSS.t627 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3458 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t11 a_n17446_n8419.t7 a_n17266_n7799.t8 VDD.t1040 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3459 VDD.t3307 mux8_6.A0.t20 mux8_6.NAND4F_3.Y.t7 VDD.t3306 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3460 a_16431_n19505.t1 Y7.t9 ZFLAG_0.nor4_1.Y.t2 VDD.t561 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X3461 a_16143_n18523.t5 Y2.t6 a_15855_n18523.t3 VDD.t1528 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X3462 VDD.t1192 mux8_3.NAND4F_3.Y.t10 mux8_3.NAND4F_8.Y.t0 VDD.t1191 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3463 VDD.t1469 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t9 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t2 VDD.t1468 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3464 a_11865_n29943.t9 mux8_8.NAND4F_8.Y.t14 VDD.t743 VDD.t742 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3465 a_4069_4914.t0 SEL3.t67 V_FLAG_0.XOR2_2.Y.t0 VSS.t921 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3466 VDD.t2469 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t22 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t5 VDD.t2468 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3467 VDD.t711 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t17 a_n15707_n4534.t6 VDD.t710 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3468 a_n12314_n31661.t3 B6.t31 VDD.t3563 VDD.t3562 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3469 a_n12316_n34281.t9 a_n12347_n33735.t7 XOR8_0.S7.t2 VDD.t1596 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3470 a_n15737_n11709.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t18 VSS.t424 VSS.t423 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3471 MULT_0.inv_13.A.t2 B2.t43 VDD.t477 VDD.t476 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3472 a_7644_n3766.t1 mux8_1.NAND4F_4.B.t14 a_7548_n3766.t1 VSS.t628 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3473 a_n17677_n16825.t5 A1.t40 OR8_0.NOT8_0.A1.t1 VDD.t4234 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3474 a_7452_n17350.t0 SEL2.t117 VSS.t1744 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3475 right_shifter_0.buffer_0.inv_1.A.t1 B2.t44 VDD.t478 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3476 a_n10884_1406.t3 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t23 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t2 VSS.t303 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3477 MULT_0.4bit_ADDER_0.B2.t3 MULT_0.NAND2_0.Y.t10 VDD.t1205 VDD.t1157 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3478 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t10 a_n8432_n6187.t0 VSS.t101 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3479 right_shifter_0.C.t3 right_shifter_0.buffer_6.inv_1.A.t7 VDD.t1704 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3480 a_n9125_n5154.t2 a_n9155_n5180.t7 VSS.t148 VSS.t147 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3481 a_n14005_n8445.t1 MULT_0.4bit_ADDER_1.A1.t11 VSS.t51 VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3482 MULT_0.NAND2_15.Y.t0 A3.t42 a_n22425_n12548.t0 VSS.t1849 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3483 mux8_1.NAND4F_0.Y.t2 MULT_0.SO.t6 a_10459_n2838.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3484 a_n18998_n8419.t3 a_n19028_n8445.t6 VSS.t664 VSS.t663 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3485 XOR8_0.S1.t2 a_n12345_n17569.t6 a_n12314_n18115.t4 VDD.t1304 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3486 a_n12314_n29052.t7 a_n12345_n28506.t7 XOR8_0.S5.t6 VDD.t1819 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3487 mux8_8.NAND4F_8.Y.t0 mux8_8.NAND4F_3.Y.t11 VDD.t3337 VDD.t3336 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3488 VDD.t2954 SEL0.t126 mux8_6.NAND4F_0.Y.t8 VDD.t2953 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3489 VDD.t3138 mux8_7.NAND4F_2.D.t13 mux8_7.NAND4F_2.Y.t7 VDD.t3137 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3490 VDD.t3197 MULT_0.4bit_ADDER_1.A0.t13 a_n10684_n7799.t10 VDD.t3196 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X3491 mux8_5.NAND4F_2.Y.t4 OR8_0.S4.t6 a_8592_n20950.t0 VSS.t87 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3492 VSS.t409 left_shifter_0.buffer_3.inv_1.A.t6 left_shifter_0.S6.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3493 VDD.t3183 mux8_2.NAND4F_2.D.t14 mux8_2.NAND4F_4.Y.t6 VDD.t3182 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3494 VSS.t1485 MULT_0.4bit_ADDER_1.A0.t14 a_n10108_n8419.t3 VSS.t1484 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3495 VSS.t923 SEL3.t68 a_n17548_3190.t0 VSS.t922 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X3496 VDD.t542 A2.t35 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t5 VDD.t541 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3497 a_11194_n34534.t1 mux8_6.NAND4F_0.Y.t9 VSS.t427 VSS.t197 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3498 a_n10684_n7799.t4 MULT_0.4bit_ADDER_1.B0.t21 VDD.t2508 VDD.t2507 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3499 a_n9125_n7799.t3 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t22 VDD.t1591 VDD.t1590 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3500 a_n12605_n6187.t1 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t22 VSS.t1883 VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3501 OR8_0.NOT8_0.A1.t0 B1.t45 VSS.t1187 VSS.t1186 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X3502 VDD.t2562 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t15 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t2 VDD.t2561 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3503 VDD.t2419 Y3.t5 a_15855_n18523.t2 VDD.t2001 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X3504 VSS.t925 SEL3.t69 a_n10786_3190.t0 VSS.t924 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3505 a_n10684_n8419.t0 a_n10714_n8445.t7 VSS.t533 VSS.t532 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3506 VDD.t1698 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t10 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t6 VDD.t1697 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3507 XOR8_0.S2.t6 a_n12345_n20814.t6 a_n12314_n21072.t9 VDD.t1236 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3508 ZFLAG_0.NAND2_0.Y.t4 ZFLAG_0.nor4_1.Y.t8 a_17528_n18777.t0 VSS.t1195 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3509 a_1857_4888.t0 B7.t29 VSS.t582 VSS.t581 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3510 MULT_0.4bit_ADDER_2.B2.t4 a_n19178_n8419.t6 a_n18998_n7799.t2 VDD.t277 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3511 mux8_7.NAND4F_3.Y.t5 mux8_7.NAND4F_4.B.t13 VDD.t206 VDD.t205 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3512 VDD.t410 OR8_0.S3.t4 mux8_4.NAND4F_2.Y.t4 VDD.t409 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3513 a_n914_3810.t11 a_n368_3164.t7 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t6 VDD.t2081 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3514 a_n23404_3164.t0 B7.t30 VSS.t584 VSS.t583 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3515 VDD.t4122 A3.t43 a_n11460_2026.t3 VDD.t4121 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X3516 VDD.t2952 SEL0.t127 mux8_7.NAND4F_4.B.t1 VDD.t2951 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3517 VDD.t2063 left_shifter_0.buffer_4.inv_1.A.t7 left_shifter_0.S5.t3 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3518 a_n17368_3810.t0 SEL3.t70 VDD.t1810 VDD.t1809 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3519 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t4 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t23 VDD.t2471 VDD.t2470 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3520 VSS.t142 a_n10714_n5180.t6 a_n10684_n5154.t1 VSS.t141 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3521 MULT_0.NAND2_8.Y.t0 A0.t39 VDD.t2237 VDD.t2236 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3522 VDD.t2105 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t10 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t6 VDD.t2104 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3523 a_n19774_2026.t1 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t17 VDD.t1124 VDD.t1123 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3524 VDD.t4268 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t9 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t5 VDD.t4267 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3525 left_shifter_0.S4.t1 left_shifter_0.buffer_5.inv_1.A.t7 VDD.t2553 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3526 a_n13975_n7799.t0 MULT_0.4bit_ADDER_1.A1.t12 VDD.t112 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3527 a_n20557_n11063.t0 MULT_0.4bit_ADDER_2.B3.t18 VDD.t4063 VDD.t4062 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3528 VDD.t1812 SEL3.t71 a_n23950_3810.t8 VDD.t1811 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3529 a_n6920_3190.t3 a_n6950_3164.t6 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t6 VSS.t1807 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3530 a_n15737_n5180.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t18 VSS.t350 VSS.t349 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3531 a_n7496_3810.t3 a_n7676_3190.t7 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t0 VDD.t3960 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3532 a_7548_n30006.t1 SEL1.t131 a_7452_n30006.t1 VSS.t1971 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3533 a_n13399_n8419.t4 MULT_0.4bit_ADDER_1.B1.t21 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t7 VSS.t1503 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3534 Y1.t3 mux8_2.inv_0.A.t10 VDD.t1524 VDD.t1523 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3535 a_n18686_n2915.t1 B0.t41 VSS.t510 VSS.t509 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3536 VDD.t1452 mux8_6.NAND4F_3.Y.t10 mux8_6.NAND4F_8.Y.t5 VDD.t1451 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3537 a_7452_762.t0 SEL2.t118 VSS.t1745 VSS.t1441 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3538 a_n22425_n11256.t0 A2.t36 VSS.t262 VSS.t261 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3539 mux8_1.inv_0.A.t0 mux8_1.NAND4F_8.Y.t14 VSS.t1947 VSS.t1946 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X3540 mux8_0.NAND4F_5.Y.t6 left_shifter_0.C.t6 a_7644_762.t0 VSS.t841 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3541 VDD.t544 A2.t37 MULT_0.inv_12.A.t1 VDD.t543 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3542 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t6 MULT_0.4bit_ADDER_1.B1.t22 VDD.t3280 VDD.t3279 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3543 AND8_0.NOT8_0.A0.t6 A0.t40 VDD.t2239 VDD.t2238 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3544 a_n13975_n4534.t6 a_n14155_n5154.t7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t6 VDD.t4164 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3545 VDD.t3229 mux8_2.NAND4F_4.B.t12 mux8_2.NAND4F_3.Y.t7 VDD.t3228 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3546 a_n17677_n25225.t0 A7.t40 OR8_0.NOT8_0.A7.t0 VDD.t3449 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3547 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t10 a_n11723_n6187.t1 VSS.t351 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3548 mux8_8.NAND4F_8.Y.t3 mux8_8.NAND4F_0.Y.t10 VDD.t167 VDD.t166 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3549 mux8_4.inv_0.A.t1 mux8_4.NAND4F_9.Y.t14 a_11865_n16359.t5 VDD.t964 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3550 VSS.t927 SEL3.t72 a_n4385_3190.t1 VSS.t926 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X3551 VSS.t270 a_n14781_1380.t7 a_n14751_1406.t2 VSS.t269 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3552 a_n12416_n5154.t3 a_n12446_n5180.t7 VSS.t1089 VSS.t1088 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3553 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t4 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t10 VDD.t1085 VDD.t1084 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3554 VSS.t1254 OR8_0.NOT8_0.A1.t10 OR8_0.S1.t3 VSS.t1253 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3555 VDD.t3847 SEL2.t119 mux8_4.NAND4F_6.Y.t1 VDD.t3846 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3556 a_11865_1753.t9 mux8_0.NAND4F_9.Y.t14 mux8_0.inv_0.A.t6 VDD.t3126 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3557 VDD.t114 MULT_0.4bit_ADDER_1.A1.t13 a_n13975_n7799.t1 VDD.t113 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X3558 mux8_4.NAND4F_7.Y.t0 SEL2.t120 VDD.t3849 VDD.t3848 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3559 VDD.t1053 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t22 a_n19178_n8419.t1 VDD.t1052 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3560 MULT_0.4bit_ADDER_2.B1.t2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t20 a_n15131_n8419.t2 VSS.t323 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3561 VDD.t568 mux8_6.NAND4F_0.C.t14 mux8_6.NAND4F_7.Y.t2 VDD.t567 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3562 a_n12314_n26419.t2 a_n12345_n25873.t7 XOR8_0.S4.t2 VDD.t629 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3563 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t4 A2.t38 VDD.t546 VDD.t545 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3564 mux8_2.NAND4F_1.Y.t1 SEL2.t121 VDD.t3851 VDD.t3850 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3565 XOR8_0.S3.t1 a_n12345_n23393.t7 a_n12314_n23651.t0 VDD.t3490 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3566 AND8_0.S7.t1 AND8_0.NOT8_0.A7.t10 VDD.t3489 VDD.t3488 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3567 VSS.t1370 a_1857_4888.t6 a_1887_4914.t1 VSS.t1369 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3568 VDD.t2757 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t15 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t3 VDD.t2756 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3569 VDD.t653 mux8_0.NAND4F_0.C.t13 mux8_0.NAND4F_1.Y.t5 VDD.t652 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3570 a_n12314_n31661.t6 a_n12345_n31115.t6 XOR8_0.S6.t11 VDD.t2641 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3571 VDD.t1995 mux8_5.NAND4F_4.B.t12 mux8_5.NAND4F_4.Y.t4 VDD.t1994 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3572 Y0.t0 mux8_1.inv_0.A.t10 VSS.t545 VSS.t544 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3573 VDD.t342 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t20 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t1 VDD.t341 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3574 VDD.t1720 mux8_1.NAND4F_2.D.t15 mux8_1.NAND4F_2.Y.t4 VDD.t1719 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3575 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t6 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t20 VDD.t3907 VDD.t3906 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3576 MULT_0.NAND2_1.Y.t4 B0.t42 VDD.t1027 VDD.t1026 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3577 mux8_4.NAND4F_1.Y.t7 mux8_4.NAND4F_4.B.t15 VDD.t3374 VDD.t3373 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3578 mux8_2.NAND4F_0.Y.t7 mux8_2.NAND4F_0.C.t13 VDD.t3213 VDD.t3212 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3579 AND8_0.S6.t2 AND8_0.NOT8_0.A6.t9 VDD.t1574 VDD.t1573 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3580 mux8_2.NAND4F_5.Y.t7 SEL2.t122 VDD.t3853 VDD.t3852 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3581 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t1 a_n14005_n11709.t6 a_n13975_n11063.t10 VDD.t1651 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3582 VDD.t2510 MULT_0.4bit_ADDER_1.B0.t22 a_n10864_n8419.t1 VDD.t2509 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3583 OR8_0.NOT8_0.A7.t6 B7.t31 VSS.t585 VSS.t177 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X3584 VDD.t788 OR8_0.NOT8_0.A7.t9 OR8_0.S7.t2 VDD.t787 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3585 VDD.t149 OR8_0.S5.t5 mux8_7.NAND4F_2.Y.t0 VDD.t148 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3586 VDD.t2950 SEL0.t128 mux8_6.NAND4F_4.B.t1 VDD.t2949 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3587 MULT_0.inv_15.Y.t0 MULT_0.NAND2_15.Y.t10 VSS.t1324 VSS.t1323 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3588 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t8 a_n21513_1406.t7 a_n21333_1406.t3 VSS.t599 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3589 a_n15707_n7799.t7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t16 VDD.t3676 VDD.t3675 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3590 a_n17266_n11063.t6 a_n17296_n11709.t7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t11 VDD.t2858 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3591 VDD.t4502 SEL1.t132 mux8_3.NAND4F_2.Y.t5 VDD.t4501 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3592 a_n19981_n11683.t3 MULT_0.inv_15.Y.t12 VSS.t1533 VSS.t1532 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3593 a_7452_n30934.t0 SEL2.t123 VSS.t1746 VSS.t738 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3594 NOT8_0.S7.t0 B7.t32 VDD.t1166 VDD.t1165 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3595 mux8_4.NAND4F_8.Y.t6 mux8_4.NAND4F_4.Y.t11 a_11386_n16422.t1 VSS.t1377 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3596 VSS.t161 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t21 a_n8350_1406.t0 VSS.t160 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X3597 mux8_7.NAND4F_7.Y.t7 SEL0.t129 VDD.t2948 VDD.t2947 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3598 mux8_5.NAND4F_0.C.t0 SEL1.t133 VSS.t1985 VSS.t1984 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3599 ZFLAG_0.NAND2_0.Y.t5 ZFLAG_0.nor4_1.Y.t9 VDD.t2390 VDD.t2389 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3600 VDD.t2131 B3.t47 a_n10786_3810.t8 VDD.t2130 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X3601 a_n1012_1406.t5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t22 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t11 VSS.t1081 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3602 mux8_0.NAND4F_7.Y.t5 VSS.t2063 VDD.t1923 VDD.t1922 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3603 a_n15131_n8419.t1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t21 MULT_0.4bit_ADDER_2.B1.t1 VSS.t324 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3604 a_n14077_3810.t9 a_n13531_3164.t7 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t3 VDD.t2729 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3605 VDD.t3855 SEL2.t124 mux8_5.NAND4F_6.Y.t7 VDD.t3854 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3606 a_11386_n20950.t1 mux8_5.NAND4F_2.Y.t11 a_11290_n20950.t1 VSS.t701 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3607 VDD.t2019 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t22 a_n12416_n11063.t6 VDD.t2018 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3608 mux8_7.A1.t0 a_n15887_n11683.t7 a_n15707_n11683.t0 VSS.t797 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3609 mux8_5.NAND4F_7.Y.t0 SEL2.t125 VDD.t3857 VDD.t3856 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3610 OR8_0.S6.t1 OR8_0.NOT8_0.A6.t9 VDD.t322 VDD.t321 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3611 left_shifter_0.S6.t1 left_shifter_0.buffer_3.inv_1.A.t7 VDD.t817 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3612 VDD.t3565 B6.t32 a_n20659_3810.t3 VDD.t3564 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3613 VSS.t625 a_n1618_1380.t6 a_n1588_1406.t5 VSS.t624 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3614 a_7644_762.t1 mux8_0.NAND4F_4.B.t13 a_7548_762.t0 VSS.t426 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3615 MULT_0.4bit_ADDER_0.B1.t0 MULT_0.NAND2_1.Y.t10 VSS.t108 VSS.t107 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3616 VDD.t4041 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t9 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t2 VDD.t4040 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3617 a_n8170_1406.t0 a_n8350_1406.t7 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t11 VSS.t747 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3618 a_5167_4886.t1 mux8_6.A0.t21 VSS.t1525 VSS.t1524 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3619 right_shifter_0.buffer_6.inv_1.A.t2 B0.t43 VDD.t1028 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3620 a_n12345_n25873.t1 A4.t25 VDD.t2200 VDD.t2199 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3621 left_shifter_0.C.t2 left_shifter_0.buffer_1.inv_1.A.t6 VDD.t138 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3622 mux8_0.NAND4F_3.Y.t6 8bit_ADDER_0.C.t9 a_9528_1690.t1 VSS.t776 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3623 mux8_5.NAND4F_1.Y.t4 mux8_5.NAND4F_4.B.t13 VDD.t1997 VDD.t1996 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3624 AND8_0.NOT8_0.A6.t1 A6.t28 VDD.t2833 VDD.t2832 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3625 a_n12347_n14753.t0 A0.t41 VSS.t1135 VSS.t1134 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3626 MULT_0.inv_12.A.t0 A2.t39 VDD.t548 VDD.t547 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3627 a_8400_n26406.t0 SEL2.t126 VSS.t1747 VSS.t1460 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3628 a_n13192_2026.t2 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t21 VDD.t352 VDD.t351 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3629 a_n11460_2026.t9 a_n11640_1406.t7 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t11 VDD.t1577 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3630 VDD.t2759 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t16 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t2 VDD.t2758 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3631 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t0 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t22 VDD.t344 VDD.t343 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3632 mux8_8.A0.t7 a_n19954_1406.t7 a_n19774_2026.t7 VDD.t1494 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3633 a_n1588_2026.t6 a_n1618_1380.t7 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t8 VDD.t1254 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3634 a_n9125_n11063.t2 a_n9155_n11709.t7 mux8_4.A1.t2 VDD.t907 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3635 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t21 VDD.t3909 VDD.t3908 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3636 a_n17677_n16825.t1 B1.t46 VDD.t2377 VDD.t2376 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3637 VDD.t550 A2.t40 a_n8170_2026.t3 VDD.t549 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3638 VDD.t1621 right_shifter_0.S3.t5 mux8_4.NAND4F_6.Y.t3 VDD.t1620 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3639 a_n15790_373.t1 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t7 VSS.t953 VSS.t952 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3640 mux8_2.NAND4F_4.Y.t1 AND8_0.S1.t5 VDD.t792 VDD.t791 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3641 NOT8_0.S7.t1 B7.t33 VDD.t1168 VDD.t1167 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3642 mux8_7.NAND4F_1.Y.t6 XOR8_0.S5.t14 a_9528_n26406.t0 VSS.t296 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3643 mux8_2.inv_0.A.t0 mux8_2.NAND4F_8.Y.t14 VSS.t14 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X3644 mux8_3.NAND4F_0.Y.t7 SEL0.t130 VDD.t2946 VDD.t2945 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3645 8bit_ADDER_0.S0.t8 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t20 a_547_1406.t3 VSS.t1145 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3646 a_n8432_n6187.t1 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t9 VSS.t1221 VSS.t101 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3647 VSS.t866 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t18 a_n9325_1406.t0 VSS.t865 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3648 a_n12314_n18115.t5 a_n12345_n17569.t7 XOR8_0.S1.t3 VDD.t1305 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3649 VSS.t1188 B1.t47 right_shifter_0.buffer_7.inv_1.A.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3650 a_n22425_n12548.t1 B3.t48 VSS.t1098 VSS.t1097 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3651 VDD.t1744 mux8_0.NAND4F_2.Y.t11 mux8_0.NAND4F_8.Y.t5 VDD.t1743 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3652 a_9432_762.t1 mux8_0.NAND4F_0.C.t14 a_9336_762.t1 VSS.t317 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3653 a_11865_n11831.t0 mux8_3.NAND4F_8.Y.t14 VDD.t3929 VDD.t3928 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3654 VDD.t79 mux8_1.NAND4F_0.C.t15 mux8_1.NAND4F_7.Y.t3 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3655 mux8_4.NAND4F_2.Y.t0 mux8_4.NAND4F_2.D.t14 VDD.t132 VDD.t131 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3656 VSS.t194 A5.t26 a_n17466_1406.t3 VSS.t193 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3657 mux8_0.NAND4F_4.B.t1 SEL0.t131 VDD.t2944 VDD.t2943 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3658 VDD.t1921 VSS.t2064 mux8_0.NAND4F_2.Y.t1 VDD.t1920 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3659 mux8_8.A0.t5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t22 a_n19198_1406.t3 VSS.t1208 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3660 a_7548_762.t1 SEL1.t134 a_7452_762.t1 VSS.t1970 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3661 VDD.t3859 SEL2.t127 mux8_2.NAND4F_5.Y.t8 VDD.t3858 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3662 VSS.t1040 a_n10714_n11709.t7 a_n10684_n11683.t3 VSS.t1039 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3663 a_9336_n30006.t1 mux8_8.NAND4F_2.D.t15 VSS.t745 VSS.t744 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3664 VDD.t4292 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t16 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t1 VDD.t4291 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3665 VDD.t3861 SEL2.t128 mux8_8.NAND4F_6.Y.t1 VDD.t3860 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3666 VDD.t4504 SEL1.t135 mux8_6.NAND4F_2.Y.t5 VDD.t4503 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3667 VDD.t1169 B7.t34 left_shifter_0.buffer_1.inv_1.A.t1 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3668 VDD.t1079 MULT_0.4bit_ADDER_2.B0.t22 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t0 VDD.t1078 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3669 a_n3659_3164.t0 B1.t48 VSS.t1190 VSS.t1189 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3670 VDD.t3245 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t22 a_n21513_1406.t1 VDD.t3244 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3671 mux8_8.NAND4F_7.Y.t0 SEL2.t129 VDD.t3863 VDD.t3862 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3672 mux8_0.NAND4F_4.Y.t1 mux8_0.NAND4F_4.B.t14 VDD.t859 VDD.t858 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3673 a_n24048_1406.t0 A7.t41 VSS.t1588 VSS.t1587 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3674 VDD.t1343 MULT_0.4bit_ADDER_0.B1.t14 a_n14155_n5154.t1 VDD.t1342 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3675 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t3 a_n14155_n8419.t6 a_n13975_n7799.t3 VDD.t3691 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3676 a_n9125_n11063.t5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t20 VDD.t3390 VDD.t3389 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3677 right_shifter_0.buffer_6.inv_1.A.t1 B0.t44 VDD.t1029 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3678 a_n17677_n15425.t5 B0.t45 VDD.t1031 VDD.t1030 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X3679 mux8_3.NAND4F_5.Y.t8 left_shifter_0.S2.t6 a_7644_n12822.t0 VSS.t208 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3680 VDD.t404 A5.t27 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t6 VDD.t403 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3681 a_2463_4914.t0 A7.t42 V_FLAG_0.XOR2_2.B.t3 VSS.t1589 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3682 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t2 a_n14155_n8419.t7 a_n13975_n8419.t0 VSS.t1691 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3683 a_n12314_n21072.t10 a_n12345_n20814.t7 XOR8_0.S2.t7 VDD.t1237 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3684 a_17528_n18777.t1 ZFLAG_0.nor4_0.Y.t9 VSS.t91 VSS.t90 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3685 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t2 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t19 VDD.t2879 VDD.t2878 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3686 MULT_0.4bit_ADDER_1.B3.t1 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t8 VDD.t721 VDD.t720 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3687 mux8_5.NAND4F_0.Y.t6 mux8_5.NAND4F_2.D.t15 VDD.t1383 VDD.t1382 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3688 a_n29_2026.t9 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t21 VDD.t2261 VDD.t2260 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3689 VDD.t175 right_shifter_0.S4.t5 mux8_5.NAND4F_6.Y.t1 VDD.t174 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3690 mux8_8.NAND4F_1.Y.t5 mux8_8.NAND4F_4.B.t15 VDD.t3166 VDD.t3165 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3691 ZFLAG_0.nor4_1.Y.t1 Y7.t10 a_16431_n19505.t0 VDD.t562 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X3692 a_15855_n18523.t1 Y3.t6 VDD.t2420 VDD.t2003 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X3693 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t1 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t17 VDD.t2761 VDD.t2760 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3694 mux8_3.NAND4F_8.Y.t1 mux8_3.NAND4F_3.Y.t11 VDD.t1194 VDD.t1193 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3695 a_8400_n35462.t0 SEL2.t130 VSS.t1748 VSS.t202 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3696 VDD.t480 B2.t45 a_n12345_n20814.t1 VDD.t479 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3697 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t1 MULT_0.4bit_ADDER_0.B0.t14 VDD.t294 VDD.t293 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3698 VSS.t12 MULT_0.4bit_ADDER_1.A2.t14 a_n16690_n8419.t3 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3699 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t3 MULT_0.4bit_ADDER_1.A1.t14 a_n13714_n9452.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3700 VDD.t3911 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t22 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t4 VDD.t3910 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3701 VDD.t3865 SEL2.t131 mux8_1.NAND4F_6.Y.t0 VDD.t3864 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3702 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t1 B7.t35 a_n23950_3190.t3 VSS.t586 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3703 mux8_0.NAND4F_0.Y.t3 VSS.t2065 VDD.t1919 VDD.t1918 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3704 a_n22176_n2915.t1 B0.t46 VSS.t512 VSS.t511 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3705 a_n15707_n7799.t3 a_n15887_n8419.t7 MULT_0.4bit_ADDER_2.B1.t7 VDD.t1440 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3706 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t23 VDD.t2021 VDD.t2020 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3707 a_n15707_n8419.t3 a_n15737_n8445.t7 VSS.t30 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3708 VDD.t31 MULT_0.4bit_ADDER_1.A2.t15 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t3 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3709 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t2 a_n17296_n5180.t7 a_n17266_n4534.t11 VDD.t2395 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3710 VDD.t3231 mux8_2.NAND4F_4.B.t13 mux8_2.NAND4F_1.Y.t8 VDD.t3230 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3711 V_FLAG_0.XOR2_2.B.t0 a_1707_4914.t7 a_1887_5534.t0 VDD.t278 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3712 VDD.t1033 B0.t47 a_n914_3810.t6 VDD.t1032 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3713 mux8_7.A0.t8 a_n16513_1380.t7 a_n16483_2026.t8 VDD.t1485 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3714 VDD.t2202 A4.t26 a_n14751_2026.t11 VDD.t2201 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X3715 a_n23065_1406.t3 a_n23245_1406.t7 mux8_6.A0.t6 VSS.t1258 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3716 a_n17677_n25225.t6 B7.t36 VDD.t1171 VDD.t1170 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3717 mux8_5.NAND4F_2.D.t0 SEL2.t132 VSS.t1750 VSS.t1749 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3718 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t11 B1.t49 a_n4205_3190.t3 VSS.t1191 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3719 VDD.t4065 mux8_1.NAND4F_2.Y.t10 mux8_1.NAND4F_8.Y.t8 VDD.t4064 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3720 MULT_0.4bit_ADDER_1.B1.t6 a_n15887_n5154.t7 a_n15707_n5154.t0 VSS.t1152 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3721 a_n11723_n6187.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t10 VSS.t1267 VSS.t351 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3722 a_9336_762.t0 SEL2.t133 VSS.t1751 VSS.t1439 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3723 mux8_1.NAND4F_2.Y.t1 OR8_0.S0.t5 VDD.t883 VDD.t882 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3724 VDD.t723 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t9 MULT_0.4bit_ADDER_1.B3.t2 VDD.t722 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3725 a_9432_n8194.t0 mux8_2.NAND4F_0.C.t14 a_9336_n8194.t1 VSS.t1486 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3726 VSS.t986 VSS.t984 a_n8549_n8419.t3 VSS.t985 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3727 mux8_6.NAND4F_1.Y.t8 XOR8_0.S7.t14 a_9528_n35462.t1 VSS.t1499 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3728 mux8_0.NAND4F_2.Y.t0 VSS.t982 a_8592_1690.t0 VSS.t983 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3729 VSS.t587 B7.t37 right_shifter_0.buffer_1.inv_1.A.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3730 mux8_2.NAND4F_7.Y.t4 NOT8_0.S1.t6 VDD.t2212 VDD.t2211 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3731 mux8_4.NAND4F_2.Y.t2 OR8_0.S3.t5 a_8592_n16422.t0 VSS.t196 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3732 VSS.t1591 A7.t43 a_5017_4912.t0 VSS.t1590 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X3733 8bit_ADDER_0.S1.t3 a_n3350_1380.t7 a_n3320_2026.t3 VDD.t178 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3734 a_n8549_n5154.t0 VSS.t979 VSS.t981 VSS.t980 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3735 a_n18422_n8419.t3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t18 VSS.t1872 VSS.t1871 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3736 a_n9125_n11063.t4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t21 VDD.t3392 VDD.t3391 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3737 VDD.t169 mux8_8.NAND4F_0.Y.t11 mux8_8.NAND4F_8.Y.t2 VDD.t168 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3738 mux8_6.NAND4F_0.Y.t7 SEL0.t132 VDD.t2942 VDD.t2941 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3739 XOR8_0.S4.t6 a_n12345_n26161.t7 a_n12314_n26419.t6 VDD.t4166 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3740 a_n12314_n23651.t6 B3.t49 VDD.t2133 VDD.t2132 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3741 a_3493_4914.t0 a_3463_4888.t7 VSS.t233 VSS.t232 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3742 mux8_7.NAND4F_2.Y.t8 mux8_7.NAND4F_2.D.t14 VDD.t3140 VDD.t3139 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3743 a_n18998_n4534.t11 a_n19028_n5180.t6 MULT_0.4bit_ADDER_1.B2.t11 VDD.t2847 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3744 VDD.t406 A5.t28 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t5 VDD.t405 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3745 VSS.t1789 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t18 a_n12616_1406.t3 VSS.t1788 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3746 mux8_1.NAND4F_7.Y.t7 SEL0.t133 VDD.t2940 VDD.t2939 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3747 VDD.t2938 SEL0.t134 mux8_5.NAND4F_4.B.t1 VDD.t2937 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3748 VSS.t929 SEL3.t73 a_n7676_3190.t0 VSS.t928 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X3749 VSS.t1063 a_n18072_1380.t6 a_n18042_1406.t0 VSS.t1062 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3750 a_n17677_n23825.t5 B6.t33 VDD.t3567 VDD.t3566 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.3968 ps=3.18 w=1.28 l=0.15
X3751 a_15855_n18523.t0 Y3.t7 VDD.t2422 VDD.t2421 sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=1.3268 ps=9.18 w=4.28 l=0.15
X3752 VDD.t173 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t17 a_n23065_2026.t3 VDD.t172 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3753 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t1 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t20 VDD.t2881 VDD.t2880 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3754 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t23 VDD.t1593 VDD.t1592 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3755 mux8_3.NAND4F_8.Y.t2 mux8_3.NAND4F_0.Y.t10 VDD.t1456 VDD.t1455 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3756 VSS.t1305 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t18 a_n2744_1406.t3 VSS.t1304 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3757 mux8_4.NAND4F_2.Y.t3 OR8_0.S3.t6 VDD.t412 VDD.t411 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3758 mux8_3.NAND4F_6.Y.t7 SEL0.t135 VDD.t2936 VDD.t2935 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3759 a_n8170_2026.t0 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t23 VDD.t346 VDD.t345 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3760 MULT_0.NAND2_2.Y.t0 B0.t48 VDD.t1035 VDD.t1034 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3761 mux8_7.NAND4F_0.Y.t3 mux8_7.A1.t13 a_10459_n25478.t0 VSS.t19 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3762 VDD.t2135 B3.t50 MULT_0.NAND2_8.Y.t5 VDD.t2134 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3763 MULT_0.NAND2_3.Y.t1 A0.t42 VDD.t2241 VDD.t2240 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3764 VDD.t1065 right_shifter_0.S6.t5 mux8_8.NAND4F_6.Y.t3 VDD.t1064 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3765 VDD.t2934 SEL0.t136 mux8_1.NAND4F_4.B.t1 VDD.t2933 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3766 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t6 a_n20737_n11683.t5 a_n20557_n11063.t3 VDD.t3455 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3767 a_7452_1690.t0 mux8_0.NAND4F_2.D.t13 VSS.t1442 VSS.t1441 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3768 MULT_0.inv_6.A.t4 A0.t43 VDD.t2243 VDD.t2242 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3769 a_8400_n8194.t0 SEL2.t134 VSS.t1752 VSS.t1472 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3770 VSS.t341 mux8_6.NAND4F_9.Y.t14 mux8_6.inv_0.A.t6 VSS.t340 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X3771 a_5773_4912.t0 A7.t44 V_FLAG_0.XOR2_0.Y.t11 VSS.t1592 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3772 a_n13501_3190.t0 a_n14257_3190.t7 VSS.t277 VSS.t276 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3773 mux8_6.NAND4F_8.Y.t6 mux8_6.NAND4F_3.Y.t11 VDD.t1454 VDD.t1453 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3774 OR8_0.NOT8_0.A2.t1 A2.t41 a_n17677_n18225.t1 VDD.t551 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3775 XOR8_0.S0.t6 a_n12347_n15041.t7 a_n12316_n15299.t6 VDD.t3687 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3776 VDD.t1210 XOR8_0.S2.t14 mux8_3.NAND4F_1.Y.t3 VDD.t1209 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3777 VDD.t296 MULT_0.4bit_ADDER_0.B0.t15 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t2 VDD.t295 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3778 MULT_0.inv_12.A.t3 B2.t46 a_n22425_n7992.t1 VSS.t220 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3779 VDD.t1814 SEL3.t74 a_n14257_3190.t1 VDD.t1813 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3780 a_n18042_2026.t8 a_n18072_1380.t7 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t8 VDD.t2047 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3781 VSS.t1935 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t17 a_n11840_n8419.t3 VSS.t1934 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3782 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t3 a_n24804_1406.t7 a_n24624_1406.t5 VSS.t1599 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3783 AND8_0.NOT8_0.A6.t4 B6.t34 VDD.t3569 VDD.t3568 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3784 VSS.t326 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t22 a_n15887_n8419.t0 VSS.t325 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X3785 a_n15014_n12716.t1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t10 VSS.t726 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3786 a_n11840_n5154.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t18 VSS.t100 VSS.t99 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3787 a_n20557_n11683.t4 a_n20737_n11683.t6 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t7 VSS.t1595 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3788 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t4 MULT_0.inv_15.Y.t13 VDD.t3321 VDD.t3320 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3789 VDD.t3933 MULT_0.NAND2_9.Y.t10 MULT_0.inv_9.Y.t1 VDD.t3930 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3790 a_8592_n21878.t1 SEL0.t137 a_8496_n21878.t1 VSS.t2003 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3791 mux8_4.NAND4F_6.Y.t0 SEL2.t135 VDD.t3867 VDD.t3866 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3792 a_n17368_3810.t3 a_n16822_3164.t7 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t3 VDD.t2856 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3793 a_n11274_n31085.t2 B6.t35 XOR8_0.S6.t0 VSS.t1638 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3794 a_10363_n21877.t0 mux8_5.NAND4F_0.C.t14 a_10267_n21877.t1 VSS.t1665 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3795 VSS.t1552 a_n4909_1380.t6 a_n4879_1406.t5 VSS.t1551 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3796 a_9528_n8194.t1 mux8_2.NAND4F_4.B.t14 a_9432_n8194.t1 VSS.t1488 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3797 mux8_6.NAND4F_7.Y.t3 mux8_6.NAND4F_0.C.t15 VDD.t570 VDD.t569 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3798 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t4 A5.t29 VDD.t408 VDD.t407 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3799 mux8_5.NAND4F_4.Y.t3 mux8_5.NAND4F_4.B.t14 VDD.t1722 VDD.t1721 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3800 a_n4205_3810.t5 a_n3659_3164.t7 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t8 VDD.t1200 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3801 V_FLAG_0.XOR2_0.Y.t3 a_5017_4912.t7 a_5197_5532.t1 VDD.t1907 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3802 VDD.t2379 B1.t50 a_n17677_n16825.t0 VDD.t2378 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3803 VDD.t2883 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t21 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t0 VDD.t2882 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3804 VSS.t264 A2.t42 a_n11274_n20496.t0 VSS.t263 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3805 mux8_2.NAND4F_5.Y.t2 left_shifter_0.S1.t6 VDD.t1251 VDD.t1250 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3806 a_n914_3190.t0 SEL3.t75 VSS.t931 VSS.t930 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3807 VDD.t3327 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t9 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t5 VDD.t3326 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3808 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t3 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t7 a_n15790_373.t0 VSS.t952 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3809 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t6 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t23 VDD.t3896 VDD.t3895 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3810 VDD.t2137 B3.t51 MULT_0.NAND2_8.Y.t4 VDD.t2136 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3811 VDD.t17 mux8_4.A1.t14 mux8_4.NAND4F_0.Y.t5 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3812 a_n13975_n11063.t9 a_n14005_n11709.t7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t2 VDD.t1652 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3813 a_7644_n8194.t1 mux8_2.NAND4F_4.B.t15 a_7548_n8194.t1 VSS.t1489 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3814 a_n11490_1380.t0 A3.t44 VSS.t1851 VSS.t1850 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3815 VDD.t1471 mux8_8.NAND4F_4.Y.t10 mux8_8.NAND4F_8.Y.t8 VDD.t1470 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3816 mux8_7.NAND4F_2.Y.t4 OR8_0.S5.t6 VDD.t2647 VDD.t2646 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3817 OR8_0.S7.t1 OR8_0.NOT8_0.A7.t10 VDD.t790 VDD.t789 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3818 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t0 MULT_0.4bit_ADDER_1.B3.t18 VDD.t2725 VDD.t2724 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3819 a_n12314_n18115.t0 B1.t51 VDD.t1832 VDD.t1831 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3820 mux8_0.NAND4F_3.Y.t8 mux8_0.NAND4F_2.D.t14 VDD.t2900 VDD.t2899 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3821 a_n16483_2026.t9 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t23 VDD.t3913 VDD.t3912 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3822 a_n20557_n4534.t11 a_n20587_n5180.t7 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t6 VDD.t2036 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3823 a_11386_n16422.t0 mux8_4.NAND4F_2.Y.t9 a_11290_n16422.t1 VSS.t103 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3824 a_n23950_3810.t11 a_n23404_3164.t7 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t11 VDD.t2413 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3825 mux8_6.NAND4F_8.Y.t0 mux8_6.NAND4F_0.Y.t10 VDD.t863 VDD.t862 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3826 VDD.t776 SEL3.t76 a_n1094_3190.t1 VDD.t775 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3827 a_n4879_2026.t11 a_n4909_1380.t7 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t11 VDD.t3380 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3828 VDD.t2392 ZFLAG_0.nor4_1.Y.t10 ZFLAG_0.NAND2_0.Y.t6 VDD.t2391 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3829 mux8_5.NAND4F_6.Y.t8 SEL2.t136 VDD.t3869 VDD.t3868 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3830 a_n12314_n23651.t9 a_n12345_n23105.t7 XOR8_0.S3.t9 VDD.t2762 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3831 a_n3320_2026.t0 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t22 VDD.t761 VDD.t760 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3832 a_n17266_n7799.t0 a_n17296_n8445.t7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t0 VDD.t3290 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3833 mux8_2.NAND4F_0.Y.t2 MULT_0.S1.t14 a_10459_n7266.t1 VSS.t1051 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3834 VSS.t1137 A0.t44 a_n11276_n14723.t0 VSS.t1136 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3835 VSS.t495 V_FLAG_0.XOR2_2.B.t19 a_4069_4914.t3 VSS.t494 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3836 VDD.t462 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t21 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t0 VDD.t461 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3837 a_n16690_n8419.t0 MULT_0.4bit_ADDER_1.B2.t21 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t8 VSS.t1821 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3838 a_n18998_n11063.t9 a_n19028_n11709.t6 mux8_8.A1.t8 VDD.t2726 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3839 mux8_1.NAND4F_6.Y.t4 right_shifter_0.S0.t6 VDD.t1063 VDD.t1062 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3840 VDD.t633 mux8_1.NAND4F_6.Y.t11 mux8_1.NAND4F_9.Y.t0 VDD.t632 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3841 VSS.t1498 left_shifter_0.buffer_7.inv_1.A.t7 left_shifter_0.S2.t0 VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3842 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t9 VDD.t869 VDD.t868 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3843 a_n13975_n11063.t7 MULT_0.4bit_ADDER_2.B1.t22 VDD.t1903 VDD.t1902 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3844 a_n11274_n29052.t0 a_n12345_n28794.t7 XOR8_0.S5.t0 VSS.t241 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3845 VSS.t1606 AND8_0.NOT8_0.A2.t10 AND8_0.S2.t0 VSS.t329 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3846 a_n20113_3164.t0 B6.t36 VSS.t1640 VSS.t1639 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3847 a_n14175_1406.t3 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t23 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t9 VSS.t702 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3848 VDD.t1206 left_shifter_0.buffer_1.inv_1.A.t7 left_shifter_0.C.t3 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3849 VDD.t2851 mux8_3.NAND4F_1.Y.t10 mux8_3.NAND4F_9.Y.t7 VDD.t2850 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3850 a_n13192_1406.t3 a_n13222_1380.t7 VSS.t384 VSS.t383 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3851 mux8_0.NAND4F_6.Y.t0 SEL2.t137 VDD.t3871 VDD.t3870 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3852 VDD.t819 mux8_4.NAND4F_2.Y.t10 mux8_4.NAND4F_8.Y.t3 VDD.t818 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3853 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t3 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t23 a_n20757_1406.t0 VSS.t1495 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3854 VDD.t4129 V_FLAG_0.XOR2_0.Y.t15 V_FLAG_0.NAND2_0.Y.t4 VDD.t4128 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3855 VDD.t2315 MULT_0.4bit_ADDER_0.A1.t14 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t1 VDD.t2314 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3856 a_n6950_3164.t0 B2.t47 VSS.t222 VSS.t221 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3857 VDD.t3652 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t22 a_n24804_1406.t1 VDD.t3651 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3858 a_n9125_n8419.t3 a_n9305_n8419.t7 MULT_0.S2.t8 VSS.t519 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3859 MULT_0.4bit_ADDER_2.B2.t11 a_n19028_n8445.t7 a_n18998_n7799.t6 VDD.t1346 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3860 VSS.t224 B2.t48 NOT8_0.S2.t0 VSS.t223 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3861 MULT_0.NAND2_9.Y.t4 B3.t52 VDD.t2139 VDD.t2138 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3862 VDD.t3491 right_shifter_0.buffer_2.inv_1.A.t5 right_shifter_0.S5.t3 VDD.t361 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3863 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t0 a_n10864_n5154.t7 a_n10684_n5154.t3 VSS.t498 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3864 MULT_0.S1.t8 a_n9305_n5154.t7 a_n9125_n5154.t3 VSS.t763 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3865 ZFLAG_0.nor4_0.Y.t5 Y1.t7 VSS.t1566 VSS.t1565 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3866 MULT_0.4bit_ADDER_2.B2.t5 a_n19178_n8419.t7 a_n18998_n8419.t0 VSS.t126 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3867 VDD.t3451 A7.t45 a_1707_4914.t1 VDD.t3450 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3868 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t6 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t10 VDD.t3329 VDD.t3328 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3869 a_n20557_n4534.t0 MULT_0.4bit_ADDER_0.A3.t14 VDD.t1612 VDD.t1611 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3870 mux8_2.inv_0.A.t1 mux8_2.NAND4F_9.Y.t13 a_11865_n7203.t9 VDD.t2117 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3871 left_shifter_0.buffer_6.inv_1.A.t1 B0.t49 VDD.t1036 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3872 VDD.t1173 B7.t38 a_n17677_n25225.t5 VDD.t1172 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3873 mux8_5.NAND4F_4.Y.t0 AND8_0.S4.t6 a_7644_n20950.t0 VSS.t328 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3874 mux8_4.NAND4F_6.Y.t4 right_shifter_0.S3.t6 VDD.t1623 VDD.t1622 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3875 a_n9155_n8445.t1 VSS.t2066 VDD.t1917 VDD.t1916 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3876 VDD.t1108 mux8_7.A1.t14 mux8_7.NAND4F_0.Y.t4 VDD.t1107 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3877 a_9528_n26406.t1 mux8_7.NAND4F_4.B.t14 a_9432_n26406.t1 VSS.t92 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3878 VDD.t3873 SEL2.t138 mux8_0.NAND4F_5.Y.t0 VDD.t3872 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3879 VDD.t501 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t23 a_n18998_n4534.t0 VDD.t500 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3880 VSS.t1374 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t17 a_n11840_n11683.t4 VSS.t1373 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3881 VDD.t947 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t18 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t4 VDD.t946 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3882 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t5 MULT_0.inv_15.Y.t14 a_n20296_n12716.t1 VSS.t1534 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3883 VDD.t4236 A1.t41 MULT_0.NAND2_5.Y.t5 VDD.t4235 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3884 a_n20659_3190.t0 SEL3.t77 VSS.t386 VSS.t385 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3885 a_n15131_n11683.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t23 mux8_7.A1.t6 VSS.t634 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3886 a_11290_n21878.t0 mux8_5.NAND4F_1.Y.t11 a_11194_n21878.t0 VSS.t1329 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3887 VDD.t3185 mux8_2.NAND4F_2.D.t15 mux8_2.NAND4F_3.Y.t3 VDD.t3184 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3888 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t2 a_n1094_3190.t7 a_n914_3810.t5 VDD.t920 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3889 a_n12416_n5154.t1 a_n12596_n5154.t6 MULT_0.4bit_ADDER_1.B0.t1 VSS.t496 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3890 a_n11460_2026.t0 a_n11490_1380.t7 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t5 VDD.t955 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3891 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t3 VSS.t978 a_n9314_n9452.t1 VSS.t290 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3892 mux8_8.NAND4F_6.Y.t0 SEL2.t139 VDD.t3875 VDD.t3874 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3893 a_n17266_n4534.t3 MULT_0.4bit_ADDER_0.B2.t15 VDD.t2922 VDD.t2921 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3894 a_n13975_n11063.t6 MULT_0.4bit_ADDER_2.B1.t23 VDD.t1905 VDD.t1904 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3895 VDD.t3394 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t22 a_n9125_n11063.t3 VDD.t3393 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3896 VSS.t1083 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t23 a_n1768_1406.t1 VSS.t1082 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.1885 ps=1.88 w=0.65 l=0.15
X3897 mux8_0.NAND4F_6.Y.t7 SEL0.t138 VDD.t2932 VDD.t2931 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3898 a_7644_n12822.t1 mux8_3.NAND4F_4.B.t15 a_7548_n12822.t0 VSS.t1269 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3899 VDD.t3323 MULT_0.inv_15.Y.t15 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t6 VDD.t3322 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3900 a_5197_5532.t9 mux8_6.A0.t22 VDD.t3309 VDD.t3308 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3901 8bit_ADDER_0.S2.t3 a_n6641_1380.t7 a_n6611_2026.t8 VDD.t886 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3902 VDD.t2701 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t8 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t4 VDD.t2700 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3903 VDD.t2426 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t10 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t6 VDD.t2425 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3904 MULT_0.NAND2_5.Y.t4 A1.t42 VDD.t4238 VDD.t4237 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3905 a_n11276_n33705.t4 B7.t39 XOR8_0.S7.t10 VSS.t588 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3906 mux8_0.NAND4F_2.Y.t6 mux8_0.NAND4F_2.D.t15 VDD.t2902 VDD.t2901 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X3907 VDD.t4264 mux8_7.NAND4F_2.Y.t11 mux8_7.NAND4F_8.Y.t7 VDD.t4263 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3908 mux8_5.NAND4F_6.Y.t2 right_shifter_0.S4.t6 VDD.t177 VDD.t176 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3909 VSS.t1299 mux8_3.NAND4F_9.Y.t14 mux8_3.inv_0.A.t6 VSS.t1298 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X3910 a_n15707_n11683.t3 a_n15737_n11709.t7 VSS.t406 VSS.t405 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3911 a_n10714_n5180.t1 MULT_0.4bit_ADDER_0.A0.t14 VSS.t698 VSS.t697 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3912 VDD.t1458 mux8_3.NAND4F_0.Y.t11 mux8_3.NAND4F_8.Y.t3 VDD.t1457 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3913 AND8_0.NOT8_0.A2.t0 B2.t49 VDD.t482 VDD.t481 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3914 a_n20587_n8445.t0 MULT_0.4bit_ADDER_1.A3.t15 VSS.t1916 VSS.t1915 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3915 MULT_0.4bit_ADDER_1.B0.t2 a_n12596_n5154.t7 a_n12416_n5154.t0 VSS.t497 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3916 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t0 MULT_0.4bit_ADDER_0.A3.t15 a_n20296_n6187.t0 VSS.t790 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3917 VDD.t3638 mux8_5.NAND4F_0.C.t15 mux8_5.NAND4F_3.Y.t0 VDD.t3637 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3918 a_n17677_n18225.t0 A2.t43 OR8_0.NOT8_0.A2.t0 VDD.t552 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3919 VDD.t4505 SEL1.t136 mux8_4.NAND4F_0.C.t1 VDD.t4448 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3920 VSS.t1358 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t18 a_n15907_1406.t5 VSS.t1357 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3921 VDD.t861 mux8_0.NAND4F_4.B.t15 mux8_0.NAND4F_5.Y.t2 VDD.t860 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3922 a_7452_n11894.t0 mux8_3.NAND4F_2.D.t15 VSS.t1385 VSS.t1384 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3923 a_n12316_n15299.t9 B0.t50 VDD.t1038 VDD.t1037 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3924 VSS.t35 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t18 a_n6035_1406.t0 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3925 a_n17266_n7799.t6 MULT_0.4bit_ADDER_1.B2.t22 VDD.t4035 VDD.t4034 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3926 a_n17296_n11709.t0 MULT_0.inv_14.Y.t15 VSS.t1245 VSS.t1244 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3927 mux8_1.NAND4F_1.Y.t4 XOR8_0.S0.t14 a_9528_n3766.t0 VSS.t1543 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3928 VSS.t1914 A1.t43 a_n11274_n17539.t3 VSS.t1913 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3929 a_9528_n35462.t0 mux8_6.NAND4F_4.B.t14 a_9432_n35462.t1 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3930 a_n11274_n28476.t1 B5.t35 XOR8_0.S5.t2 VSS.t1802 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3931 VDD.t554 A2.t44 MULT_0.NAND2_1.Y.t1 VDD.t553 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X3932 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t8 a_n20737_n8419.t7 a_n20557_n8419.t3 VSS.t1418 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3933 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t5 a_n10240_3164.t7 a_n10210_3190.t0 VSS.t334 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3934 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t18 a_n12605_n9452.t1 VSS.t1761 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3935 mux8_4.A1.t6 a_n9305_n11683.t7 a_n9125_n11063.t6 VDD.t2734 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3936 VDD.t1039 B0.t51 NOT8_0.S0.t1 VDD.t887 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3937 a_n16792_3190.t4 a_n17548_3190.t7 VSS.t566 VSS.t565 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3938 mux8_1.NAND4F_5.Y.t2 left_shifter_0.S0.t6 a_7644_n3766.t0 VSS.t275 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3939 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t6 a_n14931_1406.t7 a_n14751_2026.t3 VDD.t3376 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3940 a_n21333_1406.t0 a_n21363_1380.t7 VSS.t611 VSS.t610 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3941 VDD.t2564 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t16 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t3 VDD.t2563 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3942 VDD.t208 mux8_7.NAND4F_4.B.t15 mux8_7.NAND4F_5.Y.t6 VDD.t207 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3943 VDD.t778 SEL3.t78 a_n17548_3190.t1 VDD.t777 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3944 VSS.t86 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t18 a_n22489_1406.t1 VSS.t85 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X3945 VDD.t3678 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t17 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t3 VDD.t3677 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3946 left_shifter_0.S0.t1 VDD.t3103 VDD.t3104 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3947 VDD.t165 MULT_0.NAND2_3.Y.t10 MULT_0.SO.t1 VDD.t162 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3948 OR8_0.NOT8_0.A4.t1 A4.t27 a_n17677_n21025.t8 VDD.t2203 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X3949 VDD.t780 SEL3.t79 a_n10786_3810.t0 VDD.t779 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3950 a_n368_3164.t0 B0.t52 VSS.t514 VSS.t513 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3951 VDD.t2703 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t9 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t5 VDD.t2702 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3952 VDD.t231 mux8_4.NAND4F_6.Y.t11 mux8_4.NAND4F_9.Y.t3 VDD.t230 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3953 VDD.t2930 SEL0.t139 mux8_4.NAND4F_2.Y.t7 VDD.t2929 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3954 VDD.t4507 SEL1.t137 mux8_3.NAND4F_6.Y.t5 VDD.t4506 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3955 a_10459_n25478.t1 SEL0.t140 a_10363_n25478.t1 VSS.t1994 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3956 a_n23404_3164.t1 B7.t40 VDD.t1175 VDD.t1174 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3957 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t0 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t8 VDD.t1848 VDD.t1847 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3958 a_n14005_n5180.t0 MULT_0.4bit_ADDER_0.A1.t15 VSS.t1170 VSS.t1169 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3959 MULT_0.4bit_ADDER_1.B3.t3 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t10 a_n18305_n6187.t0 VSS.t352 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3960 a_n10684_n7799.t9 MULT_0.4bit_ADDER_1.A0.t15 VDD.t3199 VDD.t3198 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3961 a_n18998_n5154.t5 a_n19028_n5180.t7 VSS.t1409 VSS.t1408 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3962 MULT_0.4bit_ADDER_1.A3.t1 MULT_0.inv_13.A.t10 VDD.t4324 VDD.t4273 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3963 mux8_8.NAND4F_6.Y.t4 right_shifter_0.S6.t6 VDD.t1067 VDD.t1066 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3964 mux8_2.NAND4F_4.Y.t3 SEL1.t138 VDD.t4509 VDD.t4508 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3965 a_n10423_n12716.t0 MULT_0.4bit_ADDER_2.B0.t23 VSS.t529 VSS.t428 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3966 a_n7496_3810.t6 a_n6950_3164.t7 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t3 VDD.t3987 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3967 a_n10108_n8419.t0 MULT_0.4bit_ADDER_1.B0.t23 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t2 VSS.t1266 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3968 VDD.t2885 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t22 a_n18222_1406.t1 VDD.t2884 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3969 VSS.t700 MULT_0.4bit_ADDER_0.A0.t15 a_n10108_n5154.t2 VSS.t699 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3970 mux8_6.inv_0.A.t0 mux8_6.NAND4F_8.Y.t14 VSS.t1444 VSS.t1443 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X3971 a_n13381_373.t0 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t22 VSS.t164 VSS.t163 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3972 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t4 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t17 VDD.t2566 VDD.t2565 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3973 VDD.t865 mux8_6.NAND4F_0.Y.t11 mux8_6.NAND4F_8.Y.t1 VDD.t864 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3974 a_n9901_2026.t6 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t22 VDD.t1551 VDD.t1550 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3975 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t23 VDD.t3396 VDD.t3395 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3976 a_n18998_n7799.t3 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t23 VDD.t1055 VDD.t1054 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3977 a_n1588_2026.t0 A0.t45 VDD.t2245 VDD.t2244 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3978 a_n14781_1380.t0 A4.t28 VSS.t1122 VSS.t1121 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X3979 a_n10684_n5154.t0 a_n10714_n5180.t7 VSS.t320 VSS.t319 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X3980 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t10 VDD.t4270 VDD.t4269 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X3981 a_n19774_2026.t10 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t23 VDD.t2410 VDD.t2409 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X3982 VDD.t2645 mux8_3.NAND4F_4.Y.t11 mux8_3.NAND4F_8.Y.t6 VDD.t2644 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X3983 VDD.t116 MULT_0.4bit_ADDER_1.A1.t15 a_n13975_n7799.t2 VDD.t115 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3984 a_7452_n34534.t0 mux8_6.NAND4F_2.D.t15 VSS.t207 VSS.t206 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3985 Y7.t0 mux8_6.inv_0.A.t10 VSS.t843 VSS.t842 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3986 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t8 a_n20737_n11683.t7 a_n20557_n11683.t3 VSS.t1609 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3987 a_n11274_n25843.t0 B4.t36 XOR8_0.S4.t3 VSS.t1657 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3988 VSS.t1308 AND8_0.NOT8_0.A5.t10 AND8_0.S5.t0 VSS.t329 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3989 VDD.t782 SEL3.t80 a_n4385_3190.t0 VDD.t781 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X3990 a_n8170_2026.t9 a_n8200_1380.t7 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t4 VDD.t336 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3991 a_8496_n21878.t0 SEL1.t139 a_8400_n21878.t1 VSS.t1967 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3992 VDD.t2061 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t23 a_n9125_n4534.t11 VDD.t2060 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3993 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t8 MULT_0.4bit_ADDER_1.B1.t23 a_n13399_n8419.t3 VSS.t1504 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3994 VDD.t1177 B7.t41 a_n12316_n34281.t6 VDD.t1176 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3995 VDD.t4248 mux8_5.NAND4F_6.Y.t11 mux8_5.NAND4F_9.Y.t5 VDD.t4247 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3996 a_10267_n21877.t0 SEL2.t140 VSS.t1753 VSS.t679 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3997 mux8_8.NAND4F_0.Y.t4 mux8_8.A1.t14 a_10459_n30006.t0 VSS.t1157 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3998 VDD.t4037 MULT_0.4bit_ADDER_1.B2.t23 a_n17266_n7799.t5 VDD.t4036 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X3999 a_547_1406.t0 SEL3.t81 VSS.t388 VSS.t387 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4000 VDD.t1071 mux8_0.NAND4F_1.Y.t11 mux8_0.NAND4F_9.Y.t3 VDD.t1070 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4001 VSS.t650 mux8_1.NAND4F_9.Y.t14 mux8_1.inv_0.A.t6 VSS.t649 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X4002 a_n13399_n5154.t3 MULT_0.4bit_ADDER_0.B1.t15 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t0 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4003 VDD.t556 A2.t45 MULT_0.NAND2_14.Y.t0 VDD.t555 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4004 VSS.t540 Y7.t11 ZFLAG_0.nor4_1.Y.t3 VSS.t539 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X4005 V.t1 V_FLAG_0.NAND2_0.Y.t10 VDD.t3501 VDD.t3500 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4006 a_n9325_1406.t3 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t23 mux8_4.A0.t1 VSS.t2030 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4007 VDD.t4511 SEL1.t140 mux8_5.NAND4F_4.Y.t7 VDD.t4510 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4008 VDD.t2263 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t22 a_n209_1406.t1 VDD.t2262 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X4009 mux8_2.NAND4F_3.Y.t5 8bit_ADDER_0.S1.t14 VDD.t1535 VDD.t1534 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4010 VDD.t2456 mux8_6.NAND4F_4.B.t15 mux8_6.NAND4F_5.Y.t7 VDD.t2455 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4011 VDD.t4240 A1.t44 AND8_0.NOT8_0.A1.t1 VDD.t4239 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X4012 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t6 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t10 VDD.t2705 VDD.t2704 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4013 mux8_4.NAND4F_4.Y.t0 mux8_4.NAND4F_2.D.t15 VDD.t134 VDD.t133 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X4014 a_n17466_1406.t0 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t23 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t11 VSS.t1433 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4015 right_shifter_0.S5.t2 right_shifter_0.buffer_2.inv_1.A.t6 VDD.t3492 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X4016 a_9432_n12822.t1 mux8_3.NAND4F_0.C.t15 a_9336_n12822.t1 VSS.t1322 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X4017 VDD.t1850 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t9 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t1 VDD.t1849 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4018 VDD.t1915 VSS.t2067 mux8_0.NAND4F_4.Y.t4 VDD.t1914 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X4019 VDD.t4147 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t23 a_n5059_1406.t1 VDD.t4146 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X4020 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t9 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t23 a_n24048_1406.t3 VSS.t1672 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4021 a_n20557_n4534.t6 VSS.t2068 VDD.t1913 VDD.t1912 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X4022 mux8_8.NAND4F_8.Y.t7 mux8_8.NAND4F_4.Y.t11 VDD.t1473 VDD.t1472 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4023 VSS.t803 a_n23095_1380.t7 a_n23065_1406.t0 VSS.t802 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4024 a_n6611_1406.t0 a_n6791_1406.t7 8bit_ADDER_0.S2.t0 VSS.t414 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4025 a_n15131_n8419.t0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t23 MULT_0.4bit_ADDER_2.B1.t0 VSS.t327 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4026 VDD.t2928 SEL0.t141 mux8_7.NAND4F_2.Y.t5 VDD.t2927 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4027 VDD.t3876 SEL2.t141 mux8_4.NAND4F_2.D.t1 VDD.t3791 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X4028 mux8_6.A1.t0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t10 a_n18305_n12716.t0 VSS.t483 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X4029 VDD.t3878 SEL2.t142 mux8_2.NAND4F_1.Y.t0 VDD.t3877 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4030 VDD.t3879 SEL2.t143 mux8_3.NAND4F_2.D.t1 VDD.t3789 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X4031 a_n11274_n23075.t3 B3.t53 XOR8_0.S3.t6 VSS.t1099 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4032 VDD.t1179 B7.t42 AND8_0.NOT8_0.A7.t4 VDD.t1178 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4033 VSS.t590 B7.t43 a_2463_4914.t3 VSS.t589 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10725 ps=0.98 w=0.65 l=0.15
X4034 left_shifter_0.buffer_2.inv_1.A.t1 B6.t37 VDD.t3570 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X4035 mux8_1.NAND4F_2.Y.t5 SEL1.t141 VDD.t4513 VDD.t4512 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4036 MULT_0.4bit_ADDER_1.B1.t1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t22 a_n15131_n5154.t1 VSS.t217 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4037 VDD.t1911 VSS.t2069 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t4 VDD.t1910 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X4038 ZFLAG_0.NAND2_0.Y.t0 ZFLAG_0.nor4_0.Y.t10 VDD.t196 VDD.t195 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4039 VDD.t4514 SEL1.t142 mux8_0.NAND4F_0.C.t1 VDD.t4405 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X4040 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t4 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t10 VDD.t3410 VDD.t3409 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X4041 8bit_ADDER_0.S0.t3 a_n209_1406.t7 a_n29_2026.t3 VDD.t3121 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X4042 VDD.t3215 mux8_2.NAND4F_0.C.t15 mux8_2.NAND4F_0.Y.t8 VDD.t3214 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4043 VSS.t772 AND8_0.NOT8_0.A6.t10 AND8_0.S6.t3 VSS.t771 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4044 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t6 B5.t36 a_n17368_3190.t3 VSS.t1803 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4045 mux8_8.A1.t7 a_n19028_n11709.t7 a_n18998_n11063.t10 VDD.t2727 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X4046 VDD.t1181 B7.t44 a_n12347_n34023.t1 VDD.t1180 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.7975 ps=6.08 w=2.75 l=0.15
X4047 a_n12314_n21072.t3 B2.t50 VDD.t484 VDD.t483 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X4048 VDD.t3680 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t18 a_n15707_n7799.t6 VDD.t3679 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X4049 VDD.t871 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t10 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t0 VDD.t870 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4050 a_n23950_3190.t0 SEL3.t82 VSS.t390 VSS.t389 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4051 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t9 B2.t51 a_n7496_3190.t3 VSS.t225 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4052 a_n11274_n31661.t5 a_n12345_n31115.t7 VSS.t1314 VSS.t1313 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10075 ps=0.96 w=0.65 l=0.15
X4053 XOR8_0.S7.t9 B7.t45 a_n11276_n33705.t3 VSS.t591 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4054 Y3.t3 mux8_4.inv_0.A.t10 VDD.t3461 VDD.t3460 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4055 VDD.t4184 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t23 a_n12416_n4534.t6 VDD.t4183 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X4056 mux8_4.NAND4F_8.Y.t2 mux8_4.NAND4F_2.Y.t11 VDD.t821 VDD.t820 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4057 mux8_3.NAND4F_9.Y.t8 mux8_3.NAND4F_1.Y.t11 VDD.t2853 VDD.t2852 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4058 VSS.t274 OR8_0.NOT8_0.A6.t10 OR8_0.S6.t0 VSS.t273 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4059 a_1887_5534.t11 a_1857_4888.t7 V_FLAG_0.XOR2_2.B.t10 VDD.t2771 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X4060 mux8_0.NAND4F_1.Y.t4 mux8_0.NAND4F_0.C.t15 VDD.t655 VDD.t654 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4061 mux8_1.NAND4F_8.Y.t7 mux8_1.NAND4F_0.Y.t11 VDD.t3333 VDD.t3332 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X4062 VDD.t356 mux8_8.NAND4F_6.Y.t11 mux8_8.NAND4F_9.Y.t3 VDD.t355 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4063 VDD.t486 B2.t52 AND8_0.NOT8_0.A2.t1 VDD.t485 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4064 mux8_1.NAND4F_3.Y.t7 mux8_1.NAND4F_4.B.t15 VDD.t1274 VDD.t1273 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4065 a_n15131_n5154.t0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t23 MULT_0.4bit_ADDER_1.B1.t0 VSS.t218 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4066 a_n20296_n6187.t1 VSS.t976 VSS.t977 VSS.t790 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X4067 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t10 VDD.t4039 VDD.t4038 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4068 VDD.t913 mux8_6.NAND4F_4.Y.t11 mux8_6.NAND4F_8.Y.t3 VDD.t912 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X4069 right_shifter_0.S5.t1 right_shifter_0.buffer_2.inv_1.A.t7 VDD.t3493 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X4070 mux8_4.NAND4F_4.Y.t8 AND8_0.S3.t6 a_7644_n16422.t1 VSS.t957 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X4071 VSS.t516 B0.t53 a_n24013_n15316.t1 VSS.t515 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X4072 mux8_1.NAND4F_2.Y.t0 OR8_0.S0.t6 a_8592_n2838.t0 VSS.t433 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X4073 a_11386_n2838.t1 mux8_1.NAND4F_2.Y.t11 a_11290_n2838.t0 VSS.t311 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X4074 VDD.t4242 A1.t45 MULT_0.NAND2_9.Y.t1 VDD.t4241 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4075 VSS.t768 OR8_0.NOT8_0.A2.t10 OR8_0.S2.t0 VSS.t172 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4076 VSS.t792 Y2.t7 ZFLAG_0.nor4_0.Y.t6 VSS.t791 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X4077 a_n3320_2026.t9 a_n3500_1406.t7 8bit_ADDER_0.S1.t9 VDD.t1624 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X4078 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t6 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t10 a_n8432_n9452.t0 VSS.t1123 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X4079 VDD.t4019 MULT_0.inv_9.Y.t15 a_n13975_n11063.t3 VDD.t4018 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X4080 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t2 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t10 VDD.t1852 VDD.t1851 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4081 mux8_7.NAND4F_4.Y.t3 mux8_7.NAND4F_2.D.t15 VDD.t3142 VDD.t3141 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X4082 V_FLAG_0.XOR2_2.Y.t11 a_3313_4914.t7 a_3493_4914.t3 VSS.t543 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4083 a_7644_n20950.t1 mux8_5.NAND4F_4.B.t15 a_7548_n20950.t0 VSS.t857 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X4084 VDD.t2926 SEL0.t142 mux8_4.NAND4F_6.Y.t7 VDD.t2925 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4085 a_n11274_n17539.t0 B1.t52 XOR8_0.S1.t4 VSS.t943 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4086 XOR8_0.S5.t1 B5.t37 a_n11274_n28476.t0 VSS.t1804 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4087 VDD.t2568 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t18 a_n18998_n4534.t6 VDD.t2567 sky130_fd_pr__pfet_01v8 ad=0.42625 pd=3.06 as=0.45375 ps=3.08 w=2.75 l=0.15
X4088 a_n11840_n11683.t3 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t18 VSS.t1376 VSS.t1375 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4089 VDD.t2924 SEL0.t143 mux8_0.NAND4F_7.Y.t7 VDD.t2923 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4090 a_n29_2026.t8 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t23 VDD.t2265 VDD.t2264 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X4091 a_n12616_1406.t0 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t23 mux8_5.A0.t1 VSS.t165 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4092 a_n10884_1406.t0 A3.t45 VSS.t1853 VSS.t1852 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4093 VDD.t3619 B4.t37 a_n12314_n26419.t3 VDD.t3618 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X4094 a_11194_n21878.t1 mux8_5.NAND4F_7.Y.t11 VSS.t105 VSS.t104 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X4095 a_n21333_2026.t4 A6.t29 VDD.t2835 VDD.t2834 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X4096 Y4.t1 mux8_5.inv_0.A.t10 VDD.t3346 VDD.t3345 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4097 VSS.t556 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t18 a_n19198_1406.t0 VSS.t555 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4098 a_n2744_1406.t0 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t23 8bit_ADDER_0.S1.t1 VSS.t370 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4099 a_n3659_3164.t1 B1.t53 VDD.t1834 VDD.t1833 sky130_fd_pr__pfet_01v8 ad=0.7975 pd=6.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X4100 a_n11274_n20496.t3 B2.t53 XOR8_0.S2.t2 VSS.t226 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4101 VDD.t794 AND8_0.S1.t6 mux8_2.NAND4F_4.Y.t2 VDD.t793 sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
X4102 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t11 a_n14155_n11683.t7 a_n13975_n11063.t0 VDD.t2024 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.45375 ps=3.08 w=2.75 l=0.15
X4103 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t0 MULT_0.4bit_ADDER_2.B2.t23 a_n16690_n11683.t0 VSS.t932 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4104 VDD.t1059 MULT_0.NAND2_2.Y.t10 MULT_0.4bit_ADDER_0.B0.t1 VDD.t1056 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X4105 mux8_0.NAND4F_4.Y.t6 VSS.t975 a_7644_1690.t1 VSS.t841 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X4106 VSS.t1091 mux8_2.NAND4F_9.Y.t14 mux8_2.inv_0.A.t6 VSS.t1090 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X4107 a_n17677_n21025.t9 A4.t29 OR8_0.NOT8_0.A4.t0 VDD.t2204 sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.2112 ps=1.61 w=1.28 l=0.15
X4108 mux8_3.NAND4F_9.Y.t5 mux8_3.NAND4F_7.Y.t11 VDD.t3354 VDD.t3353 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X4109 a_7548_n12822.t1 SEL1.t143 a_7452_n12822.t1 VSS.t1973 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X4110 a_3493_5534.t0 SEL3.t83 VDD.t784 VDD.t783 sky130_fd_pr__pfet_01v8 ad=0.45375 pd=3.08 as=0.42625 ps=3.06 w=2.75 l=0.15
X4111 mux8_0.NAND4F_1.Y.t7 VSS.t2070 VDD.t1909 VDD.t1908 sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
R0 a_n13531_3164.n0 a_n13531_3164.t7 539.788
R1 a_n13531_3164.n1 a_n13531_3164.t5 531.496
R2 a_n13531_3164.n0 a_n13531_3164.t3 490.034
R3 a_n13531_3164.n5 a_n13531_3164.t0 283.788
R4 a_n13531_3164.t1 a_n13531_3164.n5 205.489
R5 a_n13531_3164.n2 a_n13531_3164.t6 182.625
R6 a_n13531_3164.n3 a_n13531_3164.t4 179.054
R7 a_n13531_3164.n2 a_n13531_3164.t2 139.78
R8 a_n13531_3164.n4 a_n13531_3164.n3 101.368
R9 a_n13531_3164.n5 a_n13531_3164.n4 77.9135
R10 a_n13531_3164.n4 a_n13531_3164.n1 76.1557
R11 a_n13531_3164.n1 a_n13531_3164.n0 8.29297
R12 a_n13531_3164.n3 a_n13531_3164.n2 3.57087
R13 a_n13501_3190.n3 a_n13501_3190.n2 121.353
R14 a_n13501_3190.n2 a_n13501_3190.n1 121.001
R15 a_n13501_3190.n2 a_n13501_3190.n0 120.977
R16 a_n13501_3190.n0 a_n13501_3190.t5 30.462
R17 a_n13501_3190.n0 a_n13501_3190.t3 30.462
R18 a_n13501_3190.n1 a_n13501_3190.t2 30.462
R19 a_n13501_3190.n1 a_n13501_3190.t4 30.462
R20 a_n13501_3190.n3 a_n13501_3190.t1 30.462
R21 a_n13501_3190.t0 a_n13501_3190.n3 30.462
R22 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t21 491.64
R23 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t19 491.64
R24 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t13 491.64
R25 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t22 491.64
R26 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t12 485.221
R27 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t16 367.928
R28 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t17 255.588
R29 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t14 224.478
R30 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t15 213.688
R31 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n18 209.19
R32 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t20 139.78
R33 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t23 139.78
R34 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t18 139.78
R35 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n1 120.999
R36 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n0 120.999
R37 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n13 104.489
R38 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 103.258
R39 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n3 92.5005
R40 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n8 86.2638
R41 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n9 85.8873
R42 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n6 85.724
R43 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n16 84.5046
R44 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n14 84.0545
R45 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n8 75.0672
R46 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n11 75.0672
R47 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n6 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n5 73.1255
R48 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n8 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n7 73.1255
R49 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n10 73.1255
R50 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n15 72.3005
R51 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n6 68.8946
R52 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n17 60.9816
R53 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n4 41.9827
R54 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t6 30.462
R55 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t10 30.462
R56 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t9 30.462
R57 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t11 30.462
R58 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t7 30.462
R59 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t8 30.462
R60 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n2 28.124
R61 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n19 17.8661
R62 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n20 17.8661
R63 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n21 17.1217
R64 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n23 15.6329
R65 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t4 11.8205
R66 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t5 11.8205
R67 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t3 11.8205
R68 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t1 11.8205
R69 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t0 11.8205
R70 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t2 11.8205
R71 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 10.8165
R72 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n12 9.3005
R73 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n24 2.50602
R74 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n22 1.8615
R75 VSS.n1332 VSS.n1331 7.282e+06
R76 VSS.n1632 VSS.t688 2.88729e+06
R77 VSS.n1182 VSS.n1181 1.85404e+06
R78 VSS.n1408 VSS.n107 1.63109e+06
R79 VSS.n1333 VSS.n1332 1.0076e+06
R80 VSS.t1195 VSS.t271 979097
R81 VSS.n1408 VSS.t1094 552347
R82 VSS.n363 VSS.n355 473733
R83 VSS.t837 VSS.n1408 202500
R84 VSS.n184 VSS.t192 192754
R85 VSS.n355 VSS.t209 179397
R86 VSS.n1184 VSS.n1183 52956.5
R87 VSS.n868 VSS.n867 52460.5
R88 VSS.n1210 VSS.n1209 46130.2
R89 VSS.n626 VSS.n624 43843
R90 VSS.n983 VSS.n622 43843
R91 VSS.n1019 VSS.n620 43843
R92 VSS.n881 VSS.n610 43843
R93 VSS.n735 VSS.n612 43843
R94 VSS.n915 VSS.n614 43843
R95 VSS.n1053 VSS.n616 43843
R96 VSS.n949 VSS.n618 43843
R97 VSS.n1201 VSS.n1200 40403.2
R98 VSS.n1207 VSS.n1206 39530.2
R99 VSS.n1198 VSS.n1197 39530.2
R100 VSS.n1195 VSS.n1194 39530.2
R101 VSS.n1192 VSS.n1191 39530.2
R102 VSS.n1189 VSS.n1188 39530.2
R103 VSS.n1186 VSS.n1185 39530.2
R104 VSS.n1204 VSS.n1203 38657.1
R105 VSS.n1208 VSS.n1207 37679.4
R106 VSS.n1205 VSS.n1204 37679.4
R107 VSS.n1202 VSS.n1201 37679.4
R108 VSS.n1199 VSS.n1198 37679.4
R109 VSS.n1196 VSS.n1195 37679.4
R110 VSS.n1193 VSS.n1192 37679.4
R111 VSS.n1190 VSS.n1189 37679.4
R112 VSS.n1187 VSS.n1186 37679.4
R113 VSS.n603 VSS.n573 35313.4
R114 VSS.n983 VSS.n624 28593.6
R115 VSS.n1019 VSS.n622 28593.6
R116 VSS.n867 VSS.n610 28593.6
R117 VSS.n881 VSS.n612 28593.6
R118 VSS.n735 VSS.n614 28593.6
R119 VSS.n915 VSS.n616 28593.6
R120 VSS.n1053 VSS.n618 28593.6
R121 VSS.n949 VSS.n620 28593.6
R122 VSS.n1182 VSS.n626 28575.8
R123 VSS.t1094 VSS.t1910 28160
R124 VSS.n1399 VSS.n1397 24230.8
R125 VSS.t560 VSS.n848 22188.4
R126 VSS.n1204 VSS.n612 21841.7
R127 VSS.n1192 VSS.n620 19730.8
R128 VSS.n1189 VSS.n622 19730.8
R129 VSS.n1186 VSS.n624 19730.8
R130 VSS.n1207 VSS.n610 19730.8
R131 VSS.n1198 VSS.n616 19730.8
R132 VSS.n1195 VSS.n618 19730.8
R133 VSS.n1655 VSS.t1323 18634.8
R134 VSS.n792 VSS.n757 18052.9
R135 VSS.n1201 VSS.n614 17992
R136 VSS.n870 VSS.n755 17513.7
R137 VSS.n775 VSS.n758 17513.7
R138 VSS.n809 VSS.n808 17513.7
R139 VSS.n819 VSS.n818 17513.7
R140 VSS.n829 VSS.n828 17513.7
R141 VSS.n1400 VSS.n1399 17346.2
R142 VSS.n766 VSS.n756 16974.5
R143 VSS.n1637 VSS.n104 15508.9
R144 VSS.n869 VSS.n760 15098
R145 VSS.n1401 VSS.n211 14748.5
R146 VSS.n1417 VSS.n107 14167.7
R147 VSS.n1634 VSS.n1633 13515.7
R148 VSS.n1493 VSS.n156 13488.3
R149 VSS.n487 VSS.n124 13455
R150 VSS.n1635 VSS.n107 13377.7
R151 VSS.t1780 VSS.n85 13095.2
R152 VSS.n1634 VSS.n108 12988.6
R153 VSS.n1637 VSS.n1636 12660.2
R154 VSS.t1910 VSS.t1780 12545.2
R155 VSS.t1323 VSS.t1849 12335.7
R156 VSS.n561 VSS.n560 12228.2
R157 VSS.n1401 VSS.n210 12161.6
R158 VSS.n365 VSS.n355 12097.7
R159 VSS.n1493 VSS.n155 11123.2
R160 VSS.n1636 VSS.n1635 10939.5
R161 VSS.n850 VSS.t537 10908.7
R162 VSS.n1436 VSS.n1435 10535.5
R163 VSS.n1435 VSS.n105 10529
R164 VSS.n1417 VSS.n106 10529
R165 VSS.n563 VSS.n562 10076
R166 VSS.n1436 VSS.n104 10064.5
R167 VSS.n1654 VSS.n85 10031
R168 VSS.t1849 VSS.n1654 9821.43
R169 VSS.n354 VSS.n353 9815.03
R170 VSS.n1635 VSS.n1634 9533.6
R171 VSS.n385 VSS.n84 8411.26
R172 VSS.n1494 VSS.n152 8189.68
R173 VSS.n1497 VSS.n152 8189.68
R174 VSS.n356 VSS.n327 8093.35
R175 VSS.n1332 VSS.n573 8041.05
R176 VSS.n1639 VSS.n102 7309.7
R177 VSS.n1185 VSS.n1184 7019.05
R178 VSS.n387 VSS.n386 6721.97
R179 VSS.n364 VSS.n356 6712.94
R180 VSS.n868 VSS.n606 6609.45
R181 VSS.n1400 VSS.n213 6497.02
R182 VSS.n1333 VSS.n574 6453.33
R183 VSS.n1636 VSS.n106 6374.19
R184 VSS.n1211 VSS.n1210 6327.21
R185 VSS.n606 VSS.n605 6098.06
R186 VSS.t1306 VSS.n84 6001.6
R187 VSS.n1486 VSS.n110 5953.41
R188 VSS.n1391 VSS.n108 5940.11
R189 VSS.n1336 VSS.n1335 5799.12
R190 VSS.n1338 VSS.n1337 5799.12
R191 VSS.n1339 VSS.n1338 5799.12
R192 VSS.n1340 VSS.n1339 5799.12
R193 VSS.n1340 VSS.n102 5799.12
R194 VSS.n1337 VSS.n1336 5797.36
R195 VSS.n1632 VSS.n110 5575.11
R196 VSS.n488 VSS.n487 5519.3
R197 VSS.t1687 VSS.n330 5427.65
R198 VSS.t1822 VSS.n335 5427.65
R199 VSS.t67 VSS.n339 5427.65
R200 VSS.n1509 VSS.t351 5422.48
R201 VSS.t53 VSS.n165 5422.48
R202 VSS.t352 VSS.n344 5422.48
R203 VSS.n549 VSS.n121 5387.66
R204 VSS.n1454 VSS.t525 5307.47
R205 VSS.n1401 VSS.t810 5095.85
R206 VSS.n1211 VSS.n603 5073.04
R207 VSS.t513 VSS.n574 4830.05
R208 VSS.n386 VSS.n374 4714.54
R209 VSS.t1263 VSS.n329 4626.5
R210 VSS.t52 VSS.n333 4626.5
R211 VSS.t10 VSS.n337 4626.5
R212 VSS.t1336 VSS.n372 4626.5
R213 VSS.n1517 VSS.t130 4622.1
R214 VSS.n1506 VSS.t657 4622.1
R215 VSS.n1477 VSS.t115 4622.1
R216 VSS.n368 VSS.t790 4622.1
R217 VSS.n327 VSS.t407 4585.88
R218 VSS.n1428 VSS.n199 4417.6
R219 VSS.n1424 VSS.n201 4411.73
R220 VSS.n1210 VSS.n608 4375.51
R221 VSS.t177 VSS.n109 4366.49
R222 VSS.n352 VSS.n350 4347.2
R223 VSS.n353 VSS.n352 4304.69
R224 VSS.n488 VSS.n485 4303.51
R225 VSS.n1335 VSS.n1334 4185.02
R226 VSS.n1638 VSS.n1637 4180.82
R227 VSS.n1636 VSS.n105 4154.84
R228 VSS.n1427 VSS.n1426 4124.22
R229 VSS.n1425 VSS.n1424 4117.1
R230 VSS.n1423 VSS.n85 4117.1
R231 VSS.n1429 VSS.n1428 4110.66
R232 VSS.n351 VSS.n198 4104.92
R233 VSS.n1633 VSS.n109 3979.88
R234 VSS.n367 VSS.n365 3960
R235 VSS.n1653 VSS.n1652 3766.22
R236 VSS.n362 VSS.n356 3733.33
R237 VSS.n606 VSS.n603 3711.47
R238 VSS.t290 VSS.n328 3674.36
R239 VSS.t1761 VSS.n332 3674.36
R240 VSS.t321 VSS.n336 3674.36
R241 VSS.t1138 VSS.n341 3674.36
R242 VSS.n1518 VSS.t988 3670.86
R243 VSS.n1508 VSS.t98 3670.86
R244 VSS.n1478 VSS.t215 3670.86
R245 VSS.t238 VSS.n346 3670.86
R246 VSS.n1459 VSS.n184 3553.85
R247 VSS.n1449 VSS.n1448 3309.37
R248 VSS.t537 VSS.n849 3221.13
R249 VSS.n1401 VSS.n212 3167.08
R250 VSS.n849 VSS.t560 3071.7
R251 VSS.n89 VSS.n88 3040.2
R252 VSS.n1397 VSS.n1396 2966.33
R253 VSS.n1493 VSS.n1492 2896.67
R254 VSS.n351 VSS.t557 2839.47
R255 VSS.n1427 VSS.t535 2839.47
R256 VSS.n1423 VSS.t353 2833.6
R257 VSS.t375 VSS.n102 2825.06
R258 VSS.n1340 VSS.t922 2825.06
R259 VSS.n1339 VSS.t917 2825.06
R260 VSS.n1338 VSS.t870 2825.06
R261 VSS.n1336 VSS.t926 2825.06
R262 VSS.n1335 VSS.t919 2825.06
R263 VSS.n102 VSS.t583 2822.58
R264 VSS.t1639 VSS.n1340 2822.58
R265 VSS.n1339 VSS.t1797 2822.58
R266 VSS.n1338 VSS.t1647 2822.58
R267 VSS.n1337 VSS.t1105 2822.58
R268 VSS.n1337 VSS.t928 2822.58
R269 VSS.n1336 VSS.t221 2822.58
R270 VSS.n1335 VSS.t1189 2822.58
R271 VSS.t259 VSS.n348 2798.4
R272 VSS.n1422 VSS.t1109 2792.53
R273 VSS.n1438 VSS.t831 2786.67
R274 VSS.n319 VSS.t838 2786.67
R275 VSS.n326 VSS.t220 2769.07
R276 VSS.n202 VSS.t261 2769.07
R277 VSS.t401 VSS.t1082 2761.22
R278 VSS.t1862 VSS.t38 2761.22
R279 VSS.t1782 VSS.t298 2761.22
R280 VSS.t705 VSS.t1350 2761.22
R281 VSS.t567 VSS.t1429 2761.22
R282 VSS.t1492 VSS.t958 2761.22
R283 VSS.t133 VSS.t94 2761.22
R284 VSS.t349 VSS.t655 2761.22
R285 VSS.t1279 VSS.t1446 2761.22
R286 VSS.t1261 VSS.t1928 2761.22
R287 VSS.t1501 VSS.t1685 2761.22
R288 VSS.t1816 VSS.t1867 2761.22
R289 VSS.t965 VSS.t1371 2761.22
R290 VSS.t969 VSS.t423 2761.22
R291 VSS.t73 VSS.t472 2761.22
R292 VSS.t863 VSS.t160 2755.61
R293 VSS.n1203 VSS.n1202 2723.81
R294 VSS.n1437 VSS.n1436 2722.13
R295 VSS.n318 VSS.n105 2722.13
R296 VSS.n1418 VSS.n1417 2722.13
R297 VSS.n1639 VSS.n1638 2658.62
R298 VSS.n555 VSS.n545 2623.96
R299 VSS.n869 VSS.n759 2415.69
R300 VSS.n1637 VSS.n103 2341.47
R301 VSS.n357 VSS.n198 2315.3
R302 VSS.n1426 VSS.n200 2313.85
R303 VSS.n1638 VSS.t1669 2149.49
R304 VSS.n354 VSS.t1015 2149.49
R305 VSS.t1334 VSS.n387 2149.49
R306 VSS.t1828 VSS.n1655 2149.49
R307 VSS.n486 VSS.t70 2139.63
R308 VSS.n1334 VSS.n1333 2117.97
R309 VSS.t506 VSS.t1905 2098.88
R310 VSS.n1348 VSS.t951 2062.9
R311 VSS.n1458 VSS.t509 2060.55
R312 VSS.n1334 VSS.n573 2048.36
R313 VSS.n1453 VSS.t502 1981.46
R314 VSS.n1209 VSS.n1208 1850.79
R315 VSS.n1200 VSS.n1199 1850.79
R316 VSS.n1197 VSS.n1196 1850.79
R317 VSS.n1194 VSS.n1193 1850.79
R318 VSS.n1191 VSS.n1190 1850.79
R319 VSS.n1188 VSS.n1187 1850.79
R320 VSS.n850 VSS.n830 1815.53
R321 VSS.n862 VSS.n761 1801.01
R322 VSS.t833 VSS.t1143 1790.31
R323 VSS.t367 VSS.t1895 1790.31
R324 VSS.t1248 VSS.t253 1790.31
R325 VSS.t1850 VSS.t2025 1790.31
R326 VSS.t1121 VSS.t136 1790.31
R327 VSS.t1771 VSS.t175 1790.31
R328 VSS.t1388 VSS.t412 1790.31
R329 VSS.t1603 VSS.t1571 1790.31
R330 VSS.t1069 VSS.t697 1790.31
R331 VSS.t1879 VSS.t1169 1790.31
R332 VSS.t212 VSS.t116 1790.31
R333 VSS.t235 VSS.t312 1790.31
R334 VSS.t292 VSS.t1482 1790.31
R335 VSS.t1763 VSS.t50 1790.31
R336 VSS.t325 VSS.t8 1790.31
R337 VSS.t521 VSS.t1915 1790.31
R338 VSS.t1560 VSS.t1616 1790.31
R339 VSS.t1043 VSS.t1812 1790.31
R340 VSS.t1244 VSS.t632 1790.31
R341 VSS.t1528 VSS.t1674 1790.31
R342 VSS.n1349 VSS.t1400 1758.41
R343 VSS.n1387 VSS.t1575 1758.41
R344 VSS.t777 VSS.n184 1720.14
R345 VSS.n851 VSS.n761 1592.91
R346 VSS.n605 VSS.n604 1591.74
R347 VSS.n755 VSS.t1514 1574.51
R348 VSS.n766 VSS.t544 1574.51
R349 VSS.n792 VSS.t748 1574.51
R350 VSS.n775 VSS.t1776 1574.51
R351 VSS.n808 VSS.t1539 1574.51
R352 VSS.n818 VSS.t1330 1574.51
R353 VSS.n828 VSS.t1270 1574.51
R354 VSS.n759 VSS.t1596 1574.51
R355 VSS.n830 VSS.t842 1559.22
R356 VSS.n605 VSS.t1612 1559.22
R357 VSS.n211 VSS.t415 1559.22
R358 VSS.n156 VSS.t1253 1559.22
R359 VSS.n560 VSS.t1181 1559.22
R360 VSS.t1464 VSS.n1429 1494.34
R361 VSS.n1425 VSS.t1076 1486.15
R362 VSS.n384 VSS.t1284 1467.69
R363 VSS.n377 VSS.t1292 1464.62
R364 VSS.n488 VSS.t1123 1463.87
R365 VSS.n488 VSS.t101 1462.48
R366 VSS.n1430 VSS.t1173 1454.37
R367 VSS.n361 VSS.t1183 1448.22
R368 VSS.n376 VSS.n106 1427.69
R369 VSS.n1435 VSS.n1434 1426.69
R370 VSS.t552 VSS.n1346 1396.52
R371 VSS.t960 VSS.n1386 1396.52
R372 VSS.n1226 VSS.n122 1387.3
R373 VSS.n387 VSS.n327 1375.08
R374 VSS.n1500 VSS.t1132 1365.68
R375 VSS.n385 VSS.t1920 1350.77
R376 VSS.n1404 VSS.n1403 1337.13
R377 VSS.n848 VSS.n847 1320.03
R378 VSS.n496 VSS.t453 1310.38
R379 VSS.n521 VSS.t952 1310.38
R380 VSS.n1655 VSS.n84 1288.89
R381 VSS.n1500 VSS.n152 1286.77
R382 VSS.n155 VSS.t149 1284.8
R383 VSS.n210 VSS.t670 1284.8
R384 VSS.n563 VSS.t499 1284.8
R385 VSS.n353 VSS.n104 1284.25
R386 VSS.n870 VSS.n869 1186.27
R387 VSS.n869 VSS.n756 1186.27
R388 VSS.n869 VSS.n757 1186.27
R389 VSS.n869 VSS.n758 1186.27
R390 VSS.n850 VSS.n809 1186.27
R391 VSS.n850 VSS.n819 1186.27
R392 VSS.n850 VSS.n829 1186.27
R393 VSS.n485 VSS.t428 1157.89
R394 VSS.t954 VSS.n488 1139.24
R395 VSS.t300 VSS.n493 1116.96
R396 VSS.n522 VSS.t707 1116.96
R397 VSS.n267 VSS.t192 1116.96
R398 VSS.t1178 VSS.n1612 1063.15
R399 VSS.n832 VSS.n830 1054.96
R400 VSS.t1524 VSS.n1211 1033.39
R401 VSS.n1131 VSS.t982 1032.02
R402 VSS.n1136 VSS.t1010 1032.02
R403 VSS.n1139 VSS.t975 1032.02
R404 VSS.n1128 VSS.t1001 1032.02
R405 VSS.n1126 VSS.t1003 1032.02
R406 VSS.n1035 VSS.t242 1011.19
R407 VSS.n999 VSS.t613 1011.19
R408 VSS.n1165 VSS.t167 1011.19
R409 VSS.n965 VSS.t328 1011.19
R410 VSS.n1069 VSS.t957 1011.19
R411 VSS.n931 VSS.t208 1011.19
R412 VSS.n1098 VSS.t396 1011.19
R413 VSS.n897 VSS.t275 1011.19
R414 VSS.n1122 VSS.t841 1011.19
R415 VSS.n189 VSS.n104 990.187
R416 VSS.n1039 VSS.t1050 988.638
R417 VSS.n1003 VSS.t527 988.638
R418 VSS.t127 VSS.n1163 988.638
R419 VSS.n969 VSS.t87 988.638
R420 VSS.n1073 VSS.t196 988.638
R421 VSS.n935 VSS.t562 988.638
R422 VSS.t304 VSS.n1096 988.638
R423 VSS.n901 VSS.t433 988.638
R424 VSS.t983 VSS.n1120 988.638
R425 VSS.n608 VSS.t1856 979.592
R426 VSS.n1041 VSS.t296 979.24
R427 VSS.n1005 VSS.t736 979.24
R428 VSS.t1499 VSS.n1159 979.24
R429 VSS.n971 VSS.t1541 979.24
R430 VSS.n1075 VSS.t16 979.24
R431 VSS.n937 VSS.t0 979.24
R432 VSS.t31 VSS.n1092 979.24
R433 VSS.n903 VSS.t1543 979.24
R434 VSS.t776 VSS.n1116 979.24
R435 VSS.n1206 VSS.n1205 977.779
R436 VSS.n1180 VSS.t199 971.722
R437 VSS.t19 VSS.n1023 971.529
R438 VSS.t1157 VSS.n987 971.529
R439 VSS.t674 VSS.n953 971.529
R440 VSS.t3 VSS.n1057 971.529
R441 VSS.t822 VSS.n919 971.529
R442 VSS.n737 VSS.t1051 971.529
R443 VSS.t43 VSS.n885 971.529
R444 VSS.n866 VSS.t1002 971.529
R445 VSS.t1092 VSS.t814 934.428
R446 VSS.n761 VSS.n760 927.452
R447 VSS.t860 VSS.n490 887.09
R448 VSS.n495 VSS.t163 887.09
R449 VSS.n269 VSS.t1356 887.09
R450 VSS.n355 VSS.n354 885.422
R451 VSS.n1459 VSS.t75 882.499
R452 VSS.t1651 VSS.t183 851.87
R453 VSS.t1635 VSS.t1579 843.919
R454 VSS.t1287 VSS.t1840 818.846
R455 VSS.n1575 VSS.t1392 817.013
R456 VSS.n487 VSS.n486 792.374
R457 VSS.n1183 VSS.t1443 788.635
R458 VSS.t1856 VSS.t1155 783.674
R459 VSS.n843 VSS.t340 754.973
R460 VSS.t465 VSS.n208 707.75
R461 VSS.n217 VSS.t1607 674.043
R462 VSS.n1485 VSS.t394 674.043
R463 VSS.n548 VSS.t692 674.043
R464 VSS.n362 VSS.t1300 618.029
R465 VSS.t878 VSS.n574 611.736
R466 VSS.n488 VSS.t1005 611.736
R467 VSS.n488 VSS.t1008 611.736
R468 VSS.n488 VSS.t1012 611.736
R469 VSS.n1612 VSS.t255 602.597
R470 VSS.t282 VSS.n1497 600.419
R471 VSS.n1497 VSS.t1903 600.419
R472 VSS.t1186 VSS.n1494 600.419
R473 VSS.n1494 VSS.t121 600.419
R474 VSS.n191 VSS.n190 589.682
R475 VSS.n348 VSS.n347 589.682
R476 VSS.n1439 VSS.n1438 589.682
R477 VSS.n1458 VSS.n1457 589.682
R478 VSS.n1453 VSS.n1452 589.682
R479 VSS.n187 VSS.n186 589.682
R480 VSS.n361 VSS.n360 589.682
R481 VSS.n1431 VSS.n1430 589.682
R482 VSS.n326 VSS.n325 589.682
R483 VSS.n384 VSS.n383 589.682
R484 VSS.n378 VSS.n377 589.682
R485 VSS.n203 VSS.n202 589.682
R486 VSS.n1422 VSS.n1421 589.682
R487 VSS.n1405 VSS.n1404 589.682
R488 VSS.n1411 VSS.n87 589.682
R489 VSS.n320 VSS.n319 589.682
R490 VSS.n1307 VSS.n1237 589.667
R491 VSS.n1307 VSS.n1238 589.667
R492 VSS.n1307 VSS.n1239 589.667
R493 VSS.n1307 VSS.n1240 589.667
R494 VSS.n1307 VSS.n1241 589.667
R495 VSS.n1307 VSS.n1242 589.667
R496 VSS.n1307 VSS.n1243 589.667
R497 VSS.n1307 VSS.n1306 589.667
R498 VSS.n1561 VSS.n1559 589.667
R499 VSS.n1561 VSS.n1557 589.667
R500 VSS.n1561 VSS.n1555 589.667
R501 VSS.n1561 VSS.n1553 589.667
R502 VSS.n1561 VSS.n1551 589.667
R503 VSS.n1561 VSS.n1549 589.667
R504 VSS.n1561 VSS.n1547 589.667
R505 VSS.n1565 VSS.n1564 589.667
R506 VSS.n847 VSS.n846 589.658
R507 VSS.n1307 VSS.n1228 589.654
R508 VSS.n1307 VSS.n1229 589.654
R509 VSS.n1307 VSS.n1230 589.654
R510 VSS.n1307 VSS.n1231 589.654
R511 VSS.n1307 VSS.n1232 589.654
R512 VSS.n1307 VSS.n1233 589.654
R513 VSS.n1307 VSS.n1234 589.654
R514 VSS.n1307 VSS.n1235 589.654
R515 VSS.n1562 VSS.n1561 589.654
R516 VSS.n1561 VSS.n1545 589.654
R517 VSS.n1561 VSS.n1544 589.654
R518 VSS.n1561 VSS.n1543 589.654
R519 VSS.n1561 VSS.n1542 589.654
R520 VSS.n1561 VSS.n1541 589.654
R521 VSS.n1561 VSS.n1540 589.654
R522 VSS.n1561 VSS.n1539 589.654
R523 VSS.n1307 VSS.n1236 589.65
R524 VSS.n215 VSS.n210 589.65
R525 VSS.n218 VSS.n217 589.65
R526 VSS.n227 VSS.n213 589.65
R527 VSS.n221 VSS.n211 589.65
R528 VSS.n223 VSS.n212 589.65
R529 VSS.n228 VSS.n212 589.65
R530 VSS.n225 VSS.n212 589.65
R531 VSS.n219 VSS.n212 589.65
R532 VSS.n1485 VSS.n1484 589.65
R533 VSS.n1487 VSS.n1486 589.65
R534 VSS.n1481 VSS.n155 589.65
R535 VSS.n160 VSS.n156 589.65
R536 VSS.n1492 VSS.n1491 589.65
R537 VSS.n1492 VSS.n157 589.65
R538 VSS.n1492 VSS.n159 589.65
R539 VSS.n1492 VSS.n158 589.65
R540 VSS.n678 VSS.n677 589.65
R541 VSS.n676 VSS.n675 589.65
R542 VSS.n672 VSS.n583 589.65
R543 VSS.n665 VSS.n664 589.65
R544 VSS.n667 VSS.n666 589.65
R545 VSS.n668 VSS.n584 589.65
R546 VSS.n686 VSS.n685 589.65
R547 VSS.n684 VSS.n683 589.65
R548 VSS.n680 VSS.n585 589.65
R549 VSS.n658 VSS.n657 589.65
R550 VSS.n660 VSS.n659 589.65
R551 VSS.n661 VSS.n586 589.65
R552 VSS.n694 VSS.n693 589.65
R553 VSS.n692 VSS.n691 589.65
R554 VSS.n688 VSS.n587 589.65
R555 VSS.n651 VSS.n650 589.65
R556 VSS.n653 VSS.n652 589.65
R557 VSS.n654 VSS.n588 589.65
R558 VSS.n702 VSS.n701 589.65
R559 VSS.n700 VSS.n699 589.65
R560 VSS.n696 VSS.n589 589.65
R561 VSS.n644 VSS.n643 589.65
R562 VSS.n646 VSS.n645 589.65
R563 VSS.n647 VSS.n590 589.65
R564 VSS.n710 VSS.n709 589.65
R565 VSS.n708 VSS.n707 589.65
R566 VSS.n704 VSS.n591 589.65
R567 VSS.n843 VSS.n831 589.65
R568 VSS.n843 VSS.n842 589.65
R569 VSS.n755 VSS.n754 589.65
R570 VSS.n767 VSS.n766 589.65
R571 VSS.n793 VSS.n792 589.65
R572 VSS.n776 VSS.n775 589.65
R573 VSS.n808 VSS.n807 589.65
R574 VSS.n818 VSS.n817 589.65
R575 VSS.n828 VSS.n827 589.65
R576 VSS.n784 VSS.n759 589.65
R577 VSS.n564 VSS.n563 589.65
R578 VSS.n556 VSS.n555 589.65
R579 VSS.n555 VSS.n552 589.65
R580 VSS.n555 VSS.n554 589.65
R581 VSS.n555 VSS.n553 589.65
R582 VSS.n548 VSS.n547 589.65
R583 VSS.n550 VSS.n549 589.65
R584 VSS.n560 VSS.n559 589.65
R585 VSS.n1561 VSS.n1560 589.65
R586 VSS.t649 VSS.n756 568.013
R587 VSS.t1946 VSS.n612 562.14
R588 VSS.n819 VSS.t546 553.633
R589 VSS.n829 VSS.t1505 553.633
R590 VSS.t1454 VSS.n870 553.633
R591 VSS.t1298 VSS.n758 553.633
R592 VSS.t481 VSS.n760 553.633
R593 VSS.n809 VSS.t335 553.633
R594 VSS.n1561 VSS.n122 553.595
R595 VSS.t894 VSS.n1639 549.37
R596 VSS.t359 VSS.n624 547.913
R597 VSS.t1917 VSS.n622 547.913
R598 VSS.t1614 VSS.n610 547.913
R599 VSS.t1778 VSS.n616 547.913
R600 VSS.t728 VSS.n618 547.913
R601 VSS.t1936 VSS.n620 547.913
R602 VSS.n1652 VSS.t1103 547.15
R603 VSS.n304 VSS.t987 540.38
R604 VSS.n434 VSS.t978 540.38
R605 VSS.n472 VSS.t995 540.38
R606 VSS.t1090 VSS.n757 539.962
R607 VSS.t387 VSS.t911 538.777
R608 VSS.t872 VSS.t387 538.777
R609 VSS.t1142 VSS.t872 538.777
R610 VSS.t1145 VSS.t1142 538.777
R611 VSS.t1140 VSS.t1145 538.777
R612 VSS.t1453 VSS.t1452 538.777
R613 VSS.t1451 VSS.t1453 538.777
R614 VSS.t1196 VSS.t1451 538.777
R615 VSS.t1549 VSS.t1196 538.777
R616 VSS.t1198 VSS.t1549 538.777
R617 VSS.t1127 VSS.t829 538.777
R618 VSS.t835 VSS.t1127 538.777
R619 VSS.t1081 VSS.t835 538.777
R620 VSS.t1080 VSS.t1081 538.777
R621 VSS.t1079 VSS.t1080 538.777
R622 VSS.t279 VSS.t1274 538.777
R623 VSS.t278 VSS.t279 538.777
R624 VSS.t620 VSS.t278 538.777
R625 VSS.t624 VSS.t620 538.777
R626 VSS.t622 VSS.t624 538.777
R627 VSS.t1302 VSS.t1304 538.777
R628 VSS.t403 VSS.t1302 538.777
R629 VSS.t370 VSS.t403 538.777
R630 VSS.t369 VSS.t370 538.777
R631 VSS.t366 VSS.t369 538.777
R632 VSS.t767 VSS.t765 538.777
R633 VSS.t765 VSS.t766 538.777
R634 VSS.t766 VSS.t1148 538.777
R635 VSS.t1148 VSS.t1146 538.777
R636 VSS.t1146 VSS.t1150 538.777
R637 VSS.t1911 VSS.t1899 538.777
R638 VSS.t1899 VSS.t1901 538.777
R639 VSS.t1901 VSS.t1858 538.777
R640 VSS.t1858 VSS.t1864 538.777
R641 VSS.t1864 VSS.t1861 538.777
R642 VSS.t399 VSS.t576 538.777
R643 VSS.t576 VSS.t400 538.777
R644 VSS.t400 VSS.t1225 538.777
R645 VSS.t1225 VSS.t1551 538.777
R646 VSS.t1551 VSS.t592 538.777
R647 VSS.t34 VSS.t40 538.777
R648 VSS.t40 VSS.t36 538.777
R649 VSS.t36 VSS.t1237 538.777
R650 VSS.t1237 VSS.t1250 538.777
R651 VSS.t1250 VSS.t1251 538.777
R652 VSS.t1557 VSS.t414 538.777
R653 VSS.t414 VSS.t1513 538.777
R654 VSS.t1513 VSS.t436 538.777
R655 VSS.t436 VSS.t434 538.777
R656 VSS.t434 VSS.t438 538.777
R657 VSS.t119 VSS.t257 538.777
R658 VSS.t257 VSS.t249 538.777
R659 VSS.t249 VSS.t431 538.777
R660 VSS.t431 VSS.t159 538.777
R661 VSS.t159 VSS.t432 538.777
R662 VSS.t747 VSS.t102 538.777
R663 VSS.t746 VSS.t747 538.777
R664 VSS.t157 VSS.t746 538.777
R665 VSS.t155 VSS.t157 538.777
R666 VSS.t153 VSS.t155 538.777
R667 VSS.t858 VSS.t861 538.777
R668 VSS.t865 VSS.t858 538.777
R669 VSS.t2028 VSS.t865 538.777
R670 VSS.t2027 VSS.t2028 538.777
R671 VSS.t2030 VSS.t2027 538.777
R672 VSS.t2024 VSS.t2023 538.777
R673 VSS.t2022 VSS.t2024 538.777
R674 VSS.t1117 VSS.t2022 538.777
R675 VSS.t1115 VSS.t1117 538.777
R676 VSS.t1113 VSS.t1115 538.777
R677 VSS.t1852 VSS.t1837 538.777
R678 VSS.t1846 VSS.t1852 538.777
R679 VSS.t302 VSS.t1846 538.777
R680 VSS.t297 VSS.t302 538.777
R681 VSS.t303 VSS.t297 538.777
R682 VSS.t774 VSS.t775 538.777
R683 VSS.t773 VSS.t774 538.777
R684 VSS.t474 VSS.t773 538.777
R685 VSS.t478 VSS.t474 538.777
R686 VSS.t476 VSS.t478 538.777
R687 VSS.t1784 VSS.t1786 538.777
R688 VSS.t1788 VSS.t1784 538.777
R689 VSS.t162 VSS.t1788 538.777
R690 VSS.t138 VSS.t162 538.777
R691 VSS.t165 VSS.t138 538.777
R692 VSS.t580 VSS.t1075 538.777
R693 VSS.t669 VSS.t580 538.777
R694 VSS.t383 VSS.t669 538.777
R695 VSS.t381 VSS.t383 538.777
R696 VSS.t379 VSS.t381 538.777
R697 VSS.t808 VSS.t816 538.777
R698 VSS.t1119 VSS.t808 538.777
R699 VSS.t702 VSS.t1119 538.777
R700 VSS.t703 VSS.t702 538.777
R701 VSS.t704 VSS.t703 538.777
R702 VSS.t1548 VSS.t1547 538.777
R703 VSS.t1547 VSS.t1546 538.777
R704 VSS.t1546 VSS.t265 538.777
R705 VSS.t265 VSS.t269 538.777
R706 VSS.t269 VSS.t267 538.777
R707 VSS.t1354 VSS.t1352 538.777
R708 VSS.t1352 VSS.t1357 538.777
R709 VSS.t1357 VSS.t1774 538.777
R710 VSS.t1774 VSS.t1773 538.777
R711 VSS.t1773 VSS.t1770 538.777
R712 VSS.t64 VSS.t66 538.777
R713 VSS.t66 VSS.t65 538.777
R714 VSS.t65 VSS.t730 538.777
R715 VSS.t730 VSS.t734 538.777
R716 VSS.t734 VSS.t732 538.777
R717 VSS.t193 VSS.t189 538.777
R718 VSS.t189 VSS.t179 538.777
R719 VSS.t179 VSS.t1433 538.777
R720 VSS.t1433 VSS.t1431 538.777
R721 VSS.t1431 VSS.t1428 538.777
R722 VSS.t1769 VSS.t1767 538.777
R723 VSS.t1768 VSS.t1769 538.777
R724 VSS.t1066 VSS.t1768 538.777
R725 VSS.t1062 VSS.t1066 538.777
R726 VSS.t1064 VSS.t1062 538.777
R727 VSS.t550 VSS.t553 538.777
R728 VSS.t555 VSS.t550 538.777
R729 VSS.t411 VSS.t555 538.777
R730 VSS.t1208 VSS.t411 538.777
R731 VSS.t1206 VSS.t1208 538.777
R732 VSS.t804 VSS.t227 538.777
R733 VSS.t559 VSS.t804 538.777
R734 VSS.t715 VSS.t559 538.777
R735 VSS.t719 VSS.t715 538.777
R736 VSS.t717 VSS.t719 538.777
R737 VSS.t1398 VSS.t1402 538.777
R738 VSS.t1390 VSS.t1398 538.777
R739 VSS.t1490 VSS.t1390 538.777
R740 VSS.t1495 VSS.t1490 538.777
R741 VSS.t1491 VSS.t1495 538.777
R742 VSS.t597 VSS.t598 538.777
R743 VSS.t598 VSS.t599 538.777
R744 VSS.t599 VSS.t608 538.777
R745 VSS.t608 VSS.t606 538.777
R746 VSS.t606 VSS.t610 538.777
R747 VSS.t85 VSS.t83 538.777
R748 VSS.t83 VSS.t961 538.777
R749 VSS.t961 VSS.t1600 538.777
R750 VSS.t1600 VSS.t1605 538.777
R751 VSS.t1605 VSS.t1601 538.777
R752 VSS.t1256 VSS.t1258 538.777
R753 VSS.t1258 VSS.t1257 538.777
R754 VSS.t1257 VSS.t800 538.777
R755 VSS.t800 VSS.t802 538.777
R756 VSS.t802 VSS.t798 538.777
R757 VSS.t1159 VSS.t1587 538.777
R758 VSS.t1587 VSS.t1573 538.777
R759 VSS.t1573 VSS.t1667 538.777
R760 VSS.t1667 VSS.t1672 538.777
R761 VSS.t1672 VSS.t1671 538.777
R762 VSS.t1598 VSS.t24 538.777
R763 VSS.t24 VSS.t1599 538.777
R764 VSS.t1599 VSS.t1758 538.777
R765 VSS.t1758 VSS.t1756 538.777
R766 VSS.t1756 VSS.t1754 538.777
R767 VSS.t990 VSS.t980 538.777
R768 VSS.t980 VSS.t1028 538.777
R769 VSS.t1028 VSS.t1068 538.777
R770 VSS.t1068 VSS.t1071 538.777
R771 VSS.t1071 VSS.t1072 538.777
R772 VSS.t763 VSS.t170 538.777
R773 VSS.t170 VSS.t171 538.777
R774 VSS.t171 VSS.t143 538.777
R775 VSS.t143 VSS.t145 538.777
R776 VSS.t145 VSS.t147 538.777
R777 VSS.t635 VSS.t637 538.777
R778 VSS.t637 VSS.t699 538.777
R779 VSS.t699 VSS.t129 538.777
R780 VSS.t129 VSS.t132 538.777
R781 VSS.t132 VSS.t135 538.777
R782 VSS.t498 VSS.t548 538.777
R783 VSS.t548 VSS.t549 538.777
R784 VSS.t549 VSS.t139 538.777
R785 VSS.t139 VSS.t141 538.777
R786 VSS.t141 VSS.t319 538.777
R787 VSS.t96 VSS.t99 538.777
R788 VSS.t99 VSS.t1217 538.777
R789 VSS.t1217 VSS.t1878 538.777
R790 VSS.t1878 VSS.t1881 538.777
R791 VSS.t1881 VSS.t1882 538.777
R792 VSS.t497 VSS.t496 538.777
R793 VSS.t496 VSS.t575 538.777
R794 VSS.t575 VSS.t1537 538.777
R795 VSS.t1537 VSS.t1086 538.777
R796 VSS.t1086 VSS.t1088 538.777
R797 VSS.t1165 VSS.t1163 538.777
R798 VSS.t1163 VSS.t1167 538.777
R799 VSS.t1167 VSS.t106 538.777
R800 VSS.t106 VSS.t653 538.777
R801 VSS.t653 VSS.t654 538.777
R802 VSS.t1875 VSS.t1874 538.777
R803 VSS.t1873 VSS.t1875 538.777
R804 VSS.t750 VSS.t1873 538.777
R805 VSS.t754 VSS.t750 538.777
R806 VSS.t752 VSS.t754 538.777
R807 VSS.t345 VSS.t343 538.777
R808 VSS.t347 VSS.t345 538.777
R809 VSS.t218 VSS.t347 538.777
R810 VSS.t217 VSS.t218 538.777
R811 VSS.t214 VSS.t217 538.777
R812 VSS.t1154 VSS.t1153 538.777
R813 VSS.t1153 VSS.t1152 538.777
R814 VSS.t1152 VSS.t1830 538.777
R815 VSS.t1830 VSS.t1832 538.777
R816 VSS.t1832 VSS.t462 538.777
R817 VSS.t109 VSS.t111 538.777
R818 VSS.t111 VSS.t113 538.777
R819 VSS.t113 VSS.t1449 538.777
R820 VSS.t1449 VSS.t1450 538.777
R821 VSS.t1450 VSS.t1445 538.777
R822 VSS.t1223 VSS.t1222 538.777
R823 VSS.t1224 VSS.t1223 538.777
R824 VSS.t1200 VSS.t1224 538.777
R825 VSS.t1202 VSS.t1200 538.777
R826 VSS.t1204 VSS.t1202 538.777
R827 VSS.t1275 VSS.t1281 538.777
R828 VSS.t1277 VSS.t1275 538.777
R829 VSS.t1349 VSS.t1277 538.777
R830 VSS.t237 VSS.t1349 538.777
R831 VSS.t240 VSS.t237 538.777
R832 VSS.t337 VSS.t338 538.777
R833 VSS.t338 VSS.t339 538.777
R834 VSS.t339 VSS.t1404 538.777
R835 VSS.t1404 VSS.t1406 538.777
R836 VSS.t1406 VSS.t1408 538.777
R837 VSS.t314 VSS.t786 538.777
R838 VSS.t786 VSS.t788 538.777
R839 VSS.t788 VSS.t1020 538.777
R840 VSS.t1020 VSS.t1018 538.777
R841 VSS.t1018 VSS.t997 538.777
R842 VSS.t362 VSS.t361 538.777
R843 VSS.t363 VSS.t362 538.777
R844 VSS.t1056 VSS.t363 538.777
R845 VSS.t1058 VSS.t1056 538.777
R846 VSS.t1060 VSS.t1058 538.777
R847 VSS.t999 VSS.t993 538.777
R848 VSS.t993 VSS.t985 538.777
R849 VSS.t985 VSS.t289 538.777
R850 VSS.t289 VSS.t294 538.777
R851 VSS.t294 VSS.t295 538.777
R852 VSS.t518 VSS.t519 538.777
R853 VSS.t519 VSS.t517 538.777
R854 VSS.t517 VSS.t601 538.777
R855 VSS.t601 VSS.t846 538.777
R856 VSS.t846 VSS.t946 538.777
R857 VSS.t1478 VSS.t1480 538.777
R858 VSS.t1480 VSS.t1484 538.777
R859 VSS.t1484 VSS.t1266 538.777
R860 VSS.t1266 VSS.t1260 538.777
R861 VSS.t1260 VSS.t1265 538.777
R862 VSS.t845 VSS.t342 538.777
R863 VSS.t342 VSS.t844 538.777
R864 VSS.t844 VSS.t665 538.777
R865 VSS.t665 VSS.t530 538.777
R866 VSS.t530 VSS.t532 538.777
R867 VSS.t1930 VSS.t1932 538.777
R868 VSS.t1932 VSS.t1934 538.777
R869 VSS.t1934 VSS.t1760 538.777
R870 VSS.t1760 VSS.t1765 538.777
R871 VSS.t1765 VSS.t1766 538.777
R872 VSS.t950 VSS.t949 538.777
R873 VSS.t949 VSS.t948 538.777
R874 VSS.t948 VSS.t1231 538.777
R875 VSS.t1231 VSS.t1233 538.777
R876 VSS.t1233 VSS.t1235 538.777
R877 VSS.t46 VSS.t44 538.777
R878 VSS.t44 VSS.t48 538.777
R879 VSS.t48 VSS.t1503 538.777
R880 VSS.t1503 VSS.t1504 538.777
R881 VSS.t1504 VSS.t1500 538.777
R882 VSS.t1688 VSS.t1690 538.777
R883 VSS.t1690 VSS.t1691 538.777
R884 VSS.t1691 VSS.t1658 538.777
R885 VSS.t1658 VSS.t1662 538.777
R886 VSS.t1662 VSS.t1660 538.777
R887 VSS.t1679 VSS.t1681 538.777
R888 VSS.t1681 VSS.t1683 538.777
R889 VSS.t1683 VSS.t324 538.777
R890 VSS.t324 VSS.t323 538.777
R891 VSS.t323 VSS.t327 538.777
R892 VSS.t709 VSS.t710 538.777
R893 VSS.t710 VSS.t711 538.777
R894 VSS.t711 VSS.t29 538.777
R895 VSS.t29 VSS.t25 538.777
R896 VSS.t25 VSS.t27 538.777
R897 VSS.t11 VSS.t4 538.777
R898 VSS.t4 VSS.t6 538.777
R899 VSS.t6 VSS.t1818 538.777
R900 VSS.t1818 VSS.t1819 538.777
R901 VSS.t1819 VSS.t1821 538.777
R902 VSS.t356 VSS.t357 538.777
R903 VSS.t357 VSS.t358 538.777
R904 VSS.t358 VSS.t1507 538.777
R905 VSS.t1507 VSS.t1509 538.777
R906 VSS.t1509 VSS.t1511 538.777
R907 VSS.t1869 VSS.t1871 538.777
R908 VSS.t1871 VSS.t1865 538.777
R909 VSS.t1865 VSS.t520 538.777
R910 VSS.t520 VSS.t523 538.777
R911 VSS.t523 VSS.t524 538.777
R912 VSS.t126 VSS.t124 538.777
R913 VSS.t124 VSS.t125 538.777
R914 VSS.t125 VSS.t659 538.777
R915 VSS.t659 VSS.t661 538.777
R916 VSS.t661 VSS.t663 538.777
R917 VSS.t1944 VSS.t1893 538.777
R918 VSS.t1893 VSS.t1887 538.777
R919 VSS.t1887 VSS.t1332 538.777
R920 VSS.t1332 VSS.t1333 538.777
R921 VSS.t1333 VSS.t1338 538.777
R922 VSS.t1418 VSS.t1416 538.777
R923 VSS.t1416 VSS.t1417 538.777
R924 VSS.t1417 VSS.t1419 538.777
R925 VSS.t1419 VSS.t1421 538.777
R926 VSS.t1421 VSS.t1423 538.777
R927 VSS.t1022 VSS.t1025 538.777
R928 VSS.t1025 VSS.t1031 538.777
R929 VSS.t1031 VSS.t1563 538.777
R930 VSS.t1563 VSS.t1562 538.777
R931 VSS.t1562 VSS.t1559 538.777
R932 VSS.t1055 VSS.t1054 538.777
R933 VSS.t1054 VSS.t1348 538.777
R934 VSS.t1348 VSS.t449 538.777
R935 VSS.t449 VSS.t451 538.777
R936 VSS.t451 VSS.t447 538.777
R937 VSS.t1622 VSS.t1620 538.777
R938 VSS.t1620 VSS.t1618 538.777
R939 VSS.t1618 VSS.t964 538.777
R940 VSS.t964 VSS.t963 538.777
R941 VSS.t963 VSS.t528 538.777
R942 VSS.t762 VSS.t761 538.777
R943 VSS.t761 VSS.t760 538.777
R944 VSS.t760 VSS.t1035 538.777
R945 VSS.t1035 VSS.t1039 538.777
R946 VSS.t1039 VSS.t1037 538.777
R947 VSS.t1052 VSS.t1375 538.777
R948 VSS.t1375 VSS.t1373 538.777
R949 VSS.t1373 VSS.t1046 538.777
R950 VSS.t1046 VSS.t1045 538.777
R951 VSS.t1045 VSS.t1042 538.777
R952 VSS.t616 VSS.t617 538.777
R953 VSS.t617 VSS.t615 538.777
R954 VSS.t615 VSS.t1938 538.777
R955 VSS.t1938 VSS.t1942 538.777
R956 VSS.t1942 VSS.t1940 538.777
R957 VSS.t1814 VSS.t1810 538.777
R958 VSS.t1810 VSS.t1808 538.777
R959 VSS.t1808 VSS.t972 538.777
R960 VSS.t972 VSS.t971 538.777
R961 VSS.t971 VSS.t956 538.777
R962 VSS.t1048 VSS.t1047 538.777
R963 VSS.t1047 VSS.t1049 538.777
R964 VSS.t1049 VSS.t827 538.777
R965 VSS.t827 VSS.t823 538.777
R966 VSS.t823 VSS.t825 538.777
R967 VSS.t421 VSS.t419 538.777
R968 VSS.t419 VSS.t417 538.777
R969 VSS.t417 VSS.t634 538.777
R970 VSS.t634 VSS.t630 538.777
R971 VSS.t630 VSS.t629 538.777
R972 VSS.t796 VSS.t797 538.777
R973 VSS.t795 VSS.t796 538.777
R974 VSS.t81 VSS.t795 538.777
R975 VSS.t79 VSS.t81 538.777
R976 VSS.t405 VSS.t79 538.777
R977 VSS.t1240 VSS.t1242 538.777
R978 VSS.t1238 VSS.t1240 538.777
R979 VSS.t69 VSS.t1238 538.777
R980 VSS.t932 VSS.t69 538.777
R981 VSS.t72 VSS.t932 538.777
R982 VSS.t646 VSS.t647 538.777
R983 VSS.t647 VSS.t648 538.777
R984 VSS.t648 VSS.t1414 538.777
R985 VSS.t1414 VSS.t1317 538.777
R986 VSS.t1317 VSS.t1315 538.777
R987 VSS.t468 VSS.t470 538.777
R988 VSS.t470 VSS.t466 538.777
R989 VSS.t466 VSS.t1678 538.777
R990 VSS.t1678 VSS.t1677 538.777
R991 VSS.t1677 VSS.t1676 538.777
R992 VSS.t1255 VSS.t769 538.777
R993 VSS.t770 VSS.t1255 538.777
R994 VSS.t1192 VSS.t770 538.777
R995 VSS.t1339 VSS.t1192 538.777
R996 VSS.t1341 VSS.t1339 538.777
R997 VSS.t1532 VSS.t1526 538.777
R998 VSS.t1530 VSS.t1532 538.777
R999 VSS.t1827 VSS.t1530 538.777
R1000 VSS.t1826 VSS.t1827 538.777
R1001 VSS.t1825 VSS.t1826 538.777
R1002 VSS.t1609 VSS.t1595 538.777
R1003 VSS.t1595 VSS.t1594 538.777
R1004 VSS.t1594 VSS.t1229 538.777
R1005 VSS.t1229 VSS.t1227 538.777
R1006 VSS.t1227 VSS.t391 538.777
R1007 VSS.t13 VSS.n614 534.388
R1008 VSS.t1346 VSS.n851 524.718
R1009 VSS.t1577 VSS.n574 518.669
R1010 VSS.t911 VSS.t878 516.327
R1011 VSS.t1143 VSS.t1198 516.327
R1012 VSS.t829 VSS.t833 516.327
R1013 VSS.t1082 VSS.t622 516.327
R1014 VSS.t1304 VSS.t401 516.327
R1015 VSS.t1150 VSS.t367 516.327
R1016 VSS.t1895 VSS.t1911 516.327
R1017 VSS.t592 VSS.t1862 516.327
R1018 VSS.t38 VSS.t34 516.327
R1019 VSS.t438 VSS.t1248 516.327
R1020 VSS.t253 VSS.t119 516.327
R1021 VSS.t160 VSS.t153 516.327
R1022 VSS.t861 VSS.t863 516.327
R1023 VSS.t2025 VSS.t1113 516.327
R1024 VSS.t1837 VSS.t1850 516.327
R1025 VSS.t298 VSS.t476 516.327
R1026 VSS.t1786 VSS.t1782 516.327
R1027 VSS.t136 VSS.t379 516.327
R1028 VSS.t816 VSS.t1121 516.327
R1029 VSS.t267 VSS.t705 516.327
R1030 VSS.t1350 VSS.t1354 516.327
R1031 VSS.t732 VSS.t1771 516.327
R1032 VSS.t175 VSS.t193 516.327
R1033 VSS.t1429 VSS.t1064 516.327
R1034 VSS.t553 VSS.t567 516.327
R1035 VSS.t412 VSS.t717 516.327
R1036 VSS.t1402 VSS.t1388 516.327
R1037 VSS.t610 VSS.t1492 516.327
R1038 VSS.t958 VSS.t85 516.327
R1039 VSS.t798 VSS.t1603 516.327
R1040 VSS.t1571 VSS.t1159 516.327
R1041 VSS.t1754 VSS.t1669 516.327
R1042 VSS.t1005 VSS.t990 516.327
R1043 VSS.t147 VSS.t1069 516.327
R1044 VSS.t697 VSS.t635 516.327
R1045 VSS.t319 VSS.t133 516.327
R1046 VSS.t94 VSS.t96 516.327
R1047 VSS.t1088 VSS.t1879 516.327
R1048 VSS.t1169 VSS.t1165 516.327
R1049 VSS.t655 VSS.t752 516.327
R1050 VSS.t343 VSS.t349 516.327
R1051 VSS.t462 VSS.t212 516.327
R1052 VSS.t116 VSS.t109 516.327
R1053 VSS.t1446 VSS.t1204 516.327
R1054 VSS.t1281 VSS.t1279 516.327
R1055 VSS.t1408 VSS.t235 516.327
R1056 VSS.t312 VSS.t314 516.327
R1057 VSS.t1015 VSS.t1060 516.327
R1058 VSS.t1008 VSS.t999 516.327
R1059 VSS.t946 VSS.t292 516.327
R1060 VSS.t1482 VSS.t1478 516.327
R1061 VSS.t532 VSS.t1261 516.327
R1062 VSS.t1928 VSS.t1930 516.327
R1063 VSS.t1235 VSS.t1763 516.327
R1064 VSS.t50 VSS.t46 516.327
R1065 VSS.t1660 VSS.t1501 516.327
R1066 VSS.t1685 VSS.t1679 516.327
R1067 VSS.t27 VSS.t325 516.327
R1068 VSS.t8 VSS.t11 516.327
R1069 VSS.t1511 VSS.t1816 516.327
R1070 VSS.t1867 VSS.t1869 516.327
R1071 VSS.t663 VSS.t521 516.327
R1072 VSS.t1915 VSS.t1944 516.327
R1073 VSS.t1423 VSS.t1334 516.327
R1074 VSS.t1012 VSS.t1022 516.327
R1075 VSS.t447 VSS.t1560 516.327
R1076 VSS.t1616 VSS.t1622 516.327
R1077 VSS.t1037 VSS.t965 516.327
R1078 VSS.t1371 VSS.t1052 516.327
R1079 VSS.t1940 VSS.t1043 516.327
R1080 VSS.t1812 VSS.t1814 516.327
R1081 VSS.t825 VSS.t969 516.327
R1082 VSS.t423 VSS.t421 516.327
R1083 VSS.t632 VSS.t405 516.327
R1084 VSS.t1242 VSS.t1244 516.327
R1085 VSS.t1315 VSS.t73 516.327
R1086 VSS.t472 VSS.t468 516.327
R1087 VSS.t1674 VSS.t1341 516.327
R1088 VSS.t1526 VSS.t1528 516.327
R1089 VSS.t391 VSS.t1828 516.327
R1090 VSS.n1671 VSS.t2054 491.64
R1091 VSS.n1672 VSS.t2056 491.64
R1092 VSS.n1673 VSS.t2068 491.64
R1093 VSS.n1674 VSS.t2055 491.64
R1094 VSS.n298 VSS.t2033 491.64
R1095 VSS.n298 VSS.t2043 491.64
R1096 VSS.n298 VSS.t2037 491.64
R1097 VSS.n298 VSS.t2062 491.64
R1098 VSS.n428 VSS.t2039 491.64
R1099 VSS.n428 VSS.t2050 491.64
R1100 VSS.n428 VSS.t2044 491.64
R1101 VSS.n428 VSS.t2066 491.64
R1102 VSS.n466 VSS.t2051 491.64
R1103 VSS.n466 VSS.t2045 491.64
R1104 VSS.n466 VSS.t2047 491.64
R1105 VSS.n466 VSS.t2057 491.64
R1106 VSS.t1980 VSS.n644 487.774
R1107 VSS.n645 VSS.t1710 487.774
R1108 VSS.n1667 VSS.t976 485.221
R1109 VSS.t1698 VSS.t1696 483.849
R1110 VSS.t1696 VSS.t1694 483.849
R1111 VSS.t1694 VSS.t1210 483.849
R1112 VSS.t1210 VSS.t1209 483.849
R1113 VSS.t1209 VSS.t393 483.849
R1114 VSS.t586 VSS.t696 483.849
R1115 VSS.t696 VSS.t690 483.849
R1116 VSS.t690 VSS.t389 483.849
R1117 VSS.t389 VSS.t915 483.849
R1118 VSS.t915 VSS.t881 483.849
R1119 VSS.t1922 VSS.t1924 483.849
R1120 VSS.t1926 VSS.t1922 483.849
R1121 VSS.t1326 VSS.t1926 483.849
R1122 VSS.t1325 VSS.t1326 483.849
R1123 VSS.t1327 VSS.t1325 483.849
R1124 VSS.t1634 VSS.t1632 483.849
R1125 VSS.t1632 VSS.t1630 483.849
R1126 VSS.t1630 VSS.t385 483.849
R1127 VSS.t385 VSS.t909 483.849
R1128 VSS.t909 VSS.t876 483.849
R1129 VSS.t1516 VSS.t565 483.849
R1130 VSS.t565 VSS.t563 483.849
R1131 VSS.t563 VSS.t1410 483.849
R1132 VSS.t1410 VSS.t1434 483.849
R1133 VSS.t1434 VSS.t1411 483.849
R1134 VSS.t444 VSS.t1796 483.849
R1135 VSS.t1796 VSS.t1803 483.849
R1136 VSS.t1803 VSS.t913 483.849
R1137 VSS.t913 VSS.t900 483.849
R1138 VSS.t900 VSS.t883 483.849
R1139 VSS.t758 VSS.t276 483.849
R1140 VSS.t276 VSS.t793 483.849
R1141 VSS.t793 VSS.t1344 483.849
R1142 VSS.t1344 VSS.t1345 483.849
R1143 VSS.t1345 VSS.t1343 483.849
R1144 VSS.t1649 VSS.t1643 483.849
R1145 VSS.t1643 VSS.t1654 483.849
R1146 VSS.t1654 VSS.t891 483.849
R1147 VSS.t891 VSS.t898 483.849
R1148 VSS.t898 VSS.t371 483.849
R1149 VSS.t1555 VSS.t1553 483.849
R1150 VSS.t1553 VSS.t713 483.849
R1151 VSS.t713 VSS.t332 483.849
R1152 VSS.t332 VSS.t334 483.849
R1153 VSS.t334 VSS.t333 483.849
R1154 VSS.t1107 VSS.t1100 483.849
R1155 VSS.t1100 VSS.t1112 483.849
R1156 VSS.t1112 VSS.t887 483.849
R1157 VSS.t887 VSS.t924 483.849
R1158 VSS.t924 VSS.t907 483.849
R1159 VSS.t1794 VSS.t1792 483.849
R1160 VSS.t1792 VSS.t1790 483.849
R1161 VSS.t1790 VSS.t1806 483.849
R1162 VSS.t1806 VSS.t1805 483.849
R1163 VSS.t1805 VSS.t1807 483.849
R1164 VSS.t225 VSS.t219 483.849
R1165 VSS.t219 VSS.t1286 483.849
R1166 VSS.t1286 VSS.t868 483.849
R1167 VSS.t868 VSS.t904 483.849
R1168 VSS.t904 VSS.t889 483.849
R1169 VSS.t1889 VSS.t1891 483.849
R1170 VSS.t1885 VSS.t1889 483.849
R1171 VSS.t604 VSS.t1885 483.849
R1172 VSS.t603 VSS.t604 483.849
R1173 VSS.t605 VSS.t603 483.849
R1174 VSS.t1180 VSS.t1177 483.849
R1175 VSS.t1177 VSS.t1191 483.849
R1176 VSS.t1191 VSS.t373 483.849
R1177 VSS.t373 VSS.t902 483.849
R1178 VSS.t902 VSS.t885 483.849
R1179 VSS.t455 VSS.t457 483.849
R1180 VSS.t459 VSS.t455 483.849
R1181 VSS.t821 VSS.t459 483.849
R1182 VSS.t820 VSS.t821 483.849
R1183 VSS.t1412 VSS.t820 483.849
R1184 VSS.t508 VSS.t501 483.849
R1185 VSS.t501 VSS.t284 483.849
R1186 VSS.t284 VSS.t930 483.849
R1187 VSS.t930 VSS.t896 483.849
R1188 VSS.t896 VSS.t874 483.849
R1189 VSS.t1978 VSS.n665 475.705
R1190 VSS.n666 VSS.t1734 475.705
R1191 VSS.n685 VSS.t1957 475.705
R1192 VSS.n684 VSS.t1708 475.705
R1193 VSS.t1984 VSS.n658 475.705
R1194 VSS.n659 VSS.t1749 475.705
R1195 VSS.n693 VSS.t1954 475.705
R1196 VSS.n692 VSS.t1706 475.705
R1197 VSS.t1976 VSS.n651 475.705
R1198 VSS.n652 VSS.t1732 475.705
R1199 VSS.n709 VSS.t1961 475.705
R1200 VSS.n708 VSS.t1701 475.705
R1201 VSS.n701 VSS.t1982 464.221
R1202 VSS.n700 VSS.t1714 464.221
R1203 VSS.n1401 VSS.n209 463.753
R1204 VSS.t583 VSS.t1698 463.688
R1205 VSS.t881 VSS.t894 463.688
R1206 VSS.t1924 VSS.t1639 463.688
R1207 VSS.t876 VSS.t375 463.688
R1208 VSS.t1797 VSS.t1516 463.688
R1209 VSS.t883 VSS.t922 463.688
R1210 VSS.t1647 VSS.t758 463.688
R1211 VSS.t371 VSS.t917 463.688
R1212 VSS.t1105 VSS.t1555 463.688
R1213 VSS.t907 VSS.t870 463.688
R1214 VSS.t221 VSS.t1794 463.688
R1215 VSS.t889 VSS.t928 463.688
R1216 VSS.t1891 VSS.t1189 463.688
R1217 VSS.t885 VSS.t926 463.688
R1218 VSS.t457 VSS.t513 463.688
R1219 VSS.t874 VSS.t919 463.688
R1220 VSS.n89 VSS.t1645 442.212
R1221 VSS.n1396 VSS.t441 440
R1222 VSS.t1103 VSS.t1839 437.721
R1223 VSS.t1534 VSS.n1401 427.397
R1224 VSS.t1590 VSS.t488 424.45
R1225 VSS.n1653 VSS.n87 420.933
R1226 VSS.n677 VSS.t1974 415.024
R1227 VSS.n676 VSS.t1728 415.024
R1228 VSS.n1191 VSS.n621 400.342
R1229 VSS.n1188 VSS.n623 400.342
R1230 VSS.n1185 VSS.n625 400.342
R1231 VSS.n1194 VSS.n619 400.342
R1232 VSS.n1197 VSS.n617 400.342
R1233 VSS.n1200 VSS.n615 400.342
R1234 VSS.n1203 VSS.n613 400.342
R1235 VSS.n1206 VSS.n611 400.342
R1236 VSS.n1209 VSS.n609 400.342
R1237 VSS.n487 VSS.t1134 395.522
R1238 VSS.n1496 VSS.n1495 390
R1239 VSS.n1499 VSS.n1498 390
R1240 VSS.n252 VSS.n154 390
R1241 VSS.n250 VSS.n154 390
R1242 VSS.n254 VSS.n154 390
R1243 VSS.n178 VSS.n153 390
R1244 VSS.n180 VSS.n153 390
R1245 VSS.n182 VSS.n153 390
R1246 VSS.n839 VSS.n838 390
R1247 VSS.n814 VSS.n813 390
R1248 VSS.n824 VSS.n823 390
R1249 VSS.n872 VSS.n871 390
R1250 VSS.n764 VSS.n763 390
R1251 VSS.n790 VSS.n789 390
R1252 VSS.n773 VSS.n772 390
R1253 VSS.n782 VSS.n781 390
R1254 VSS.n804 VSS.n803 390
R1255 VSS.n1501 VSS.n151 389.536
R1256 VSS.n1535 VSS.t211 387.267
R1257 VSS.n1633 VSS.n1632 379.269
R1258 VSS.n1404 VSS.t1097 378.113
R1259 VSS.n1502 VSS.n1501 370.646
R1260 VSS.n1665 VSS.t2058 367.928
R1261 VSS.n302 VSS.t2069 367.928
R1262 VSS.n432 VSS.t2041 367.928
R1263 VSS.n470 VSS.t2060 367.928
R1264 VSS.t280 VSS.t1848 357.361
R1265 VSS.t1645 VSS.t805 353.769
R1266 VSS.n869 VSS.n868 353.735
R1267 VSS.t441 VSS.t191 352
R1268 VSS.n1131 VSS.t2064 336.962
R1269 VSS.n1136 VSS.t2052 336.962
R1270 VSS.n1139 VSS.t2067 336.962
R1271 VSS.n1128 VSS.t2042 336.962
R1272 VSS.n1126 VSS.t2049 336.962
R1273 VSS.t234 VSS.n626 336.438
R1274 VSS.t243 VSS.n1019 336.295
R1275 VSS.t727 VSS.n983 336.295
R1276 VSS.t577 VSS.n949 336.295
R1277 VSS.t1377 VSS.n1053 336.295
R1278 VSS.t461 VSS.n915 336.295
R1279 VSS.t454 VSS.n735 336.295
R1280 VSS.t785 VSS.n881 336.295
R1281 VSS.n867 VSS.t626 336.295
R1282 VSS.n1448 VSS.n1447 335.543
R1283 VSS.n212 VSS.t329 334.584
R1284 VSS.n1492 VSS.t172 334.584
R1285 VSS.n555 VSS.t223 334.584
R1286 VSS.t118 VSS.n448 330.106
R1287 VSS.n1131 VSS.t2036 326.154
R1288 VSS.n1136 VSS.t2065 326.154
R1289 VSS.n1139 VSS.t2040 326.154
R1290 VSS.n1128 VSS.t2063 326.154
R1291 VSS.n1126 VSS.t2070 326.154
R1292 VSS.t1859 VSS.n122 325.317
R1293 VSS.n862 VSS.t1219 320.356
R1294 VSS.t1522 VSS.t1520 305.644
R1295 VSS.t1518 VSS.t1522 305.644
R1296 VSS.t1592 VSS.t1518 305.644
R1297 VSS.t1162 VSS.t1592 305.644
R1298 VSS.t1584 VSS.t1162 305.644
R1299 VSS.t974 VSS.t1085 305.644
R1300 VSS.n1654 VSS.n86 298.127
R1301 VSS.n1654 VSS.n1653 294.896
R1302 VSS.t1520 VSS.t1524 292.909
R1303 VSS.n851 VSS.n850 288.707
R1304 VSS.t1452 VSS.n1259 280.613
R1305 VSS.t1274 VSS.n1268 280.613
R1306 VSS.n1278 VSS.t767 280.613
R1307 VSS.n1277 VSS.t399 280.613
R1308 VSS.n1525 VSS.t1557 280.613
R1309 VSS.n1524 VSS.t102 280.613
R1310 VSS.t2023 VSS.n281 280.613
R1311 VSS.t775 VSS.n502 280.613
R1312 VSS.t1075 VSS.n511 280.613
R1313 VSS.n512 VSS.t1548 280.613
R1314 VSS.n1467 VSS.t64 280.613
R1315 VSS.n1466 VSS.t1767 280.613
R1316 VSS.t227 VSS.n1355 280.613
R1317 VSS.n1377 VSS.t597 280.613
R1318 VSS.n1376 VSS.t1256 280.613
R1319 VSS.n1367 VSS.t1598 280.613
R1320 VSS.n316 VSS.t763 280.613
R1321 VSS.n296 VSS.t498 280.613
R1322 VSS.n1719 VSS.t497 280.613
R1323 VSS.n1718 VSS.t1874 280.613
R1324 VSS.n1699 VSS.t1154 280.613
R1325 VSS.n1698 VSS.t1222 280.613
R1326 VSS.n1679 VSS.t337 280.613
R1327 VSS.n1678 VSS.t361 280.613
R1328 VSS.n446 VSS.t518 280.613
R1329 VSS.n426 VSS.t845 280.613
R1330 VSS.n417 VSS.t950 280.613
R1331 VSS.n412 VSS.t1688 280.613
R1332 VSS.n407 VSS.t709 280.613
R1333 VSS.n402 VSS.t356 280.613
R1334 VSS.n397 VSS.t126 280.613
R1335 VSS.n392 VSS.t1418 280.613
R1336 VSS.n484 VSS.t1055 280.613
R1337 VSS.n464 VSS.t762 280.613
R1338 VSS.n455 VSS.t616 280.613
R1339 VSS.n1709 VSS.t1048 280.613
R1340 VSS.n1708 VSS.t797 280.613
R1341 VSS.n1689 VSS.t646 280.613
R1342 VSS.n1688 VSS.t769 280.613
R1343 VSS.n1656 VSS.t1609 280.613
R1344 VSS.n190 VSS.n189 275.466
R1345 VSS.n1331 VSS.n575 263.452
R1346 VSS.n1298 VSS.t364 262.168
R1347 VSS.n1391 VSS.t686 259.205
R1348 VSS.n1647 VSS.n87 258.538
R1349 VSS.n1259 VSS.t1140 258.163
R1350 VSS.n1268 VSS.t1079 258.163
R1351 VSS.n1278 VSS.t366 258.163
R1352 VSS.t1861 VSS.n1277 258.163
R1353 VSS.n1525 VSS.t1251 258.163
R1354 VSS.t432 VSS.n1524 258.163
R1355 VSS.n281 VSS.t2030 258.163
R1356 VSS.n502 VSS.t303 258.163
R1357 VSS.n511 VSS.t165 258.163
R1358 VSS.n512 VSS.t704 258.163
R1359 VSS.n1467 VSS.t1770 258.163
R1360 VSS.t1428 VSS.n1466 258.163
R1361 VSS.n1355 VSS.t1206 258.163
R1362 VSS.n1377 VSS.t1491 258.163
R1363 VSS.t1601 VSS.n1376 258.163
R1364 VSS.t1671 VSS.n1367 258.163
R1365 VSS.t1072 VSS.n316 258.163
R1366 VSS.t135 VSS.n296 258.163
R1367 VSS.n1719 VSS.t1882 258.163
R1368 VSS.t654 VSS.n1718 258.163
R1369 VSS.n1699 VSS.t214 258.163
R1370 VSS.t1445 VSS.n1698 258.163
R1371 VSS.n1679 VSS.t240 258.163
R1372 VSS.t997 VSS.n1678 258.163
R1373 VSS.t295 VSS.n446 258.163
R1374 VSS.t1265 VSS.n426 258.163
R1375 VSS.t1766 VSS.n417 258.163
R1376 VSS.t1500 VSS.n412 258.163
R1377 VSS.t327 VSS.n407 258.163
R1378 VSS.t1821 VSS.n402 258.163
R1379 VSS.t524 VSS.n397 258.163
R1380 VSS.t1338 VSS.n392 258.163
R1381 VSS.t1559 VSS.n484 258.163
R1382 VSS.t528 VSS.n464 258.163
R1383 VSS.t1042 VSS.n455 258.163
R1384 VSS.n1709 VSS.t956 258.163
R1385 VSS.t629 VSS.n1708 258.163
R1386 VSS.n1689 VSS.t72 258.163
R1387 VSS.t1676 VSS.n1688 258.163
R1388 VSS.n1656 VSS.t1825 258.163
R1389 VSS.n1640 VSS.t393 257.046
R1390 VSS.n1341 VSS.t1327 257.046
R1391 VSS.t1411 VSS.n262 257.046
R1392 VSS.t1343 VSS.n531 257.046
R1393 VSS.t333 VSS.n540 257.046
R1394 VSS.t1807 VSS.n572 257.046
R1395 VSS.n1291 VSS.t605 257.046
R1396 VSS.n1317 VSS.t1412 257.046
R1397 VSS.n1675 VSS.t1014 255.588
R1398 VSS.n1225 VSS.n1224 252.06
R1399 VSS.t672 VSS.t168 241.638
R1400 VSS.n1205 VSS.t2020 236.631
R1401 VSS.n450 VSS.n449 236.256
R1402 VSS.n1406 VSS.n86 235.869
R1403 VSS.n204 VSS.n201 235.869
R1404 VSS.n381 VSS.n200 235.869
R1405 VSS.n323 VSS.n199 235.869
R1406 VSS.n358 VSS.n357 235.869
R1407 VSS.n1455 VSS.n1454 235.869
R1408 VSS.n189 VSS.n188 235.869
R1409 VSS.n350 VSS.n349 235.869
R1410 VSS.n1437 VSS.n196 235.869
R1411 VSS.n1450 VSS.n1449 235.869
R1412 VSS.n1447 VSS.n1446 235.869
R1413 VSS.n1434 VSS.n1433 235.869
R1414 VSS.n318 VSS.n317 235.869
R1415 VSS.n376 VSS.n375 235.869
R1416 VSS.n1419 VSS.n1418 235.869
R1417 VSS.n1410 VSS.n1409 235.869
R1418 VSS VSS.n844 235.867
R1419 VSS.n1513 VSS.n142 235.861
R1420 VSS.n1514 VSS.n1513 235.861
R1421 VSS.n448 VSS.n447 235.861
R1422 VSS.n1534 VSS.n1533 235.861
R1423 VSS.n1536 VSS.n1535 235.861
R1424 VSS.n1297 VSS.n1296 235.861
R1425 VSS.n1299 VSS.n1298 235.861
R1426 VSS.n1309 VSS.n1308 235.861
R1427 VSS.n1323 VSS.n1322 235.861
R1428 VSS.n1325 VSS.n1324 235.861
R1429 VSS.n1392 VSS.n1391 235.861
R1430 VSS.n1391 VSS.n1390 235.861
R1431 VSS.n1396 VSS.n1395 235.861
R1432 VSS.n90 VSS.n89 235.861
R1433 VSS.n1652 VSS.n1651 235.861
R1434 VSS.n1403 VSS.n1402 235.861
R1435 VSS.n342 VSS.n209 235.861
R1436 VSS.n208 VSS.n207 235.861
R1437 VSS.n94 VSS.n93 235.861
R1438 VSS.n1646 VSS.n1645 235.861
R1439 VSS.n1648 VSS.n1647 235.861
R1440 VSS.n374 VSS.n373 235.861
R1441 VSS.n372 VSS.n371 235.861
R1442 VSS.n341 VSS.n340 235.861
R1443 VSS.n339 VSS.n338 235.861
R1444 VSS.n337 VSS.n167 235.861
R1445 VSS.n336 VSS.n162 235.861
R1446 VSS.n335 VSS.n334 235.861
R1447 VSS.n333 VSS.n147 235.861
R1448 VSS.n332 VSS.n331 235.861
R1449 VSS.n330 VSS.n145 235.861
R1450 VSS.n329 VSS.n140 235.861
R1451 VSS.n328 VSS.n136 235.861
R1452 VSS.n367 VSS.n366 235.861
R1453 VSS.n369 VSS.n368 235.861
R1454 VSS.n346 VSS.n345 235.861
R1455 VSS.n344 VSS.n343 235.861
R1456 VSS.n1477 VSS.n1476 235.861
R1457 VSS.n1479 VSS.n1478 235.861
R1458 VSS.n165 VSS.n164 235.861
R1459 VSS.n1506 VSS.n1505 235.861
R1460 VSS.n1508 VSS.n1507 235.861
R1461 VSS.n1510 VSS.n1509 235.861
R1462 VSS.n1517 VSS.n1516 235.861
R1463 VSS.n1519 VSS.n1518 235.861
R1464 VSS.n1362 VSS.n103 235.861
R1465 VSS.n1388 VSS.n1387 235.861
R1466 VSS.n1386 VSS.n1385 235.861
R1467 VSS.n1348 VSS.n1347 235.861
R1468 VSS.n1350 VSS.n1349 235.861
R1469 VSS.n1346 VSS.n1345 235.861
R1470 VSS.n1461 VSS.n1460 235.861
R1471 VSS.n267 VSS.n266 235.861
R1472 VSS.n269 VSS.n268 235.861
R1473 VSS.n521 VSS.n520 235.861
R1474 VSS.n523 VSS.n522 235.861
R1475 VSS.n495 VSS.n494 235.861
R1476 VSS.n497 VSS.n496 235.861
R1477 VSS.n493 VSS.n492 235.861
R1478 VSS.n490 VSS.n489 235.861
R1479 VSS.n151 VSS.n149 235.861
R1480 VSS.n1474 VSS.n151 235.861
R1481 VSS.n163 VSS.n151 235.861
R1482 VSS.n151 VSS.n150 235.861
R1483 VSS.n1503 VSS.n1502 235.861
R1484 VSS.n608 VSS.n607 235.861
R1485 VSS.n485 VSS.n138 235.861
R1486 VSS.n1513 VSS.n1512 235.861
R1487 VSS.t810 VSS.n153 234.464
R1488 VSS.n154 VSS.t177 234.34
R1489 VSS.n1187 VSS.t1995 230.778
R1490 VSS.n1190 VSS.t2010 230.778
R1491 VSS.n1193 VSS.t2004 230.778
R1492 VSS.n1196 VSS.t2012 230.778
R1493 VSS.n1199 VSS.t1992 230.778
R1494 VSS.n1208 VSS.t2016 230.778
R1495 VSS.n1041 VSS.t1458 229.304
R1496 VSS.t1462 VSS.n1039 229.304
R1497 VSS.t1460 VSS.n1035 229.304
R1498 VSS.t1456 VSS.n621 229.304
R1499 VSS.n1005 VSS.t740 229.304
R1500 VSS.t744 VSS.n1003 229.304
R1501 VSS.t742 VSS.n999 229.304
R1502 VSS.t738 VSS.n623 229.304
R1503 VSS.t197 VSS.n1180 229.304
R1504 VSS.n1159 VSS.t200 229.304
R1505 VSS.n1163 VSS.t204 229.304
R1506 VSS.n1165 VSS.t202 229.304
R1507 VSS.t206 VSS.n625 229.304
R1508 VSS.n971 VSS.t679 229.304
R1509 VSS.t675 VSS.n969 229.304
R1510 VSS.t681 VSS.n965 229.304
R1511 VSS.t677 VSS.n619 229.304
R1512 VSS.n1075 VSS.t58 229.304
R1513 VSS.t54 VSS.n1073 229.304
R1514 VSS.t60 VSS.n1069 229.304
R1515 VSS.t56 VSS.n617 229.304
R1516 VSS.n937 VSS.t1378 229.304
R1517 VSS.t1382 VSS.n935 229.304
R1518 VSS.t1380 VSS.n931 229.304
R1519 VSS.t1384 VSS.n615 229.304
R1520 VSS.n1092 VSS.t1474 229.304
R1521 VSS.n1096 VSS.t1470 229.304
R1522 VSS.n1098 VSS.t1472 229.304
R1523 VSS.t1476 VSS.n613 229.304
R1524 VSS.n903 VSS.t853 229.304
R1525 VSS.t849 VSS.n901 229.304
R1526 VSS.t851 VSS.n897 229.304
R1527 VSS.t855 VSS.n611 229.304
R1528 VSS.n1116 VSS.t1437 229.304
R1529 VSS.n1120 VSS.t1439 229.304
R1530 VSS.n1122 VSS.t1435 229.304
R1531 VSS.t1441 VSS.n609 229.304
R1532 VSS.n1023 VSS.t17 229.207
R1533 VSS.n987 VSS.t77 229.207
R1534 VSS.n953 VSS.t104 229.207
R1535 VSS.n1057 VSS.t397 229.207
R1536 VSS.n919 VSS.t722 229.207
R1537 VSS.n737 VSS.t667 229.207
R1538 VSS.n885 VSS.t651 229.207
R1539 VSS.t618 VSS.n866 229.207
R1540 VSS.n1323 VSS.t840 228.032
R1541 VSS.n303 VSS.t2035 227.356
R1542 VSS.n433 VSS.t2048 227.356
R1543 VSS.n471 VSS.t2053 227.356
R1544 VSS.n1640 VSS.t586 226.804
R1545 VSS.n1341 VSS.t1634 226.804
R1546 VSS.n262 VSS.t444 226.804
R1547 VSS.n531 VSS.t1649 226.804
R1548 VSS.n540 VSS.t1107 226.804
R1549 VSS.n572 VSS.t225 226.804
R1550 VSS.n1291 VSS.t1180 226.804
R1551 VSS.n1317 VSS.t508 226.804
R1552 VSS.n1202 VSS.t2018 225.206
R1553 VSS.n1666 VSS.t2038 224.478
R1554 VSS.n1224 VSS.n590 221.006
R1555 VSS.n1565 VSS.n122 219.048
R1556 VSS.t939 VSS.n1226 216.869
R1557 VSS.n1224 VSS.n584 215.537
R1558 VSS.n1224 VSS.n585 215.537
R1559 VSS.n1224 VSS.n586 215.537
R1560 VSS.n1224 VSS.n587 215.537
R1561 VSS.n1224 VSS.n588 215.537
R1562 VSS.n1224 VSS.n591 215.537
R1563 VSS.n1665 VSS.t2061 213.688
R1564 VSS.n302 VSS.t2034 213.688
R1565 VSS.n432 VSS.t2046 213.688
R1566 VSS.n470 VSS.t2059 213.688
R1567 VSS.n869 VSS.n862 212.206
R1568 VSS.n1224 VSS.n589 210.333
R1569 VSS.n1671 VSS.n1670 209.19
R1570 VSS.n365 VSS.n364 207.804
R1571 VSS.t686 VSS.t1158 207.364
R1572 VSS.n1534 VSS.n124 204.708
R1573 VSS.n1184 VSS.t1986 201.339
R1574 VSS.n1448 VSS.n104 195.733
R1575 VSS.t511 VSS.t252 191.739
R1576 VSS.n1460 VSS.n1459 191.393
R1577 VSS.n1210 VSS.n606 190.877
R1578 VSS.n1224 VSS.n583 188.042
R1579 VSS.n1501 VSS.n1500 186.94
R1580 VSS.n1324 VSS.t880 181.102
R1581 VSS.t1994 VSS.t19 180.436
R1582 VSS.t89 VSS.t1994 180.436
R1583 VSS.t1458 VSS.t89 180.436
R1584 VSS.t296 VSS.t92 180.436
R1585 VSS.t92 VSS.t88 180.436
R1586 VSS.t88 VSS.t1462 180.436
R1587 VSS.t1050 VSS.t1989 180.436
R1588 VSS.t1989 VSS.t1951 180.436
R1589 VSS.t1951 VSS.t1460 180.436
R1590 VSS.t242 VSS.t93 180.436
R1591 VSS.t93 VSS.t1963 180.436
R1592 VSS.t1963 VSS.t1456 180.436
R1593 VSS.t1988 VSS.t1157 180.436
R1594 VSS.t1319 VSS.t1988 180.436
R1595 VSS.t740 VSS.t1319 180.436
R1596 VSS.t736 VSS.t1467 180.436
R1597 VSS.t1467 VSS.t1320 180.436
R1598 VSS.t1320 VSS.t744 180.436
R1599 VSS.t527 VSS.t1991 180.436
R1600 VSS.t1991 VSS.t1956 180.436
R1601 VSS.t1956 VSS.t742 180.436
R1602 VSS.t613 VSS.t1466 180.436
R1603 VSS.t1466 VSS.t1971 180.436
R1604 VSS.t1971 VSS.t738 180.436
R1605 VSS.t123 VSS.t234 180.436
R1606 VSS.t721 VSS.t123 180.436
R1607 VSS.t1990 VSS.t199 180.436
R1608 VSS.t151 VSS.t1990 180.436
R1609 VSS.t200 VSS.t151 180.436
R1610 VSS.t2 VSS.t1499 180.436
R1611 VSS.t152 VSS.t2 180.436
R1612 VSS.t204 VSS.t152 180.436
R1613 VSS.t2009 VSS.t127 180.436
R1614 VSS.t1972 VSS.t2009 180.436
R1615 VSS.t202 VSS.t1972 180.436
R1616 VSS.t167 VSS.t1 180.436
R1617 VSS.t1 VSS.t1964 180.436
R1618 VSS.t1964 VSS.t206 180.436
R1619 VSS.t2000 VSS.t674 180.436
R1620 VSS.t1665 VSS.t2000 180.436
R1621 VSS.t679 VSS.t1665 180.436
R1622 VSS.t1541 VSS.t1033 180.436
R1623 VSS.t1033 VSS.t1664 180.436
R1624 VSS.t1664 VSS.t675 180.436
R1625 VSS.t87 VSS.t2003 180.436
R1626 VSS.t2003 VSS.t1967 180.436
R1627 VSS.t1967 VSS.t681 180.436
R1628 VSS.t328 VSS.t857 180.436
R1629 VSS.t857 VSS.t1950 180.436
R1630 VSS.t1950 VSS.t677 180.436
R1631 VSS.t2001 VSS.t3 180.436
R1632 VSS.t1497 VSS.t2001 180.436
R1633 VSS.t58 VSS.t1497 180.436
R1634 VSS.t16 VSS.t1545 180.436
R1635 VSS.t1545 VSS.t1496 180.436
R1636 VSS.t1496 VSS.t54 180.436
R1637 VSS.t196 VSS.t2002 180.436
R1638 VSS.t2002 VSS.t1969 180.436
R1639 VSS.t1969 VSS.t60 180.436
R1640 VSS.t957 VSS.t1544 180.436
R1641 VSS.t1544 VSS.t1953 180.436
R1642 VSS.t1953 VSS.t56 180.436
R1643 VSS.t2015 VSS.t822 180.436
R1644 VSS.t1321 VSS.t2015 180.436
R1645 VSS.t1378 VSS.t1321 180.436
R1646 VSS.t0 VSS.t1268 180.436
R1647 VSS.t1268 VSS.t1322 180.436
R1648 VSS.t1322 VSS.t1382 180.436
R1649 VSS.t562 VSS.t1999 180.436
R1650 VSS.t1999 VSS.t1965 180.436
R1651 VSS.t1965 VSS.t1380 180.436
R1652 VSS.t208 VSS.t1269 180.436
R1653 VSS.t1269 VSS.t1973 180.436
R1654 VSS.t1973 VSS.t1384 180.436
R1655 VSS.t1051 VSS.t1998 180.436
R1656 VSS.t1998 VSS.t1487 180.436
R1657 VSS.t1487 VSS.t1474 180.436
R1658 VSS.t1488 VSS.t31 180.436
R1659 VSS.t1486 VSS.t1488 180.436
R1660 VSS.t1470 VSS.t1486 180.436
R1661 VSS.t2008 VSS.t304 180.436
R1662 VSS.t1966 VSS.t2008 180.436
R1663 VSS.t1472 VSS.t1966 180.436
R1664 VSS.t396 VSS.t1489 180.436
R1665 VSS.t1489 VSS.t1959 180.436
R1666 VSS.t1959 VSS.t1476 180.436
R1667 VSS.t1997 VSS.t43 180.436
R1668 VSS.t32 VSS.t1997 180.436
R1669 VSS.t853 VSS.t32 180.436
R1670 VSS.t1543 VSS.t627 180.436
R1671 VSS.t627 VSS.t33 180.436
R1672 VSS.t33 VSS.t849 180.436
R1673 VSS.t433 VSS.t2006 180.436
R1674 VSS.t2006 VSS.t1960 180.436
R1675 VSS.t1960 VSS.t851 180.436
R1676 VSS.t275 VSS.t628 180.436
R1677 VSS.t628 VSS.t1952 180.436
R1678 VSS.t1952 VSS.t855 180.436
R1679 VSS.t1002 VSS.t2014 180.436
R1680 VSS.t2014 VSS.t316 180.436
R1681 VSS.t316 VSS.t1437 180.436
R1682 VSS.t425 VSS.t776 180.436
R1683 VSS.t317 VSS.t425 180.436
R1684 VSS.t1439 VSS.t317 180.436
R1685 VSS.t2007 VSS.t983 180.436
R1686 VSS.t1968 VSS.t2007 180.436
R1687 VSS.t1435 VSS.t1968 180.436
R1688 VSS.t841 VSS.t426 180.436
R1689 VSS.t426 VSS.t1970 180.436
R1690 VSS.t1970 VSS.t1441 180.436
R1691 VSS.t1084 VSS.t243 180.359
R1692 VSS.t1272 VSS.t1084 180.359
R1693 VSS.t17 VSS.t1272 180.359
R1694 VSS.t166 VSS.t727 180.359
R1695 VSS.t712 VSS.t166 180.359
R1696 VSS.t77 VSS.t712 180.359
R1697 VSS.t701 VSS.t577 180.359
R1698 VSS.t1329 VSS.t701 180.359
R1699 VSS.t104 VSS.t1329 180.359
R1700 VSS.t103 VSS.t1377 180.359
R1701 VSS.t967 VSS.t103 180.359
R1702 VSS.t397 VSS.t967 180.359
R1703 VSS.t612 VSS.t461 180.359
R1704 VSS.t596 VSS.t612 180.359
R1705 VSS.t722 VSS.t596 180.359
R1706 VSS.t764 VSS.t454 180.359
R1707 VSS.t318 VSS.t764 180.359
R1708 VSS.t667 VSS.t318 180.359
R1709 VSS.t311 VSS.t785 180.359
R1710 VSS.t464 VSS.t311 180.359
R1711 VSS.t651 VSS.t464 180.359
R1712 VSS.t626 VSS.t867 180.359
R1713 VSS.t867 VSS.t174 180.359
R1714 VSS.t174 VSS.t618 180.359
R1715 VSS.n1677 VSS.n1676 179.369
R1716 VSS.n486 VSS.n143 179.054
R1717 VSS.n190 VSS.t280 171.236
R1718 VSS.n1226 VSS.n1225 170.826
R1719 VSS.t483 VSS.n152 167.243
R1720 VSS.n562 VSS.n124 165.24
R1721 VSS.n1132 VSS.n1131 162.952
R1722 VSS.n1137 VSS.n1136 162.952
R1723 VSS.n1129 VSS.n1128 162.952
R1724 VSS.n1127 VSS.n1126 162.946
R1725 VSS.n1140 VSS.n1139 162.945
R1726 VSS.n301 VSS.n300 162.852
R1727 VSS.n431 VSS.n430 162.852
R1728 VSS.n469 VSS.n468 162.852
R1729 VSS.n304 VSS.n303 160.439
R1730 VSS.n434 VSS.n433 160.439
R1731 VSS.n472 VSS.n471 160.439
R1732 VSS.n1212 VSS.t974 159.19
R1733 VSS.n352 VSS.n351 158.4
R1734 VSS.n844 VSS.t90 158.037
R1735 VSS.n182 VSS.t1295 156.332
R1736 VSS.n182 VSS.t122 156.332
R1737 VSS.n180 VSS.t1108 156.332
R1738 VSS.n180 VSS.t1834 156.332
R1739 VSS.n178 VSS.t1655 156.332
R1740 VSS.n178 VSS.t811 156.332
R1741 VSS.n254 VSS.t445 156.332
R1742 VSS.n254 VSS.t178 156.332
R1743 VSS.n250 VSS.t1629 156.332
R1744 VSS.n250 VSS.t1401 156.332
R1745 VSS.n252 VSS.t585 156.332
R1746 VSS.n252 VSS.t1576 156.332
R1747 VSS.n1498 VSS.t283 156.332
R1748 VSS.n1498 VSS.t1133 156.332
R1749 VSS.n1495 VSS.t1187 156.332
R1750 VSS.n1495 VSS.t1904 156.332
R1751 VSS.n804 VSS.t336 156.332
R1752 VSS.n804 VSS.t1937 156.332
R1753 VSS.n838 VSS.t341 156.332
R1754 VSS.n838 VSS.t1444 156.332
R1755 VSS.n814 VSS.t547 156.332
R1756 VSS.n814 VSS.t360 156.332
R1757 VSS.n824 VSS.t1506 156.332
R1758 VSS.n824 VSS.t1918 156.332
R1759 VSS.n872 VSS.t1455 156.332
R1760 VSS.n872 VSS.t1615 156.332
R1761 VSS.n764 VSS.t650 156.332
R1762 VSS.n764 VSS.t1947 156.332
R1763 VSS.n790 VSS.t1091 156.332
R1764 VSS.n790 VSS.t14 156.332
R1765 VSS.n773 VSS.t1299 156.332
R1766 VSS.n773 VSS.t1779 156.332
R1767 VSS.n782 VSS.t482 156.332
R1768 VSS.n782 VSS.t729 156.332
R1769 VSS.n1493 VSS.n153 155.143
R1770 VSS.n1493 VSS.n154 155.061
R1771 VSS.n859 VSS.t1220 150.175
R1772 VSS.n799 VSS.t1347 150.175
R1773 VSS.n860 VSS.t272 149.728
R1774 VSS.n853 VSS.t540 149.728
R1775 VSS.n1447 VSS.n186 147.798
R1776 VSS.n1212 VSS.t1584 146.454
R1777 VSS.n1670 VSS.t1017 139.78
R1778 VSS.n1670 VSS.t1019 139.78
R1779 VSS.n1670 VSS.t996 139.78
R1780 VSS.n299 VSS.t979 139.78
R1781 VSS.n299 VSS.t1004 139.78
R1782 VSS.n299 VSS.t989 139.78
R1783 VSS.n299 VSS.t1027 139.78
R1784 VSS.n429 VSS.t992 139.78
R1785 VSS.n429 VSS.t1007 139.78
R1786 VSS.n429 VSS.t998 139.78
R1787 VSS.n429 VSS.t984 139.78
R1788 VSS.n467 VSS.t1024 139.78
R1789 VSS.n467 VSS.t1011 139.78
R1790 VSS.n467 VSS.t1021 139.78
R1791 VSS.n467 VSS.t1030 139.78
R1792 VSS.n1041 VSS.n1040 128.913
R1793 VSS.n1039 VSS.n1038 128.913
R1794 VSS.n1035 VSS.n1034 128.913
R1795 VSS.n1025 VSS.n621 128.913
R1796 VSS.n1023 VSS.n1022 128.913
R1797 VSS.n1005 VSS.n1004 128.913
R1798 VSS.n1003 VSS.n1002 128.913
R1799 VSS.n999 VSS.n998 128.913
R1800 VSS.n989 VSS.n623 128.913
R1801 VSS.n987 VSS.n986 128.913
R1802 VSS.n1180 VSS.n1179 128.913
R1803 VSS.n1159 VSS.n1158 128.913
R1804 VSS.n1163 VSS.n1162 128.913
R1805 VSS.n1165 VSS.n1164 128.913
R1806 VSS.n1168 VSS.n625 128.913
R1807 VSS.n971 VSS.n970 128.913
R1808 VSS.n969 VSS.n968 128.913
R1809 VSS.n965 VSS.n964 128.913
R1810 VSS.n955 VSS.n619 128.913
R1811 VSS.n953 VSS.n952 128.913
R1812 VSS.n1075 VSS.n1074 128.913
R1813 VSS.n1073 VSS.n1072 128.913
R1814 VSS.n1069 VSS.n1068 128.913
R1815 VSS.n1059 VSS.n617 128.913
R1816 VSS.n1057 VSS.n1056 128.913
R1817 VSS.n937 VSS.n936 128.913
R1818 VSS.n935 VSS.n934 128.913
R1819 VSS.n931 VSS.n930 128.913
R1820 VSS.n921 VSS.n615 128.913
R1821 VSS.n919 VSS.n918 128.913
R1822 VSS.n1092 VSS.n1091 128.913
R1823 VSS.n1096 VSS.n1095 128.913
R1824 VSS.n1098 VSS.n1097 128.913
R1825 VSS.n1101 VSS.n613 128.913
R1826 VSS.n737 VSS.n736 128.913
R1827 VSS.n903 VSS.n902 128.913
R1828 VSS.n901 VSS.n900 128.913
R1829 VSS.n897 VSS.n896 128.913
R1830 VSS.n887 VSS.n611 128.913
R1831 VSS.n885 VSS.n884 128.913
R1832 VSS.n1116 VSS.n1115 128.913
R1833 VSS.n1120 VSS.n1119 128.913
R1834 VSS.n1122 VSS.n1121 128.913
R1835 VSS.n1133 VSS.n609 128.913
R1836 VSS.n866 VSS.n865 128.913
R1837 VSS.n1042 VSS.n1041 128.855
R1838 VSS.n1039 VSS.n1036 128.855
R1839 VSS.n1035 VSS.n1024 128.855
R1840 VSS.n1026 VSS.n621 128.855
R1841 VSS.n1023 VSS.n1020 128.855
R1842 VSS.n1006 VSS.n1005 128.855
R1843 VSS.n1003 VSS.n1000 128.855
R1844 VSS.n999 VSS.n988 128.855
R1845 VSS.n990 VSS.n623 128.855
R1846 VSS.n987 VSS.n984 128.855
R1847 VSS.n1180 VSS.n627 128.855
R1848 VSS.n1159 VSS.n1157 128.855
R1849 VSS.n1163 VSS.n1160 128.855
R1850 VSS.n1166 VSS.n1165 128.855
R1851 VSS.n1169 VSS.n625 128.855
R1852 VSS.n972 VSS.n971 128.855
R1853 VSS.n969 VSS.n966 128.855
R1854 VSS.n965 VSS.n954 128.855
R1855 VSS.n956 VSS.n619 128.855
R1856 VSS.n953 VSS.n950 128.855
R1857 VSS.n1076 VSS.n1075 128.855
R1858 VSS.n1073 VSS.n1070 128.855
R1859 VSS.n1069 VSS.n1058 128.855
R1860 VSS.n1060 VSS.n617 128.855
R1861 VSS.n1057 VSS.n1054 128.855
R1862 VSS.n938 VSS.n937 128.855
R1863 VSS.n935 VSS.n932 128.855
R1864 VSS.n931 VSS.n920 128.855
R1865 VSS.n922 VSS.n615 128.855
R1866 VSS.n919 VSS.n916 128.855
R1867 VSS.n1092 VSS.n734 128.855
R1868 VSS.n1096 VSS.n1093 128.855
R1869 VSS.n1099 VSS.n1098 128.855
R1870 VSS.n1102 VSS.n613 128.855
R1871 VSS.n738 VSS.n737 128.855
R1872 VSS.n904 VSS.n903 128.855
R1873 VSS.n901 VSS.n898 128.855
R1874 VSS.n897 VSS.n886 128.855
R1875 VSS.n888 VSS.n611 128.855
R1876 VSS.n885 VSS.n882 128.855
R1877 VSS.n1116 VSS.n719 128.855
R1878 VSS.n1120 VSS.n1117 128.855
R1879 VSS.n1123 VSS.n1122 128.855
R1880 VSS.n866 VSS.n863 128.855
R1881 VSS.n1147 VSS.n609 128.823
R1882 VSS.t1897 VSS.t1908 127.922
R1883 VSS.t1908 VSS.t1913 127.922
R1884 VSS.t1913 VSS.t943 127.922
R1885 VSS.t943 VSS.t1175 127.922
R1886 VSS.t1175 VSS.t1176 127.922
R1887 VSS.t1247 VSS.t128 127.922
R1888 VSS.t128 VSS.t1246 127.922
R1889 VSS.t1246 VSS.t639 127.922
R1890 VSS.t639 VSS.t641 127.922
R1891 VSS.t641 VSS.t643 127.922
R1892 VSS.t1125 VSS.t1129 127.846
R1893 VSS.t1129 VSS.t1136 127.846
R1894 VSS.t1136 VSS.t287 127.846
R1895 VSS.t287 VSS.t288 127.846
R1896 VSS.t288 VSS.t505 127.846
R1897 VSS.t1693 VSS.t1689 127.846
R1898 VSS.t1689 VSS.t1692 127.846
R1899 VSS.t1692 VSS.t569 127.846
R1900 VSS.t569 VSS.t571 127.846
R1901 VSS.t571 VSS.t573 127.846
R1902 VSS.n848 VSS.t539 123.335
R1903 VSS.t1905 VSS.t1897 122.593
R1904 VSS.t643 VSS.t1178 122.593
R1905 VSS.t1134 VSS.t1125 122.519
R1906 VSS.t573 VSS.t506 122.519
R1907 VSS.n1626 VSS.n1624 120.757
R1908 VSS.n120 VSS.n118 120.757
R1909 VSS.n1618 VSS.n1616 120.757
R1910 VSS.n1615 VSS.n1613 120.757
R1911 VSS.n1608 VSS.n1606 120.757
R1912 VSS.n1605 VSS.n1603 120.757
R1913 VSS.n1599 VSS.n1597 120.757
R1914 VSS.n1596 VSS.n1594 120.757
R1915 VSS.n1590 VSS.n1588 120.757
R1916 VSS.n1587 VSS.n1585 120.757
R1917 VSS.n1581 VSS.n1579 120.757
R1918 VSS.n1578 VSS.n1576 120.757
R1919 VSS.n1571 VSS.n1569 120.757
R1920 VSS.n1568 VSS.n1566 120.757
R1921 VSS.n116 VSS.n114 120.757
R1922 VSS.n113 VSS.n111 120.757
R1923 VSS.n578 VSS.n576 120.757
R1924 VSS.n581 VSS.n579 120.757
R1925 VSS.n594 VSS.n592 120.757
R1926 VSS.n597 VSS.n595 120.757
R1927 VSS.n1287 VSS.n1285 120.757
R1928 VSS.n1290 VSS.n1288 120.757
R1929 VSS.n543 VSS.n541 120.757
R1930 VSS.n570 VSS.n568 120.757
R1931 VSS.n534 VSS.n532 120.757
R1932 VSS.n538 VSS.n536 120.757
R1933 VSS.n265 VSS.n263 120.757
R1934 VSS.n529 VSS.n527 120.757
R1935 VSS.n249 VSS.n247 120.757
R1936 VSS.n260 VSS.n258 120.757
R1937 VSS.n243 VSS.n241 120.757
R1938 VSS.n246 VSS.n244 120.757
R1939 VSS.n98 VSS.n96 120.757
R1940 VSS.n101 VSS.n99 120.757
R1941 VSS.n1358 VSS.n1356 120.757
R1942 VSS.n1361 VSS.n1359 120.757
R1943 VSS.n1370 VSS.n1368 120.757
R1944 VSS.n1373 VSS.n1371 120.757
R1945 VSS.n233 VSS.n231 120.757
R1946 VSS.n1381 VSS.n1379 120.757
R1947 VSS.n236 VSS.n234 120.757
R1948 VSS.n239 VSS.n237 120.757
R1949 VSS.n174 VSS.n172 120.757
R1950 VSS.n177 VSS.n175 120.757
R1951 VSS.n171 VSS.n169 120.757
R1952 VSS.n1471 VSS.n1469 120.757
R1953 VSS.n272 VSS.n270 120.757
R1954 VSS.n516 VSS.n514 120.757
R1955 VSS.n505 VSS.n503 120.757
R1956 VSS.n508 VSS.n506 120.757
R1957 VSS.n284 VSS.n282 120.757
R1958 VSS.n287 VSS.n285 120.757
R1959 VSS.n275 VSS.n273 120.757
R1960 VSS.n278 VSS.n276 120.757
R1961 VSS.n131 VSS.n129 120.757
R1962 VSS.n134 VSS.n132 120.757
R1963 VSS.n128 VSS.n126 120.757
R1964 VSS.n1529 VSS.n1527 120.757
R1965 VSS.n1271 VSS.n1269 120.757
R1966 VSS.n1274 VSS.n1272 120.757
R1967 VSS.n1250 VSS.n1248 120.757
R1968 VSS.n1282 VSS.n1280 120.757
R1969 VSS.n1262 VSS.n1260 120.757
R1970 VSS.n1265 VSS.n1263 120.757
R1971 VSS.n1253 VSS.n1251 120.757
R1972 VSS.n1256 VSS.n1254 120.757
R1973 VSS.n72 VSS.n70 120.757
R1974 VSS.n75 VSS.n73 120.757
R1975 VSS.n69 VSS.n67 120.757
R1976 VSS.n1683 VSS.n1681 120.757
R1977 VSS.n42 VSS.n40 120.757
R1978 VSS.n45 VSS.n43 120.757
R1979 VSS.n39 VSS.n37 120.757
R1980 VSS.n1703 VSS.n1701 120.757
R1981 VSS.n15 VSS.n13 120.757
R1982 VSS.n18 VSS.n16 120.757
R1983 VSS.n12 VSS.n10 120.757
R1984 VSS.n1723 VSS.n1721 120.757
R1985 VSS.n290 VSS.n288 120.757
R1986 VSS.n293 VSS.n291 120.757
R1987 VSS.n310 VSS.n297 120.757
R1988 VSS.n313 VSS.n311 120.757
R1989 VSS.n390 VSS.n388 120.757
R1990 VSS.n79 VSS.n77 120.757
R1991 VSS.n395 VSS.n393 120.757
R1992 VSS.n64 VSS.n62 120.757
R1993 VSS.n400 VSS.n398 120.757
R1994 VSS.n49 VSS.n47 120.757
R1995 VSS.n405 VSS.n403 120.757
R1996 VSS.n35 VSS.n33 120.757
R1997 VSS.n410 VSS.n408 120.757
R1998 VSS.n22 VSS.n20 120.757
R1999 VSS.n415 VSS.n413 120.757
R2000 VSS.n3 VSS.n1 120.757
R2001 VSS.n420 VSS.n418 120.757
R2002 VSS.n423 VSS.n421 120.757
R2003 VSS.n440 VSS.n427 120.757
R2004 VSS.n443 VSS.n441 120.757
R2005 VSS.n83 VSS.n81 120.757
R2006 VSS.n1660 VSS.n1658 120.757
R2007 VSS.n57 VSS.n55 120.757
R2008 VSS.n60 VSS.n58 120.757
R2009 VSS.n54 VSS.n52 120.757
R2010 VSS.n1693 VSS.n1691 120.757
R2011 VSS.n29 VSS.n27 120.757
R2012 VSS.n32 VSS.n30 120.757
R2013 VSS.n26 VSS.n24 120.757
R2014 VSS.n1713 VSS.n1711 120.757
R2015 VSS.n453 VSS.n451 120.757
R2016 VSS.n8 VSS.n6 120.757
R2017 VSS.n458 VSS.n456 120.757
R2018 VSS.n461 VSS.n459 120.757
R2019 VSS.n481 VSS.n479 120.757
R2020 VSS.n1313 VSS.n1311 120.757
R2021 VSS.n1316 VSS.n1314 120.757
R2022 VSS.n602 VSS.n600 120.757
R2023 VSS.n1216 VSS.n1214 120.757
R2024 VSS.n478 VSS.n465 120.754
R2025 VSS.n859 VSS.n858 119.644
R2026 VSS.n799 VSS.n798 119.644
R2027 VSS.n853 VSS.n852 117.001
R2028 VSS.n861 VSS.n860 117.001
R2029 VSS.n151 VSS.t70 110.507
R2030 VSS.n1424 VSS.n1423 99.7338
R2031 VSS.n1181 VSS.t197 97.7365
R2032 VSS.n120 VSS.n119 97.6833
R2033 VSS.n1615 VSS.n1614 97.6833
R2034 VSS.n1605 VSS.n1604 97.6833
R2035 VSS.n1596 VSS.n1595 97.6833
R2036 VSS.n1587 VSS.n1586 97.6833
R2037 VSS.n1578 VSS.n1577 97.6833
R2038 VSS.n1568 VSS.n1567 97.6833
R2039 VSS.n113 VSS.n112 97.6833
R2040 VSS.n578 VSS.n577 97.6833
R2041 VSS.n594 VSS.n593 97.6833
R2042 VSS.n1290 VSS.n1289 97.6833
R2043 VSS.n570 VSS.n569 97.6833
R2044 VSS.n538 VSS.n537 97.6833
R2045 VSS.n529 VSS.n528 97.6833
R2046 VSS.n260 VSS.n259 97.6833
R2047 VSS.n246 VSS.n245 97.6833
R2048 VSS.n101 VSS.n100 97.6833
R2049 VSS.n1358 VSS.n1357 97.6833
R2050 VSS.n1370 VSS.n1369 97.6833
R2051 VSS.n233 VSS.n232 97.6833
R2052 VSS.n236 VSS.n235 97.6833
R2053 VSS.n174 VSS.n173 97.6833
R2054 VSS.n171 VSS.n170 97.6833
R2055 VSS.n272 VSS.n271 97.6833
R2056 VSS.n505 VSS.n504 97.6833
R2057 VSS.n284 VSS.n283 97.6833
R2058 VSS.n275 VSS.n274 97.6833
R2059 VSS.n131 VSS.n130 97.6833
R2060 VSS.n128 VSS.n127 97.6833
R2061 VSS.n1271 VSS.n1270 97.6833
R2062 VSS.n1250 VSS.n1249 97.6833
R2063 VSS.n1262 VSS.n1261 97.6833
R2064 VSS.n1253 VSS.n1252 97.6833
R2065 VSS.n72 VSS.n71 97.6833
R2066 VSS.n69 VSS.n68 97.6833
R2067 VSS.n42 VSS.n41 97.6833
R2068 VSS.n39 VSS.n38 97.6833
R2069 VSS.n15 VSS.n14 97.6833
R2070 VSS.n12 VSS.n11 97.6833
R2071 VSS.n290 VSS.n289 97.6833
R2072 VSS.n390 VSS.n389 97.6833
R2073 VSS.n395 VSS.n394 97.6833
R2074 VSS.n400 VSS.n399 97.6833
R2075 VSS.n405 VSS.n404 97.6833
R2076 VSS.n410 VSS.n409 97.6833
R2077 VSS.n415 VSS.n414 97.6833
R2078 VSS.n420 VSS.n419 97.6833
R2079 VSS.n83 VSS.n82 97.6833
R2080 VSS.n57 VSS.n56 97.6833
R2081 VSS.n54 VSS.n53 97.6833
R2082 VSS.n29 VSS.n28 97.6833
R2083 VSS.n26 VSS.n25 97.6833
R2084 VSS.n453 VSS.n452 97.6833
R2085 VSS.n458 VSS.n457 97.6833
R2086 VSS.n1316 VSS.n1315 97.6833
R2087 VSS.n602 VSS.n601 97.6833
R2088 VSS.n1626 VSS.n1625 97.6819
R2089 VSS.n1618 VSS.n1617 97.6819
R2090 VSS.n1608 VSS.n1607 97.6819
R2091 VSS.n1599 VSS.n1598 97.6819
R2092 VSS.n1590 VSS.n1589 97.6819
R2093 VSS.n1581 VSS.n1580 97.6819
R2094 VSS.n1571 VSS.n1570 97.6819
R2095 VSS.n116 VSS.n115 97.6819
R2096 VSS.n581 VSS.n580 97.6819
R2097 VSS.n597 VSS.n596 97.6819
R2098 VSS.n1287 VSS.n1286 97.6819
R2099 VSS.n543 VSS.n542 97.6819
R2100 VSS.n534 VSS.n533 97.6819
R2101 VSS.n265 VSS.n264 97.6819
R2102 VSS.n249 VSS.n248 97.6819
R2103 VSS.n243 VSS.n242 97.6819
R2104 VSS.n98 VSS.n97 97.6819
R2105 VSS.n1361 VSS.n1360 97.6819
R2106 VSS.n1373 VSS.n1372 97.6819
R2107 VSS.n1381 VSS.n1380 97.6819
R2108 VSS.n239 VSS.n238 97.6819
R2109 VSS.n177 VSS.n176 97.6819
R2110 VSS.n1471 VSS.n1470 97.6819
R2111 VSS.n516 VSS.n515 97.6819
R2112 VSS.n508 VSS.n507 97.6819
R2113 VSS.n287 VSS.n286 97.6819
R2114 VSS.n278 VSS.n277 97.6819
R2115 VSS.n134 VSS.n133 97.6819
R2116 VSS.n1529 VSS.n1528 97.6819
R2117 VSS.n1274 VSS.n1273 97.6819
R2118 VSS.n1282 VSS.n1281 97.6819
R2119 VSS.n1265 VSS.n1264 97.6819
R2120 VSS.n1256 VSS.n1255 97.6819
R2121 VSS.n75 VSS.n74 97.6819
R2122 VSS.n1683 VSS.n1682 97.6819
R2123 VSS.n45 VSS.n44 97.6819
R2124 VSS.n1703 VSS.n1702 97.6819
R2125 VSS.n18 VSS.n17 97.6819
R2126 VSS.n1723 VSS.n1722 97.6819
R2127 VSS.n293 VSS.n292 97.6819
R2128 VSS.n313 VSS.n312 97.6819
R2129 VSS.n79 VSS.n78 97.6819
R2130 VSS.n64 VSS.n63 97.6819
R2131 VSS.n49 VSS.n48 97.6819
R2132 VSS.n35 VSS.n34 97.6819
R2133 VSS.n22 VSS.n21 97.6819
R2134 VSS.n3 VSS.n2 97.6819
R2135 VSS.n423 VSS.n422 97.6819
R2136 VSS.n443 VSS.n442 97.6819
R2137 VSS.n1660 VSS.n1659 97.6819
R2138 VSS.n60 VSS.n59 97.6819
R2139 VSS.n1693 VSS.n1692 97.6819
R2140 VSS.n32 VSS.n31 97.6819
R2141 VSS.n1713 VSS.n1712 97.6819
R2142 VSS.n8 VSS.n7 97.6819
R2143 VSS.n461 VSS.n460 97.6819
R2144 VSS.n481 VSS.n480 97.6819
R2145 VSS.n1313 VSS.n1312 97.6819
R2146 VSS.n1216 VSS.n1215 97.6819
R2147 VSS.n309 VSS.n308 97.6215
R2148 VSS.n1561 VSS.t285 97.6148
R2149 VSS.n477 VSS.n476 97.5878
R2150 VSS.n439 VSS.n438 97.5611
R2151 VSS.t724 VSS.t1195 97.4563
R2152 VSS.n303 VSS.n302 94.4341
R2153 VSS.n433 VSS.n432 94.4341
R2154 VSS.n471 VSS.n470 94.4341
R2155 VSS.n1428 VSS.n1427 93.8672
R2156 VSS.t1289 VSS.n93 92.1048
R2157 VSS.n186 VSS.t511 91.8752
R2158 VSS.n1676 VSS 89.5858
R2159 VSS.t973 VSS.t22 87.8175
R2160 VSS.t22 VSS.t20 87.8175
R2161 VSS.t20 VSS.t1854 87.8175
R2162 VSS.t490 VSS.t492 87.8175
R2163 VSS.t492 VSS.t494 87.8175
R2164 VSS.t494 VSS.t893 87.8175
R2165 VSS.t893 VSS.t906 87.8175
R2166 VSS.t906 VSS.t921 87.8175
R2167 VSS.t543 VSS.t541 87.8175
R2168 VSS.t541 VSS.t542 87.8175
R2169 VSS.t542 VSS.t232 87.8175
R2170 VSS.t232 VSS.t228 87.8175
R2171 VSS.t228 VSS.t230 87.8175
R2172 VSS.t589 VSS.t683 87.8175
R2173 VSS.t683 VSS.t694 87.8175
R2174 VSS.t694 VSS.t1589 87.8175
R2175 VSS.t1589 VSS.t1161 87.8175
R2176 VSS.t1161 VSS.t1583 87.8175
R2177 VSS.t410 VSS.t945 87.8175
R2178 VSS.t945 VSS.t1413 87.8175
R2179 VSS.t1413 VSS.t1367 87.8175
R2180 VSS.t1367 VSS.t1369 87.8175
R2181 VSS.t1369 VSS.t1365 87.8175
R2182 VSS.n1513 VSS.n143 84.9212
R2183 VSS.n1667 VSS.n1666 84.5046
R2184 VSS.t1854 VSS.t1590 84.1585
R2185 VSS.t488 VSS.t490 84.1585
R2186 VSS.t230 VSS.t377 84.1585
R2187 VSS.t581 VSS.t589 84.1585
R2188 VSS.t1365 VSS.t1577 84.1585
R2189 VSS.n223 VSS.t1606 83.8604
R2190 VSS.n219 VSS.t1308 83.8604
R2191 VSS.n1236 VSS.t2031 83.7809
R2192 VSS.n215 VSS.t671 83.7809
R2193 VSS.n218 VSS.t772 83.7809
R2194 VSS.n227 VSS.t1608 83.7809
R2195 VSS.n221 VSS.t416 83.7809
R2196 VSS.n228 VSS.t1194 83.7809
R2197 VSS.n225 VSS.t330 83.7809
R2198 VSS.n1484 VSS.t274 83.7809
R2199 VSS.n1487 VSS.t395 83.7809
R2200 VSS.n1481 VSS.t150 83.7809
R2201 VSS.n160 VSS.t1254 83.7809
R2202 VSS.n1491 VSS.t768 83.7809
R2203 VSS.n157 VSS.t355 83.7809
R2204 VSS.n159 VSS.t173 83.7809
R2205 VSS.n158 VSS.t1156 83.7809
R2206 VSS.n678 VSS.t1987 83.7809
R2207 VSS.n672 VSS.t1729 83.7809
R2208 VSS.n675 VSS.t1975 83.7809
R2209 VSS.n664 VSS.t1996 83.7809
R2210 VSS.n668 VSS.t1735 83.7809
R2211 VSS.n667 VSS.t1979 83.7809
R2212 VSS.n686 VSS.t2011 83.7809
R2213 VSS.n680 VSS.t1709 83.7809
R2214 VSS.n683 VSS.t1958 83.7809
R2215 VSS.n657 VSS.t2005 83.7809
R2216 VSS.n661 VSS.t1750 83.7809
R2217 VSS.n660 VSS.t1985 83.7809
R2218 VSS.n694 VSS.t2013 83.7809
R2219 VSS.n688 VSS.t1707 83.7809
R2220 VSS.n691 VSS.t1955 83.7809
R2221 VSS.n650 VSS.t1993 83.7809
R2222 VSS.n654 VSS.t1733 83.7809
R2223 VSS.n653 VSS.t1977 83.7809
R2224 VSS.n702 VSS.t2019 83.7809
R2225 VSS.n696 VSS.t1715 83.7809
R2226 VSS.n699 VSS.t1983 83.7809
R2227 VSS.n643 VSS.t2021 83.7809
R2228 VSS.n647 VSS.t1711 83.7809
R2229 VSS.n646 VSS.t1981 83.7809
R2230 VSS.n710 VSS.t2017 83.7809
R2231 VSS.n704 VSS.t1702 83.7809
R2232 VSS.n707 VSS.t1962 83.7809
R2233 VSS.n604 VSS.t1613 83.7809
R2234 VSS.n564 VSS.t500 83.7809
R2235 VSS.n556 VSS.t224 83.7809
R2236 VSS.n552 VSS.t1111 83.7809
R2237 VSS.n554 VSS.t1653 83.7809
R2238 VSS.n553 VSS.t446 83.7809
R2239 VSS.n547 VSS.t1628 83.7809
R2240 VSS.n550 VSS.t693 83.7809
R2241 VSS.n559 VSS.t1182 83.7809
R2242 VSS.n1560 VSS.t2032 83.7809
R2243 VSS.n846 VSS.t725 83.774
R2244 VSS.n840 VSS.t561 83.7659
R2245 VSS.n841 VSS.t538 83.7659
R2246 VSS.n1306 VSS.t848 83.7653
R2247 VSS.n1243 VSS.t169 83.7653
R2248 VSS.n1242 VSS.t1034 83.7653
R2249 VSS.n1241 VSS.t1259 83.7653
R2250 VSS.n1240 VSS.t195 83.7653
R2251 VSS.n1239 VSS.t331 83.7653
R2252 VSS.n1238 VSS.t1884 83.7653
R2253 VSS.n1237 VSS.t594 83.7653
R2254 VSS.n1559 VSS.t614 83.7653
R2255 VSS.n1557 VSS.t1498 83.7653
R2256 VSS.n1555 VSS.t595 83.7653
R2257 VSS.n1553 VSS.t1273 83.7653
R2258 VSS.n1551 VSS.t1074 83.7653
R2259 VSS.n1549 VSS.t409 83.7653
R2260 VSS.n1547 VSS.t645 83.7653
R2261 VSS.n1564 VSS.t63 83.7653
R2262 VSS.n1411 VSS.t1781 83.7497
R2263 VSS.n1405 VSS.t1324 83.7497
R2264 VSS.n1421 VSS.t354 83.7497
R2265 VSS.n203 VSS.t1307 83.7497
R2266 VSS.n378 VSS.t1077 83.7497
R2267 VSS.n383 VSS.t1921 83.7497
R2268 VSS.n325 VSS.t408 83.7497
R2269 VSS.n1431 VSS.t1465 83.7497
R2270 VSS.n360 VSS.t1301 83.7497
R2271 VSS.n1452 VSS.t526 83.7497
R2272 VSS.n1457 VSS.t76 83.7497
R2273 VSS.n191 VSS.t579 83.7497
R2274 VSS.n187 VSS.t108 83.7497
R2275 VSS.n1439 VSS.t558 83.7497
R2276 VSS.n347 VSS.t210 83.7497
R2277 VSS.n320 VSS.t536 83.7495
R2278 VSS VSS.t1540 83.7183
R2279 VSS VSS.t843 83.7183
R2280 VSS VSS.t1331 83.7183
R2281 VSS VSS.t1271 83.7183
R2282 VSS VSS.t1515 83.7183
R2283 VSS VSS.t545 83.7183
R2284 VSS VSS.t749 83.7183
R2285 VSS VSS.t1777 83.7183
R2286 VSS VSS.t1597 83.7183
R2287 VSS.n1228 VSS.t504 83.7172
R2288 VSS.n1229 VSS.t1188 83.7172
R2289 VSS.n1230 VSS.t1294 83.7172
R2290 VSS.n1231 VSS.t1102 83.7172
R2291 VSS.n1232 VSS.t1656 83.7172
R2292 VSS.n1233 VSS.t440 83.7172
R2293 VSS.n1234 VSS.t1637 83.7172
R2294 VSS.n1235 VSS.t587 83.7172
R2295 VSS.n1539 VSS.t286 83.7172
R2296 VSS.n1540 VSS.t1185 83.7172
R2297 VSS.n1541 VSS.t1291 83.7172
R2298 VSS.n1542 VSS.t1096 83.7172
R2299 VSS.n1543 VSS.t1644 83.7172
R2300 VSS.n1544 VSS.t1801 83.7172
R2301 VSS.n1545 VSS.t1633 83.7172
R2302 VSS.n1562 VSS.t691 83.7172
R2303 VSS.n1181 VSS.t721 82.7002
R2304 VSS.n1224 VSS.t973 79.5847
R2305 VSS.n1225 VSS.n575 79.5698
R2306 VSS.t340 VSS.n839 76.9404
R2307 VSS.n839 VSS.t1443 76.9404
R2308 VSS.n1666 VSS.n1665 72.3005
R2309 VSS.n1331 VSS.t581 70.4371
R2310 VSS.n1623 VSS.n1622 69.4053
R2311 VSS.n1621 VSS.n1620 69.4053
R2312 VSS.n1611 VSS.n1610 69.4053
R2313 VSS.n1602 VSS.n1601 69.4053
R2314 VSS.n1593 VSS.n1592 69.4053
R2315 VSS.n1584 VSS.n1583 69.4053
R2316 VSS.n1574 VSS.n1573 69.4053
R2317 VSS.n1631 VSS.n1630 69.4053
R2318 VSS.n1330 VSS.n1329 69.4053
R2319 VSS.n1223 VSS.n1222 69.4053
R2320 VSS.n1292 VSS.n1291 69.4053
R2321 VSS.n572 VSS.n571 69.4053
R2322 VSS.n540 VSS.n539 69.4053
R2323 VSS.n531 VSS.n530 69.4053
R2324 VSS.n262 VSS.n261 69.4053
R2325 VSS.n1342 VSS.n1341 69.4053
R2326 VSS.n1641 VSS.n1640 69.4053
R2327 VSS.n1367 VSS.n1366 69.4053
R2328 VSS.n1376 VSS.n1375 69.4053
R2329 VSS.n1378 VSS.n1377 69.4053
R2330 VSS.n1355 VSS.n1354 69.4053
R2331 VSS.n1466 VSS.n1465 69.4053
R2332 VSS.n1468 VSS.n1467 69.4053
R2333 VSS.n513 VSS.n512 69.4053
R2334 VSS.n511 VSS.n510 69.4053
R2335 VSS.n502 VSS.n501 69.4053
R2336 VSS.n281 VSS.n280 69.4053
R2337 VSS.n1524 VSS.n1523 69.4053
R2338 VSS.n1526 VSS.n1525 69.4053
R2339 VSS.n1277 VSS.n1276 69.4053
R2340 VSS.n1279 VSS.n1278 69.4053
R2341 VSS.n1268 VSS.n1267 69.4053
R2342 VSS.n1259 VSS.n1258 69.4053
R2343 VSS.n1680 VSS.n1679 69.4053
R2344 VSS.n1698 VSS.n1697 69.4053
R2345 VSS.n1700 VSS.n1699 69.4053
R2346 VSS.n1718 VSS.n1717 69.4053
R2347 VSS.n1720 VSS.n1719 69.4053
R2348 VSS.n296 VSS.n295 69.4053
R2349 VSS.n316 VSS.n315 69.4053
R2350 VSS.n392 VSS.n391 69.4053
R2351 VSS.n397 VSS.n396 69.4053
R2352 VSS.n402 VSS.n401 69.4053
R2353 VSS.n407 VSS.n406 69.4053
R2354 VSS.n412 VSS.n411 69.4053
R2355 VSS.n417 VSS.n416 69.4053
R2356 VSS.n426 VSS.n425 69.4053
R2357 VSS.n446 VSS.n445 69.4053
R2358 VSS.n1657 VSS.n1656 69.4053
R2359 VSS.n1688 VSS.n1687 69.4053
R2360 VSS.n1690 VSS.n1689 69.4053
R2361 VSS.n1708 VSS.n1707 69.4053
R2362 VSS.n1710 VSS.n1709 69.4053
R2363 VSS.n455 VSS.n454 69.4053
R2364 VSS.n464 VSS.n463 69.4053
R2365 VSS.n484 VSS.n483 69.4053
R2366 VSS.n1318 VSS.n1317 69.4053
R2367 VSS.n1213 VSS.n1212 69.4053
R2368 VSS.n1678 VSS.n1677 68.824
R2369 VSS.n1621 VSS.t1247 66.6268
R2370 VSS.n1622 VSS.t1693 66.5865
R2371 VSS.n1308 VSS.n1307 64.0892
R2372 VSS.t263 VSS.t244 62.9607
R2373 VSS.t244 VSS.t246 62.9607
R2374 VSS.t246 VSS.t1296 62.9607
R2375 VSS.t1296 VSS.t1297 62.9607
R2376 VSS.t1297 VSS.t226 62.9607
R2377 VSS.t1425 VSS.t1426 62.9607
R2378 VSS.t1426 VSS.t1427 62.9607
R2379 VSS.t1427 VSS.t1215 62.9607
R2380 VSS.t1215 VSS.t1211 62.9607
R2381 VSS.t1211 VSS.t1213 62.0747
R2382 VSS.t1176 VSS.n1621 61.2967
R2383 VSS.n1622 VSS.t505 61.2596
R2384 VSS.n1668 VSS.n1667 60.9816
R2385 VSS.t255 VSS.t263 60.3374
R2386 VSS.t1835 VSS.t1842 58.7079
R2387 VSS.t1842 VSS.t1844 58.7079
R2388 VSS.t1844 VSS.t1099 58.7079
R2389 VSS.t1099 VSS.t1101 58.7079
R2390 VSS.t1101 VSS.t1110 58.7079
R2391 VSS.t1610 VSS.t1593 58.7079
R2392 VSS.t1593 VSS.t15 58.7079
R2393 VSS.t15 VSS.t1361 58.7079
R2394 VSS.t1361 VSS.t1363 58.7079
R2395 VSS.t1363 VSS.t1359 58.7079
R2396 VSS.t806 VSS.t812 58.7079
R2397 VSS.t812 VSS.t818 58.7079
R2398 VSS.t818 VSS.t1657 58.7079
R2399 VSS.t1657 VSS.t1642 58.7079
R2400 VSS.t1642 VSS.t1650 58.7079
R2401 VSS.t1877 VSS.t1624 58.7079
R2402 VSS.t1624 VSS.t1876 58.7079
R2403 VSS.t1876 VSS.t305 58.7079
R2404 VSS.t305 VSS.t307 58.7079
R2405 VSS.t307 VSS.t309 58.7079
R2406 VSS.t181 VSS.t185 58.7079
R2407 VSS.t185 VSS.t187 58.7079
R2408 VSS.t187 VSS.t1802 58.7079
R2409 VSS.t1802 VSS.t1804 58.7079
R2410 VSS.t1804 VSS.t443 58.7079
R2411 VSS.t944 VSS.t241 58.7079
R2412 VSS.t241 VSS.t600 58.7079
R2413 VSS.t600 VSS.t935 58.7079
R2414 VSS.t935 VSS.t937 58.7079
R2415 VSS.t937 VSS.t933 58.7079
R2416 VSS.t1386 VSS.t1394 58.7079
R2417 VSS.t1394 VSS.t1396 58.7079
R2418 VSS.t1396 VSS.t1638 58.7079
R2419 VSS.t1638 VSS.t1626 58.7079
R2420 VSS.t1626 VSS.t1631 58.7079
R2421 VSS.t941 VSS.t942 58.7079
R2422 VSS.t942 VSS.t940 58.7079
R2423 VSS.t940 VSS.t1309 58.7079
R2424 VSS.t1309 VSS.t1311 58.7079
R2425 VSS.t1311 VSS.t1313 58.7079
R2426 VSS.t1569 VSS.t1581 58.7079
R2427 VSS.t1581 VSS.t1585 58.7079
R2428 VSS.t1585 VSS.t588 58.7079
R2429 VSS.t588 VSS.t591 58.7079
R2430 VSS.t591 VSS.t685 58.7079
R2431 VSS.t487 VSS.t486 58.7079
R2432 VSS.t485 VSS.t487 58.7079
R2433 VSS.t779 VSS.t485 58.7079
R2434 VSS.t781 VSS.t779 58.7079
R2435 VSS.t783 VSS.t781 58.7079
R2436 VSS.t42 VSS.n124 57.4621
R2437 VSS.t1213 VSS.t1287 56.2618
R2438 VSS.t1840 VSS.t1835 56.2618
R2439 VSS.t1359 VSS.t1092 56.2618
R2440 VSS.t814 VSS.t806 56.2618
R2441 VSS.t309 VSS.t1651 56.2618
R2442 VSS.t183 VSS.t181 56.2618
R2443 VSS.t933 VSS.t1799 56.2618
R2444 VSS.t1392 VSS.t1386 56.2618
R2445 VSS.t1313 VSS.t1635 56.2618
R2446 VSS.t1579 VSS.t1569 56.2618
R2447 VSS.t688 VSS.t783 56.2618
R2448 VSS.n1397 VSS.n88 55.2769
R2449 VSS.n763 VSS.t649 54.8434
R2450 VSS.n763 VSS.t1946 54.8434
R2451 VSS.n813 VSS.t546 53.4553
R2452 VSS.n813 VSS.t359 53.4553
R2453 VSS.n823 VSS.t1505 53.4553
R2454 VSS.n823 VSS.t1917 53.4553
R2455 VSS.n871 VSS.t1454 53.4553
R2456 VSS.n871 VSS.t1614 53.4553
R2457 VSS.n772 VSS.t1298 53.4553
R2458 VSS.n772 VSS.t1778 53.4553
R2459 VSS.n781 VSS.t481 53.4553
R2460 VSS.n781 VSS.t728 53.4553
R2461 VSS.n803 VSS.t335 53.4553
R2462 VSS.n803 VSS.t1936 53.4553
R2463 VSS.n789 VSS.t1090 52.1358
R2464 VSS.n789 VSS.t13 52.1358
R2465 VSS.t428 VSS.n143 50.7962
R2466 VSS.n386 VSS.n385 49.2313
R2467 VSS.n1426 VSS.n1425 49.2313
R2468 VSS.n1398 VSS.n109 46.6115
R2469 VSS.n1429 VSS.n198 46.1221
R2470 VSS.n1223 VSS.t543 45.7385
R2471 VSS.n1330 VSS.t410 45.7385
R2472 VSS.t1132 VSS.n1499 44.2031
R2473 VSS.n1499 VSS.t282 44.2031
R2474 VSS.t1903 VSS.n1496 44.2031
R2475 VSS.n1496 VSS.t1186 44.2031
R2476 VSS.n1409 VSS.t251 43.6289
R2477 VSS.t121 VSS.n1493 43.2822
R2478 VSS.n363 VSS.n362 43.0473
R2479 VSS VSS.t1857 42.6224
R2480 VSS VSS.t1567 42.6029
R2481 VSS VSS.t1558 42.6029
R2482 VSS VSS.t1252 42.6029
R2483 VSS VSS.t1535 42.6029
R2484 VSS VSS.t365 42.6029
R2485 VSS VSS.t673 42.6029
R2486 VSS VSS.t1141 42.6029
R2487 VSS VSS.t1564 42.6029
R2488 VSS VSS.t1625 42.6029
R2489 VSS VSS.t687 42.6029
R2490 VSS VSS.t442 42.6029
R2491 VSS VSS.t1646 42.6029
R2492 VSS VSS.t1104 42.6029
R2493 VSS VSS.t1098 42.6029
R2494 VSS VSS.t1095 42.6029
R2495 VSS VSS.t1673 42.6029
R2496 VSS VSS.t484 42.6029
R2497 VSS VSS.t516 42.6029
R2498 VSS VSS.t1172 42.6029
R2499 VSS VSS.t1290 42.6029
R2500 VSS VSS.t262 42.6029
R2501 VSS VSS.t1131 42.6029
R2502 VSS VSS.t1285 42.6029
R2503 VSS VSS.t1293 42.6029
R2504 VSS VSS.t1139 42.6029
R2505 VSS VSS.t68 42.6029
R2506 VSS VSS.t322 42.6029
R2507 VSS VSS.t1823 42.6029
R2508 VSS VSS.t1762 42.6029
R2509 VSS VSS.t1919 42.6029
R2510 VSS VSS.t291 42.6029
R2511 VSS VSS.t1124 42.6029
R2512 VSS VSS.t248 42.6029
R2513 VSS VSS.t839 42.6029
R2514 VSS VSS.t1184 42.6029
R2515 VSS VSS.t1174 42.6029
R2516 VSS VSS.t239 42.6029
R2517 VSS VSS.t1948 42.6029
R2518 VSS VSS.t216 42.6029
R2519 VSS VSS.t534 42.6029
R2520 VSS VSS.t1883 42.6029
R2521 VSS VSS.t1267 42.6029
R2522 VSS VSS.t1073 42.6029
R2523 VSS VSS.t1221 42.6029
R2524 VSS VSS.t510 42.6029
R2525 VSS VSS.t503 42.6029
R2526 VSS VSS.t1602 42.6029
R2527 VSS VSS.t1328 42.6029
R2528 VSS VSS.t1207 42.6029
R2529 VSS VSS.t778 42.6029
R2530 VSS VSS.t281 42.6029
R2531 VSS VSS.t512 42.6029
R2532 VSS VSS.t260 42.6029
R2533 VSS VSS.t832 42.6029
R2534 VSS VSS.t1775 42.6029
R2535 VSS VSS.t953 42.6029
R2536 VSS VSS.t164 42.6029
R2537 VSS VSS.t1666 42.6029
R2538 VSS VSS.t2029 42.6029
R2539 VSS VSS.t955 42.6029
R2540 VSS VSS.t631 42.6029
R2541 VSS VSS.t726 42.6029
R2542 VSS VSS.t1041 42.6029
R2543 VSS VSS.t429 42.6029
R2544 VSS VSS.t529 42.5938
R2545 VSS VSS.t430 42.5938
R2546 VSS VSS.t1860 42.5938
R2547 VSS VSS.t1078 42.5938
R2548 VSS VSS.t1824 42.5938
R2549 VSS VSS.t1337 42.5938
R2550 VSS VSS.t1820 42.5938
R2551 VSS VSS.t1611 42.5938
R2552 VSS VSS.t1264 42.5938
R2553 VSS VSS.t977 42.5938
R2554 VSS VSS.t1448 42.5938
R2555 VSS VSS.t658 42.5938
R2556 VSS VSS.t131 42.5938
R2557 VSS VSS.t1668 42.5938
R2558 VSS VSS.t1494 42.5938
R2559 VSS VSS.t1432 42.5938
R2560 VSS VSS.t708 42.5938
R2561 VSS VSS.t301 42.5938
R2562 VSS VSS.t71 42.5938
R2563 VSS VSS.t968 42.5938
R2564 VSS VSS.t91 42.5938
R2565 VSS.t921 VSS.n1223 42.0795
R2566 VSS.t1583 VSS.n1330 42.0795
R2567 VSS.n488 VSS.n450 38.8103
R2568 VSS.n300 VSS.n299 38.6833
R2569 VSS.n430 VSS.n429 38.6833
R2570 VSS.n468 VSS.n467 38.6833
R2571 VSS.t62 VSS.n1565 38.6248
R2572 VSS.n1575 VSS.t62 37.3021
R2573 VSS.n849 VSS.n843 35.2646
R2574 VSS.n350 VSS.t259 35.2005
R2575 VSS.t831 VSS.n1437 35.2005
R2576 VSS.t220 VSS.n199 35.2005
R2577 VSS.t838 VSS.n318 35.2005
R2578 VSS.t261 VSS.n201 35.2005
R2579 VSS.n1418 VSS.t1109 35.2005
R2580 VSS.n1611 VSS.t1425 32.7923
R2581 VSS.n1602 VSS.t1610 30.5773
R2582 VSS.n1593 VSS.t1877 30.5773
R2583 VSS.n1584 VSS.t944 30.5773
R2584 VSS.n1574 VSS.t941 30.5773
R2585 VSS.t486 VSS.n1631 30.5773
R2586 VSS.n1625 VSS.t574 30.462
R2587 VSS.n1624 VSS.t570 30.462
R2588 VSS.n1624 VSS.t572 30.462
R2589 VSS.n118 VSS.t1130 30.462
R2590 VSS.n118 VSS.t1137 30.462
R2591 VSS.n119 VSS.t1126 30.462
R2592 VSS.n1617 VSS.t644 30.462
R2593 VSS.n1616 VSS.t640 30.462
R2594 VSS.n1616 VSS.t642 30.462
R2595 VSS.n1613 VSS.t1909 30.462
R2596 VSS.n1613 VSS.t1914 30.462
R2597 VSS.n1614 VSS.t1898 30.462
R2598 VSS.n1607 VSS.t1214 30.462
R2599 VSS.n1606 VSS.t1216 30.462
R2600 VSS.n1606 VSS.t1212 30.462
R2601 VSS.n1603 VSS.t245 30.462
R2602 VSS.n1603 VSS.t247 30.462
R2603 VSS.n1604 VSS.t264 30.462
R2604 VSS.n1598 VSS.t1360 30.462
R2605 VSS.n1597 VSS.t1362 30.462
R2606 VSS.n1597 VSS.t1364 30.462
R2607 VSS.n1594 VSS.t1843 30.462
R2608 VSS.n1594 VSS.t1845 30.462
R2609 VSS.n1595 VSS.t1836 30.462
R2610 VSS.n1589 VSS.t310 30.462
R2611 VSS.n1588 VSS.t306 30.462
R2612 VSS.n1588 VSS.t308 30.462
R2613 VSS.n1585 VSS.t813 30.462
R2614 VSS.n1585 VSS.t819 30.462
R2615 VSS.n1586 VSS.t807 30.462
R2616 VSS.n1580 VSS.t934 30.462
R2617 VSS.n1579 VSS.t936 30.462
R2618 VSS.n1579 VSS.t938 30.462
R2619 VSS.n1576 VSS.t186 30.462
R2620 VSS.n1576 VSS.t188 30.462
R2621 VSS.n1577 VSS.t182 30.462
R2622 VSS.n1570 VSS.t1314 30.462
R2623 VSS.n1569 VSS.t1310 30.462
R2624 VSS.n1569 VSS.t1312 30.462
R2625 VSS.n1566 VSS.t1395 30.462
R2626 VSS.n1566 VSS.t1397 30.462
R2627 VSS.n1567 VSS.t1387 30.462
R2628 VSS.n115 VSS.t784 30.462
R2629 VSS.n114 VSS.t780 30.462
R2630 VSS.n114 VSS.t782 30.462
R2631 VSS.n111 VSS.t1582 30.462
R2632 VSS.n111 VSS.t1586 30.462
R2633 VSS.n112 VSS.t1570 30.462
R2634 VSS.n577 VSS.t590 30.462
R2635 VSS.n576 VSS.t684 30.462
R2636 VSS.n576 VSS.t695 30.462
R2637 VSS.n579 VSS.t1368 30.462
R2638 VSS.n579 VSS.t1370 30.462
R2639 VSS.n580 VSS.t1366 30.462
R2640 VSS.n593 VSS.t491 30.462
R2641 VSS.n592 VSS.t493 30.462
R2642 VSS.n592 VSS.t495 30.462
R2643 VSS.n595 VSS.t233 30.462
R2644 VSS.n595 VSS.t229 30.462
R2645 VSS.n596 VSS.t231 30.462
R2646 VSS.n1286 VSS.t1892 30.462
R2647 VSS.n1285 VSS.t1890 30.462
R2648 VSS.n1285 VSS.t1886 30.462
R2649 VSS.n1288 VSS.t374 30.462
R2650 VSS.n1288 VSS.t903 30.462
R2651 VSS.n1289 VSS.t886 30.462
R2652 VSS.n542 VSS.t1795 30.462
R2653 VSS.n541 VSS.t1793 30.462
R2654 VSS.n541 VSS.t1791 30.462
R2655 VSS.n568 VSS.t869 30.462
R2656 VSS.n568 VSS.t905 30.462
R2657 VSS.n569 VSS.t890 30.462
R2658 VSS.n533 VSS.t1556 30.462
R2659 VSS.n532 VSS.t1554 30.462
R2660 VSS.n532 VSS.t714 30.462
R2661 VSS.n536 VSS.t888 30.462
R2662 VSS.n536 VSS.t925 30.462
R2663 VSS.n537 VSS.t908 30.462
R2664 VSS.n264 VSS.t759 30.462
R2665 VSS.n263 VSS.t277 30.462
R2666 VSS.n263 VSS.t794 30.462
R2667 VSS.n527 VSS.t892 30.462
R2668 VSS.n527 VSS.t899 30.462
R2669 VSS.n528 VSS.t372 30.462
R2670 VSS.n248 VSS.t1517 30.462
R2671 VSS.n247 VSS.t566 30.462
R2672 VSS.n247 VSS.t564 30.462
R2673 VSS.n258 VSS.t914 30.462
R2674 VSS.n258 VSS.t901 30.462
R2675 VSS.n259 VSS.t884 30.462
R2676 VSS.n242 VSS.t1925 30.462
R2677 VSS.n241 VSS.t1923 30.462
R2678 VSS.n241 VSS.t1927 30.462
R2679 VSS.n244 VSS.t386 30.462
R2680 VSS.n244 VSS.t910 30.462
R2681 VSS.n245 VSS.t877 30.462
R2682 VSS.n97 VSS.t1699 30.462
R2683 VSS.n96 VSS.t1697 30.462
R2684 VSS.n96 VSS.t1695 30.462
R2685 VSS.n99 VSS.t390 30.462
R2686 VSS.n99 VSS.t916 30.462
R2687 VSS.n100 VSS.t882 30.462
R2688 VSS.n1357 VSS.t1160 30.462
R2689 VSS.n1356 VSS.t1588 30.462
R2690 VSS.n1356 VSS.t1574 30.462
R2691 VSS.n1359 VSS.t1759 30.462
R2692 VSS.n1359 VSS.t1757 30.462
R2693 VSS.n1360 VSS.t1755 30.462
R2694 VSS.n1369 VSS.t86 30.462
R2695 VSS.n1368 VSS.t84 30.462
R2696 VSS.n1368 VSS.t962 30.462
R2697 VSS.n1371 VSS.t801 30.462
R2698 VSS.n1371 VSS.t803 30.462
R2699 VSS.n1372 VSS.t799 30.462
R2700 VSS.n232 VSS.t1403 30.462
R2701 VSS.n231 VSS.t1399 30.462
R2702 VSS.n231 VSS.t1391 30.462
R2703 VSS.n1379 VSS.t609 30.462
R2704 VSS.n1379 VSS.t607 30.462
R2705 VSS.n1380 VSS.t611 30.462
R2706 VSS.n235 VSS.t554 30.462
R2707 VSS.n234 VSS.t551 30.462
R2708 VSS.n234 VSS.t556 30.462
R2709 VSS.n237 VSS.t716 30.462
R2710 VSS.n237 VSS.t720 30.462
R2711 VSS.n238 VSS.t718 30.462
R2712 VSS.n173 VSS.t194 30.462
R2713 VSS.n172 VSS.t190 30.462
R2714 VSS.n172 VSS.t180 30.462
R2715 VSS.n175 VSS.t1067 30.462
R2716 VSS.n175 VSS.t1063 30.462
R2717 VSS.n176 VSS.t1065 30.462
R2718 VSS.n170 VSS.t1355 30.462
R2719 VSS.n169 VSS.t1353 30.462
R2720 VSS.n169 VSS.t1358 30.462
R2721 VSS.n1469 VSS.t731 30.462
R2722 VSS.n1469 VSS.t735 30.462
R2723 VSS.n1470 VSS.t733 30.462
R2724 VSS.n271 VSS.t817 30.462
R2725 VSS.n270 VSS.t809 30.462
R2726 VSS.n270 VSS.t1120 30.462
R2727 VSS.n514 VSS.t266 30.462
R2728 VSS.n514 VSS.t270 30.462
R2729 VSS.n515 VSS.t268 30.462
R2730 VSS.n504 VSS.t1787 30.462
R2731 VSS.n503 VSS.t1785 30.462
R2732 VSS.n503 VSS.t1789 30.462
R2733 VSS.n506 VSS.t384 30.462
R2734 VSS.n506 VSS.t382 30.462
R2735 VSS.n507 VSS.t380 30.462
R2736 VSS.n283 VSS.t1838 30.462
R2737 VSS.n282 VSS.t1853 30.462
R2738 VSS.n282 VSS.t1847 30.462
R2739 VSS.n285 VSS.t475 30.462
R2740 VSS.n285 VSS.t479 30.462
R2741 VSS.n286 VSS.t477 30.462
R2742 VSS.n274 VSS.t862 30.462
R2743 VSS.n273 VSS.t859 30.462
R2744 VSS.n273 VSS.t866 30.462
R2745 VSS.n276 VSS.t1118 30.462
R2746 VSS.n276 VSS.t1116 30.462
R2747 VSS.n277 VSS.t1114 30.462
R2748 VSS.n130 VSS.t120 30.462
R2749 VSS.n129 VSS.t258 30.462
R2750 VSS.n129 VSS.t250 30.462
R2751 VSS.n132 VSS.t158 30.462
R2752 VSS.n132 VSS.t156 30.462
R2753 VSS.n133 VSS.t154 30.462
R2754 VSS.n127 VSS.t35 30.462
R2755 VSS.n126 VSS.t41 30.462
R2756 VSS.n126 VSS.t37 30.462
R2757 VSS.n1527 VSS.t437 30.462
R2758 VSS.n1527 VSS.t435 30.462
R2759 VSS.n1528 VSS.t439 30.462
R2760 VSS.n1270 VSS.t1912 30.462
R2761 VSS.n1269 VSS.t1900 30.462
R2762 VSS.n1269 VSS.t1902 30.462
R2763 VSS.n1272 VSS.t1226 30.462
R2764 VSS.n1272 VSS.t1552 30.462
R2765 VSS.n1273 VSS.t593 30.462
R2766 VSS.n1249 VSS.t1305 30.462
R2767 VSS.n1248 VSS.t1303 30.462
R2768 VSS.n1248 VSS.t404 30.462
R2769 VSS.n1280 VSS.t1149 30.462
R2770 VSS.n1280 VSS.t1147 30.462
R2771 VSS.n1281 VSS.t1151 30.462
R2772 VSS.n1261 VSS.t830 30.462
R2773 VSS.n1260 VSS.t1128 30.462
R2774 VSS.n1260 VSS.t836 30.462
R2775 VSS.n1263 VSS.t621 30.462
R2776 VSS.n1263 VSS.t625 30.462
R2777 VSS.n1264 VSS.t623 30.462
R2778 VSS.n1252 VSS.t912 30.462
R2779 VSS.n1251 VSS.t388 30.462
R2780 VSS.n1251 VSS.t873 30.462
R2781 VSS.n1254 VSS.t1197 30.462
R2782 VSS.n1254 VSS.t1550 30.462
R2783 VSS.n1255 VSS.t1199 30.462
R2784 VSS.n71 VSS.t315 30.462
R2785 VSS.n70 VSS.t787 30.462
R2786 VSS.n70 VSS.t789 30.462
R2787 VSS.n73 VSS.t1057 30.462
R2788 VSS.n73 VSS.t1059 30.462
R2789 VSS.n74 VSS.t1061 30.462
R2790 VSS.n68 VSS.t1282 30.462
R2791 VSS.n67 VSS.t1276 30.462
R2792 VSS.n67 VSS.t1278 30.462
R2793 VSS.n1681 VSS.t1405 30.462
R2794 VSS.n1681 VSS.t1407 30.462
R2795 VSS.n1682 VSS.t1409 30.462
R2796 VSS.n41 VSS.t110 30.462
R2797 VSS.n40 VSS.t112 30.462
R2798 VSS.n40 VSS.t114 30.462
R2799 VSS.n43 VSS.t1201 30.462
R2800 VSS.n43 VSS.t1203 30.462
R2801 VSS.n44 VSS.t1205 30.462
R2802 VSS.n38 VSS.t344 30.462
R2803 VSS.n37 VSS.t346 30.462
R2804 VSS.n37 VSS.t348 30.462
R2805 VSS.n1701 VSS.t1831 30.462
R2806 VSS.n1701 VSS.t1833 30.462
R2807 VSS.n1702 VSS.t463 30.462
R2808 VSS.n14 VSS.t1166 30.462
R2809 VSS.n13 VSS.t1164 30.462
R2810 VSS.n13 VSS.t1168 30.462
R2811 VSS.n16 VSS.t751 30.462
R2812 VSS.n16 VSS.t755 30.462
R2813 VSS.n17 VSS.t753 30.462
R2814 VSS.n11 VSS.t97 30.462
R2815 VSS.n10 VSS.t100 30.462
R2816 VSS.n10 VSS.t1218 30.462
R2817 VSS.n1721 VSS.t1538 30.462
R2818 VSS.n1721 VSS.t1087 30.462
R2819 VSS.n1722 VSS.t1089 30.462
R2820 VSS.n289 VSS.t636 30.462
R2821 VSS.n288 VSS.t638 30.462
R2822 VSS.n288 VSS.t700 30.462
R2823 VSS.n291 VSS.t140 30.462
R2824 VSS.n291 VSS.t142 30.462
R2825 VSS.n292 VSS.t320 30.462
R2826 VSS.n308 VSS.t991 30.462
R2827 VSS.n297 VSS.t981 30.462
R2828 VSS.n297 VSS.t1029 30.462
R2829 VSS.n311 VSS.t144 30.462
R2830 VSS.n311 VSS.t146 30.462
R2831 VSS.n312 VSS.t148 30.462
R2832 VSS.n389 VSS.t1945 30.462
R2833 VSS.n388 VSS.t1894 30.462
R2834 VSS.n388 VSS.t1888 30.462
R2835 VSS.n77 VSS.t1420 30.462
R2836 VSS.n77 VSS.t1422 30.462
R2837 VSS.n78 VSS.t1424 30.462
R2838 VSS.n394 VSS.t1870 30.462
R2839 VSS.n393 VSS.t1872 30.462
R2840 VSS.n393 VSS.t1866 30.462
R2841 VSS.n62 VSS.t660 30.462
R2842 VSS.n62 VSS.t662 30.462
R2843 VSS.n63 VSS.t664 30.462
R2844 VSS.n399 VSS.t12 30.462
R2845 VSS.n398 VSS.t5 30.462
R2846 VSS.n398 VSS.t7 30.462
R2847 VSS.n47 VSS.t1508 30.462
R2848 VSS.n47 VSS.t1510 30.462
R2849 VSS.n48 VSS.t1512 30.462
R2850 VSS.n404 VSS.t1680 30.462
R2851 VSS.n403 VSS.t1682 30.462
R2852 VSS.n403 VSS.t1684 30.462
R2853 VSS.n33 VSS.t30 30.462
R2854 VSS.n33 VSS.t26 30.462
R2855 VSS.n34 VSS.t28 30.462
R2856 VSS.n409 VSS.t47 30.462
R2857 VSS.n408 VSS.t45 30.462
R2858 VSS.n408 VSS.t49 30.462
R2859 VSS.n20 VSS.t1659 30.462
R2860 VSS.n20 VSS.t1663 30.462
R2861 VSS.n21 VSS.t1661 30.462
R2862 VSS.n414 VSS.t1931 30.462
R2863 VSS.n413 VSS.t1933 30.462
R2864 VSS.n413 VSS.t1935 30.462
R2865 VSS.n1 VSS.t1232 30.462
R2866 VSS.n1 VSS.t1234 30.462
R2867 VSS.n2 VSS.t1236 30.462
R2868 VSS.n419 VSS.t1479 30.462
R2869 VSS.n418 VSS.t1481 30.462
R2870 VSS.n418 VSS.t1485 30.462
R2871 VSS.n421 VSS.t666 30.462
R2872 VSS.n421 VSS.t531 30.462
R2873 VSS.n422 VSS.t533 30.462
R2874 VSS.n438 VSS.t1000 30.462
R2875 VSS.n427 VSS.t994 30.462
R2876 VSS.n427 VSS.t986 30.462
R2877 VSS.n441 VSS.t602 30.462
R2878 VSS.n441 VSS.t847 30.462
R2879 VSS.n442 VSS.t947 30.462
R2880 VSS.n82 VSS.t1527 30.462
R2881 VSS.n81 VSS.t1533 30.462
R2882 VSS.n81 VSS.t1531 30.462
R2883 VSS.n1658 VSS.t1230 30.462
R2884 VSS.n1658 VSS.t1228 30.462
R2885 VSS.n1659 VSS.t392 30.462
R2886 VSS.n56 VSS.t469 30.462
R2887 VSS.n55 VSS.t471 30.462
R2888 VSS.n55 VSS.t467 30.462
R2889 VSS.n58 VSS.t1193 30.462
R2890 VSS.n58 VSS.t1340 30.462
R2891 VSS.n59 VSS.t1342 30.462
R2892 VSS.n53 VSS.t1243 30.462
R2893 VSS.n52 VSS.t1241 30.462
R2894 VSS.n52 VSS.t1239 30.462
R2895 VSS.n1691 VSS.t1415 30.462
R2896 VSS.n1691 VSS.t1318 30.462
R2897 VSS.n1692 VSS.t1316 30.462
R2898 VSS.n28 VSS.t422 30.462
R2899 VSS.n27 VSS.t420 30.462
R2900 VSS.n27 VSS.t418 30.462
R2901 VSS.n30 VSS.t82 30.462
R2902 VSS.n30 VSS.t80 30.462
R2903 VSS.n31 VSS.t406 30.462
R2904 VSS.n25 VSS.t1815 30.462
R2905 VSS.n24 VSS.t1811 30.462
R2906 VSS.n24 VSS.t1809 30.462
R2907 VSS.n1711 VSS.t828 30.462
R2908 VSS.n1711 VSS.t824 30.462
R2909 VSS.n1712 VSS.t826 30.462
R2910 VSS.n452 VSS.t1053 30.462
R2911 VSS.n451 VSS.t1376 30.462
R2912 VSS.n451 VSS.t1374 30.462
R2913 VSS.n6 VSS.t1939 30.462
R2914 VSS.n6 VSS.t1943 30.462
R2915 VSS.n7 VSS.t1941 30.462
R2916 VSS.n457 VSS.t1623 30.462
R2917 VSS.n456 VSS.t1621 30.462
R2918 VSS.n456 VSS.t1619 30.462
R2919 VSS.n459 VSS.t1036 30.462
R2920 VSS.n459 VSS.t1040 30.462
R2921 VSS.n460 VSS.t1038 30.462
R2922 VSS.n476 VSS.t1023 30.462
R2923 VSS.n465 VSS.t1026 30.462
R2924 VSS.n465 VSS.t1032 30.462
R2925 VSS.n479 VSS.t450 30.462
R2926 VSS.n479 VSS.t452 30.462
R2927 VSS.n480 VSS.t448 30.462
R2928 VSS.n1312 VSS.t458 30.462
R2929 VSS.n1311 VSS.t456 30.462
R2930 VSS.n1311 VSS.t460 30.462
R2931 VSS.n1314 VSS.t931 30.462
R2932 VSS.n1314 VSS.t897 30.462
R2933 VSS.n1315 VSS.t875 30.462
R2934 VSS.n601 VSS.t1521 30.462
R2935 VSS.n600 VSS.t1523 30.462
R2936 VSS.n600 VSS.t1519 30.462
R2937 VSS.n1214 VSS.t23 30.462
R2938 VSS.n1214 VSS.t21 30.462
R2939 VSS.n1215 VSS.t1855 30.462
R2940 VSS.n1307 VSS.t168 30.1842
R2941 VSS.t226 VSS.n1611 30.1689
R2942 VSS.t90 VSS.t724 28.9739
R2943 VSS.n300 VSS.n298 28.3986
R2944 VSS.n430 VSS.n428 28.3986
R2945 VSS.n468 VSS.n466 28.3986
R2946 VSS.t1110 VSS.n1602 28.1311
R2947 VSS.t1650 VSS.n1593 28.1311
R2948 VSS.t443 VSS.n1584 28.1311
R2949 VSS.t1631 VSS.n1574 28.1311
R2950 VSS.n1631 VSS.t685 28.1311
R2951 VSS.n1401 VSS.n1400 28.0856
R2952 VSS.n545 VSS.n121 28.0856
R2953 VSS.n1625 VSS.t507 26.7697
R2954 VSS.n119 VSS.t1135 26.7697
R2955 VSS.n1617 VSS.t1179 26.7697
R2956 VSS.n1614 VSS.t1906 26.7697
R2957 VSS.n1607 VSS.t1288 26.7697
R2958 VSS.n1604 VSS.t256 26.7697
R2959 VSS.n1598 VSS.t1093 26.7697
R2960 VSS.n1595 VSS.t1841 26.7697
R2961 VSS.n1589 VSS.t1652 26.7697
R2962 VSS.n1586 VSS.t815 26.7697
R2963 VSS.n1580 VSS.t1800 26.7697
R2964 VSS.n1577 VSS.t184 26.7697
R2965 VSS.n1570 VSS.t1636 26.7697
R2966 VSS.n1567 VSS.t1393 26.7697
R2967 VSS.n115 VSS.t689 26.7697
R2968 VSS.n112 VSS.t1580 26.7697
R2969 VSS.n577 VSS.t582 26.7697
R2970 VSS.n580 VSS.t1578 26.7697
R2971 VSS.n593 VSS.t489 26.7697
R2972 VSS.n596 VSS.t378 26.7697
R2973 VSS.n1286 VSS.t1190 26.7697
R2974 VSS.n1289 VSS.t927 26.7697
R2975 VSS.n542 VSS.t222 26.7697
R2976 VSS.n569 VSS.t929 26.7697
R2977 VSS.n533 VSS.t1106 26.7697
R2978 VSS.n537 VSS.t871 26.7697
R2979 VSS.n264 VSS.t1648 26.7697
R2980 VSS.n528 VSS.t918 26.7697
R2981 VSS.n248 VSS.t1798 26.7697
R2982 VSS.n259 VSS.t923 26.7697
R2983 VSS.n242 VSS.t1640 26.7697
R2984 VSS.n245 VSS.t376 26.7697
R2985 VSS.n97 VSS.t584 26.7697
R2986 VSS.n100 VSS.t895 26.7697
R2987 VSS.n1357 VSS.t1572 26.7697
R2988 VSS.n1360 VSS.t1670 26.7697
R2989 VSS.n1369 VSS.t959 26.7697
R2990 VSS.n1372 VSS.t1604 26.7697
R2991 VSS.n232 VSS.t1389 26.7697
R2992 VSS.n1380 VSS.t1493 26.7697
R2993 VSS.n235 VSS.t568 26.7697
R2994 VSS.n238 VSS.t413 26.7697
R2995 VSS.n173 VSS.t176 26.7697
R2996 VSS.n176 VSS.t1430 26.7697
R2997 VSS.n170 VSS.t1351 26.7697
R2998 VSS.n1470 VSS.t1772 26.7697
R2999 VSS.n271 VSS.t1122 26.7697
R3000 VSS.n515 VSS.t706 26.7697
R3001 VSS.n504 VSS.t1783 26.7697
R3002 VSS.n507 VSS.t137 26.7697
R3003 VSS.n283 VSS.t1851 26.7697
R3004 VSS.n286 VSS.t299 26.7697
R3005 VSS.n274 VSS.t864 26.7697
R3006 VSS.n277 VSS.t2026 26.7697
R3007 VSS.n130 VSS.t254 26.7697
R3008 VSS.n133 VSS.t161 26.7697
R3009 VSS.n127 VSS.t39 26.7697
R3010 VSS.n1528 VSS.t1249 26.7697
R3011 VSS.n1270 VSS.t1896 26.7697
R3012 VSS.n1273 VSS.t1863 26.7697
R3013 VSS.n1249 VSS.t402 26.7697
R3014 VSS.n1281 VSS.t368 26.7697
R3015 VSS.n1261 VSS.t834 26.7697
R3016 VSS.n1264 VSS.t1083 26.7697
R3017 VSS.n1252 VSS.t879 26.7697
R3018 VSS.n1255 VSS.t1144 26.7697
R3019 VSS.n71 VSS.t313 26.7697
R3020 VSS.n74 VSS.t1016 26.7697
R3021 VSS.n68 VSS.t1280 26.7697
R3022 VSS.n1682 VSS.t236 26.7697
R3023 VSS.n41 VSS.t117 26.7697
R3024 VSS.n44 VSS.t1447 26.7697
R3025 VSS.n38 VSS.t350 26.7697
R3026 VSS.n1702 VSS.t213 26.7697
R3027 VSS.n14 VSS.t1170 26.7697
R3028 VSS.n17 VSS.t656 26.7697
R3029 VSS.n11 VSS.t95 26.7697
R3030 VSS.n1722 VSS.t1880 26.7697
R3031 VSS.n289 VSS.t698 26.7697
R3032 VSS.n292 VSS.t134 26.7697
R3033 VSS.n308 VSS.t1006 26.7697
R3034 VSS.n312 VSS.t1070 26.7697
R3035 VSS.n389 VSS.t1916 26.7697
R3036 VSS.n78 VSS.t1335 26.7697
R3037 VSS.n394 VSS.t1868 26.7697
R3038 VSS.n63 VSS.t522 26.7697
R3039 VSS.n399 VSS.t9 26.7697
R3040 VSS.n48 VSS.t1817 26.7697
R3041 VSS.n404 VSS.t1686 26.7697
R3042 VSS.n34 VSS.t326 26.7697
R3043 VSS.n409 VSS.t51 26.7697
R3044 VSS.n21 VSS.t1502 26.7697
R3045 VSS.n414 VSS.t1929 26.7697
R3046 VSS.n2 VSS.t1764 26.7697
R3047 VSS.n419 VSS.t1483 26.7697
R3048 VSS.n422 VSS.t1262 26.7697
R3049 VSS.n438 VSS.t1009 26.7697
R3050 VSS.n442 VSS.t293 26.7697
R3051 VSS.n82 VSS.t1529 26.7697
R3052 VSS.n1659 VSS.t1829 26.7697
R3053 VSS.n56 VSS.t473 26.7697
R3054 VSS.n59 VSS.t1675 26.7697
R3055 VSS.n53 VSS.t1245 26.7697
R3056 VSS.n1692 VSS.t74 26.7697
R3057 VSS.n28 VSS.t424 26.7697
R3058 VSS.n31 VSS.t633 26.7697
R3059 VSS.n25 VSS.t1813 26.7697
R3060 VSS.n1712 VSS.t970 26.7697
R3061 VSS.n452 VSS.t1372 26.7697
R3062 VSS.n7 VSS.t1044 26.7697
R3063 VSS.n457 VSS.t1617 26.7697
R3064 VSS.n460 VSS.t966 26.7697
R3065 VSS.n476 VSS.t1013 26.7697
R3066 VSS.n480 VSS.t1561 26.7697
R3067 VSS.n1312 VSS.t514 26.7697
R3068 VSS.n1315 VSS.t920 26.7697
R3069 VSS.n601 VSS.t1525 26.7697
R3070 VSS.n1215 VSS.t1591 26.7697
R3071 VSS.t539 VSS.t1468 26.3117
R3072 VSS.t756 VSS.t1346 26.3117
R3073 VSS.n328 VSS.t1123 25.1673
R3074 VSS.n329 VSS.t290 25.1673
R3075 VSS.n330 VSS.t1263 25.1673
R3076 VSS.n332 VSS.t1687 25.1673
R3077 VSS.n333 VSS.t1761 25.1673
R3078 VSS.n335 VSS.t52 25.1673
R3079 VSS.n336 VSS.t1822 25.1673
R3080 VSS.n337 VSS.t321 25.1673
R3081 VSS.n339 VSS.t10 25.1673
R3082 VSS.n341 VSS.t67 25.1673
R3083 VSS.n372 VSS.t1138 25.1673
R3084 VSS.n374 VSS.t1336 25.1673
R3085 VSS.n1518 VSS.t101 25.1434
R3086 VSS.t988 VSS.n1517 25.1434
R3087 VSS.n1509 VSS.t130 25.1434
R3088 VSS.t351 VSS.n1508 25.1434
R3089 VSS.t98 VSS.n1506 25.1434
R3090 VSS.n165 VSS.t657 25.1434
R3091 VSS.n1478 VSS.t53 25.1434
R3092 VSS.t215 VSS.n1477 25.1434
R3093 VSS.n344 VSS.t115 25.1434
R3094 VSS.n346 VSS.t352 25.1434
R3095 VSS.n368 VSS.t238 25.1434
R3096 VSS.t790 VSS.n367 25.1434
R3097 VSS.n1454 VSS.t509 24.9768
R3098 VSS.n1449 VSS.t502 24.9768
R3099 VSS.t1094 VSS.t515 24.2385
R3100 VSS.n1026 VSS.t1727 21.7959
R3101 VSS.n1024 VSS.t1747 21.7959
R3102 VSS.n1036 VSS.t1713 21.7959
R3103 VSS.n1020 VSS.t18 21.7959
R3104 VSS.n1042 VSS.t1723 21.7959
R3105 VSS.n990 VSS.t1746 21.7959
R3106 VSS.n988 VSS.t1705 21.7959
R3107 VSS.n1000 VSS.t1725 21.7959
R3108 VSS.n984 VSS.t1283 21.7959
R3109 VSS.n1006 VSS.t1741 21.7959
R3110 VSS.n1169 VSS.t1730 21.7959
R3111 VSS.n1166 VSS.t1748 21.7959
R3112 VSS.n1160 VSS.t1716 21.7959
R3113 VSS.n1157 VSS.t1724 21.7959
R3114 VSS.n627 VSS.t198 21.7959
R3115 VSS.n956 VSS.t1703 21.7959
R3116 VSS.n954 VSS.t1718 21.7959
R3117 VSS.n966 VSS.t1740 21.7959
R3118 VSS.n950 VSS.t105 21.7959
R3119 VSS.n972 VSS.t1753 21.7959
R3120 VSS.n1060 VSS.t1744 21.7959
R3121 VSS.n1058 VSS.t1704 21.7959
R3122 VSS.n1070 VSS.t1722 21.7959
R3123 VSS.n1054 VSS.t1641 21.7959
R3124 VSS.n1076 VSS.t1738 21.7959
R3125 VSS.n922 VSS.t1719 21.7959
R3126 VSS.n920 VSS.t1731 21.7959
R3127 VSS.n932 VSS.t1700 21.7959
R3128 VSS.n916 VSS.t1542 21.7959
R3129 VSS.n938 VSS.t1712 21.7959
R3130 VSS.n1102 VSS.t1721 21.7959
R3131 VSS.n1099 VSS.t1752 21.7959
R3132 VSS.n1093 VSS.t1742 21.7959
R3133 VSS.n738 VSS.t668 21.7959
R3134 VSS.n734 VSS.t1737 21.7959
R3135 VSS.n888 VSS.t1720 21.7959
R3136 VSS.n886 VSS.t1743 21.7959
R3137 VSS.n898 VSS.t1739 21.7959
R3138 VSS.n882 VSS.t652 21.7959
R3139 VSS.n904 VSS.t1726 21.7959
R3140 VSS.n1123 VSS.t1717 21.7959
R3141 VSS.n1117 VSS.t1751 21.7959
R3142 VSS.n863 VSS.t737 21.7959
R3143 VSS.n719 VSS.t1736 21.7959
R3144 VSS.n1040 VSS.t1459 21.7687
R3145 VSS.n1025 VSS.t1457 21.7687
R3146 VSS.n1034 VSS.t1461 21.7687
R3147 VSS.n1038 VSS.t1463 21.7687
R3148 VSS.n1022 VSS.t480 21.7687
R3149 VSS.n1004 VSS.t741 21.7687
R3150 VSS.n989 VSS.t739 21.7687
R3151 VSS.n998 VSS.t743 21.7687
R3152 VSS.n1002 VSS.t745 21.7687
R3153 VSS.n986 VSS.t78 21.7687
R3154 VSS.n1179 VSS.t427 21.7687
R3155 VSS.n1168 VSS.t207 21.7687
R3156 VSS.n1164 VSS.t203 21.7687
R3157 VSS.n1162 VSS.t205 21.7687
R3158 VSS.n1158 VSS.t201 21.7687
R3159 VSS.n970 VSS.t680 21.7687
R3160 VSS.n955 VSS.t678 21.7687
R3161 VSS.n964 VSS.t682 21.7687
R3162 VSS.n968 VSS.t676 21.7687
R3163 VSS.n952 VSS.t1568 21.7687
R3164 VSS.n1074 VSS.t59 21.7687
R3165 VSS.n1059 VSS.t57 21.7687
R3166 VSS.n1068 VSS.t61 21.7687
R3167 VSS.n1072 VSS.t55 21.7687
R3168 VSS.n1056 VSS.t398 21.7687
R3169 VSS.n936 VSS.t1379 21.7687
R3170 VSS.n921 VSS.t1385 21.7687
R3171 VSS.n930 VSS.t1381 21.7687
R3172 VSS.n934 VSS.t1383 21.7687
R3173 VSS.n918 VSS.t723 21.7687
R3174 VSS.n1091 VSS.t1475 21.7687
R3175 VSS.n1101 VSS.t1477 21.7687
R3176 VSS.n1097 VSS.t1473 21.7687
R3177 VSS.n1095 VSS.t1471 21.7687
R3178 VSS.n736 VSS.t1949 21.7687
R3179 VSS.n902 VSS.t854 21.7687
R3180 VSS.n887 VSS.t856 21.7687
R3181 VSS.n896 VSS.t852 21.7687
R3182 VSS.n900 VSS.t850 21.7687
R3183 VSS.n884 VSS.t1536 21.7687
R3184 VSS.n1115 VSS.t1438 21.7687
R3185 VSS.n1133 VSS.t1442 21.7687
R3186 VSS.n1148 VSS.t1745 21.7687
R3187 VSS.n1121 VSS.t1436 21.7687
R3188 VSS.n1119 VSS.t1440 21.7687
R3189 VSS.n865 VSS.t619 21.7687
R3190 VSS.n183 VSS.n182 20.508
R3191 VSS.n181 VSS.n180 20.337
R3192 VSS.t1799 VSS.n1575 20.1812
R3193 VSS.n179 VSS.n178 20.1096
R3194 VSS.n1498 VSS.n51 20.0737
R3195 VSS.n1495 VSS.n51 20.0088
R3196 VSS.n858 VSS.t1566 19.8005
R3197 VSS.n858 VSS.t792 19.8005
R3198 VSS.n798 VSS.t1469 19.8005
R3199 VSS.n798 VSS.t757 19.8005
R3200 VSS.n1493 VSS.n110 19.1083
R3201 VSS.t1284 VSS.n200 18.462
R3202 VSS.t1292 VSS.n376 18.462
R3203 VSS.n357 VSS.t1183 18.4491
R3204 VSS.n1434 VSS.t1173 18.4491
R3205 VSS.n1672 VSS.n1671 17.8661
R3206 VSS.n1673 VSS.n1672 17.8661
R3207 VSS.n1183 VSS.n1182 17.7999
R3208 VSS.n348 VSS.t209 17.6005
R3209 VSS.n1438 VSS.t557 17.6005
R3210 VSS.t407 VSS.n326 17.6005
R3211 VSS.n319 VSS.t535 17.6005
R3212 VSS.n202 VSS.t1306 17.6005
R3213 VSS.t353 VSS.n1422 17.6005
R3214 VSS.n1674 VSS.n1673 17.1217
R3215 VSS.t271 VSS.t1565 17.1052
R3216 VSS.t1219 VSS.t791 17.1052
R3217 VSS.n1502 VSS.t70 16.848
R3218 VSS.n91 VSS.n90 16.7948
R3219 VSS.n1649 VSS.n1648 16.7775
R3220 VSS.n1645 VSS.n1644 16.7725
R3221 VSS.n1651 VSS.n1650 16.7688
R3222 VSS.n1395 VSS.n1394 16.7676
R3223 VSS.n1393 VSS.n1392 16.7651
R3224 VSS.n95 VSS.n94 16.7205
R3225 VSS.n1390 VSS.n92 16.7156
R3226 VSS.n220 VSS.n218 16.6847
R3227 VSS.n1484 VSS.n1483 16.6847
R3228 VSS.n547 VSS.n544 16.6847
R3229 VSS.n229 VSS.n227 16.6735
R3230 VSS.n1488 VSS.n1487 16.6735
R3231 VSS.n551 VSS.n550 16.6735
R3232 VSS.n216 VSS 16.6585
R3233 VSS.n1482 VSS 16.6585
R3234 VSS.n565 VSS 16.6585
R3235 VSS.n220 VSS 16.6501
R3236 VSS.n1483 VSS 16.6501
R3237 VSS VSS.n544 16.6501
R3238 VSS.n222 VSS 16.6473
R3239 VSS.n224 VSS 16.6473
R3240 VSS.n161 VSS 16.6473
R3241 VSS VSS.n1490 16.6473
R3242 VSS.n557 VSS 16.6473
R3243 VSS VSS.n558 16.6473
R3244 VSS.n226 VSS 16.6431
R3245 VSS.n1489 VSS 16.6431
R3246 VSS VSS.n546 16.6431
R3247 VSS.n229 VSS 16.6417
R3248 VSS.n1488 VSS 16.6417
R3249 VSS VSS.n551 16.6417
R3250 VSS.n253 VSS 16.5096
R3251 VSS.n251 VSS 16.496
R3252 VSS.n1305 VSS.n1304 16.4945
R3253 VSS.n1304 VSS.n1244 16.4945
R3254 VSS.n1304 VSS.n1303 16.4945
R3255 VSS.n1304 VSS.n1245 16.4945
R3256 VSS.n1304 VSS.n1302 16.4945
R3257 VSS.n1304 VSS.n1246 16.4945
R3258 VSS.n1304 VSS.n1301 16.4945
R3259 VSS.n1304 VSS.n1247 16.4945
R3260 VSS.n840 VSS.n742 16.4945
R3261 VSS.n1558 VSS.n1538 16.4943
R3262 VSS.n1556 VSS.n1538 16.4943
R3263 VSS.n1554 VSS.n1538 16.4943
R3264 VSS.n1552 VSS.n1538 16.4943
R3265 VSS.n1550 VSS.n1538 16.4943
R3266 VSS.n1548 VSS.n1538 16.4943
R3267 VSS.n1546 VSS.n1538 16.4943
R3268 VSS.n1563 VSS.n1538 16.4943
R3269 VSS.n255 VSS 16.479
R3270 VSS.n1304 VSS 16.4313
R3271 VSS VSS.n1538 16.4312
R3272 VSS.n142 VSS.n0 16.2301
R3273 VSS.n1533 VSS.n1532 16.2301
R3274 VSS.n1300 VSS.n1299 16.2301
R3275 VSS.n1326 VSS.n1325 16.2301
R3276 VSS.n207 VSS.n61 16.2301
R3277 VSS.n340 VSS.n61 16.2301
R3278 VSS.n1480 VSS.n162 16.2301
R3279 VSS.n331 VSS.n0 16.2301
R3280 VSS.n1520 VSS.n136 16.2301
R3281 VSS.n345 VSS.n61 16.2301
R3282 VSS.n1480 VSS.n1479 16.2301
R3283 VSS.n1507 VSS.n0 16.2301
R3284 VSS.n1520 VSS.n1519 16.2301
R3285 VSS.n1385 VSS.n1384 16.2301
R3286 VSS.n1345 VSS.n66 16.2301
R3287 VSS.n268 VSS.n166 16.2301
R3288 VSS.n494 VSS.n5 16.2301
R3289 VSS.n489 VSS.n139 16.2301
R3290 VSS.n1480 VSS.n163 16.2301
R3291 VSS.n1520 VSS.n138 16.2301
R3292 VSS.n1515 VSS.n1514 16.2064
R3293 VSS.n447 VSS.n125 16.2064
R3294 VSS.n1296 VSS.n1295 16.2064
R3295 VSS.n1322 VSS.n1321 16.2064
R3296 VSS.n370 VSS.n342 16.2064
R3297 VSS.n371 VSS.n370 16.2064
R3298 VSS.n1475 VSS.n167 16.2064
R3299 VSS.n1504 VSS.n147 16.2064
R3300 VSS.n1515 VSS.n140 16.2064
R3301 VSS.n370 VSS.n369 16.2064
R3302 VSS.n1476 VSS.n1475 16.2064
R3303 VSS.n1505 VSS.n1504 16.2064
R3304 VSS.n1516 VSS.n1515 16.2064
R3305 VSS.n1389 VSS.n1388 16.2064
R3306 VSS.n1351 VSS.n1350 16.2064
R3307 VSS.n266 VSS.n168 16.2064
R3308 VSS.n524 VSS.n523 16.2064
R3309 VSS.n492 VSS.n491 16.2064
R3310 VSS.n1475 VSS.n1474 16.2064
R3311 VSS.n1504 VSS.n1503 16.2064
R3312 VSS.n845 VSS 16.2013
R3313 VSS.n1629 VSS.n1628 16.2005
R3314 VSS.n1572 VSS.n117 16.2005
R3315 VSS.n1582 VSS.n117 16.2005
R3316 VSS.n1591 VSS.n117 16.2005
R3317 VSS.n1600 VSS.n117 16.2005
R3318 VSS.n1609 VSS.n117 16.2005
R3319 VSS.n1619 VSS.n117 16.2005
R3320 VSS.n1628 VSS.n1627 16.2005
R3321 VSS.n482 VSS.n137 16.2005
R3322 VSS.n462 VSS.n146 16.2005
R3323 VSS.n1725 VSS.n9 16.2005
R3324 VSS.n1715 VSS.n1714 16.2005
R3325 VSS.n1706 VSS.n1705 16.2005
R3326 VSS.n1695 VSS.n1694 16.2005
R3327 VSS.n1686 VSS.n1685 16.2005
R3328 VSS.n1662 VSS.n1661 16.2005
R3329 VSS.n444 VSS.n137 16.2005
R3330 VSS.n424 VSS.n146 16.2005
R3331 VSS.n1725 VSS.n4 16.2005
R3332 VSS.n1715 VSS.n23 16.2005
R3333 VSS.n1705 VSS.n36 16.2005
R3334 VSS.n1695 VSS.n50 16.2005
R3335 VSS.n1685 VSS.n65 16.2005
R3336 VSS.n1662 VSS.n80 16.2005
R3337 VSS.n314 VSS.n137 16.2005
R3338 VSS.n294 VSS.n146 16.2005
R3339 VSS.n1725 VSS.n1724 16.2005
R3340 VSS.n1716 VSS.n1715 16.2005
R3341 VSS.n1705 VSS.n1704 16.2005
R3342 VSS.n1696 VSS.n1695 16.2005
R3343 VSS.n1685 VSS.n1684 16.2005
R3344 VSS.n1663 VSS.n1662 16.2005
R3345 VSS.n1257 VSS.n582 16.2005
R3346 VSS.n1266 VSS.n1227 16.2005
R3347 VSS.n1284 VSS.n1283 16.2005
R3348 VSS.n1275 VSS.n123 16.2005
R3349 VSS.n1531 VSS.n1530 16.2005
R3350 VSS.n1522 VSS.n1521 16.2005
R3351 VSS.n279 VSS.n141 16.2005
R3352 VSS.n500 VSS.n499 16.2005
R3353 VSS.n509 VSS.n148 16.2005
R3354 VSS.n518 VSS.n517 16.2005
R3355 VSS.n1473 VSS.n1472 16.2005
R3356 VSS.n1464 VSS.n1463 16.2005
R3357 VSS.n1353 VSS.n1352 16.2005
R3358 VSS.n1383 VSS.n1382 16.2005
R3359 VSS.n1374 VSS.n193 16.2005
R3360 VSS.n1365 VSS.n1364 16.2005
R3361 VSS.n1320 VSS.n1319 16.2005
R3362 VSS.n1294 VSS.n1293 16.2005
R3363 VSS.n567 VSS.n566 16.2005
R3364 VSS.n535 VSS.n144 16.2005
R3365 VSS.n526 VSS.n525 16.2005
R3366 VSS.n257 VSS.n256 16.2005
R3367 VSS.n1344 VSS.n1343 16.2005
R3368 VSS.n1643 VSS.n1642 16.2005
R3369 VSS.n1221 VSS.n1220 16.2005
R3370 VSS.n1328 VSS.n1327 16.2005
R3371 VSS.n673 VSS.n672 15.8647
R3372 VSS.n669 VSS.n668 15.8647
R3373 VSS.n681 VSS.n680 15.8647
R3374 VSS.n662 VSS.n661 15.8647
R3375 VSS.n689 VSS.n688 15.8647
R3376 VSS.n655 VSS.n654 15.8647
R3377 VSS.n697 VSS.n696 15.8647
R3378 VSS.n648 VSS.n647 15.8647
R3379 VSS.n705 VSS.n704 15.8647
R3380 VSS.n675 VSS.n674 15.8449
R3381 VSS.n670 VSS.n667 15.8449
R3382 VSS.n683 VSS.n682 15.8449
R3383 VSS.n663 VSS.n660 15.8449
R3384 VSS.n691 VSS.n690 15.8449
R3385 VSS.n656 VSS.n653 15.8449
R3386 VSS.n699 VSS.n698 15.8449
R3387 VSS.n649 VSS.n646 15.8449
R3388 VSS.n707 VSS.n706 15.8449
R3389 VSS.n679 VSS.n678 15.8355
R3390 VSS.n664 VSS.n642 15.8355
R3391 VSS.n687 VSS.n686 15.8355
R3392 VSS.n657 VSS.n641 15.8355
R3393 VSS.n695 VSS.n694 15.8355
R3394 VSS.n650 VSS.n640 15.8355
R3395 VSS.n703 VSS.n702 15.8355
R3396 VSS.n643 VSS.n639 15.8355
R3397 VSS.n711 VSS.n710 15.8355
R3398 VSS.n1130 VSS.n1129 15.6691
R3399 VSS VSS.n1675 15.6329
R3400 VSS.n1138 VSS.n1137 15.5706
R3401 VSS.n852 VSS.t756 15.3487
R3402 VSS.t1848 VSS.t578 14.8905
R3403 VSS.n1676 VSS.n1669 13.6732
R3404 VSS.n1145 VSS.n1127 13.5081
R3405 VSS.t75 VSS.n1458 12.4887
R3406 VSS.t525 VSS.n1453 12.4887
R3407 VSS.n1135 VSS.n1132 11.6937
R3408 VSS.n852 VSS.t1468 10.9635
R3409 VSS.n1669 VSS.n1668 10.8165
R3410 VSS.n437 VSS.n436 10.6145
R3411 VSS.n475 VSS.n474 10.587
R3412 VSS.n307 VSS.n306 10.5541
R3413 VSS.n1141 VSS.n1140 10.4475
R3414 VSS.t791 VSS.n861 9.97823
R3415 VSS.n604 VSS.n599 9.59666
R3416 VSS.n1346 VSS.t777 9.56572
R3417 VSS.n1349 VSS.t552 9.56572
R3418 VSS.t1400 VSS.n1348 9.56572
R3419 VSS.n1386 VSS.t951 9.56572
R3420 VSS.n1387 VSS.t960 9.56572
R3421 VSS.t1575 VSS.n103 9.56572
R3422 VSS.n1146 VSS.n1145 9.48445
R3423 VSS.n1135 VSS.n1134 9.46423
R3424 VSS.n217 VSS.n213 9.3622
R3425 VSS.t1607 VSS.t771 9.3622
R3426 VSS.n1486 VSS.n1485 9.3622
R3427 VSS.t394 VSS.t273 9.3622
R3428 VSS.n549 VSS.n548 9.3622
R3429 VSS.t692 VSS.t1627 9.3622
R3430 VSS.t1920 VSS.n384 9.23127
R3431 VSS.n377 VSS.t1076 9.23127
R3432 VSS.n364 VSS.n363 9.22482
R3433 VSS.t1300 VSS.n361 9.22482
R3434 VSS.n1430 VSS.t1464 9.22482
R3435 VSS.n607 VSS.n599 9.0566
R3436 VSS.n1218 VSS.n1217 9.0005
R3437 VSS.n562 VSS.n561 8.8005
R3438 VSS.t252 VSS.t107 7.98961
R3439 VSS.n383 VSS.n382 7.96007
R3440 VSS.n347 VSS.n195 7.96007
R3441 VSS.n1457 VSS.n1456 7.95966
R3442 VSS.n205 VSS.n203 7.95956
R3443 VSS.n325 VSS.n324 7.95956
R3444 VSS.n360 VSS.n359 7.95945
R3445 VSS.n1445 VSS.n187 7.95811
R3446 VSS.n1407 VSS.n1405 7.9581
R3447 VSS.n1412 VSS.n1411 7.9105
R3448 VSS.n1421 VSS.n1420 7.9105
R3449 VSS.n379 VSS.n378 7.9105
R3450 VSS.n321 VSS.n320 7.9105
R3451 VSS.n1432 VSS.n1431 7.9105
R3452 VSS.n1452 VSS.n1451 7.9105
R3453 VSS.n192 VSS.n191 7.9105
R3454 VSS.n1440 VSS.n1439 7.9105
R3455 VSS.n1219 VSS.n1218 7.2005
R3456 VSS.n861 VSS.t1565 7.12745
R3457 VSS.n1224 VSS.t1085 6.39585
R3458 VSS.n490 VSS.t954 6.07645
R3459 VSS.n493 VSS.t860 6.07645
R3460 VSS.n496 VSS.t300 6.07645
R3461 VSS.t453 VSS.n495 6.07645
R3462 VSS.n522 VSS.t163 6.07645
R3463 VSS.t707 VSS.n521 6.07645
R3464 VSS.t952 VSS.n269 6.07645
R3465 VSS.t1356 VSS.n267 6.07645
R3466 VSS.n1460 VSS.t192 6.07645
R3467 VSS.n847 VSS.n844 5.26838
R3468 VSS.n306 VSS.n301 5.09176
R3469 VSS.n436 VSS.n431 5.09176
R3470 VSS.n474 VSS.n469 5.09176
R3471 VSS.n208 VSS.t483 4.84809
R3472 VSS.n209 VSS.t465 4.84809
R3473 VSS.n1403 VSS.t1534 4.84809
R3474 VSS.t1097 VSS.n86 4.84809
R3475 VSS.n1409 VSS.t1094 4.84809
R3476 VSS.n1297 VSS.n122 4.78896
R3477 VSS.n1653 VSS.n88 4.56009
R3478 VSS.n306 VSS.n305 4.19292
R3479 VSS.n436 VSS.n435 4.19292
R3480 VSS.n474 VSS.n473 4.19292
R3481 VSS.n1647 VSS.n1646 4.04016
R3482 VSS.t1171 VSS.t1289 4.04016
R3483 VSS.t251 VSS.t1907 4.04016
R3484 VSS.n449 VSS.n135 3.88674
R3485 VSS.n1537 VSS.n1536 3.88674
R3486 VSS.n1310 VSS.n1309 3.88674
R3487 VSS.n1402 VSS.n76 3.88674
R3488 VSS.n373 VSS.n76 3.88674
R3489 VSS.n338 VSS.n46 3.88674
R3490 VSS.n334 VSS.n19 3.88674
R3491 VSS.n1511 VSS.n145 3.88674
R3492 VSS.n366 VSS.n76 3.88674
R3493 VSS.n343 VSS.n46 3.88674
R3494 VSS.n164 VSS.n19 3.88674
R3495 VSS.n1511 VSS.n1510 3.88674
R3496 VSS.n1363 VSS.n1362 3.88674
R3497 VSS.n1347 VSS.n230 3.88674
R3498 VSS.n1462 VSS.n1461 3.88674
R3499 VSS.n520 VSS.n519 3.88674
R3500 VSS.n498 VSS.n497 3.88674
R3501 VSS.n149 VSS.n46 3.88674
R3502 VSS.n150 VSS.n19 3.88674
R3503 VSS.n1512 VSS.n1511 3.88674
R3504 VSS.n1420 VSS.n1419 3.55497
R3505 VSS.n379 VSS.n375 3.55497
R3506 VSS.n1440 VSS.n196 3.55487
R3507 VSS.n192 VSS.n188 3.55483
R3508 VSS.n321 VSS.n317 3.55476
R3509 VSS.n1433 VSS.n1432 3.55466
R3510 VSS.n1412 VSS.n1410 3.55391
R3511 VSS.n1451 VSS.n1450 3.55279
R3512 VSS.n1407 VSS.n1406 3.5055
R3513 VSS.n205 VSS.n204 3.5055
R3514 VSS.n382 VSS.n381 3.5055
R3515 VSS.n324 VSS.n323 3.5055
R3516 VSS.n359 VSS.n358 3.5055
R3517 VSS.n1456 VSS.n1455 3.5055
R3518 VSS.n1446 VSS.n1445 3.5055
R3519 VSS.n349 VSS.n195 3.5055
R3520 VSS.n802 VSS.n745 3.41065
R3521 VSS.n836 VSS.n747 3.41065
R3522 VSS.n812 VSS.n746 3.41065
R3523 VSS.n822 VSS.n748 3.41065
R3524 VSS.n875 VSS.n874 3.41065
R3525 VSS.n762 VSS.n743 3.41065
R3526 VSS.n788 VSS.n750 3.41065
R3527 VSS.n771 VSS.n744 3.41065
R3528 VSS.n780 VSS.n749 3.41065
R3529 VSS.n801 VSS.n800 3.4105
R3530 VSS.n806 VSS.n801 3.4105
R3531 VSS.n805 VSS.n802 3.4105
R3532 VSS.n835 VSS.n834 3.4105
R3533 VSS.n835 VSS.n833 3.4105
R3534 VSS.n837 VSS.n836 3.4105
R3535 VSS.n811 VSS.n810 3.4105
R3536 VSS.n816 VSS.n811 3.4105
R3537 VSS.n815 VSS.n812 3.4105
R3538 VSS.n821 VSS.n820 3.4105
R3539 VSS.n826 VSS.n821 3.4105
R3540 VSS.n825 VSS.n822 3.4105
R3541 VSS.n752 VSS.n751 3.4105
R3542 VSS.n874 VSS.n873 3.4105
R3543 VSS.n753 VSS.n752 3.4105
R3544 VSS.n770 VSS.n769 3.4105
R3545 VSS.n765 VSS.n762 3.4105
R3546 VSS.n769 VSS.n768 3.4105
R3547 VSS.n796 VSS.n795 3.4105
R3548 VSS.n791 VSS.n788 3.4105
R3549 VSS.n795 VSS.n794 3.4105
R3550 VSS.n779 VSS.n778 3.4105
R3551 VSS.n774 VSS.n771 3.4105
R3552 VSS.n778 VSS.n777 3.4105
R3553 VSS.n787 VSS.n786 3.4105
R3554 VSS.n786 VSS.n785 3.4105
R3555 VSS.n783 VSS.n780 3.4105
R3556 VSS.n644 VSS.t2020 3.34905
R3557 VSS.n645 VSS.t1980 3.34905
R3558 VSS.t1710 VSS.n590 3.34905
R3559 VSS.n665 VSS.t1995 3.26621
R3560 VSS.n666 VSS.t1978 3.26621
R3561 VSS.t1734 VSS.n584 3.26621
R3562 VSS.n685 VSS.t2010 3.26621
R3563 VSS.t1957 VSS.n684 3.26621
R3564 VSS.t1708 VSS.n585 3.26621
R3565 VSS.n658 VSS.t2004 3.26621
R3566 VSS.n659 VSS.t1984 3.26621
R3567 VSS.t1749 VSS.n586 3.26621
R3568 VSS.n693 VSS.t2012 3.26621
R3569 VSS.t1954 VSS.n692 3.26621
R3570 VSS.t1706 VSS.n587 3.26621
R3571 VSS.n651 VSS.t1992 3.26621
R3572 VSS.n652 VSS.t1976 3.26621
R3573 VSS.t1732 VSS.n588 3.26621
R3574 VSS.n709 VSS.t2016 3.26621
R3575 VSS.t1961 VSS.n708 3.26621
R3576 VSS.t1701 VSS.n591 3.26621
R3577 VSS.n701 VSS.t2018 3.18737
R3578 VSS.t1982 VSS.n700 3.18737
R3579 VSS.t1714 VSS.n589 3.18737
R3580 VSS VSS.n252 3.163
R3581 VSS VSS.n250 3.15979
R3582 VSS VSS.n254 3.12124
R3583 VSS VSS.n804 3.11598
R3584 VSS.n838 VSS 3.11598
R3585 VSS VSS.n872 3.11598
R3586 VSS VSS.n764 3.11598
R3587 VSS VSS.n790 3.11598
R3588 VSS VSS.n814 3.10254
R3589 VSS VSS.n824 3.10254
R3590 VSS VSS.n773 3.10254
R3591 VSS VSS.n782 3.10254
R3592 VSS.n677 VSS.t1986 2.84963
R3593 VSS.t1974 VSS.n676 2.84963
R3594 VSS.t1728 VSS.n583 2.84963
R3595 VSS.n561 VSS.n545 2.29217
R3596 VSS.n807 VSS.n806 2.27663
R3597 VSS.n833 VSS.n832 2.27663
R3598 VSS.n817 VSS.n816 2.27663
R3599 VSS.n827 VSS.n826 2.27663
R3600 VSS.n754 VSS.n753 2.27663
R3601 VSS.n768 VSS.n767 2.27663
R3602 VSS.n794 VSS.n793 2.27663
R3603 VSS.n777 VSS.n776 2.27663
R3604 VSS.n785 VSS.n784 2.27663
R3605 VSS.n805 VSS 2.2624
R3606 VSS VSS.n837 2.2624
R3607 VSS.n873 VSS 2.2624
R3608 VSS.n765 VSS 2.2624
R3609 VSS.n791 VSS 2.2624
R3610 VSS.n815 VSS 2.25356
R3611 VSS.n825 VSS 2.25356
R3612 VSS.n774 VSS 2.25356
R3613 VSS.n783 VSS 2.25356
R3614 VSS.n1021 VSS.n1017 2.2505
R3615 VSS.n1037 VSS.n1018 2.2505
R3616 VSS.n1033 VSS.n1032 2.2505
R3617 VSS.n1028 VSS.n1027 2.2505
R3618 VSS.n1044 VSS.n1043 2.2505
R3619 VSS.n985 VSS.n981 2.2505
R3620 VSS.n1001 VSS.n982 2.2505
R3621 VSS.n997 VSS.n996 2.2505
R3622 VSS.n992 VSS.n991 2.2505
R3623 VSS.n1008 VSS.n1007 2.2505
R3624 VSS.n1176 VSS.n629 2.2505
R3625 VSS.n1161 VSS.n630 2.2505
R3626 VSS.n1172 VSS.n1167 2.2505
R3627 VSS.n1171 VSS.n1170 2.2505
R3628 VSS.n1178 VSS.n1177 2.2505
R3629 VSS.n951 VSS.n947 2.2505
R3630 VSS.n967 VSS.n948 2.2505
R3631 VSS.n963 VSS.n962 2.2505
R3632 VSS.n958 VSS.n957 2.2505
R3633 VSS.n974 VSS.n973 2.2505
R3634 VSS.n1055 VSS.n1051 2.2505
R3635 VSS.n1071 VSS.n1052 2.2505
R3636 VSS.n1067 VSS.n1066 2.2505
R3637 VSS.n1062 VSS.n1061 2.2505
R3638 VSS.n1078 VSS.n1077 2.2505
R3639 VSS.n917 VSS.n913 2.2505
R3640 VSS.n933 VSS.n914 2.2505
R3641 VSS.n929 VSS.n928 2.2505
R3642 VSS.n924 VSS.n923 2.2505
R3643 VSS.n940 VSS.n939 2.2505
R3644 VSS.n740 VSS.n739 2.2505
R3645 VSS.n1094 VSS.n733 2.2505
R3646 VSS.n1105 VSS.n1100 2.2505
R3647 VSS.n1104 VSS.n1103 2.2505
R3648 VSS.n1090 VSS.n1089 2.2505
R3649 VSS.n883 VSS.n879 2.2505
R3650 VSS.n899 VSS.n880 2.2505
R3651 VSS.n895 VSS.n894 2.2505
R3652 VSS.n890 VSS.n889 2.2505
R3653 VSS.n906 VSS.n905 2.2505
R3654 VSS.n864 VSS.n720 2.2505
R3655 VSS.n1118 VSS.n718 2.2505
R3656 VSS.n1125 VSS.n1124 2.2505
R3657 VSS.n1151 VSS.n1150 2.2505
R3658 VSS.n1114 VSS.n1113 2.2505
R3659 VSS.n1399 VSS.n1398 2.14536
R3660 VSS.n1218 VSS.n599 2.0027
R3661 VSS.n1144 VSS.n1143 1.96262
R3662 VSS.n1675 VSS.n1674 1.8615
R3663 VSS.n1298 VSS.t672 1.79617
R3664 VSS.t364 VSS.n1297 1.79617
R3665 VSS.n1535 VSS.t1859 1.79617
R3666 VSS.t211 VSS.n1534 1.79617
R3667 VSS.n448 VSS.t42 1.79617
R3668 VSS.n1144 VSS 1.71641
R3669 VSS.n1130 VSS 1.71262
R3670 VSS.n855 VSS.n854 1.7029
R3671 VSS.n857 VSS.n856 1.70078
R3672 VSS.n1142 VSS 1.6426
R3673 VSS.n1138 VSS 1.64065
R3674 VSS.n1141 VSS 1.63497
R3675 VSS.n450 VSS.t118 1.38705
R3676 VSS.n1324 VSS.t939 1.24093
R3677 VSS.t880 VSS.n1323 1.24093
R3678 VSS.n1308 VSS.t840 1.24093
R3679 VSS.n1147 VSS.n1146 0.990274
R3680 VSS.n854 VSS.n853 0.931911
R3681 VSS.n860 VSS.n857 0.931904
R3682 VSS.t377 VSS.n575 0.915261
R3683 VSS.n1669 VSS 0.862278
R3684 VSS.n1046 VSS.n1045 0.853
R3685 VSS.n1048 VSS.n1015 0.853
R3686 VSS.n1016 VSS.n728 0.853
R3687 VSS.n1031 VSS.n1029 0.853
R3688 VSS.n1030 VSS.n713 0.853
R3689 VSS.n1045 VSS.n1044 0.853
R3690 VSS.n1017 VSS.n1015 0.853
R3691 VSS.n1018 VSS.n1016 0.853
R3692 VSS.n1032 VSS.n1031 0.853
R3693 VSS.n1030 VSS.n1028 0.853
R3694 VSS.n1010 VSS.n1009 0.853
R3695 VSS.n1012 VSS.n979 0.853
R3696 VSS.n980 VSS.n727 0.853
R3697 VSS.n995 VSS.n993 0.853
R3698 VSS.n994 VSS.n638 0.853
R3699 VSS.n1009 VSS.n1008 0.853
R3700 VSS.n981 VSS.n979 0.853
R3701 VSS.n982 VSS.n980 0.853
R3702 VSS.n996 VSS.n995 0.853
R3703 VSS.n994 VSS.n992 0.853
R3704 VSS.n1175 VSS.n631 0.853
R3705 VSS.n1014 VSS.n628 0.853
R3706 VSS.n1174 VSS.n632 0.853
R3707 VSS.n1173 VSS.n633 0.853
R3708 VSS.n1156 VSS.n1155 0.853
R3709 VSS.n1176 VSS.n1175 0.853
R3710 VSS.n1177 VSS.n628 0.853
R3711 VSS.n1174 VSS.n630 0.853
R3712 VSS.n1173 VSS.n1172 0.853
R3713 VSS.n1171 VSS.n1156 0.853
R3714 VSS.n976 VSS.n975 0.853
R3715 VSS.n978 VSS.n945 0.853
R3716 VSS.n946 VSS.n726 0.853
R3717 VSS.n961 VSS.n959 0.853
R3718 VSS.n960 VSS.n637 0.853
R3719 VSS.n975 VSS.n974 0.853
R3720 VSS.n947 VSS.n945 0.853
R3721 VSS.n948 VSS.n946 0.853
R3722 VSS.n962 VSS.n961 0.853
R3723 VSS.n960 VSS.n958 0.853
R3724 VSS.n1080 VSS.n1079 0.853
R3725 VSS.n1082 VSS.n1049 0.853
R3726 VSS.n1050 VSS.n729 0.853
R3727 VSS.n1065 VSS.n1063 0.853
R3728 VSS.n1064 VSS.n714 0.853
R3729 VSS.n1079 VSS.n1078 0.853
R3730 VSS.n1051 VSS.n1049 0.853
R3731 VSS.n1052 VSS.n1050 0.853
R3732 VSS.n1066 VSS.n1065 0.853
R3733 VSS.n1064 VSS.n1062 0.853
R3734 VSS.n942 VSS.n941 0.853
R3735 VSS.n944 VSS.n911 0.853
R3736 VSS.n912 VSS.n725 0.853
R3737 VSS.n927 VSS.n925 0.853
R3738 VSS.n926 VSS.n636 0.853
R3739 VSS.n941 VSS.n940 0.853
R3740 VSS.n913 VSS.n911 0.853
R3741 VSS.n914 VSS.n912 0.853
R3742 VSS.n928 VSS.n927 0.853
R3743 VSS.n926 VSS.n924 0.853
R3744 VSS.n1088 VSS.n730 0.853
R3745 VSS.n1087 VSS.n1086 0.853
R3746 VSS.n1108 VSS.n731 0.853
R3747 VSS.n1107 VSS.n1106 0.853
R3748 VSS.n732 VSS.n715 0.853
R3749 VSS.n1089 VSS.n1088 0.853
R3750 VSS.n1087 VSS.n740 0.853
R3751 VSS.n733 VSS.n731 0.853
R3752 VSS.n1106 VSS.n1105 0.853
R3753 VSS.n1104 VSS.n732 0.853
R3754 VSS.n908 VSS.n907 0.853
R3755 VSS.n910 VSS.n877 0.853
R3756 VSS.n878 VSS.n724 0.853
R3757 VSS.n893 VSS.n891 0.853
R3758 VSS.n892 VSS.n635 0.853
R3759 VSS.n907 VSS.n906 0.853
R3760 VSS.n879 VSS.n877 0.853
R3761 VSS.n880 VSS.n878 0.853
R3762 VSS.n894 VSS.n893 0.853
R3763 VSS.n892 VSS.n890 0.853
R3764 VSS.n1112 VSS.n722 0.853
R3765 VSS.n1084 VSS.n721 0.853
R3766 VSS.n1111 VSS.n1110 0.853
R3767 VSS.n717 VSS.n716 0.853
R3768 VSS.n1153 VSS.n1152 0.853
R3769 VSS.n1113 VSS.n1112 0.853
R3770 VSS.n721 VSS.n720 0.853
R3771 VSS.n1111 VSS.n718 0.853
R3772 VSS.n1125 VSS.n717 0.853
R3773 VSS.n1152 VSS.n1151 0.853
R3774 VSS.n1149 VSS.n1148 0.845955
R3775 VSS.n1646 VSS.n93 0.808432
R3776 VSS.t515 VSS.t1171 0.808432
R3777 VSS.t1907 VSS.t837 0.808432
R3778 VSS.n305 VSS.n304 0.794268
R3779 VSS.n435 VSS.n434 0.794268
R3780 VSS.n473 VSS.n472 0.794268
R3781 VSS VSS.n1025 0.684563
R3782 VSS.n1034 VSS 0.684563
R3783 VSS.n1038 VSS 0.684563
R3784 VSS.n1022 VSS 0.684563
R3785 VSS.n1040 VSS 0.684563
R3786 VSS VSS.n989 0.684563
R3787 VSS.n998 VSS 0.684563
R3788 VSS.n1002 VSS 0.684563
R3789 VSS.n986 VSS 0.684563
R3790 VSS.n1004 VSS 0.684563
R3791 VSS VSS.n1168 0.684563
R3792 VSS.n1164 VSS 0.684563
R3793 VSS.n1162 VSS 0.684563
R3794 VSS.n1158 VSS 0.684563
R3795 VSS.n1179 VSS 0.684563
R3796 VSS VSS.n955 0.684563
R3797 VSS.n964 VSS 0.684563
R3798 VSS.n968 VSS 0.684563
R3799 VSS.n952 VSS 0.684563
R3800 VSS.n970 VSS 0.684563
R3801 VSS VSS.n1059 0.684563
R3802 VSS.n1068 VSS 0.684563
R3803 VSS.n1072 VSS 0.684563
R3804 VSS.n1056 VSS 0.684563
R3805 VSS.n1074 VSS 0.684563
R3806 VSS VSS.n921 0.684563
R3807 VSS.n930 VSS 0.684563
R3808 VSS.n934 VSS 0.684563
R3809 VSS.n918 VSS 0.684563
R3810 VSS.n936 VSS 0.684563
R3811 VSS VSS.n1101 0.684563
R3812 VSS.n1097 VSS 0.684563
R3813 VSS.n1095 VSS 0.684563
R3814 VSS.n736 VSS 0.684563
R3815 VSS.n1091 VSS 0.684563
R3816 VSS VSS.n887 0.684563
R3817 VSS.n896 VSS 0.684563
R3818 VSS.n900 VSS 0.684563
R3819 VSS.n884 VSS 0.684563
R3820 VSS.n902 VSS 0.684563
R3821 VSS.n1121 VSS 0.684563
R3822 VSS.n1119 VSS 0.684563
R3823 VSS.n865 VSS 0.684563
R3824 VSS.n1115 VSS 0.684563
R3825 VSS.n1143 VSS.n1135 0.659647
R3826 VSS VSS.n1026 0.653922
R3827 VSS VSS.n1024 0.653922
R3828 VSS VSS.n1036 0.653922
R3829 VSS VSS.n1020 0.653922
R3830 VSS VSS.n1042 0.653922
R3831 VSS VSS.n990 0.653922
R3832 VSS VSS.n988 0.653922
R3833 VSS VSS.n1000 0.653922
R3834 VSS VSS.n984 0.653922
R3835 VSS VSS.n1006 0.653922
R3836 VSS VSS.n1169 0.653922
R3837 VSS VSS.n1166 0.653922
R3838 VSS VSS.n1160 0.653922
R3839 VSS.n1157 VSS 0.653922
R3840 VSS VSS.n627 0.653922
R3841 VSS VSS.n956 0.653922
R3842 VSS VSS.n954 0.653922
R3843 VSS VSS.n966 0.653922
R3844 VSS VSS.n950 0.653922
R3845 VSS VSS.n972 0.653922
R3846 VSS VSS.n1060 0.653922
R3847 VSS VSS.n1058 0.653922
R3848 VSS VSS.n1070 0.653922
R3849 VSS VSS.n1054 0.653922
R3850 VSS VSS.n1076 0.653922
R3851 VSS VSS.n922 0.653922
R3852 VSS VSS.n920 0.653922
R3853 VSS VSS.n932 0.653922
R3854 VSS VSS.n916 0.653922
R3855 VSS VSS.n938 0.653922
R3856 VSS VSS.n1102 0.653922
R3857 VSS VSS.n1099 0.653922
R3858 VSS VSS.n1093 0.653922
R3859 VSS VSS.n738 0.653922
R3860 VSS VSS.n734 0.653922
R3861 VSS VSS.n888 0.653922
R3862 VSS VSS.n886 0.653922
R3863 VSS VSS.n898 0.653922
R3864 VSS VSS.n882 0.653922
R3865 VSS VSS.n904 0.653922
R3866 VSS VSS.n1123 0.653922
R3867 VSS VSS.n1117 0.653922
R3868 VSS VSS.n863 0.653922
R3869 VSS VSS.n719 0.653922
R3870 VSS.n1145 VSS.n1144 0.636864
R3871 VSS.n1677 VSS.n1664 0.58175
R3872 VSS.n1623 VSS.n120 0.523852
R3873 VSS.n1620 VSS.n1615 0.523852
R3874 VSS.n1610 VSS.n1605 0.523852
R3875 VSS.n1601 VSS.n1596 0.523852
R3876 VSS.n1592 VSS.n1587 0.523852
R3877 VSS.n1583 VSS.n1578 0.523852
R3878 VSS.n1573 VSS.n1568 0.523852
R3879 VSS.n1630 VSS.n113 0.523852
R3880 VSS.n1329 VSS.n578 0.523852
R3881 VSS.n1222 VSS.n594 0.523852
R3882 VSS.n1292 VSS.n1290 0.523852
R3883 VSS.n571 VSS.n570 0.523852
R3884 VSS.n539 VSS.n538 0.523852
R3885 VSS.n530 VSS.n529 0.523852
R3886 VSS.n261 VSS.n260 0.523852
R3887 VSS.n1342 VSS.n246 0.523852
R3888 VSS.n1641 VSS.n101 0.523852
R3889 VSS.n1366 VSS.n1358 0.523852
R3890 VSS.n1375 VSS.n1370 0.523852
R3891 VSS.n1378 VSS.n233 0.523852
R3892 VSS.n1354 VSS.n236 0.523852
R3893 VSS.n1465 VSS.n174 0.523852
R3894 VSS.n1468 VSS.n171 0.523852
R3895 VSS.n513 VSS.n272 0.523852
R3896 VSS.n510 VSS.n505 0.523852
R3897 VSS.n501 VSS.n284 0.523852
R3898 VSS.n280 VSS.n275 0.523852
R3899 VSS.n1523 VSS.n131 0.523852
R3900 VSS.n1526 VSS.n128 0.523852
R3901 VSS.n1276 VSS.n1271 0.523852
R3902 VSS.n1279 VSS.n1250 0.523852
R3903 VSS.n1267 VSS.n1262 0.523852
R3904 VSS.n1258 VSS.n1253 0.523852
R3905 VSS.n1664 VSS.n72 0.523852
R3906 VSS.n1680 VSS.n69 0.523852
R3907 VSS.n1697 VSS.n42 0.523852
R3908 VSS.n1700 VSS.n39 0.523852
R3909 VSS.n1717 VSS.n15 0.523852
R3910 VSS.n1720 VSS.n12 0.523852
R3911 VSS.n295 VSS.n290 0.523852
R3912 VSS.n315 VSS.n310 0.523852
R3913 VSS.n391 VSS.n390 0.523852
R3914 VSS.n396 VSS.n395 0.523852
R3915 VSS.n401 VSS.n400 0.523852
R3916 VSS.n406 VSS.n405 0.523852
R3917 VSS.n411 VSS.n410 0.523852
R3918 VSS.n416 VSS.n415 0.523852
R3919 VSS.n425 VSS.n420 0.523852
R3920 VSS.n445 VSS.n440 0.523852
R3921 VSS.n1657 VSS.n83 0.523852
R3922 VSS.n1687 VSS.n57 0.523852
R3923 VSS.n1690 VSS.n54 0.523852
R3924 VSS.n1707 VSS.n29 0.523852
R3925 VSS.n1710 VSS.n26 0.523852
R3926 VSS.n454 VSS.n453 0.523852
R3927 VSS.n463 VSS.n458 0.523852
R3928 VSS.n1318 VSS.n1316 0.523852
R3929 VSS.n1213 VSS.n602 0.523852
R3930 VSS.n483 VSS.n478 0.523374
R3931 VSS.n860 VSS.n859 0.447662
R3932 VSS.n853 VSS.n799 0.447662
R3933 VSS.n1134 VSS.n1133 0.443357
R3934 VSS.n800 VSS.n797 0.380713
R3935 VSS.n834 VSS.n797 0.380713
R3936 VSS.n810 VSS.n797 0.380713
R3937 VSS.n820 VSS.n797 0.380713
R3938 VSS.n797 VSS.n751 0.380713
R3939 VSS.n797 VSS.n770 0.380713
R3940 VSS.n797 VSS.n796 0.380713
R3941 VSS.n797 VSS.n779 0.380713
R3942 VSS.n797 VSS.n787 0.380713
R3943 VSS.n876 VSS.n747 0.3805
R3944 VSS.n712 VSS.n679 0.3805
R3945 VSS.n674 VSS.n671 0.3805
R3946 VSS.n673 VSS.n598 0.3805
R3947 VSS.n876 VSS.n746 0.3805
R3948 VSS.n712 VSS.n642 0.3805
R3949 VSS.n671 VSS.n670 0.3805
R3950 VSS.n669 VSS.n598 0.3805
R3951 VSS.n876 VSS.n748 0.3805
R3952 VSS.n712 VSS.n687 0.3805
R3953 VSS.n682 VSS.n671 0.3805
R3954 VSS.n681 VSS.n598 0.3805
R3955 VSS.n876 VSS.n745 0.3805
R3956 VSS.n712 VSS.n641 0.3805
R3957 VSS.n671 VSS.n663 0.3805
R3958 VSS.n662 VSS.n598 0.3805
R3959 VSS.n876 VSS.n749 0.3805
R3960 VSS.n712 VSS.n695 0.3805
R3961 VSS.n690 VSS.n671 0.3805
R3962 VSS.n689 VSS.n598 0.3805
R3963 VSS.n876 VSS.n744 0.3805
R3964 VSS.n712 VSS.n640 0.3805
R3965 VSS.n671 VSS.n656 0.3805
R3966 VSS.n655 VSS.n598 0.3805
R3967 VSS.n876 VSS.n750 0.3805
R3968 VSS.n712 VSS.n703 0.3805
R3969 VSS.n698 VSS.n671 0.3805
R3970 VSS.n697 VSS.n598 0.3805
R3971 VSS.n876 VSS.n743 0.3805
R3972 VSS.n712 VSS.n639 0.3805
R3973 VSS.n671 VSS.n649 0.3805
R3974 VSS.n648 VSS.n598 0.3805
R3975 VSS.n876 VSS.n875 0.3805
R3976 VSS.n712 VSS.n711 0.3805
R3977 VSS.n706 VSS.n671 0.3805
R3978 VSS.n705 VSS.n598 0.3805
R3979 VSS.n1013 VSS.n723 0.3805
R3980 VSS.n1085 VSS.n1014 0.3805
R3981 VSS.n1109 VSS.n632 0.3805
R3982 VSS.n634 VSS.n633 0.3805
R3983 VSS.n1155 VSS.n1154 0.3805
R3984 VSS.n1011 VSS.n723 0.3805
R3985 VSS.n1085 VSS.n1012 0.3805
R3986 VSS.n1109 VSS.n727 0.3805
R3987 VSS.n993 VSS.n634 0.3805
R3988 VSS.n1154 VSS.n638 0.3805
R3989 VSS.n1047 VSS.n723 0.3805
R3990 VSS.n1085 VSS.n1048 0.3805
R3991 VSS.n1109 VSS.n728 0.3805
R3992 VSS.n1029 VSS.n634 0.3805
R3993 VSS.n1154 VSS.n713 0.3805
R3994 VSS.n977 VSS.n723 0.3805
R3995 VSS.n1085 VSS.n978 0.3805
R3996 VSS.n1109 VSS.n726 0.3805
R3997 VSS.n959 VSS.n634 0.3805
R3998 VSS.n1154 VSS.n637 0.3805
R3999 VSS.n1081 VSS.n723 0.3805
R4000 VSS.n1085 VSS.n1082 0.3805
R4001 VSS.n1109 VSS.n729 0.3805
R4002 VSS.n1063 VSS.n634 0.3805
R4003 VSS.n1154 VSS.n714 0.3805
R4004 VSS.n943 VSS.n723 0.3805
R4005 VSS.n1085 VSS.n944 0.3805
R4006 VSS.n1109 VSS.n725 0.3805
R4007 VSS.n925 VSS.n634 0.3805
R4008 VSS.n1154 VSS.n636 0.3805
R4009 VSS.n741 VSS.n723 0.3805
R4010 VSS.n1086 VSS.n1085 0.3805
R4011 VSS.n1109 VSS.n1108 0.3805
R4012 VSS.n1107 VSS.n634 0.3805
R4013 VSS.n1154 VSS.n715 0.3805
R4014 VSS.n909 VSS.n723 0.3805
R4015 VSS.n1085 VSS.n910 0.3805
R4016 VSS.n1109 VSS.n724 0.3805
R4017 VSS.n891 VSS.n634 0.3805
R4018 VSS.n1154 VSS.n635 0.3805
R4019 VSS.n1083 VSS.n723 0.3805
R4020 VSS.n1085 VSS.n1084 0.3805
R4021 VSS.n1110 VSS.n1109 0.3805
R4022 VSS.n716 VSS.n634 0.3805
R4023 VSS.n1154 VSS.n1153 0.3805
R4024 VSS.n1032 VSS.n1018 0.364986
R4025 VSS.n996 VSS.n982 0.364986
R4026 VSS.n1172 VSS.n630 0.364986
R4027 VSS.n962 VSS.n948 0.364986
R4028 VSS.n1066 VSS.n1052 0.364986
R4029 VSS.n928 VSS.n914 0.364986
R4030 VSS.n1105 VSS.n733 0.364986
R4031 VSS.n894 VSS.n880 0.364986
R4032 VSS.n1125 VSS.n718 0.364986
R4033 VSS.n1032 VSS.n1028 0.364597
R4034 VSS.n996 VSS.n992 0.364597
R4035 VSS.n1172 VSS.n1171 0.364597
R4036 VSS.n962 VSS.n958 0.364597
R4037 VSS.n1066 VSS.n1062 0.364597
R4038 VSS.n928 VSS.n924 0.364597
R4039 VSS.n1105 VSS.n1104 0.364597
R4040 VSS.n894 VSS.n890 0.364597
R4041 VSS.n1151 VSS.n1125 0.364597
R4042 VSS.n1044 VSS.n1018 0.36265
R4043 VSS.n1008 VSS.n982 0.36265
R4044 VSS.n1176 VSS.n630 0.36265
R4045 VSS.n974 VSS.n948 0.36265
R4046 VSS.n1078 VSS.n1052 0.36265
R4047 VSS.n940 VSS.n914 0.36265
R4048 VSS.n1089 VSS.n733 0.36265
R4049 VSS.n906 VSS.n880 0.36265
R4050 VSS.n1113 VSS.n718 0.36265
R4051 VSS.n1044 VSS.n1017 0.361871
R4052 VSS.n1008 VSS.n981 0.361871
R4053 VSS.n1177 VSS.n1176 0.361871
R4054 VSS.n974 VSS.n947 0.361871
R4055 VSS.n1078 VSS.n1051 0.361871
R4056 VSS.n940 VSS.n913 0.361871
R4057 VSS.n1089 VSS.n740 0.361871
R4058 VSS.n906 VSS.n879 0.361871
R4059 VSS.n1113 VSS.n720 0.361871
R4060 VSS.n845 VSS 0.351639
R4061 VSS.n1627 VSS 0.282093
R4062 VSS.n1619 VSS 0.282093
R4063 VSS.n1609 VSS 0.282093
R4064 VSS.n1600 VSS 0.282093
R4065 VSS.n1591 VSS 0.282093
R4066 VSS.n1582 VSS 0.282093
R4067 VSS.n1572 VSS 0.282093
R4068 VSS.n1629 VSS 0.282093
R4069 VSS.n1328 VSS 0.282093
R4070 VSS.n1221 VSS 0.282093
R4071 VSS.n1365 VSS 0.282093
R4072 VSS.n1374 VSS 0.282093
R4073 VSS.n1382 VSS 0.282093
R4074 VSS.n1353 VSS 0.282093
R4075 VSS.n1464 VSS 0.282093
R4076 VSS.n1472 VSS 0.282093
R4077 VSS.n517 VSS 0.282093
R4078 VSS.n509 VSS 0.282093
R4079 VSS.n500 VSS 0.282093
R4080 VSS.n279 VSS 0.282093
R4081 VSS.n1522 VSS 0.282093
R4082 VSS.n1530 VSS 0.282093
R4083 VSS.n1275 VSS 0.282093
R4084 VSS.n1283 VSS 0.282093
R4085 VSS.n1266 VSS 0.282093
R4086 VSS.n1257 VSS 0.282093
R4087 VSS.n1663 VSS 0.282093
R4088 VSS.n1684 VSS 0.282093
R4089 VSS.n1696 VSS 0.282093
R4090 VSS.n1704 VSS 0.282093
R4091 VSS.n1716 VSS 0.282093
R4092 VSS.n1724 VSS 0.282093
R4093 VSS.n294 VSS 0.282093
R4094 VSS.n314 VSS 0.282093
R4095 VSS.n80 VSS 0.282093
R4096 VSS.n65 VSS 0.282093
R4097 VSS.n50 VSS 0.282093
R4098 VSS.n36 VSS 0.282093
R4099 VSS.n23 VSS 0.282093
R4100 VSS.n4 VSS 0.282093
R4101 VSS.n424 VSS 0.282093
R4102 VSS.n444 VSS 0.282093
R4103 VSS.n1661 VSS 0.282093
R4104 VSS.n1686 VSS 0.282093
R4105 VSS.n1694 VSS 0.282093
R4106 VSS.n1706 VSS 0.282093
R4107 VSS.n1714 VSS 0.282093
R4108 VSS.n9 VSS 0.282093
R4109 VSS.n462 VSS 0.282093
R4110 VSS.n482 VSS 0.282093
R4111 VSS.n1217 VSS 0.282093
R4112 VSS VSS.n1287 0.277973
R4113 VSS VSS.n543 0.277973
R4114 VSS VSS.n534 0.277973
R4115 VSS VSS.n265 0.277973
R4116 VSS VSS.n249 0.277973
R4117 VSS VSS.n243 0.277973
R4118 VSS VSS.n98 0.277973
R4119 VSS VSS.n1313 0.277973
R4120 VSS.n806 VSS.n805 0.255642
R4121 VSS.n837 VSS.n833 0.255642
R4122 VSS.n816 VSS.n815 0.255642
R4123 VSS.n826 VSS.n825 0.255642
R4124 VSS.n873 VSS.n753 0.255642
R4125 VSS.n768 VSS.n765 0.255642
R4126 VSS.n794 VSS.n791 0.255642
R4127 VSS.n777 VSS.n774 0.255642
R4128 VSS.n785 VSS.n783 0.255642
R4129 VSS.n1134 VSS 0.241706
R4130 VSS VSS.n1149 0.210927
R4131 VSS.n1293 VSS 0.152973
R4132 VSS.n567 VSS 0.152973
R4133 VSS.n535 VSS 0.152973
R4134 VSS.n526 VSS 0.152973
R4135 VSS.n257 VSS 0.152973
R4136 VSS.n1343 VSS 0.152973
R4137 VSS.n1642 VSS 0.152973
R4138 VSS.n1319 VSS 0.152973
R4139 VSS.n307 VSS 0.151599
R4140 VSS VSS.n1626 0.150225
R4141 VSS VSS.n1618 0.150225
R4142 VSS VSS.n1608 0.150225
R4143 VSS VSS.n1599 0.150225
R4144 VSS VSS.n1590 0.150225
R4145 VSS VSS.n1581 0.150225
R4146 VSS VSS.n1571 0.150225
R4147 VSS VSS.n116 0.150225
R4148 VSS VSS.n581 0.150225
R4149 VSS VSS.n597 0.150225
R4150 VSS VSS.n1361 0.150225
R4151 VSS VSS.n1373 0.150225
R4152 VSS VSS.n1381 0.150225
R4153 VSS VSS.n239 0.150225
R4154 VSS VSS.n177 0.150225
R4155 VSS VSS.n1471 0.150225
R4156 VSS VSS.n516 0.150225
R4157 VSS VSS.n508 0.150225
R4158 VSS VSS.n287 0.150225
R4159 VSS VSS.n278 0.150225
R4160 VSS VSS.n134 0.150225
R4161 VSS VSS.n1529 0.150225
R4162 VSS VSS.n1274 0.150225
R4163 VSS VSS.n1282 0.150225
R4164 VSS VSS.n1265 0.150225
R4165 VSS VSS.n1256 0.150225
R4166 VSS VSS.n75 0.150225
R4167 VSS VSS.n1683 0.150225
R4168 VSS VSS.n45 0.150225
R4169 VSS VSS.n1703 0.150225
R4170 VSS VSS.n18 0.150225
R4171 VSS VSS.n1723 0.150225
R4172 VSS VSS.n293 0.150225
R4173 VSS VSS.n313 0.150225
R4174 VSS VSS.n79 0.150225
R4175 VSS VSS.n64 0.150225
R4176 VSS VSS.n49 0.150225
R4177 VSS VSS.n35 0.150225
R4178 VSS VSS.n22 0.150225
R4179 VSS VSS.n3 0.150225
R4180 VSS VSS.n423 0.150225
R4181 VSS VSS.n443 0.150225
R4182 VSS VSS.n1660 0.150225
R4183 VSS VSS.n60 0.150225
R4184 VSS VSS.n1693 0.150225
R4185 VSS VSS.n32 0.150225
R4186 VSS VSS.n1713 0.150225
R4187 VSS VSS.n8 0.150225
R4188 VSS VSS.n461 0.150225
R4189 VSS VSS.n481 0.150225
R4190 VSS VSS.n1216 0.150225
R4191 VSS.n846 VSS.n845 0.148387
R4192 VSS.n840 VSS 0.143357
R4193 VSS.n1029 VSS.n728 0.137547
R4194 VSS.n1031 VSS.n1016 0.137547
R4195 VSS.n993 VSS.n727 0.137547
R4196 VSS.n995 VSS.n980 0.137547
R4197 VSS.n633 VSS.n632 0.137547
R4198 VSS.n1174 VSS.n1173 0.137547
R4199 VSS.n959 VSS.n726 0.137547
R4200 VSS.n961 VSS.n946 0.137547
R4201 VSS.n1063 VSS.n729 0.137547
R4202 VSS.n1065 VSS.n1050 0.137547
R4203 VSS.n925 VSS.n725 0.137547
R4204 VSS.n927 VSS.n912 0.137547
R4205 VSS.n1108 VSS.n1107 0.137547
R4206 VSS.n1106 VSS.n731 0.137547
R4207 VSS.n891 VSS.n724 0.137547
R4208 VSS.n893 VSS.n878 0.137547
R4209 VSS.n1110 VSS.n716 0.137547
R4210 VSS.n1111 VSS.n717 0.137547
R4211 VSS.n1029 VSS.n713 0.1374
R4212 VSS.n1031 VSS.n1030 0.1374
R4213 VSS.n993 VSS.n638 0.1374
R4214 VSS.n995 VSS.n994 0.1374
R4215 VSS.n1155 VSS.n633 0.1374
R4216 VSS.n1173 VSS.n1156 0.1374
R4217 VSS.n959 VSS.n637 0.1374
R4218 VSS.n961 VSS.n960 0.1374
R4219 VSS.n1063 VSS.n714 0.1374
R4220 VSS.n1065 VSS.n1064 0.1374
R4221 VSS.n925 VSS.n636 0.1374
R4222 VSS.n927 VSS.n926 0.1374
R4223 VSS.n1107 VSS.n715 0.1374
R4224 VSS.n1106 VSS.n732 0.1374
R4225 VSS.n891 VSS.n635 0.1374
R4226 VSS.n893 VSS.n892 0.1374
R4227 VSS.n1153 VSS.n716 0.1374
R4228 VSS.n1152 VSS.n717 0.1374
R4229 VSS.n1046 VSS.n728 0.136668
R4230 VSS.n1045 VSS.n1016 0.136668
R4231 VSS.n1010 VSS.n727 0.136668
R4232 VSS.n1009 VSS.n980 0.136668
R4233 VSS.n632 VSS.n631 0.136668
R4234 VSS.n1175 VSS.n1174 0.136668
R4235 VSS.n976 VSS.n726 0.136668
R4236 VSS.n975 VSS.n946 0.136668
R4237 VSS.n1080 VSS.n729 0.136668
R4238 VSS.n1079 VSS.n1050 0.136668
R4239 VSS.n942 VSS.n725 0.136668
R4240 VSS.n941 VSS.n912 0.136668
R4241 VSS.n1108 VSS.n730 0.136668
R4242 VSS.n1088 VSS.n731 0.136668
R4243 VSS.n908 VSS.n724 0.136668
R4244 VSS.n907 VSS.n878 0.136668
R4245 VSS.n1110 VSS.n722 0.136668
R4246 VSS.n1112 VSS.n1111 0.136668
R4247 VSS.n1045 VSS.n1015 0.136375
R4248 VSS.n1009 VSS.n979 0.136375
R4249 VSS.n1175 VSS.n628 0.136375
R4250 VSS.n975 VSS.n945 0.136375
R4251 VSS.n1079 VSS.n1049 0.136375
R4252 VSS.n941 VSS.n911 0.136375
R4253 VSS.n1088 VSS.n1087 0.136375
R4254 VSS.n907 VSS.n877 0.136375
R4255 VSS.n1112 VSS.n721 0.136375
R4256 VSS.n1048 VSS.n1047 0.136229
R4257 VSS.n1012 VSS.n1011 0.136229
R4258 VSS.n1014 VSS.n1013 0.136229
R4259 VSS.n978 VSS.n977 0.136229
R4260 VSS.n1082 VSS.n1081 0.136229
R4261 VSS.n944 VSS.n943 0.136229
R4262 VSS.n1086 VSS.n741 0.136229
R4263 VSS.n910 VSS.n909 0.136229
R4264 VSS.n1084 VSS.n1083 0.136229
R4265 VSS.n1305 VSS.n1228 0.13538
R4266 VSS.n1244 VSS.n1229 0.13538
R4267 VSS.n1303 VSS.n1230 0.13538
R4268 VSS.n1245 VSS.n1231 0.13538
R4269 VSS.n1302 VSS.n1232 0.13538
R4270 VSS.n1246 VSS.n1233 0.13538
R4271 VSS.n1301 VSS.n1234 0.13538
R4272 VSS.n1247 VSS.n1235 0.13538
R4273 VSS.n1558 VSS.n1539 0.13538
R4274 VSS.n1556 VSS.n1540 0.13538
R4275 VSS.n1554 VSS.n1541 0.13538
R4276 VSS.n1552 VSS.n1542 0.13538
R4277 VSS.n1550 VSS.n1543 0.13538
R4278 VSS.n1548 VSS.n1544 0.13538
R4279 VSS.n1546 VSS.n1545 0.13538
R4280 VSS.n1563 VSS.n1562 0.13538
R4281 VSS.n440 VSS.n439 0.122753
R4282 VSS.n475 VSS 0.118632
R4283 VSS.n305 VSS 0.107118
R4284 VSS.n435 VSS 0.107118
R4285 VSS.n473 VSS 0.107118
R4286 VSS.n1144 VSS.n1130 0.106561
R4287 VSS.n1293 VSS.n1292 0.0994011
R4288 VSS.n571 VSS.n567 0.0994011
R4289 VSS.n539 VSS.n535 0.0994011
R4290 VSS.n530 VSS.n526 0.0994011
R4291 VSS.n261 VSS.n257 0.0994011
R4292 VSS.n1343 VSS.n1342 0.0994011
R4293 VSS.n1642 VSS.n1641 0.0994011
R4294 VSS.n1319 VSS.n1318 0.0994011
R4295 VSS.n1627 VSS.n1623 0.0980275
R4296 VSS.n1620 VSS.n1619 0.0980275
R4297 VSS.n1610 VSS.n1609 0.0980275
R4298 VSS.n1601 VSS.n1600 0.0980275
R4299 VSS.n1592 VSS.n1591 0.0980275
R4300 VSS.n1583 VSS.n1582 0.0980275
R4301 VSS.n1573 VSS.n1572 0.0980275
R4302 VSS.n1630 VSS.n1629 0.0980275
R4303 VSS.n1329 VSS.n1328 0.0980275
R4304 VSS.n1222 VSS.n1221 0.0980275
R4305 VSS.n1366 VSS.n1365 0.0980275
R4306 VSS.n1375 VSS.n1374 0.0980275
R4307 VSS.n1382 VSS.n1378 0.0980275
R4308 VSS.n1354 VSS.n1353 0.0980275
R4309 VSS.n1465 VSS.n1464 0.0980275
R4310 VSS.n1472 VSS.n1468 0.0980275
R4311 VSS.n517 VSS.n513 0.0980275
R4312 VSS.n510 VSS.n509 0.0980275
R4313 VSS.n501 VSS.n500 0.0980275
R4314 VSS.n280 VSS.n279 0.0980275
R4315 VSS.n1523 VSS.n1522 0.0980275
R4316 VSS.n1530 VSS.n1526 0.0980275
R4317 VSS.n1276 VSS.n1275 0.0980275
R4318 VSS.n1283 VSS.n1279 0.0980275
R4319 VSS.n1267 VSS.n1266 0.0980275
R4320 VSS.n1258 VSS.n1257 0.0980275
R4321 VSS.n1664 VSS.n1663 0.0980275
R4322 VSS.n1684 VSS.n1680 0.0980275
R4323 VSS.n1697 VSS.n1696 0.0980275
R4324 VSS.n1704 VSS.n1700 0.0980275
R4325 VSS.n1717 VSS.n1716 0.0980275
R4326 VSS.n1724 VSS.n1720 0.0980275
R4327 VSS.n295 VSS.n294 0.0980275
R4328 VSS.n315 VSS.n314 0.0980275
R4329 VSS.n391 VSS.n80 0.0980275
R4330 VSS.n396 VSS.n65 0.0980275
R4331 VSS.n401 VSS.n50 0.0980275
R4332 VSS.n406 VSS.n36 0.0980275
R4333 VSS.n411 VSS.n23 0.0980275
R4334 VSS.n416 VSS.n4 0.0980275
R4335 VSS.n425 VSS.n424 0.0980275
R4336 VSS.n445 VSS.n444 0.0980275
R4337 VSS.n1661 VSS.n1657 0.0980275
R4338 VSS.n1687 VSS.n1686 0.0980275
R4339 VSS.n1694 VSS.n1690 0.0980275
R4340 VSS.n1707 VSS.n1706 0.0980275
R4341 VSS.n1714 VSS.n1710 0.0980275
R4342 VSS.n454 VSS.n9 0.0980275
R4343 VSS.n463 VSS.n462 0.0980275
R4344 VSS.n483 VSS.n482 0.0980275
R4345 VSS.n1217 VSS.n1213 0.0980275
R4346 VSS.n874 VSS.n752 0.0964335
R4347 VSS.n769 VSS.n762 0.0964335
R4348 VSS.n795 VSS.n788 0.0964335
R4349 VSS.n778 VSS.n771 0.0964335
R4350 VSS.n802 VSS.n801 0.0964334
R4351 VSS.n836 VSS.n835 0.0964334
R4352 VSS.n812 VSS.n811 0.0964334
R4353 VSS.n822 VSS.n821 0.0964334
R4354 VSS.n786 VSS.n780 0.0964334
R4355 VSS.n800 VSS.n745 0.0962852
R4356 VSS.n834 VSS.n747 0.0962852
R4357 VSS.n810 VSS.n746 0.0962852
R4358 VSS.n820 VSS.n748 0.0962852
R4359 VSS.n875 VSS.n751 0.0962852
R4360 VSS.n770 VSS.n743 0.0962852
R4361 VSS.n796 VSS.n750 0.0962852
R4362 VSS.n779 VSS.n744 0.0962852
R4363 VSS.n787 VSS.n749 0.0962852
R4364 VSS.n478 VSS.n477 0.09425
R4365 VSS.n437 VSS 0.0911593
R4366 VSS.n1445 VSS.n1444 0.0891315
R4367 VSS.n1027 VSS 0.0815302
R4368 VSS.n1033 VSS 0.0815302
R4369 VSS.n1037 VSS 0.0815302
R4370 VSS.n1021 VSS 0.0815302
R4371 VSS.n991 VSS 0.0815302
R4372 VSS.n997 VSS 0.0815302
R4373 VSS.n1001 VSS 0.0815302
R4374 VSS.n985 VSS 0.0815302
R4375 VSS.n1170 VSS 0.0815302
R4376 VSS.n1167 VSS 0.0815302
R4377 VSS.n1161 VSS 0.0815302
R4378 VSS.n1178 VSS 0.0815302
R4379 VSS.n957 VSS 0.0815302
R4380 VSS.n963 VSS 0.0815302
R4381 VSS.n967 VSS 0.0815302
R4382 VSS.n951 VSS 0.0815302
R4383 VSS.n1061 VSS 0.0815302
R4384 VSS.n1067 VSS 0.0815302
R4385 VSS.n1071 VSS 0.0815302
R4386 VSS.n1055 VSS 0.0815302
R4387 VSS.n923 VSS 0.0815302
R4388 VSS.n929 VSS 0.0815302
R4389 VSS.n933 VSS 0.0815302
R4390 VSS.n917 VSS 0.0815302
R4391 VSS.n1103 VSS 0.0815302
R4392 VSS.n1100 VSS 0.0815302
R4393 VSS.n1094 VSS 0.0815302
R4394 VSS.n739 VSS 0.0815302
R4395 VSS.n889 VSS 0.0815302
R4396 VSS.n895 VSS 0.0815302
R4397 VSS.n899 VSS 0.0815302
R4398 VSS.n883 VSS 0.0815302
R4399 VSS.n1150 VSS 0.0815302
R4400 VSS.n1124 VSS 0.0815302
R4401 VSS.n1118 VSS 0.0815302
R4402 VSS.n864 VSS 0.0815302
R4403 VSS.n1043 VSS 0.080902
R4404 VSS.n1007 VSS 0.080902
R4405 VSS VSS.n629 0.080902
R4406 VSS.n973 VSS 0.080902
R4407 VSS.n1077 VSS 0.080902
R4408 VSS.n939 VSS 0.080902
R4409 VSS.n1090 VSS 0.080902
R4410 VSS.n905 VSS 0.080902
R4411 VSS.n1114 VSS 0.080902
R4412 VSS.n1141 VSS.n1138 0.0762576
R4413 VSS.n1143 VSS.n1142 0.0758676
R4414 VSS.n1668 VSS 0.0755
R4415 VSS.n1612 VSS.n121 0.0748565
R4416 VSS.n309 VSS.n307 0.0733022
R4417 VSS.n439 VSS.n437 0.0733022
R4418 VSS.n477 VSS.n475 0.0733022
R4419 VSS.n301 VSS 0.0730524
R4420 VSS.n431 VSS 0.0730524
R4421 VSS.n469 VSS 0.0730524
R4422 VSS.n382 VSS.n380 0.0722856
R4423 VSS.n324 VSS.n322 0.0709486
R4424 VSS.n1444 VSS.n192 0.0688728
R4425 VSS.n1142 VSS.n1141 0.0686818
R4426 VSS.n1416 VSS.n205 0.0680689
R4427 VSS.n1413 VSS.n1407 0.0677291
R4428 VSS.n359 VSS.n197 0.0669376
R4429 VSS.n1441 VSS.n195 0.0668348
R4430 VSS.n1451 VSS.n185 0.0648054
R4431 VSS.n1432 VSS.n197 0.0634409
R4432 VSS.n1441 VSS.n1440 0.0633381
R4433 VSS.n310 VSS.n309 0.0623132
R4434 VSS.n1420 VSS.n1416 0.0621039
R4435 VSS.n1456 VSS.n185 0.061954
R4436 VSS.n1148 VSS.n1147 0.0602153
R4437 VSS.n1413 VSS.n1412 0.0596777
R4438 VSS.n322 VSS.n321 0.05943
R4439 VSS.n380 VSS.n379 0.0577845
R4440 VSS.n1140 VSS 0.0573182
R4441 VSS.n679 VSS.n674 0.0568488
R4442 VSS.n670 VSS.n642 0.0568488
R4443 VSS.n687 VSS.n682 0.0568488
R4444 VSS.n663 VSS.n641 0.0568488
R4445 VSS.n695 VSS.n690 0.0568488
R4446 VSS.n656 VSS.n640 0.0568488
R4447 VSS.n703 VSS.n698 0.0568488
R4448 VSS.n649 VSS.n639 0.0568488
R4449 VSS.n711 VSS.n706 0.0568488
R4450 VSS.n674 VSS.n673 0.0565926
R4451 VSS.n670 VSS.n669 0.0565926
R4452 VSS.n682 VSS.n681 0.0565926
R4453 VSS.n663 VSS.n662 0.0565926
R4454 VSS.n690 VSS.n689 0.0565926
R4455 VSS.n656 VSS.n655 0.0565926
R4456 VSS.n698 VSS.n697 0.0565926
R4457 VSS.n649 VSS.n648 0.0565926
R4458 VSS.n706 VSS.n705 0.0565926
R4459 VSS.n1127 VSS 0.0554242
R4460 VSS.n1414 VSS.n1413 0.0547857
R4461 VSS.n1416 VSS.n1415 0.0547857
R4462 VSS.n380 VSS.n214 0.0547857
R4463 VSS.n322 VSS.n206 0.0547857
R4464 VSS.n197 VSS.n194 0.0547857
R4465 VSS.n1442 VSS.n1441 0.0547857
R4466 VSS.n240 VSS.n185 0.0547857
R4467 VSS.n1444 VSS.n1443 0.0547857
R4468 VSS.n1306 VSS.n1305 0.0546237
R4469 VSS.n1244 VSS.n1243 0.0546237
R4470 VSS.n1303 VSS.n1242 0.0546237
R4471 VSS.n1245 VSS.n1241 0.0546237
R4472 VSS.n1302 VSS.n1240 0.0546237
R4473 VSS.n1246 VSS.n1239 0.0546237
R4474 VSS.n1301 VSS.n1238 0.0546237
R4475 VSS.n1247 VSS.n1237 0.0546237
R4476 VSS.n1559 VSS.n1558 0.0546237
R4477 VSS.n1557 VSS.n1556 0.0546237
R4478 VSS.n1555 VSS.n1554 0.0546237
R4479 VSS.n1553 VSS.n1552 0.0546237
R4480 VSS.n1551 VSS.n1550 0.0546237
R4481 VSS.n1549 VSS.n1548 0.0546237
R4482 VSS.n1547 VSS.n1546 0.0546237
R4483 VSS.n1564 VSS.n1563 0.0546237
R4484 VSS.n841 VSS.n840 0.0520464
R4485 VSS.n1027 VSS 0.0507513
R4486 VSS VSS.n1033 0.0507513
R4487 VSS VSS.n1037 0.0507513
R4488 VSS VSS.n1021 0.0507513
R4489 VSS.n1043 VSS 0.0507513
R4490 VSS.n991 VSS 0.0507513
R4491 VSS VSS.n997 0.0507513
R4492 VSS VSS.n1001 0.0507513
R4493 VSS VSS.n985 0.0507513
R4494 VSS.n1007 VSS 0.0507513
R4495 VSS.n1170 VSS 0.0507513
R4496 VSS.n1167 VSS 0.0507513
R4497 VSS VSS.n1161 0.0507513
R4498 VSS VSS.n629 0.0507513
R4499 VSS VSS.n1178 0.0507513
R4500 VSS.n957 VSS 0.0507513
R4501 VSS VSS.n963 0.0507513
R4502 VSS VSS.n967 0.0507513
R4503 VSS VSS.n951 0.0507513
R4504 VSS.n973 VSS 0.0507513
R4505 VSS.n1061 VSS 0.0507513
R4506 VSS VSS.n1067 0.0507513
R4507 VSS VSS.n1071 0.0507513
R4508 VSS VSS.n1055 0.0507513
R4509 VSS.n1077 VSS 0.0507513
R4510 VSS.n923 VSS 0.0507513
R4511 VSS VSS.n929 0.0507513
R4512 VSS VSS.n933 0.0507513
R4513 VSS VSS.n917 0.0507513
R4514 VSS.n939 VSS 0.0507513
R4515 VSS.n1103 VSS 0.0507513
R4516 VSS.n1100 VSS 0.0507513
R4517 VSS VSS.n1094 0.0507513
R4518 VSS.n739 VSS 0.0507513
R4519 VSS VSS.n1090 0.0507513
R4520 VSS.n889 VSS 0.0507513
R4521 VSS VSS.n895 0.0507513
R4522 VSS VSS.n899 0.0507513
R4523 VSS VSS.n883 0.0507513
R4524 VSS.n905 VSS 0.0507513
R4525 VSS.n1150 VSS 0.0507513
R4526 VSS.n1124 VSS 0.0507513
R4527 VSS VSS.n1118 0.0507513
R4528 VSS VSS.n864 0.0507513
R4529 VSS VSS.n1114 0.0507513
R4530 VSS.n1132 VSS 0.0497424
R4531 VSS.n1137 VSS 0.0497424
R4532 VSS.n1129 VSS 0.0497424
R4533 VSS.n607 VSS 0.0428228
R4534 VSS VSS.n223 0.0342079
R4535 VSS VSS.n219 0.0342079
R4536 VSS.n857 VSS 0.017073
R4537 VSS.n854 VSS 0.0168657
R4538 VSS.n1398 VSS.n108 0.0159873
R4539 VSS VSS.n1236 0.0155
R4540 VSS VSS.n215 0.0155
R4541 VSS VSS.n221 0.0155
R4542 VSS VSS.n228 0.0155
R4543 VSS VSS.n225 0.0155
R4544 VSS VSS.n1481 0.0155
R4545 VSS VSS.n160 0.0155
R4546 VSS.n1491 VSS 0.0155
R4547 VSS VSS.n157 0.0155
R4548 VSS VSS.n159 0.0155
R4549 VSS VSS.n158 0.0155
R4550 VSS.n842 VSS.n841 0.0155
R4551 VSS.n842 VSS 0.0155
R4552 VSS.n840 VSS.n831 0.0155
R4553 VSS.n831 VSS 0.0155
R4554 VSS VSS.n564 0.0155
R4555 VSS VSS.n556 0.0155
R4556 VSS.n552 VSS 0.0155
R4557 VSS.n554 VSS 0.0155
R4558 VSS.n553 VSS 0.0155
R4559 VSS.n559 VSS 0.0155
R4560 VSS.n1560 VSS 0.0155
R4561 VSS.n142 VSS 0.0139375
R4562 VSS.n1514 VSS 0.0139375
R4563 VSS.n447 VSS 0.0139375
R4564 VSS.n1533 VSS 0.0139375
R4565 VSS.n1296 VSS 0.0139375
R4566 VSS.n1299 VSS 0.0139375
R4567 VSS.n1322 VSS 0.0139375
R4568 VSS.n1325 VSS 0.0139375
R4569 VSS.n1392 VSS 0.0139375
R4570 VSS.n1390 VSS 0.0139375
R4571 VSS.n1395 VSS 0.0139375
R4572 VSS.n90 VSS 0.0139375
R4573 VSS.n1651 VSS 0.0139375
R4574 VSS.n342 VSS 0.0139375
R4575 VSS.n207 VSS 0.0139375
R4576 VSS.n94 VSS 0.0139375
R4577 VSS.n1645 VSS 0.0139375
R4578 VSS.n1648 VSS 0.0139375
R4579 VSS.n371 VSS 0.0139375
R4580 VSS.n340 VSS 0.0139375
R4581 VSS.n167 VSS 0.0139375
R4582 VSS.n162 VSS 0.0139375
R4583 VSS.n147 VSS 0.0139375
R4584 VSS.n331 VSS 0.0139375
R4585 VSS.n140 VSS 0.0139375
R4586 VSS.n136 VSS 0.0139375
R4587 VSS.n369 VSS 0.0139375
R4588 VSS.n345 VSS 0.0139375
R4589 VSS.n1476 VSS 0.0139375
R4590 VSS.n1479 VSS 0.0139375
R4591 VSS.n1505 VSS 0.0139375
R4592 VSS.n1507 VSS 0.0139375
R4593 VSS.n1516 VSS 0.0139375
R4594 VSS.n1519 VSS 0.0139375
R4595 VSS.n1388 VSS 0.0139375
R4596 VSS.n1385 VSS 0.0139375
R4597 VSS.n1350 VSS 0.0139375
R4598 VSS.n1345 VSS 0.0139375
R4599 VSS.n266 VSS 0.0139375
R4600 VSS.n268 VSS 0.0139375
R4601 VSS.n523 VSS 0.0139375
R4602 VSS.n494 VSS 0.0139375
R4603 VSS.n492 VSS 0.0139375
R4604 VSS.n489 VSS 0.0139375
R4605 VSS.n1474 VSS 0.0139375
R4606 VSS.n163 VSS 0.0139375
R4607 VSS.n1503 VSS 0.0139375
R4608 VSS.n138 VSS 0.0139375
R4609 VSS.n449 VSS 0.00589568
R4610 VSS.n1536 VSS 0.00589568
R4611 VSS.n1309 VSS 0.00589568
R4612 VSS.n1402 VSS 0.00589568
R4613 VSS.n373 VSS 0.00589568
R4614 VSS.n338 VSS 0.00589568
R4615 VSS.n334 VSS 0.00589568
R4616 VSS.n145 VSS 0.00589568
R4617 VSS.n366 VSS 0.00589568
R4618 VSS.n343 VSS 0.00589568
R4619 VSS.n164 VSS 0.00589568
R4620 VSS.n1510 VSS 0.00589568
R4621 VSS.n1362 VSS 0.00589568
R4622 VSS.n1347 VSS 0.00589568
R4623 VSS.n1461 VSS 0.00589568
R4624 VSS.n520 VSS 0.00589568
R4625 VSS.n497 VSS 0.00589568
R4626 VSS.n149 VSS 0.00589568
R4627 VSS.n150 VSS 0.00589568
R4628 VSS.n1512 VSS 0.00589568
R4629 VSS.n1410 VSS 0.0045625
R4630 VSS.n1406 VSS 0.0045625
R4631 VSS.n1419 VSS 0.0045625
R4632 VSS.n204 VSS 0.0045625
R4633 VSS.n375 VSS 0.0045625
R4634 VSS.n381 VSS 0.0045625
R4635 VSS.n317 VSS 0.0045625
R4636 VSS.n323 VSS 0.0045625
R4637 VSS.n1433 VSS 0.0045625
R4638 VSS.n358 VSS 0.0045625
R4639 VSS.n1450 VSS 0.0045625
R4640 VSS.n1455 VSS 0.0045625
R4641 VSS.n1446 VSS 0.0045625
R4642 VSS.n188 VSS 0.0045625
R4643 VSS.n196 VSS 0.0045625
R4644 VSS.n349 VSS 0.0045625
R4645 VSS.n855 VSS.n797 0.00268719
R4646 VSS.n1220 VSS.n1219 0.0016172
R4647 VSS.n1327 VSS.n1326 0.00148476
R4648 VSS.n1085 VSS.n876 0.00131823
R4649 VSS VSS.n1300 0.0012271
R4650 VSS.n1532 VSS 0.0012271
R4651 VSS.n1384 VSS 0.0012271
R4652 VSS.n1149 VSS.n1146 0.00112814
R4653 VSS.n1154 VSS.n634 0.00111302
R4654 VSS.n1109 VSS.n723 0.00111039
R4655 VSS.n1085 VSS.n723 0.00110777
R4656 VSS.n807 VSS 0.00106561
R4657 VSS.n832 VSS 0.00106561
R4658 VSS.n817 VSS 0.00106561
R4659 VSS.n827 VSS 0.00106561
R4660 VSS.n754 VSS 0.00106561
R4661 VSS.n767 VSS 0.00106561
R4662 VSS.n793 VSS 0.00106561
R4663 VSS.n776 VSS 0.00106561
R4664 VSS.n784 VSS 0.00106561
R4665 VSS.n1220 VSS 0.001035
R4666 VSS.n1363 VSS.n95 0.0010232
R4667 VSS.n1327 VSS 0.00101795
R4668 VSS VSS.n634 0.000979268
R4669 VSS.n1320 VSS 0.00097599
R4670 VSS.n1154 VSS.n712 0.00094452
R4671 VSS.n856 VSS 0.000911738
R4672 VSS.n498 VSS 0.000864532
R4673 VSS.n519 VSS 0.000864532
R4674 VSS.n1462 VSS 0.000864532
R4675 VSS.n551 VSS.n135 0.000856009
R4676 VSS.n1538 VSS.n1537 0.000806837
R4677 VSS.n1321 VSS.n582 0.000793724
R4678 VSS.n1295 VSS.n1284 0.000793724
R4679 VSS.n1531 VSS.n125 0.000793724
R4680 VSS.n491 VSS.n141 0.000793724
R4681 VSS.n524 VSS.n148 0.000793724
R4682 VSS.n1473 VSS.n168 0.000793724
R4683 VSS.n1352 VSS.n1351 0.000793724
R4684 VSS.n712 VSS.n671 0.000788479
R4685 VSS.n671 VSS.n598 0.000787168
R4686 VSS.n1326 VSS.n582 0.000771432
R4687 VSS.n1300 VSS.n1284 0.000771432
R4688 VSS.n1532 VSS.n1531 0.000771432
R4689 VSS.n1520 VSS.n137 0.000771432
R4690 VSS.n1685 VSS.n61 0.000771432
R4691 VSS.n1384 VSS.n193 0.000771432
R4692 VSS VSS.n0 0.000741929
R4693 VSS.n139 VSS.n137 0.000737339
R4694 VSS.n1725 VSS.n5 0.000737339
R4695 VSS.n1685 VSS.n66 0.000737339
R4696 VSS VSS.n742 0.000734061
R4697 VSS VSS.n0 0.000718326
R4698 VSS VSS.n61 0.000718326
R4699 VSS VSS.n1520 0.00071767
R4700 VSS.n1515 VSS.n141 0.000715048
R4701 VSS.n1504 VSS.n148 0.000715048
R4702 VSS.n1475 VSS.n1473 0.000715048
R4703 VSS.n876 VSS.n742 0.000699968
R4704 VSS.n1321 VSS.n1320 0.000696035
R4705 VSS.n1295 VSS.n1294 0.000696035
R4706 VSS.n566 VSS.n125 0.000696035
R4707 VSS.n491 VSS.n144 0.000696035
R4708 VSS.n525 VSS.n524 0.000696035
R4709 VSS.n1351 VSS.n1344 0.000696035
R4710 VSS.n166 VSS 0.000677021
R4711 VSS.n230 VSS.n229 0.000675054
R4712 VSS.n1443 VSS.n193 0.000651451
R4713 VSS.n1047 VSS.n1046 0.000646417
R4714 VSS.n1011 VSS.n1010 0.000646417
R4715 VSS.n1013 VSS.n631 0.000646417
R4716 VSS.n977 VSS.n976 0.000646417
R4717 VSS.n1081 VSS.n1080 0.000646417
R4718 VSS.n943 VSS.n942 0.000646417
R4719 VSS.n741 VSS.n730 0.000646417
R4720 VSS.n909 VSS.n908 0.000646417
R4721 VSS.n1083 VSS.n722 0.000646417
R4722 VSS.n1352 VSS.n240 0.000642928
R4723 VSS.n1394 VSS.n1389 0.000637683
R4724 VSS VSS.n123 0.000637027
R4725 VSS.n1521 VSS 0.000637027
R4726 VSS VSS.n146 0.000637027
R4727 VSS.n1715 VSS 0.000637027
R4728 VSS.n518 VSS 0.000637027
R4729 VSS.n1463 VSS 0.000637027
R4730 VSS.n1662 VSS 0.000637027
R4731 VSS VSS.n1383 0.000637027
R4732 VSS.n1364 VSS 0.000637027
R4733 VSS.n1109 VSS 0.000634405
R4734 VSS.n1705 VSS 0.000626537
R4735 VSS.n1538 VSS 0.000619325
R4736 VSS.n1628 VSS 0.00061408
R4737 VSS.n251 VSS.n168 0.000606213
R4738 VSS VSS.n565 0.000605557
R4739 VSS.n216 VSS 0.000605557
R4740 VSS.n1482 VSS.n1480 0.000604246
R4741 VSS.n1294 VSS 0.000599001
R4742 VSS.n1389 VSS.n214 0.000594411
R4743 VSS.n1219 VSS.n598 0.00057802
R4744 VSS.n183 VSS.n181 0.000575398
R4745 VSS.n1304 VSS 0.000574087
R4746 VSS.n370 VSS.n240 0.00057212
R4747 VSS.n1304 VSS.n1227 0.000562941
R4748 VSS.n1705 VSS 0.000560318
R4749 VSS.n256 VSS.n255 0.000560318
R4750 VSS.n1515 VSS.n139 0.000556385
R4751 VSS.n1504 VSS.n5 0.000556385
R4752 VSS.n1475 VSS.n166 0.000556385
R4753 VSS.n370 VSS.n66 0.000556385
R4754 VSS.n566 VSS 0.000555729
R4755 VSS VSS.n1310 0.000549173
R4756 VSS.n797 VSS 0.000542616
R4757 VSS.n856 VSS.n855 0.000538027
R4758 VSS.n1695 VSS.n51 0.000537371
R4759 VSS.n1488 VSS 0.00053147
R4760 VSS VSS.n1725 0.000529504
R4761 VSS.n255 VSS.n253 0.000528192
R4762 VSS.n1644 VSS.n1643 0.000526225
R4763 VSS.n499 VSS.n117 0.000521636
R4764 VSS.n1511 VSS.n144 0.000516391
R4765 VSS.n525 VSS.n19 0.000516391
R4766 VSS.n256 VSS.n46 0.000516391
R4767 VSS.n1344 VSS.n76 0.000516391
R4768 VSS.n1650 VSS.n91 0.00051508
R4769 VSS VSS.n183 0.000513768
R4770 VSS.n1443 VSS.n1442 0.000513113
R4771 VSS.n1414 VSS.n206 0.000511146
R4772 VSS.n214 VSS.n206 0.000509179
R4773 VSS.n1310 VSS.n1227 0.000507212
R4774 VSS.n1537 VSS.n123 0.000507212
R4775 VSS.n1521 VSS.n135 0.000507212
R4776 VSS.n1511 VSS.n146 0.000507212
R4777 VSS.n499 VSS.n498 0.000507212
R4778 VSS.n1715 VSS.n19 0.000507212
R4779 VSS.n519 VSS.n518 0.000507212
R4780 VSS.n1695 VSS.n46 0.000507212
R4781 VSS.n1463 VSS.n1462 0.000507212
R4782 VSS.n1662 VSS.n76 0.000507212
R4783 VSS.n1383 VSS.n230 0.000507212
R4784 VSS.n1415 VSS.n1414 0.000507212
R4785 VSS.n1364 VSS.n1363 0.000507212
R4786 VSS.n181 VSS.n179 0.000506556
R4787 VSS.n1415 VSS.n194 0.000506556
R4788 VSS.n1650 VSS.n1649 0.000505245
R4789 VSS.n565 VSS.n544 0.000503934
R4790 VSS.n1483 VSS.n1482 0.000503934
R4791 VSS.n179 VSS.n51 0.000503934
R4792 VSS.n220 VSS.n216 0.000503934
R4793 VSS.n1393 VSS.n91 0.000503934
R4794 VSS.n1644 VSS.n92 0.000503934
R4795 VSS.n557 VSS.n546 0.000501967
R4796 VSS.n1490 VSS.n1489 0.000501967
R4797 VSS.n226 VSS.n224 0.000501967
R4798 VSS.n1394 VSS.n1393 0.000501967
R4799 VSS.n1649 VSS.n92 0.000501967
R4800 VSS.n1643 VSS.n95 0.000501967
R4801 VSS.n1628 VSS.n117 0.000501311
R4802 VSS.n1480 VSS 0.000501311
R4803 VSS.n253 VSS.n251 0.000501311
R4804 VSS.n558 VSS.n544 0.000500656
R4805 VSS.n558 VSS.n557 0.000500656
R4806 VSS.n551 VSS.n546 0.000500656
R4807 VSS.n1483 VSS.n161 0.000500656
R4808 VSS.n1490 VSS.n161 0.000500656
R4809 VSS.n1489 VSS.n1488 0.000500656
R4810 VSS.n222 VSS.n220 0.000500656
R4811 VSS.n224 VSS.n222 0.000500656
R4812 VSS.n229 VSS.n226 0.000500656
R4813 VSS.n1442 VSS.n194 0.000500656
R4814 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t22 491.64
R4815 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t21 491.64
R4816 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t19 491.64
R4817 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t18 491.64
R4818 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t14 485.221
R4819 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t17 367.928
R4820 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t12 255.588
R4821 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t15 224.478
R4822 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t16 213.688
R4823 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n0 209.19
R4824 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t13 139.78
R4825 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t20 139.78
R4826 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t23 139.78
R4827 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n10 120.999
R4828 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n9 120.999
R4829 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n22 104.489
R4830 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n12 92.5005
R4831 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n18 86.2638
R4832 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n17 85.8873
R4833 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n15 85.724
R4834 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n7 84.5046
R4835 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n23 83.8907
R4836 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n20 75.0672
R4837 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n17 75.0672
R4838 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n19 73.1255
R4839 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n17 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n16 73.1255
R4840 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n15 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n14 73.1255
R4841 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n6 72.3005
R4842 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n15 68.8946
R4843 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n8 60.9797
R4844 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n13 41.9827
R4845 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t2 30.462
R4846 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t10 30.462
R4847 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t8 30.462
R4848 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t7 30.462
R4849 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t1 30.462
R4850 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t0 30.462
R4851 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n11 28.124
R4852 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n5 19.963
R4853 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n1 17.8661
R4854 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n2 17.8661
R4855 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n3 17.1217
R4856 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t5 11.8205
R4857 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t4 11.8205
R4858 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t11 11.8205
R4859 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t9 11.8205
R4860 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t3 11.8205
R4861 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t6 11.8205
R4862 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n21 9.3005
R4863 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n4 1.8615
R4864 a_n10081_1406.n0 a_n10081_1406.t3 539.788
R4865 a_n10081_1406.n1 a_n10081_1406.t5 531.496
R4866 a_n10081_1406.n0 a_n10081_1406.t6 490.034
R4867 a_n10081_1406.n5 a_n10081_1406.t0 283.788
R4868 a_n10081_1406.t1 a_n10081_1406.n5 205.489
R4869 a_n10081_1406.n2 a_n10081_1406.t7 182.625
R4870 a_n10081_1406.n3 a_n10081_1406.t2 179.054
R4871 a_n10081_1406.n2 a_n10081_1406.t4 139.78
R4872 a_n10081_1406.n4 a_n10081_1406.n3 101.368
R4873 a_n10081_1406.n5 a_n10081_1406.n4 77.9135
R4874 a_n10081_1406.n4 a_n10081_1406.n1 76.1557
R4875 a_n10081_1406.n1 a_n10081_1406.n0 8.29297
R4876 a_n10081_1406.n3 a_n10081_1406.n2 3.57087
R4877 SEL0.n176 SEL0.t93 933.563
R4878 SEL0.n173 SEL0.t103 933.563
R4879 SEL0.n183 SEL0.t51 933.563
R4880 SEL0.n180 SEL0.t18 933.563
R4881 SEL0.n154 SEL0.t100 933.563
R4882 SEL0.n151 SEL0.t118 933.563
R4883 SEL0.n161 SEL0.t61 933.563
R4884 SEL0.n158 SEL0.t30 933.563
R4885 SEL0.n132 SEL0.t106 933.563
R4886 SEL0.n129 SEL0.t101 933.563
R4887 SEL0.n139 SEL0.t36 933.563
R4888 SEL0.n136 SEL0.t116 933.563
R4889 SEL0.n110 SEL0.t48 933.563
R4890 SEL0.n107 SEL0.t41 933.563
R4891 SEL0.n117 SEL0.t95 933.563
R4892 SEL0.n114 SEL0.t45 933.563
R4893 SEL0.n88 SEL0.t43 933.563
R4894 SEL0.n85 SEL0.t34 933.563
R4895 SEL0.n95 SEL0.t137 933.563
R4896 SEL0.n92 SEL0.t81 933.563
R4897 SEL0.n66 SEL0.t2 933.563
R4898 SEL0.n63 SEL0.t140 933.563
R4899 SEL0.n73 SEL0.t73 933.563
R4900 SEL0.n70 SEL0.t10 933.563
R4901 SEL0.n45 SEL0.t14 933.563
R4902 SEL0.n42 SEL0.t6 933.563
R4903 SEL0.n52 SEL0.t98 933.563
R4904 SEL0.n49 SEL0.t52 933.563
R4905 SEL0.n24 SEL0.t109 933.563
R4906 SEL0.n21 SEL0.t102 933.563
R4907 SEL0.n31 SEL0.t75 933.563
R4908 SEL0.n28 SEL0.t15 933.563
R4909 SEL0.n4 SEL0.t64 933.563
R4910 SEL0.n1 SEL0.t94 933.563
R4911 SEL0.n11 SEL0.t50 933.563
R4912 SEL0.n8 SEL0.t99 933.563
R4913 SEL0.n189 SEL0.t114 385.697
R4914 SEL0.n167 SEL0.t117 385.697
R4915 SEL0.n145 SEL0.t13 385.697
R4916 SEL0.n123 SEL0.t86 385.697
R4917 SEL0.n101 SEL0.t53 385.697
R4918 SEL0.n79 SEL0.t88 385.697
R4919 SEL0.n58 SEL0.t19 385.697
R4920 SEL0.n37 SEL0.t7 385.697
R4921 SEL0.n17 SEL0.t110 385.697
R4922 SEL0.n176 SEL0.t112 367.635
R4923 SEL0.n173 SEL0.t54 367.635
R4924 SEL0.n183 SEL0.t119 367.635
R4925 SEL0.n180 SEL0.t4 367.635
R4926 SEL0.n154 SEL0.t89 367.635
R4927 SEL0.n151 SEL0.t22 367.635
R4928 SEL0.n161 SEL0.t91 367.635
R4929 SEL0.n158 SEL0.t113 367.635
R4930 SEL0.n132 SEL0.t71 367.635
R4931 SEL0.n129 SEL0.t123 367.635
R4932 SEL0.n139 SEL0.t79 367.635
R4933 SEL0.n136 SEL0.t47 367.635
R4934 SEL0.n110 SEL0.t139 367.635
R4935 SEL0.n107 SEL0.t59 367.635
R4936 SEL0.n117 SEL0.t142 367.635
R4937 SEL0.n114 SEL0.t9 367.635
R4938 SEL0.n88 SEL0.t96 367.635
R4939 SEL0.n85 SEL0.t17 367.635
R4940 SEL0.n95 SEL0.t1 367.635
R4941 SEL0.n92 SEL0.t11 367.635
R4942 SEL0.n66 SEL0.t141 367.635
R4943 SEL0.n63 SEL0.t63 367.635
R4944 SEL0.n73 SEL0.t105 367.635
R4945 SEL0.n70 SEL0.t122 367.635
R4946 SEL0.n45 SEL0.t67 367.635
R4947 SEL0.n42 SEL0.t111 367.635
R4948 SEL0.n52 SEL0.t3 367.635
R4949 SEL0.n49 SEL0.t16 367.635
R4950 SEL0.n24 SEL0.t74 367.635
R4951 SEL0.n21 SEL0.t126 367.635
R4952 SEL0.n31 SEL0.t107 367.635
R4953 SEL0.n28 SEL0.t85 367.635
R4954 SEL0.n4 SEL0.t55 367.635
R4955 SEL0.n1 SEL0.t25 367.635
R4956 SEL0.n11 SEL0.t49 367.635
R4957 SEL0.n8 SEL0.t143 367.635
R4958 SEL0.n177 SEL0.t72 308.481
R4959 SEL0.n174 SEL0.t39 308.481
R4960 SEL0.n184 SEL0.t76 308.481
R4961 SEL0.n181 SEL0.t133 308.481
R4962 SEL0.n155 SEL0.t38 308.481
R4963 SEL0.n152 SEL0.t0 308.481
R4964 SEL0.n162 SEL0.t44 308.481
R4965 SEL0.n159 SEL0.t97 308.481
R4966 SEL0.n133 SEL0.t121 308.481
R4967 SEL0.n130 SEL0.t130 308.481
R4968 SEL0.n140 SEL0.t135 308.481
R4969 SEL0.n137 SEL0.t56 308.481
R4970 SEL0.n111 SEL0.t58 308.481
R4971 SEL0.n108 SEL0.t69 308.481
R4972 SEL0.n118 SEL0.t62 308.481
R4973 SEL0.n115 SEL0.t21 308.481
R4974 SEL0.n89 SEL0.t12 308.481
R4975 SEL0.n86 SEL0.t28 308.481
R4976 SEL0.n96 SEL0.t66 308.481
R4977 SEL0.n93 SEL0.t24 308.481
R4978 SEL0.n67 SEL0.t60 308.481
R4979 SEL0.n64 SEL0.t70 308.481
R4980 SEL0.n74 SEL0.t29 308.481
R4981 SEL0.n71 SEL0.t129 308.481
R4982 SEL0.n46 SEL0.t108 308.481
R4983 SEL0.n43 SEL0.t125 308.481
R4984 SEL0.n53 SEL0.t68 308.481
R4985 SEL0.n50 SEL0.t27 308.481
R4986 SEL0.n25 SEL0.t124 308.481
R4987 SEL0.n22 SEL0.t132 308.481
R4988 SEL0.n32 SEL0.t32 308.481
R4989 SEL0.n29 SEL0.t90 308.481
R4990 SEL0.n5 SEL0.t115 308.481
R4991 SEL0.n2 SEL0.t57 308.481
R4992 SEL0.n12 SEL0.t138 308.481
R4993 SEL0.n9 SEL0.t23 308.481
R4994 SEL0.n172 SEL0.t136 291.829
R4995 SEL0.n172 SEL0.t46 291.829
R4996 SEL0.n150 SEL0.t104 291.829
R4997 SEL0.n150 SEL0.t26 291.829
R4998 SEL0.n128 SEL0.t31 291.829
R4999 SEL0.n128 SEL0.t82 291.829
R5000 SEL0.n106 SEL0.t5 291.829
R5001 SEL0.n106 SEL0.t65 291.829
R5002 SEL0.n84 SEL0.t33 291.829
R5003 SEL0.n84 SEL0.t134 291.829
R5004 SEL0.n62 SEL0.t77 291.829
R5005 SEL0.n62 SEL0.t127 291.829
R5006 SEL0.n41 SEL0.t37 291.829
R5007 SEL0.n41 SEL0.t92 291.829
R5008 SEL0.n20 SEL0.t78 291.829
R5009 SEL0.n20 SEL0.t128 291.829
R5010 SEL0.n0 SEL0.t40 291.829
R5011 SEL0.n0 SEL0.t87 291.829
R5012 SEL0.n172 SEL0.t42 221.72
R5013 SEL0.n150 SEL0.t20 221.72
R5014 SEL0.n128 SEL0.t35 221.72
R5015 SEL0.n106 SEL0.t8 221.72
R5016 SEL0.n84 SEL0.t80 221.72
R5017 SEL0.n62 SEL0.t120 221.72
R5018 SEL0.n41 SEL0.t83 221.72
R5019 SEL0.n20 SEL0.t84 221.72
R5020 SEL0.n0 SEL0.t131 221.72
R5021 SEL0.n182 SEL0.n181 161.607
R5022 SEL0.n160 SEL0.n159 161.607
R5023 SEL0.n138 SEL0.n137 161.607
R5024 SEL0.n116 SEL0.n115 161.607
R5025 SEL0.n94 SEL0.n93 161.607
R5026 SEL0.n72 SEL0.n71 161.607
R5027 SEL0.n51 SEL0.n50 161.607
R5028 SEL0.n30 SEL0.n29 161.607
R5029 SEL0.n10 SEL0.n9 161.607
R5030 SEL0.n185 SEL0.n184 161.606
R5031 SEL0.n163 SEL0.n162 161.606
R5032 SEL0.n141 SEL0.n140 161.606
R5033 SEL0.n119 SEL0.n118 161.606
R5034 SEL0.n97 SEL0.n96 161.606
R5035 SEL0.n75 SEL0.n74 161.606
R5036 SEL0.n54 SEL0.n53 161.606
R5037 SEL0.n33 SEL0.n32 161.606
R5038 SEL0.n13 SEL0.n12 161.606
R5039 SEL0.n178 SEL0.n177 161.599
R5040 SEL0.n156 SEL0.n155 161.599
R5041 SEL0.n134 SEL0.n133 161.599
R5042 SEL0.n112 SEL0.n111 161.599
R5043 SEL0.n90 SEL0.n89 161.599
R5044 SEL0.n68 SEL0.n67 161.599
R5045 SEL0.n47 SEL0.n46 161.599
R5046 SEL0.n26 SEL0.n25 161.599
R5047 SEL0.n6 SEL0.n5 161.599
R5048 SEL0.n175 SEL0.n174 161.579
R5049 SEL0.n153 SEL0.n152 161.579
R5050 SEL0.n131 SEL0.n130 161.579
R5051 SEL0.n109 SEL0.n108 161.579
R5052 SEL0.n87 SEL0.n86 161.579
R5053 SEL0.n65 SEL0.n64 161.579
R5054 SEL0.n44 SEL0.n43 161.579
R5055 SEL0.n23 SEL0.n22 161.579
R5056 SEL0.n3 SEL0.n2 161.579
R5057 SEL0.n190 SEL0.n189 89.6005
R5058 SEL0.n168 SEL0.n167 89.6005
R5059 SEL0.n146 SEL0.n145 89.6005
R5060 SEL0.n124 SEL0.n123 89.6005
R5061 SEL0.n102 SEL0.n101 89.6005
R5062 SEL0.n80 SEL0.n79 89.6005
R5063 SEL0.n59 SEL0.n58 89.6005
R5064 SEL0.n38 SEL0.n37 89.6005
R5065 SEL0.n18 SEL0.n17 89.6005
R5066 SEL0.n190 SEL0.n172 50.6672
R5067 SEL0.n168 SEL0.n150 50.6672
R5068 SEL0.n146 SEL0.n128 50.6672
R5069 SEL0.n124 SEL0.n106 50.6672
R5070 SEL0.n102 SEL0.n84 50.6672
R5071 SEL0.n80 SEL0.n62 50.6672
R5072 SEL0.n59 SEL0.n41 50.6672
R5073 SEL0.n38 SEL0.n20 50.6672
R5074 SEL0.n18 SEL0.n0 50.6672
R5075 SEL0.n186 SEL0.n182 13.8557
R5076 SEL0.n164 SEL0.n160 13.8557
R5077 SEL0.n142 SEL0.n138 13.8557
R5078 SEL0.n120 SEL0.n116 13.8557
R5079 SEL0.n98 SEL0.n94 13.8557
R5080 SEL0.n76 SEL0.n72 13.8557
R5081 SEL0.n55 SEL0.n51 13.8557
R5082 SEL0.n34 SEL0.n30 13.8557
R5083 SEL0.n14 SEL0.n10 13.8557
R5084 SEL0.n188 SEL0.n187 13.8507
R5085 SEL0.n166 SEL0.n165 13.8507
R5086 SEL0.n144 SEL0.n143 13.8507
R5087 SEL0.n122 SEL0.n121 13.8507
R5088 SEL0.n100 SEL0.n99 13.8507
R5089 SEL0.n78 SEL0.n77 13.8507
R5090 SEL0.n57 SEL0.n56 13.8507
R5091 SEL0.n36 SEL0.n35 13.8507
R5092 SEL0.n16 SEL0.n15 13.8507
R5093 SEL0.n179 SEL0.n175 13.6141
R5094 SEL0.n157 SEL0.n153 13.6141
R5095 SEL0.n135 SEL0.n131 13.6141
R5096 SEL0.n113 SEL0.n109 13.6141
R5097 SEL0.n91 SEL0.n87 13.6141
R5098 SEL0.n69 SEL0.n65 13.6141
R5099 SEL0.n48 SEL0.n44 13.6141
R5100 SEL0.n27 SEL0.n23 13.6141
R5101 SEL0.n7 SEL0.n3 13.6141
R5102 SEL0.n179 SEL0.n178 12.6478
R5103 SEL0.n157 SEL0.n156 12.6478
R5104 SEL0.n135 SEL0.n134 12.6478
R5105 SEL0.n113 SEL0.n112 12.6478
R5106 SEL0.n91 SEL0.n90 12.6478
R5107 SEL0.n69 SEL0.n68 12.6478
R5108 SEL0.n48 SEL0.n47 12.6478
R5109 SEL0.n27 SEL0.n26 12.6478
R5110 SEL0.n7 SEL0.n6 12.6478
R5111 SEL0.n186 SEL0.n185 12.4772
R5112 SEL0.n164 SEL0.n163 12.4772
R5113 SEL0.n142 SEL0.n141 12.4772
R5114 SEL0.n120 SEL0.n119 12.4772
R5115 SEL0.n98 SEL0.n97 12.4772
R5116 SEL0.n76 SEL0.n75 12.4772
R5117 SEL0.n55 SEL0.n54 12.4772
R5118 SEL0.n34 SEL0.n33 12.4772
R5119 SEL0.n14 SEL0.n13 12.4772
R5120 SEL0.n177 SEL0.n176 10.955
R5121 SEL0.n174 SEL0.n173 10.955
R5122 SEL0.n184 SEL0.n183 10.955
R5123 SEL0.n181 SEL0.n180 10.955
R5124 SEL0.n155 SEL0.n154 10.955
R5125 SEL0.n152 SEL0.n151 10.955
R5126 SEL0.n162 SEL0.n161 10.955
R5127 SEL0.n159 SEL0.n158 10.955
R5128 SEL0.n133 SEL0.n132 10.955
R5129 SEL0.n130 SEL0.n129 10.955
R5130 SEL0.n140 SEL0.n139 10.955
R5131 SEL0.n137 SEL0.n136 10.955
R5132 SEL0.n111 SEL0.n110 10.955
R5133 SEL0.n108 SEL0.n107 10.955
R5134 SEL0.n118 SEL0.n117 10.955
R5135 SEL0.n115 SEL0.n114 10.955
R5136 SEL0.n89 SEL0.n88 10.955
R5137 SEL0.n86 SEL0.n85 10.955
R5138 SEL0.n96 SEL0.n95 10.955
R5139 SEL0.n93 SEL0.n92 10.955
R5140 SEL0.n67 SEL0.n66 10.955
R5141 SEL0.n64 SEL0.n63 10.955
R5142 SEL0.n74 SEL0.n73 10.955
R5143 SEL0.n71 SEL0.n70 10.955
R5144 SEL0.n46 SEL0.n45 10.955
R5145 SEL0.n43 SEL0.n42 10.955
R5146 SEL0.n53 SEL0.n52 10.955
R5147 SEL0.n50 SEL0.n49 10.955
R5148 SEL0.n25 SEL0.n24 10.955
R5149 SEL0.n22 SEL0.n21 10.955
R5150 SEL0.n32 SEL0.n31 10.955
R5151 SEL0.n29 SEL0.n28 10.955
R5152 SEL0.n5 SEL0.n4 10.955
R5153 SEL0.n2 SEL0.n1 10.955
R5154 SEL0.n12 SEL0.n11 10.955
R5155 SEL0.n9 SEL0.n8 10.955
R5156 SEL0 SEL0.n60 9.59074
R5157 SEL0.n126 SEL0.n125 9.56176
R5158 SEL0.n40 SEL0.n39 9.54908
R5159 SEL0.n194 SEL0.n19 9.5364
R5160 SEL0.n82 SEL0.n81 9.52224
R5161 SEL0.n192 SEL0.n191 9.5219
R5162 SEL0.n104 SEL0.n103 9.5219
R5163 SEL0.n148 SEL0.n147 9.51647
R5164 SEL0.n170 SEL0.n169 9.51103
R5165 SEL0.n189 SEL0.n188 9.3005
R5166 SEL0.n167 SEL0.n166 9.3005
R5167 SEL0.n145 SEL0.n144 9.3005
R5168 SEL0.n123 SEL0.n122 9.3005
R5169 SEL0.n101 SEL0.n100 9.3005
R5170 SEL0.n79 SEL0.n78 9.3005
R5171 SEL0.n58 SEL0.n57 9.3005
R5172 SEL0.n37 SEL0.n36 9.3005
R5173 SEL0.n17 SEL0.n16 9.3005
R5174 SEL0.n61 SEL0.n40 6.81149
R5175 SEL0.n194 SEL0.n193 6.80812
R5176 SEL0.n171 SEL0.n149 3.42946
R5177 SEL0.n61 SEL0 3.41775
R5178 SEL0.n83 SEL0.n82 3.4105
R5179 SEL0.n105 SEL0.n104 3.4105
R5180 SEL0.n127 SEL0.n126 3.4105
R5181 SEL0.n149 SEL0.n148 3.4105
R5182 SEL0.n171 SEL0.n170 3.4105
R5183 SEL0.n193 SEL0.n192 3.4105
R5184 SEL0.n127 SEL0.n105 3.38859
R5185 SEL0.n83 SEL0.n61 3.36815
R5186 SEL0.n149 SEL0.n127 3.34499
R5187 SEL0.n105 SEL0.n83 3.34227
R5188 SEL0.n193 SEL0.n171 3.29391
R5189 SEL0.n191 SEL0.n190 3.1005
R5190 SEL0.n169 SEL0.n168 3.1005
R5191 SEL0.n147 SEL0.n146 3.1005
R5192 SEL0.n125 SEL0.n124 3.1005
R5193 SEL0.n103 SEL0.n102 3.1005
R5194 SEL0.n81 SEL0.n80 3.1005
R5195 SEL0.n60 SEL0.n59 3.1005
R5196 SEL0.n39 SEL0.n38 3.1005
R5197 SEL0.n19 SEL0.n18 3.1005
R5198 SEL0.n187 SEL0.n186 3.01361
R5199 SEL0.n165 SEL0.n164 3.01361
R5200 SEL0.n143 SEL0.n142 3.01361
R5201 SEL0.n121 SEL0.n120 3.01361
R5202 SEL0.n99 SEL0.n98 3.01361
R5203 SEL0.n77 SEL0.n76 3.01361
R5204 SEL0.n56 SEL0.n55 3.01361
R5205 SEL0.n35 SEL0.n34 3.01361
R5206 SEL0.n15 SEL0.n14 3.01361
R5207 SEL0.n187 SEL0.n179 1.42612
R5208 SEL0.n165 SEL0.n157 1.42612
R5209 SEL0.n143 SEL0.n135 1.42612
R5210 SEL0.n121 SEL0.n113 1.42612
R5211 SEL0.n99 SEL0.n91 1.42612
R5212 SEL0.n77 SEL0.n69 1.42612
R5213 SEL0.n56 SEL0.n48 1.42612
R5214 SEL0.n35 SEL0.n27 1.42612
R5215 SEL0.n15 SEL0.n7 1.42612
R5216 SEL0.n175 SEL0 0.593405
R5217 SEL0.n153 SEL0 0.593405
R5218 SEL0.n131 SEL0 0.593405
R5219 SEL0.n109 SEL0 0.593405
R5220 SEL0.n87 SEL0 0.593405
R5221 SEL0.n65 SEL0 0.593405
R5222 SEL0.n44 SEL0 0.593405
R5223 SEL0.n23 SEL0 0.593405
R5224 SEL0.n3 SEL0 0.593405
R5225 SEL0.n178 SEL0 0.574824
R5226 SEL0.n156 SEL0 0.574824
R5227 SEL0.n134 SEL0 0.574824
R5228 SEL0.n112 SEL0 0.574824
R5229 SEL0.n90 SEL0 0.574824
R5230 SEL0.n68 SEL0 0.574824
R5231 SEL0.n47 SEL0 0.574824
R5232 SEL0.n26 SEL0 0.574824
R5233 SEL0.n6 SEL0 0.574824
R5234 SEL0.n185 SEL0 0.568068
R5235 SEL0.n163 SEL0 0.568068
R5236 SEL0.n141 SEL0 0.568068
R5237 SEL0.n119 SEL0 0.568068
R5238 SEL0.n97 SEL0 0.568068
R5239 SEL0.n75 SEL0 0.568068
R5240 SEL0.n54 SEL0 0.568068
R5241 SEL0.n33 SEL0 0.568068
R5242 SEL0.n13 SEL0 0.568068
R5243 SEL0.n182 SEL0 0.567223
R5244 SEL0.n160 SEL0 0.567223
R5245 SEL0.n138 SEL0 0.567223
R5246 SEL0.n116 SEL0 0.567223
R5247 SEL0.n94 SEL0 0.567223
R5248 SEL0.n72 SEL0 0.567223
R5249 SEL0.n51 SEL0 0.567223
R5250 SEL0.n30 SEL0 0.567223
R5251 SEL0.n10 SEL0 0.567223
R5252 SEL0.n188 SEL0 0.397239
R5253 SEL0.n166 SEL0 0.397239
R5254 SEL0.n144 SEL0 0.397239
R5255 SEL0.n122 SEL0 0.397239
R5256 SEL0.n100 SEL0 0.397239
R5257 SEL0.n78 SEL0 0.397239
R5258 SEL0.n57 SEL0 0.397239
R5259 SEL0.n36 SEL0 0.397239
R5260 SEL0.n16 SEL0 0.397239
R5261 SEL0.n191 SEL0 0.237819
R5262 SEL0.n169 SEL0 0.237819
R5263 SEL0.n147 SEL0 0.237819
R5264 SEL0.n125 SEL0 0.237819
R5265 SEL0.n103 SEL0 0.237819
R5266 SEL0.n81 SEL0 0.237819
R5267 SEL0.n60 SEL0 0.237819
R5268 SEL0.n39 SEL0 0.237819
R5269 SEL0.n19 SEL0 0.237819
R5270 SEL0.n170 SEL0 0.0802101
R5271 SEL0.n148 SEL0 0.0747754
R5272 SEL0.n192 SEL0 0.0693406
R5273 SEL0.n104 SEL0 0.0693406
R5274 SEL0.n40 SEL0 0.0421667
R5275 SEL0.n126 SEL0 0.0294855
R5276 SEL0 SEL0.n194 0.0276739
R5277 SEL0.n82 SEL0 0.0149928
R5278 VDD.n1063 VDD.t1519 15549.3
R5279 VDD.n934 VDD.t3918 15549.3
R5280 VDD.n805 VDD.t3456 15549.3
R5281 VDD.n654 VDD.t1316 15549.3
R5282 VDD.n525 VDD.t2545 15549.3
R5283 VDD.n396 VDD.t2706 15549.3
R5284 VDD.n267 VDD.t1691 15549.3
R5285 VDD.n129 VDD.t1101 15549.3
R5286 VDD.n2913 VDD.t3292 15549.3
R5287 VDD.t1026 VDD.n2400 2135.7
R5288 VDD.t2300 VDD.t3568 1823.03
R5289 VDD.t2318 VDD.t269 1811.88
R5290 VDD.t889 VDD.t2830 1806.46
R5291 VDD.t4194 VDD.t595 1663.3
R5292 VDD.n2382 VDD.t1021 1648.11
R5293 VDD.t989 VDD.n2407 1613.92
R5294 VDD.t2199 VDD.t2153 1612.38
R5295 VDD.t2320 VDD.t257 1596.32
R5296 VDD.t1633 VDD.t2126 1564.05
R5297 VDD.t4239 VDD.t1024 1547.34
R5298 VDD.t4004 VDD.t1076 1498.08
R5299 VDD.t1695 VDD.t1892 1498.08
R5300 VDD.t2074 VDD.t152 1498.08
R5301 VDD.t2503 VDD.t3681 1498.08
R5302 VDD.t3279 VDD.t4040 1498.08
R5303 VDD.t4030 VDD.t573 1498.08
R5304 VDD.t712 VDD.t283 1498.08
R5305 VDD.t1336 VDD.t117 1498.08
R5306 VDD.t2909 VDD.t722 1498.08
R5307 VDD.t1327 VDD.t2084 1498.08
R5308 VDD.t447 VDD.t4138 1498.08
R5309 VDD.t908 VDD.t611 1498.08
R5310 VDD.t1435 VDD.t2700 1498.08
R5311 VDD.t2472 VDD.t2880 1498.08
R5312 VDD.t3240 VDD.t1840 1498.08
R5313 VDD.t337 VDD.t2189 1496.25
R5314 VDD.t3592 VDD.t397 1493.96
R5315 VDD.t3579 VDD.t376 1469.88
R5316 VDD.t2288 VDD.t3539 1456.41
R5317 VDD.t897 VDD.t2843 1444.55
R5318 VDD.t479 VDD.t4073 1412.88
R5319 VDD.t2592 VDD.t4116 1366.39
R5320 VDD.t3524 VDD.t3395 1149.13
R5321 VDD.t2020 VDD.t4008 1149.13
R5322 VDD.t1283 VDD.t2443 1149.13
R5323 VDD.t3322 VDD.t3659 1149.13
R5324 VDD.t1592 VDD.t3192 1149.13
R5325 VDD.t3895 VDD.t103 1149.13
R5326 VDD.t668 VDD.t20 1149.13
R5327 VDD.t2250 VDD.t4243 1149.13
R5328 VDD.t2056 VDD.t1293 1149.13
R5329 VDD.t4181 VDD.t2314 1149.13
R5330 VDD.t243 VDD.t449 1149.13
R5331 VDD.t496 VDD.t1609 1149.13
R5332 VDD.t2256 VDD.t2223 1149.13
R5333 VDD.t748 VDD.t4206 1149.13
R5334 VDD.t2466 VDD.t265 1149.13
R5335 VDD.t1562 VDD.t4105 1149.13
R5336 VDD.t299 VDD.t1625 1149.13
R5337 VDD.t3908 VDD.t403 1149.13
R5338 VDD.t2405 VDD.t2836 1149.13
R5339 VDD.t3475 VDD.t3432 1149.13
R5340 VDD.t2982 VDD.n1021 858.129
R5341 VDD.n1017 VDD.t4353 858.129
R5342 VDD.t3001 VDD.n892 858.129
R5343 VDD.n888 VDD.t4373 858.129
R5344 VDD.t3026 VDD.n763 858.129
R5345 VDD.n759 VDD.t4448 858.129
R5346 VDD.t2937 VDD.n612 858.129
R5347 VDD.n608 VDD.t4355 858.129
R5348 VDD.t2951 VDD.n483 858.129
R5349 VDD.n479 VDD.t4345 858.129
R5350 VDD.t2988 VDD.n354 858.129
R5351 VDD.n350 VDD.t4357 858.129
R5352 VDD.t2949 VDD.n225 858.129
R5353 VDD.n221 VDD.t4347 858.129
R5354 VDD.t2933 VDD.n87 858.129
R5355 VDD.n83 VDD.t4409 858.129
R5356 VDD.t2943 VDD.n25 858.129
R5357 VDD.n21 VDD.t4405 858.129
R5358 VDD.t560 VDD.t2423 851.116
R5359 VDD.n1136 VDD.t3496 769.712
R5360 VDD.t868 VDD.t1928 734.423
R5361 VDD.t3409 VDD.t2784 734.423
R5362 VDD.t836 VDD.t1464 734.423
R5363 VDD.t965 VDD.t944 734.423
R5364 VDD.t1966 VDD.t2215 734.423
R5365 VDD.t4269 VDD.t4291 734.423
R5366 VDD.t4048 VDD.t3669 734.423
R5367 VDD.t142 VDD.t4148 734.423
R5368 VDD.t1910 VDD.t2246 734.423
R5369 VDD.t217 VDD.t2519 734.423
R5370 VDD.t1082 VDD.t700 734.423
R5371 VDD.t2561 VDD.t4329 734.423
R5372 VDD.t1775 VDD.t3401 734.423
R5373 VDD.t805 VDD.t1358 734.423
R5374 VDD.t94 VDD.t3324 734.423
R5375 VDD.t1858 VDD.t1733 734.423
R5376 VDD.t3940 VDD.t3994 734.423
R5377 VDD.t1847 VDD.t2756 734.423
R5378 VDD.t1119 VDD.t1584 734.423
R5379 VDD.t170 VDD.t2692 734.423
R5380 VDD.t4273 VDD.t4081 711.524
R5381 VDD.t2077 VDD.t4223 709.568
R5382 VDD.t162 VDD.t2234 687.312
R5383 VDD.t1157 VDD.t4087 663.92
R5384 VDD.n2219 VDD.t3558 662.178
R5385 VDD.t321 VDD.n2242 662.178
R5386 VDD.n1881 VDD.t1573 662.178
R5387 VDD.t824 VDD.n1859 656
R5388 VDD.t4210 VDD.t1056 653.125
R5389 VDD.n1062 VDD.n1061 651.75
R5390 VDD.n933 VDD.n932 651.75
R5391 VDD.n804 VDD.n803 651.75
R5392 VDD.n653 VDD.n652 651.75
R5393 VDD.n524 VDD.n523 651.75
R5394 VDD.n395 VDD.n394 651.75
R5395 VDD.n266 VDD.n265 651.75
R5396 VDD.n128 VDD.n127 651.75
R5397 VDD.n2912 VDD.n2911 651.75
R5398 VDD.t2368 VDD.t439 638.008
R5399 VDD.t3930 VDD.t4186 636.255
R5400 VDD.t725 VDD.t2136 636.255
R5401 VDD.n675 VDD.t1475 636.122
R5402 VDD.t1086 VDD.t2598 634.503
R5403 VDD.t553 VDD.t236 633.333
R5404 VDD.t3147 VDD.t4217 630.996
R5405 VDD.t2632 VDD.t2174 629.245
R5406 VDD.t811 VDD.t2585 629.245
R5407 VDD.t2620 VDD.t4068 627.491
R5408 VDD.t2683 VDD.t4111 622.232
R5409 VDD.t1125 VDD.t2335 616.308
R5410 VDD.n1886 VDD.t1354 607.301
R5411 VDD.t1165 VDD.n2217 591.591
R5412 VDD.t785 VDD.n2239 591.591
R5413 VDD.t3484 VDD.n1883 591.591
R5414 VDD.t291 VDD.t215 513.063
R5415 VDD.t1342 VDD.t3988 513.063
R5416 VDD.t2911 VDD.t2559 513.063
R5417 VDD.t1074 VDD.t2780 513.063
R5418 VDD.t1898 VDD.t832 513.063
R5419 VDD.t940 VDD.t150 513.063
R5420 VDD.t4289 VDD.t2509 513.063
R5421 VDD.t3667 VDD.t3494 513.063
R5422 VDD.t4032 VDD.t4160 513.063
R5423 VDD.t2086 VDD.t2626 513.063
R5424 VDD.t4146 VDD.t92 513.063
R5425 VDD.t619 VDD.t3948 513.063
R5426 VDD.t2752 VDD.t1425 513.063
R5427 VDD.t2884 VDD.t1115 513.063
R5428 VDD.t1876 VDD.t3244 513.063
R5429 VDD.t1727 VDD.t876 512.02
R5430 VDD.t3423 VDD.t978 489.522
R5431 VDD.t872 VDD.t1376 456
R5432 VDD.t2382 VDD.t3834 455.209
R5433 VDD.t1248 VDD.t3783 455.209
R5434 VDD.t3397 VDD.t3755 455.209
R5435 VDD.t1864 VDD.t3866 455.209
R5436 VDD.t1486 VDD.t3868 455.209
R5437 VDD.t1567 VDD.t3805 455.209
R5438 VDD.t1860 VDD.t3874 455.209
R5439 VDD.t357 VDD.t3809 455.209
R5440 VDD.t1683 VDD.t3870 455.209
R5441 VDD.t793 VDD.t3174 449.49
R5442 VDD.t435 VDD.t2804 449.49
R5443 VDD.t2792 VDD.t131 449.49
R5444 VDD.t502 VDD.t3139 449.49
R5445 VDD.t1232 VDD.t1509 449.49
R5446 VDD.t506 VDD.t427 449.49
R5447 VDD.t579 VDD.t1717 449.49
R5448 VDD.t1914 VDD.t2901 449.49
R5449 VDD.t1372 VDD.t2041 436.175
R5450 VDD.t3710 VDD.t1060 435.418
R5451 VDD.t3850 VDD.t625 435.418
R5452 VDD.t3742 VDD.t1138 435.418
R5453 VDD.t3823 VDD.t1620 435.418
R5454 VDD.t3825 VDD.t174 435.418
R5455 VDD.t3772 VDD.t2111 435.418
R5456 VDD.t3829 VDD.t1064 435.418
R5457 VDD.t3778 VDD.t279 435.418
R5458 VDD.t3819 VDD.t2511 435.418
R5459 VDD.t3178 VDD.t950 434.663
R5460 VDD.t2800 VDD.t1490 434.663
R5461 VDD.t127 VDD.t409 434.663
R5462 VDD.t3135 VDD.t148 434.663
R5463 VDD.t1505 VDD.t3143 434.663
R5464 VDD.t423 VDD.t1222 434.663
R5465 VDD.t1705 VDD.t880 434.663
R5466 VDD.t2899 VDD.t1920 434.663
R5467 VDD.t3347 VDD.t1382 427.913
R5468 VDD.t3695 VDD.t3746 427.171
R5469 VDD.t64 VDD.t3718 427.171
R5470 VDD.t1209 VDD.t3716 427.171
R5471 VDD.t43 VDD.t3848 427.171
R5472 VDD.t4130 VDD.t3856 427.171
R5473 VDD.t1201 VDD.t3799 427.171
R5474 VDD.t3990 VDD.t3862 427.171
R5475 VDD.t3265 VDD.t3748 427.171
R5476 VDD.t1950 VDD.t3785 427.171
R5477 VDD.t1532 VDD.t3170 426.43
R5478 VDD.t2 VDD.t2810 426.43
R5479 VDD.t239 VDD.t121 426.43
R5480 VDD.t605 VDD.t3129 426.43
R5481 VDD.t1497 VDD.t1515 426.43
R5482 VDD.t3306 VDD.t433 426.43
R5483 VDD.t3357 VDD.t1713 426.43
R5484 VDD.t1580 VDD.t2891 426.43
R5485 VDD.t3413 VDD.t1366 421.305
R5486 VDD.t1323 VDD.t809 420.978
R5487 VDD.t1350 VDD.t2209 420.978
R5488 VDD.t3353 VDD.t1725 420.978
R5489 VDD.t4167 VDD.t3573 420.978
R5490 VDD.t232 VDD.t3956 420.978
R5491 VDD.t47 VDD.t51 420.978
R5492 VDD.t2569 VDD.t2282 420.978
R5493 VDD.t2064 VDD.t415 420.978
R5494 VDD.t1501 VDD.t1964 420.978
R5495 VDD.t4333 VDD.t2031 420.498
R5496 VDD.t1455 VDD.t1646 420.498
R5497 VDD.t795 VDD.t16 420.498
R5498 VDD.t956 VDD.t1107 420.498
R5499 VDD.t166 VDD.t2490 420.498
R5500 VDD.t862 VDD.t3338 420.498
R5501 VDD.t3332 VDD.t98 420.498
R5502 VDD.t1246 VDD.t1944 420.498
R5503 VDD.n2189 VDD.t4516 394.37
R5504 VDD.n2081 VDD.t4515 394.37
R5505 VDD.t1781 VDD.t1391 385.906
R5506 VDD.n1264 VDD.t2077 381.257
R5507 VDD.n1276 VDD.t4273 381.257
R5508 VDD.n1022 VDD.t2982 381.255
R5509 VDD.n893 VDD.t3001 381.255
R5510 VDD.n764 VDD.t3026 381.255
R5511 VDD.n613 VDD.t2937 381.255
R5512 VDD.n484 VDD.t2951 381.255
R5513 VDD.n355 VDD.t2988 381.255
R5514 VDD.n226 VDD.t2949 381.255
R5515 VDD.n88 VDD.t2933 381.255
R5516 VDD.n26 VDD.t2943 381.255
R5517 VDD.n2371 VDD.t162 381.101
R5518 VDD.n1240 VDD.t1086 381.055
R5519 VDD.n1312 VDD.t3930 381.055
R5520 VDD.n1324 VDD.t2683 381.055
R5521 VDD.n1288 VDD.t725 381.055
R5522 VDD.n1300 VDD.t2632 381.055
R5523 VDD.n1252 VDD.t811 381.055
R5524 VDD.n1216 VDD.t3147 381.055
R5525 VDD.n1228 VDD.t2620 381.055
R5526 VDD.t439 VDD.n1185 381.055
R5527 VDD.n1203 VDD.t1125 381.005
R5528 VDD.n148 VDD.n147 379.366
R5529 VDD.n2400 VDD.n2399 379.301
R5530 VDD.n2407 VDD.n2406 379.301
R5531 VDD.n2382 VDD.n2381 379.301
R5532 VDD.n2230 VDD.n2229 379.3
R5533 VDD.n2228 VDD.n2204 379.3
R5534 VDD.n2228 VDD.n2224 379.3
R5535 VDD.n2228 VDD.n2207 379.3
R5536 VDD.n2228 VDD.n2210 379.3
R5537 VDD.n2228 VDD.n2227 379.3
R5538 VDD.n2193 VDD.n2192 379.3
R5539 VDD.n2192 VDD.n2185 379.3
R5540 VDD.n2192 VDD.n2180 379.3
R5541 VDD.n2192 VDD.n2150 379.3
R5542 VDD.n2192 VDD.n2149 379.3
R5543 VDD.n2192 VDD.n2148 379.3
R5544 VDD.n2192 VDD.n2147 379.3
R5545 VDD.n2192 VDD.n2146 379.3
R5546 VDD.n2192 VDD.n2145 379.3
R5547 VDD.n2192 VDD.n2142 379.3
R5548 VDD.n2192 VDD.n2139 379.3
R5549 VDD.n2192 VDD.n2136 379.3
R5550 VDD.n2192 VDD.n2133 379.3
R5551 VDD.n2192 VDD.n2130 379.3
R5552 VDD.n2192 VDD.n2127 379.3
R5553 VDD.n2192 VDD.n2124 379.3
R5554 VDD.n2192 VDD.n2191 379.3
R5555 VDD.n2115 VDD.n2114 379.3
R5556 VDD.n2114 VDD.n2053 379.3
R5557 VDD.n2114 VDD.n2057 379.3
R5558 VDD.n2114 VDD.n2061 379.3
R5559 VDD.n2114 VDD.n2065 379.3
R5560 VDD.n2114 VDD.n2069 379.3
R5561 VDD.n2114 VDD.n2073 379.3
R5562 VDD.n2114 VDD.n2077 379.3
R5563 VDD.n2114 VDD.n2074 379.3
R5564 VDD.n2114 VDD.n2070 379.3
R5565 VDD.n2114 VDD.n2066 379.3
R5566 VDD.n2114 VDD.n2062 379.3
R5567 VDD.n2114 VDD.n2058 379.3
R5568 VDD.n2114 VDD.n2054 379.3
R5569 VDD.n2114 VDD.n2046 379.3
R5570 VDD.n2114 VDD.n2045 379.3
R5571 VDD.n2114 VDD.n2113 379.3
R5572 VDD.n2263 VDD.n2247 379.3
R5573 VDD.n2255 VDD.n2244 379.3
R5574 VDD.n2263 VDD.n2250 379.3
R5575 VDD.n2263 VDD.n2259 379.3
R5576 VDD.n2264 VDD.n2263 379.3
R5577 VDD.n2263 VDD.n2262 379.3
R5578 VDD.n1876 VDD.n1875 379.3
R5579 VDD.n1876 VDD.n1867 379.3
R5580 VDD.n1876 VDD.n1870 379.3
R5581 VDD.n1877 VDD.n1876 379.3
R5582 VDD.n1018 VDD.n1017 379.3
R5583 VDD.n1021 VDD.n1020 379.3
R5584 VDD.n889 VDD.n888 379.3
R5585 VDD.n892 VDD.n891 379.3
R5586 VDD.n760 VDD.n759 379.3
R5587 VDD.n763 VDD.n762 379.3
R5588 VDD.n609 VDD.n608 379.3
R5589 VDD.n612 VDD.n611 379.3
R5590 VDD.n480 VDD.n479 379.3
R5591 VDD.n483 VDD.n482 379.3
R5592 VDD.n351 VDD.n350 379.3
R5593 VDD.n354 VDD.n353 379.3
R5594 VDD.n222 VDD.n221 379.3
R5595 VDD.n225 VDD.n224 379.3
R5596 VDD.n147 VDD.n144 379.3
R5597 VDD.n84 VDD.n83 379.3
R5598 VDD.n87 VDD.n86 379.3
R5599 VDD.n22 VDD.n21 379.3
R5600 VDD.n25 VDD.n24 379.3
R5601 VDD.t1289 VDD.t2054 332.656
R5602 VDD.t2306 VDD.t4179 332.656
R5603 VDD.t453 VDD.t255 332.656
R5604 VDD.t494 VDD.t638 332.656
R5605 VDD.t3387 VDD.t3518 332.656
R5606 VDD.t2014 VDD.t4014 332.656
R5607 VDD.t1287 VDD.t2439 332.656
R5608 VDD.t3665 VDD.t3318 332.656
R5609 VDD.t3188 VDD.t603 332.656
R5610 VDD.t109 VDD.t3893 332.656
R5611 VDD.t28 VDD.t666 332.656
R5612 VDD.t1052 VDD.t4310 332.656
R5613 VDD.t2262 VDD.t2227 332.656
R5614 VDD.t758 VDD.t4221 332.656
R5615 VDD.t261 VDD.t2464 332.656
R5616 VDD.t1556 VDD.t4099 332.656
R5617 VDD.t1638 VDD.t349 332.656
R5618 VDD.t3902 VDD.t391 332.656
R5619 VDD.t2823 VDD.t2403 332.656
R5620 VDD.t3440 VDD.t3467 332.656
R5621 VDD.n1135 VDD.t2275 326.818
R5622 VDD.n2188 VDD.t3103 291.829
R5623 VDD.n2188 VDD.t3111 291.829
R5624 VDD.n2080 VDD.t3105 291.829
R5625 VDD.n2080 VDD.t3107 291.829
R5626 VDD.n1130 VDD.t3497 258.021
R5627 VDD.n2398 VDD.t1159 258.021
R5628 VDD.n2384 VDD.t1329 258.021
R5629 VDD.n2380 VDD.t1057 258.021
R5630 VDD.n2370 VDD.t163 258.021
R5631 VDD.n2201 VDD.t2340 258.021
R5632 VDD.n2203 VDD.t2581 258.021
R5633 VDD.n2212 VDD.t2118 258.021
R5634 VDD.n2206 VDD.t3610 258.021
R5635 VDD.n2209 VDD.t3970 258.021
R5636 VDD.n2216 VDD.t1166 258.021
R5637 VDD.n2214 VDD.t3559 258.021
R5638 VDD.n2226 VDD.t1012 258.021
R5639 VDD.n2043 VDD.t1703 258.021
R5640 VDD.n2041 VDD.t1028 258.021
R5641 VDD.n2048 VDD.t364 258.021
R5642 VDD.n2052 VDD.t2331 258.021
R5643 VDD.n2083 VDD.t1999 258.021
R5644 VDD.n2056 VDD.t475 258.021
R5645 VDD.n2088 VDD.t2495 258.021
R5646 VDD.n2060 VDD.t2164 258.021
R5647 VDD.n2093 VDD.t952 258.021
R5648 VDD.n2064 VDD.t3588 258.021
R5649 VDD.n2098 VDD.t681 258.021
R5650 VDD.n2068 VDD.t902 258.021
R5651 VDD.n2103 VDD.t3492 258.021
R5652 VDD.n2072 VDD.t3531 258.021
R5653 VDD.n2108 VDD.t1188 258.021
R5654 VDD.n2076 VDD.t1389 258.021
R5655 VDD.n2079 VDD.t3108 258.021
R5656 VDD.n2246 VDD.t312 258.021
R5657 VDD.n2254 VDD.t2479 258.021
R5658 VDD.n2249 VDD.t1545 258.021
R5659 VDD.n2252 VDD.t730 258.021
R5660 VDD.n2236 VDD.t2277 258.021
R5661 VDD.n2238 VDD.t786 258.021
R5662 VDD.n2241 VDD.t322 258.021
R5663 VDD.n2261 VDD.t369 258.021
R5664 VDD.n1872 VDD.t3481 258.021
R5665 VDD.n1866 VDD.t2385 258.021
R5666 VDD.n1869 VDD.t675 258.021
R5667 VDD.n1864 VDD.t2636 258.021
R5668 VDD.n1856 VDD.t1355 258.021
R5669 VDD.n1858 VDD.t825 258.021
R5670 VDD.n1880 VDD.t1574 258.021
R5671 VDD.n1861 VDD.t3485 258.021
R5672 VDD.n1311 VDD.t3931 258.021
R5673 VDD.n1323 VDD.t2684 258.021
R5674 VDD.n1287 VDD.t726 258.021
R5675 VDD.n1299 VDD.t2634 258.021
R5676 VDD.n1263 VDD.t2080 258.021
R5677 VDD.n1275 VDD.t4275 258.021
R5678 VDD.n1239 VDD.t1087 258.021
R5679 VDD.n1251 VDD.t812 258.021
R5680 VDD.n1215 VDD.t3150 258.021
R5681 VDD.n1227 VDD.t2622 258.021
R5682 VDD.n1202 VDD.t1126 258.021
R5683 VDD.n1184 VDD.t440 258.021
R5684 VDD.n1016 VDD.t3734 258.021
R5685 VDD.n1014 VDD.t4478 258.021
R5686 VDD.n1011 VDD.t2983 258.021
R5687 VDD.n1058 VDD.t1522 258.021
R5688 VDD.n887 VDD.t3790 258.021
R5689 VDD.n885 VDD.t4374 258.021
R5690 VDD.n882 VDD.t3064 258.021
R5691 VDD.n929 VDD.t3915 258.021
R5692 VDD.n758 VDD.t3792 258.021
R5693 VDD.n756 VDD.t4449 258.021
R5694 VDD.n753 VDD.t3094 258.021
R5695 VDD.n800 VDD.t3459 258.021
R5696 VDD.n607 VDD.t3831 258.021
R5697 VDD.n605 VDD.t4481 258.021
R5698 VDD.n602 VDD.t3061 258.021
R5699 VDD.n649 VDD.t3344 258.021
R5700 VDD.n478 VDD.t3709 258.021
R5701 VDD.n476 VDD.t4346 258.021
R5702 VDD.n473 VDD.t3007 258.021
R5703 VDD.n520 VDD.t2542 258.021
R5704 VDD.n349 VDD.t3836 258.021
R5705 VDD.n347 VDD.t4482 258.021
R5706 VDD.n344 VDD.t3059 258.021
R5707 VDD.n391 VDD.t2709 258.021
R5708 VDD.n220 VDD.t3715 258.021
R5709 VDD.n218 VDD.t4348 258.021
R5710 VDD.n215 VDD.t3006 258.021
R5711 VDD.n262 VDD.t1688 258.021
R5712 VDD.n673 VDD.t1476 258.021
R5713 VDD.n82 VDD.t3730 258.021
R5714 VDD.n80 VDD.t4410 258.021
R5715 VDD.n77 VDD.t2934 258.021
R5716 VDD.n124 VDD.t1104 258.021
R5717 VDD.n20 VDD.t3761 258.021
R5718 VDD.n18 VDD.t4457 258.021
R5719 VDD.n15 VDD.t3054 258.021
R5720 VDD.n2908 VDD.t3297 258.021
R5721 VDD.n2460 VDD.t4207 257.805
R5722 VDD.n2681 VDD.t3433 257.805
R5723 VDD.n2699 VDD.t2837 257.805
R5724 VDD.n1368 VDD.t1294 257.805
R5725 VDD.n1772 VDD.t2315 257.805
R5726 VDD.n1722 VDD.t244 257.805
R5727 VDD.n1337 VDD.t2444 257.805
R5728 VDD.n1686 VDD.t3525 257.805
R5729 VDD.n1343 VDD.t4009 257.805
R5730 VDD.n1328 VDD.t3323 257.805
R5731 VDD.n1500 VDD.t21 257.805
R5732 VDD.n1548 VDD.t3193 257.805
R5733 VDD.n1524 VDD.t104 257.805
R5734 VDD.n1476 VDD.t4244 257.805
R5735 VDD.n1732 VDD.t1610 257.805
R5736 VDD.n2420 VDD.t404 257.805
R5737 VDD.n2432 VDD.t1626 257.805
R5738 VDD.n2440 VDD.t4106 257.805
R5739 VDD.n2452 VDD.t266 257.805
R5740 VDD.n2468 VDD.t2224 257.805
R5741 VDD.n2676 VDD.t1841 257.798
R5742 VDD.n2415 VDD.t2473 257.798
R5743 VDD.n1726 VDD.t723 257.798
R5744 VDD.n1715 VDD.t713 257.798
R5745 VDD.n1765 VDD.t118 257.798
R5746 VDD.n1333 VDD.t2075 257.798
R5747 VDD.n1819 VDD.t1696 257.798
R5748 VDD.n1415 VDD.t4005 257.798
R5749 VDD.n1493 VDD.t574 257.798
R5750 VDD.n1517 VDD.t4041 257.798
R5751 VDD.n1541 VDD.t3682 257.798
R5752 VDD.n2619 VDD.t2701 257.798
R5753 VDD.n2435 VDD.t909 257.798
R5754 VDD.n2555 VDD.t2190 257.798
R5755 VDD.n2455 VDD.t448 257.798
R5756 VDD.n2463 VDD.t1328 257.798
R5757 VDD.n1128 VDD.t2276 257.767
R5758 VDD.n2466 VDD.t749 257.757
R5759 VDD.n2679 VDD.t3476 257.757
R5760 VDD.n2418 VDD.t2406 257.757
R5761 VDD.n2394 VDD.t1018 257.757
R5762 VDD.n2391 VDD.t4088 257.757
R5763 VDD.n2389 VDD.t1027 257.757
R5764 VDD.n2387 VDD.t554 257.757
R5765 VDD.n1168 VDD.t990 257.757
R5766 VDD.n1166 VDD.t4211 257.757
R5767 VDD.n2376 VDD.t1022 257.757
R5768 VDD.n1170 VDD.t2235 257.757
R5769 VDD.n1897 VDD.t2226 257.757
R5770 VDD.n1893 VDD.t4240 257.757
R5771 VDD.n1895 VDD.t2321 257.757
R5772 VDD.n1940 VDD.t258 257.757
R5773 VDD.n1942 VDD.t2593 257.757
R5774 VDD.n1901 VDD.t4117 257.757
R5775 VDD.n1935 VDD.t2127 257.757
R5776 VDD.n1904 VDD.t1634 257.757
R5777 VDD.n1930 VDD.t3593 257.757
R5778 VDD.n1921 VDD.t398 257.757
R5779 VDD.n1923 VDD.t890 257.757
R5780 VDD.n1906 VDD.t2831 257.757
R5781 VDD.n1916 VDD.t3569 257.757
R5782 VDD.n1908 VDD.t2301 257.757
R5783 VDD.n1912 VDD.t1403 257.757
R5784 VDD.n1889 VDD.t1025 257.757
R5785 VDD.n1307 VDD.t2173 257.757
R5786 VDD.n1304 VDD.t4187 257.757
R5787 VDD.n1319 VDD.t2125 257.757
R5788 VDD.n1316 VDD.t4112 257.757
R5789 VDD.n1283 VDD.t1675 257.757
R5790 VDD.n1280 VDD.t2137 257.757
R5791 VDD.n1295 VDD.t534 257.757
R5792 VDD.n1292 VDD.t2175 257.757
R5793 VDD.n1259 VDD.t2608 257.757
R5794 VDD.n1256 VDD.t4224 257.757
R5795 VDD.n1271 VDD.t477 257.757
R5796 VDD.n1268 VDD.t4082 257.757
R5797 VDD.n1235 VDD.t1670 257.757
R5798 VDD.n1232 VDD.t2599 257.757
R5799 VDD.n1247 VDD.t548 257.757
R5800 VDD.n1244 VDD.t2586 257.757
R5801 VDD.n1211 VDD.t2352 257.757
R5802 VDD.n1208 VDD.t4218 257.757
R5803 VDD.n1223 VDD.t2373 257.757
R5804 VDD.n1220 VDD.t4069 257.757
R5805 VDD.n1198 VDD.t1664 257.757
R5806 VDD.n1195 VDD.t2336 257.757
R5807 VDD.n1189 VDD.t524 257.757
R5808 VDD.n1187 VDD.t2369 257.757
R5809 VDD.n1730 VDD.t497 257.757
R5810 VDD.n1393 VDD.t2057 257.757
R5811 VDD.n1366 VDD.t4182 257.757
R5812 VDD.n1761 VDD.t450 257.757
R5813 VDD.n1847 VDD.t3660 257.757
R5814 VDD.n1341 VDD.t1284 257.757
R5815 VDD.n1682 VDD.t3396 257.757
R5816 VDD.n1696 VDD.t2021 257.757
R5817 VDD.n1489 VDD.t2251 257.757
R5818 VDD.n1513 VDD.t669 257.757
R5819 VDD.n1470 VDD.t1593 257.757
R5820 VDD.n1537 VDD.t3896 257.757
R5821 VDD.n2615 VDD.t3909 257.757
R5822 VDD.n2438 VDD.t300 257.757
R5823 VDD.n2551 VDD.t1563 257.757
R5824 VDD.n2458 VDD.t2467 257.757
R5825 VDD.n2473 VDD.t2257 257.757
R5826 VDD.n680 VDD.t2424 257.757
R5827 VDD.n2695 VDD.t2693 257.755
R5828 VDD.n2672 VDD.t1585 257.755
R5829 VDD.n1747 VDD.t4330 257.755
R5830 VDD.n1718 VDD.t2520 257.755
R5831 VDD.n1768 VDD.t1083 257.755
R5832 VDD.n1335 VDD.t966 257.755
R5833 VDD.n1822 VDD.t1465 257.755
R5834 VDD.n1417 VDD.t3410 257.755
R5835 VDD.n1421 VDD.t869 257.755
R5836 VDD.n1496 VDD.t143 257.755
R5837 VDD.n1520 VDD.t4049 257.755
R5838 VDD.n1544 VDD.t4270 257.755
R5839 VDD.n1472 VDD.t2216 257.755
R5840 VDD.n1395 VDD.t2247 257.755
R5841 VDD.n2622 VDD.t1848 257.755
R5842 VDD.n2608 VDD.t3995 257.755
R5843 VDD.n2558 VDD.t1859 257.755
R5844 VDD.n2544 VDD.t3325 257.755
R5845 VDD.n2528 VDD.t1359 257.755
R5846 VDD.n2475 VDD.t3402 257.755
R5847 VDD.n2540 VDD.t4139 257.755
R5848 VDD.n2684 VDD.t3648 257.755
R5849 VDD.n2702 VDD.t3241 257.755
R5850 VDD.n1711 VDD.t284 257.755
R5851 VDD.n1775 VDD.t1337 257.755
R5852 VDD.n1724 VDD.t2910 257.755
R5853 VDD.n1835 VDD.t153 257.755
R5854 VDD.n1689 VDD.t1077 257.755
R5855 VDD.n1815 VDD.t1893 257.755
R5856 VDD.n1330 VDD.t4053 257.755
R5857 VDD.n1503 VDD.t4031 257.755
R5858 VDD.n1551 VDD.t2504 257.755
R5859 VDD.n1527 VDD.t3280 257.755
R5860 VDD.n1479 VDD.t2717 257.755
R5861 VDD.n1735 VDD.t1973 257.755
R5862 VDD.n2668 VDD.t2881 257.755
R5863 VDD.n2626 VDD.t1436 257.755
R5864 VDD.n2604 VDD.t612 257.755
R5865 VDD.n2562 VDD.t338 257.755
R5866 VDD.n2524 VDD.t2085 257.755
R5867 VDD.n1419 VDD.t2105 257.755
R5868 VDD.n1467 VDD.t2742 257.755
R5869 VDD.n1390 VDD.t222 257.755
R5870 VDD.n2470 VDD.t1825 257.755
R5871 VDD.n2535 VDD.t806 257.705
R5872 VDD.n2691 VDD.t171 257.705
R5873 VDD.n2709 VDD.t1120 257.705
R5874 VDD.n1742 VDD.t2562 257.705
R5875 VDD.n1402 VDD.t1911 257.705
R5876 VDD.n1782 VDD.t218 257.705
R5877 VDD.n1757 VDD.t701 257.705
R5878 VDD.n1843 VDD.t945 257.705
R5879 VDD.n1829 VDD.t837 257.705
R5880 VDD.n1678 VDD.t1929 257.705
R5881 VDD.n1692 VDD.t2785 257.705
R5882 VDD.n1485 VDD.t4149 257.705
R5883 VDD.n1509 VDD.t3670 257.705
R5884 VDD.n1558 VDD.t1967 257.705
R5885 VDD.n1533 VDD.t4292 257.705
R5886 VDD.n2611 VDD.t2757 257.705
R5887 VDD.n2633 VDD.t3941 257.705
R5888 VDD.n2547 VDD.t1734 257.705
R5889 VDD.n2569 VDD.t95 257.705
R5890 VDD.n2482 VDD.t1776 257.705
R5891 VDD.n1126 VDD.t4125 257.683
R5892 VDD.n2123 VDD.t1001 257.644
R5893 VDD.n2121 VDD.t1239 257.644
R5894 VDD.n2126 VDD.t2326 257.644
R5895 VDD.n2182 VDD.t3262 257.644
R5896 VDD.n2129 VDD.t465 257.644
R5897 VDD.n2152 VDD.t1185 257.644
R5898 VDD.n2132 VDD.t2149 257.644
R5899 VDD.n2173 VDD.t2551 257.644
R5900 VDD.n2135 VDD.t3612 257.644
R5901 VDD.n2168 VDD.t2062 257.644
R5902 VDD.n2138 VDD.t899 257.644
R5903 VDD.n2163 VDD.t815 257.644
R5904 VDD.n2141 VDD.t3570 257.644
R5905 VDD.n2158 VDD.t1310 257.644
R5906 VDD.n2144 VDD.t1418 257.644
R5907 VDD.n2154 VDD.t138 257.644
R5908 VDD.n2187 VDD.t3104 257.644
R5909 VDD.n146 VDD.t1137 257.644
R5910 VDD.n143 VDD.t1095 257.644
R5911 VDD.n676 VDD.t2388 257.644
R5912 VDD.n674 VDD.t2387 248.495
R5913 VDD.n1130 VDD.n1129 227.905
R5914 VDD.n2398 VDD.n2397 227.905
R5915 VDD.n2384 VDD.n2383 227.905
R5916 VDD.n2380 VDD.n2379 227.905
R5917 VDD.n2370 VDD.n2369 227.905
R5918 VDD.n2201 VDD.n2200 227.905
R5919 VDD.n2203 VDD.n2202 227.905
R5920 VDD.n2212 VDD.n2211 227.905
R5921 VDD.n2206 VDD.n2205 227.905
R5922 VDD.n2209 VDD.n2208 227.905
R5923 VDD.n2216 VDD.n2215 227.905
R5924 VDD.n2214 VDD.n2213 227.905
R5925 VDD.n2226 VDD.n2225 227.905
R5926 VDD.n2043 VDD.n2042 227.905
R5927 VDD.n2041 VDD.n2040 227.905
R5928 VDD.n2048 VDD.n2047 227.905
R5929 VDD.n2052 VDD.n2051 227.905
R5930 VDD.n2083 VDD.n2082 227.905
R5931 VDD.n2056 VDD.n2055 227.905
R5932 VDD.n2088 VDD.n2087 227.905
R5933 VDD.n2060 VDD.n2059 227.905
R5934 VDD.n2093 VDD.n2092 227.905
R5935 VDD.n2064 VDD.n2063 227.905
R5936 VDD.n2098 VDD.n2097 227.905
R5937 VDD.n2068 VDD.n2067 227.905
R5938 VDD.n2103 VDD.n2102 227.905
R5939 VDD.n2072 VDD.n2071 227.905
R5940 VDD.n2108 VDD.n2107 227.905
R5941 VDD.n2076 VDD.n2075 227.905
R5942 VDD.n2079 VDD.n2078 227.905
R5943 VDD.n2246 VDD.n2245 227.905
R5944 VDD.n2254 VDD.n2253 227.905
R5945 VDD.n2249 VDD.n2248 227.905
R5946 VDD.n2252 VDD.n2251 227.905
R5947 VDD.n2236 VDD.n2235 227.905
R5948 VDD.n2238 VDD.n2237 227.905
R5949 VDD.n2241 VDD.n2240 227.905
R5950 VDD.n2261 VDD.n2260 227.905
R5951 VDD.n1872 VDD.n1871 227.905
R5952 VDD.n1866 VDD.n1865 227.905
R5953 VDD.n1869 VDD.n1868 227.905
R5954 VDD.n1864 VDD.n1863 227.905
R5955 VDD.n1856 VDD.n1855 227.905
R5956 VDD.n1858 VDD.n1857 227.905
R5957 VDD.n1880 VDD.n1879 227.905
R5958 VDD.n1861 VDD.n1860 227.905
R5959 VDD.n1311 VDD.n1310 227.905
R5960 VDD.n1323 VDD.n1322 227.905
R5961 VDD.n1287 VDD.n1286 227.905
R5962 VDD.n1299 VDD.n1298 227.905
R5963 VDD.n1263 VDD.n1262 227.905
R5964 VDD.n1275 VDD.n1274 227.905
R5965 VDD.n1239 VDD.n1238 227.905
R5966 VDD.n1251 VDD.n1250 227.905
R5967 VDD.n1215 VDD.n1214 227.905
R5968 VDD.n1227 VDD.n1226 227.905
R5969 VDD.n1202 VDD.n1201 227.905
R5970 VDD.n1184 VDD.n1183 227.905
R5971 VDD.n1016 VDD.n1015 227.905
R5972 VDD.n1014 VDD.n1013 227.905
R5973 VDD.n1011 VDD.n1010 227.905
R5974 VDD.n1058 VDD.n1057 227.905
R5975 VDD.n887 VDD.n886 227.905
R5976 VDD.n885 VDD.n884 227.905
R5977 VDD.n882 VDD.n881 227.905
R5978 VDD.n929 VDD.n928 227.905
R5979 VDD.n758 VDD.n757 227.905
R5980 VDD.n756 VDD.n755 227.905
R5981 VDD.n753 VDD.n752 227.905
R5982 VDD.n800 VDD.n799 227.905
R5983 VDD.n607 VDD.n606 227.905
R5984 VDD.n605 VDD.n604 227.905
R5985 VDD.n602 VDD.n601 227.905
R5986 VDD.n649 VDD.n648 227.905
R5987 VDD.n478 VDD.n477 227.905
R5988 VDD.n476 VDD.n475 227.905
R5989 VDD.n473 VDD.n472 227.905
R5990 VDD.n520 VDD.n519 227.905
R5991 VDD.n349 VDD.n348 227.905
R5992 VDD.n347 VDD.n346 227.905
R5993 VDD.n344 VDD.n343 227.905
R5994 VDD.n391 VDD.n390 227.905
R5995 VDD.n220 VDD.n219 227.905
R5996 VDD.n218 VDD.n217 227.905
R5997 VDD.n215 VDD.n214 227.905
R5998 VDD.n262 VDD.n261 227.905
R5999 VDD.n673 VDD.n672 227.905
R6000 VDD.n82 VDD.n81 227.905
R6001 VDD.n80 VDD.n79 227.905
R6002 VDD.n77 VDD.n76 227.905
R6003 VDD.n124 VDD.n123 227.905
R6004 VDD.n20 VDD.n19 227.905
R6005 VDD.n18 VDD.n17 227.905
R6006 VDD.n15 VDD.n14 227.905
R6007 VDD.n2908 VDD.n2907 227.905
R6008 VDD.n2123 VDD.n2122 227.529
R6009 VDD.n2121 VDD.n2120 227.529
R6010 VDD.n2126 VDD.n2125 227.529
R6011 VDD.n2182 VDD.n2181 227.529
R6012 VDD.n2129 VDD.n2128 227.529
R6013 VDD.n2152 VDD.n2151 227.529
R6014 VDD.n2132 VDD.n2131 227.529
R6015 VDD.n2173 VDD.n2172 227.529
R6016 VDD.n2135 VDD.n2134 227.529
R6017 VDD.n2168 VDD.n2167 227.529
R6018 VDD.n2138 VDD.n2137 227.529
R6019 VDD.n2163 VDD.n2162 227.529
R6020 VDD.n2141 VDD.n2140 227.529
R6021 VDD.n2158 VDD.n2157 227.529
R6022 VDD.n2144 VDD.n2143 227.529
R6023 VDD.n2154 VDD.n2153 227.529
R6024 VDD.n2187 VDD.n2186 227.529
R6025 VDD.n146 VDD.n145 227.529
R6026 VDD.n143 VDD.n142 227.529
R6027 VDD.n1132 VDD.n1131 227.266
R6028 VDD.n1128 VDD.n1127 227.266
R6029 VDD.n2528 VDD.n2527 227.266
R6030 VDD.n2463 VDD.n2462 227.266
R6031 VDD.n2534 VDD.n2533 227.266
R6032 VDD.n2466 VDD.n2465 227.266
R6033 VDD.n2540 VDD.n2539 227.266
R6034 VDD.n2460 VDD.n2459 227.266
R6035 VDD.n2690 VDD.n2689 227.266
R6036 VDD.n2679 VDD.n2678 227.266
R6037 VDD.n2695 VDD.n2694 227.266
R6038 VDD.n2676 VDD.n2675 227.266
R6039 VDD.n2684 VDD.n2683 227.266
R6040 VDD.n2681 VDD.n2680 227.266
R6041 VDD.n2708 VDD.n2707 227.266
R6042 VDD.n2418 VDD.n2417 227.266
R6043 VDD.n2672 VDD.n2671 227.266
R6044 VDD.n2415 VDD.n2414 227.266
R6045 VDD.n2702 VDD.n2701 227.266
R6046 VDD.n2699 VDD.n2698 227.266
R6047 VDD.n2394 VDD.n2393 227.266
R6048 VDD.n2391 VDD.n2390 227.266
R6049 VDD.n2389 VDD.n2388 227.266
R6050 VDD.n2387 VDD.n2386 227.266
R6051 VDD.n1168 VDD.n1167 227.266
R6052 VDD.n1166 VDD.n1165 227.266
R6053 VDD.n2376 VDD.n2375 227.266
R6054 VDD.n1170 VDD.n1169 227.266
R6055 VDD.n1893 VDD.n1892 227.266
R6056 VDD.n1895 VDD.n1894 227.266
R6057 VDD.n1940 VDD.n1939 227.266
R6058 VDD.n1942 VDD.n1941 227.266
R6059 VDD.n1901 VDD.n1900 227.266
R6060 VDD.n1935 VDD.n1934 227.266
R6061 VDD.n1904 VDD.n1903 227.266
R6062 VDD.n1930 VDD.n1929 227.266
R6063 VDD.n1921 VDD.n1920 227.266
R6064 VDD.n1923 VDD.n1922 227.266
R6065 VDD.n1906 VDD.n1905 227.266
R6066 VDD.n1916 VDD.n1915 227.266
R6067 VDD.n1908 VDD.n1907 227.266
R6068 VDD.n1912 VDD.n1911 227.266
R6069 VDD.n1897 VDD.n1896 227.266
R6070 VDD.n1889 VDD.n1888 227.266
R6071 VDD.n1307 VDD.n1306 227.266
R6072 VDD.n1304 VDD.n1303 227.266
R6073 VDD.n1319 VDD.n1318 227.266
R6074 VDD.n1316 VDD.n1315 227.266
R6075 VDD.n1283 VDD.n1282 227.266
R6076 VDD.n1280 VDD.n1279 227.266
R6077 VDD.n1295 VDD.n1294 227.266
R6078 VDD.n1292 VDD.n1291 227.266
R6079 VDD.n1259 VDD.n1258 227.266
R6080 VDD.n1256 VDD.n1255 227.266
R6081 VDD.n1271 VDD.n1270 227.266
R6082 VDD.n1268 VDD.n1267 227.266
R6083 VDD.n1235 VDD.n1234 227.266
R6084 VDD.n1232 VDD.n1231 227.266
R6085 VDD.n1247 VDD.n1246 227.266
R6086 VDD.n1244 VDD.n1243 227.266
R6087 VDD.n1211 VDD.n1210 227.266
R6088 VDD.n1208 VDD.n1207 227.266
R6089 VDD.n1223 VDD.n1222 227.266
R6090 VDD.n1220 VDD.n1219 227.266
R6091 VDD.n1198 VDD.n1197 227.266
R6092 VDD.n1195 VDD.n1194 227.266
R6093 VDD.n1189 VDD.n1188 227.266
R6094 VDD.n1187 VDD.n1186 227.266
R6095 VDD.n1730 VDD.n1729 227.266
R6096 VDD.n1741 VDD.n1740 227.266
R6097 VDD.n1747 VDD.n1746 227.266
R6098 VDD.n1726 VDD.n1725 227.266
R6099 VDD.n1395 VDD.n1394 227.266
R6100 VDD.n1390 VDD.n1389 227.266
R6101 VDD.n1401 VDD.n1400 227.266
R6102 VDD.n1393 VDD.n1392 227.266
R6103 VDD.n1711 VDD.n1710 227.266
R6104 VDD.n1368 VDD.n1367 227.266
R6105 VDD.n1781 VDD.n1780 227.266
R6106 VDD.n1366 VDD.n1365 227.266
R6107 VDD.n1718 VDD.n1717 227.266
R6108 VDD.n1715 VDD.n1714 227.266
R6109 VDD.n1775 VDD.n1774 227.266
R6110 VDD.n1772 VDD.n1771 227.266
R6111 VDD.n1759 VDD.n1758 227.266
R6112 VDD.n1761 VDD.n1760 227.266
R6113 VDD.n1768 VDD.n1767 227.266
R6114 VDD.n1765 VDD.n1764 227.266
R6115 VDD.n1724 VDD.n1723 227.266
R6116 VDD.n1722 VDD.n1721 227.266
R6117 VDD.n1847 VDD.n1846 227.266
R6118 VDD.n1845 VDD.n1844 227.266
R6119 VDD.n1335 VDD.n1334 227.266
R6120 VDD.n1333 VDD.n1332 227.266
R6121 VDD.n1822 VDD.n1821 227.266
R6122 VDD.n1819 VDD.n1818 227.266
R6123 VDD.n1828 VDD.n1827 227.266
R6124 VDD.n1341 VDD.n1340 227.266
R6125 VDD.n1835 VDD.n1834 227.266
R6126 VDD.n1337 VDD.n1336 227.266
R6127 VDD.n1421 VDD.n1420 227.266
R6128 VDD.n1419 VDD.n1418 227.266
R6129 VDD.n1680 VDD.n1679 227.266
R6130 VDD.n1682 VDD.n1681 227.266
R6131 VDD.n1689 VDD.n1688 227.266
R6132 VDD.n1686 VDD.n1685 227.266
R6133 VDD.n1694 VDD.n1693 227.266
R6134 VDD.n1696 VDD.n1695 227.266
R6135 VDD.n1417 VDD.n1416 227.266
R6136 VDD.n1415 VDD.n1414 227.266
R6137 VDD.n1815 VDD.n1814 227.266
R6138 VDD.n1343 VDD.n1342 227.266
R6139 VDD.n1330 VDD.n1329 227.266
R6140 VDD.n1328 VDD.n1327 227.266
R6141 VDD.n1489 VDD.n1488 227.266
R6142 VDD.n1487 VDD.n1486 227.266
R6143 VDD.n1496 VDD.n1495 227.266
R6144 VDD.n1493 VDD.n1492 227.266
R6145 VDD.n1520 VDD.n1519 227.266
R6146 VDD.n1517 VDD.n1516 227.266
R6147 VDD.n1511 VDD.n1510 227.266
R6148 VDD.n1513 VDD.n1512 227.266
R6149 VDD.n1503 VDD.n1502 227.266
R6150 VDD.n1500 VDD.n1499 227.266
R6151 VDD.n1472 VDD.n1471 227.266
R6152 VDD.n1467 VDD.n1466 227.266
R6153 VDD.n1557 VDD.n1556 227.266
R6154 VDD.n1470 VDD.n1469 227.266
R6155 VDD.n1551 VDD.n1550 227.266
R6156 VDD.n1548 VDD.n1547 227.266
R6157 VDD.n1535 VDD.n1534 227.266
R6158 VDD.n1537 VDD.n1536 227.266
R6159 VDD.n1544 VDD.n1543 227.266
R6160 VDD.n1541 VDD.n1540 227.266
R6161 VDD.n1527 VDD.n1526 227.266
R6162 VDD.n1524 VDD.n1523 227.266
R6163 VDD.n1479 VDD.n1478 227.266
R6164 VDD.n1476 VDD.n1475 227.266
R6165 VDD.n1735 VDD.n1734 227.266
R6166 VDD.n1732 VDD.n1731 227.266
R6167 VDD.n2613 VDD.n2612 227.266
R6168 VDD.n2615 VDD.n2614 227.266
R6169 VDD.n2622 VDD.n2621 227.266
R6170 VDD.n2619 VDD.n2618 227.266
R6171 VDD.n2668 VDD.n2667 227.266
R6172 VDD.n2420 VDD.n2419 227.266
R6173 VDD.n2632 VDD.n2631 227.266
R6174 VDD.n2438 VDD.n2437 227.266
R6175 VDD.n2608 VDD.n2607 227.266
R6176 VDD.n2435 VDD.n2434 227.266
R6177 VDD.n2626 VDD.n2625 227.266
R6178 VDD.n2432 VDD.n2431 227.266
R6179 VDD.n2549 VDD.n2548 227.266
R6180 VDD.n2551 VDD.n2550 227.266
R6181 VDD.n2558 VDD.n2557 227.266
R6182 VDD.n2555 VDD.n2554 227.266
R6183 VDD.n2604 VDD.n2603 227.266
R6184 VDD.n2440 VDD.n2439 227.266
R6185 VDD.n2568 VDD.n2567 227.266
R6186 VDD.n2458 VDD.n2457 227.266
R6187 VDD.n2544 VDD.n2543 227.266
R6188 VDD.n2455 VDD.n2454 227.266
R6189 VDD.n2562 VDD.n2561 227.266
R6190 VDD.n2452 VDD.n2451 227.266
R6191 VDD.n2473 VDD.n2472 227.266
R6192 VDD.n2481 VDD.n2480 227.266
R6193 VDD.n2475 VDD.n2474 227.266
R6194 VDD.n2470 VDD.n2469 227.266
R6195 VDD.n2524 VDD.n2523 227.266
R6196 VDD.n2468 VDD.n2467 227.266
R6197 VDD.n680 VDD.n679 227.266
R6198 VDD.n678 VDD.n677 227.266
R6199 VDD.t3560 VDD.t3545 226.304
R6200 VDD.t317 VDD.t319 226.304
R6201 VDD.t1569 VDD.t1571 226.304
R6202 VDD.t1521 VDD.t1523 223.53
R6203 VDD.t1523 VDD.t1519 223.53
R6204 VDD.t3914 VDD.t3916 223.53
R6205 VDD.t3916 VDD.t3918 223.53
R6206 VDD.t3458 VDD.t3460 223.53
R6207 VDD.t3460 VDD.t3456 223.53
R6208 VDD.t3343 VDD.t3345 223.53
R6209 VDD.t3345 VDD.t1316 223.53
R6210 VDD.t2541 VDD.t2543 223.53
R6211 VDD.t2543 VDD.t2545 223.53
R6212 VDD.t2708 VDD.t2710 223.53
R6213 VDD.t2710 VDD.t2706 223.53
R6214 VDD.t1687 VDD.t1689 223.53
R6215 VDD.t1689 VDD.t1691 223.53
R6216 VDD.t1103 VDD.t1099 223.53
R6217 VDD.t1099 VDD.t1101 223.53
R6218 VDD.t3296 VDD.t3294 223.53
R6219 VDD.t3294 VDD.t3292 223.53
R6220 VDD.n2188 VDD.t3113 221.72
R6221 VDD.n2080 VDD.t3109 221.72
R6222 VDD.t826 VDD.t828 221.359
R6223 VDD.n1959 VDD.t1031 220.395
R6224 VDD.n2335 VDD.t2363 220.395
R6225 VDD.n2325 VDD.t2597 220.395
R6226 VDD.n2315 VDD.t2148 220.395
R6227 VDD.n2304 VDD.t3599 220.395
R6228 VDD.n2294 VDD.t896 220.395
R6229 VDD.n2284 VDD.t3567 220.395
R6230 VDD.n2274 VDD.t1417 220.395
R6231 VDD.n1070 VDD.t33 220.395
R6232 VDD.n941 VDD.t3927 220.395
R6233 VDD.n812 VDD.t1229 220.395
R6234 VDD.n661 VDD.t4304 220.395
R6235 VDD.n532 VDD.t4260 220.395
R6236 VDD.n403 VDD.t741 220.395
R6237 VDD.n274 VDD.t2908 220.395
R6238 VDD.n136 VDD.t4317 220.395
R6239 VDD.n2920 VDD.t3505 220.395
R6240 VDD.t2275 VDD.t2271 211.112
R6241 VDD.t2271 VDD.t2273 211.112
R6242 VDD.t4126 VDD.t4128 211.112
R6243 VDD.t4128 VDD.t4124 211.112
R6244 VDD.t2830 VDD.t2832 211.112
R6245 VDD.t2832 VDD.t2819 211.112
R6246 VDD.t3556 VDD.t3543 211.112
R6247 VDD.t3568 VDD.t3556 211.112
R6248 VDD.t3419 VDD.t2300 211.112
R6249 VDD.t3434 VDD.t3419 211.112
R6250 VDD.t1414 VDD.t1178 211.112
R6251 VDD.t1178 VDD.t1402 211.112
R6252 VDD.t397 VDD.t381 211.112
R6253 VDD.t381 VDD.t393 211.112
R6254 VDD.t903 VDD.t3974 211.112
R6255 VDD.t1640 VDD.t1633 211.112
R6256 VDD.t2197 VDD.t1640 211.112
R6257 VDD.t3600 VDD.t3613 211.112
R6258 VDD.t4116 VDD.t4066 211.112
R6259 VDD.t4066 VDD.t4070 211.112
R6260 VDD.t2162 VDD.t2157 211.112
R6261 VDD.t257 VDD.t519 211.112
R6262 VDD.t519 VDD.t531 211.112
R6263 VDD.t481 VDD.t485 211.112
R6264 VDD.t4188 VDD.t4239 211.112
R6265 VDD.t4208 VDD.t4188 211.112
R6266 VDD.t2364 VDD.t2370 211.112
R6267 VDD.t2238 VDD.t2225 211.112
R6268 VDD.t1661 VDD.t2238 211.112
R6269 VDD.t1019 VDD.t997 211.112
R6270 VDD.t2387 VDD.t2389 211.112
R6271 VDD.t2389 VDD.t2391 211.112
R6272 VDD.t1820 VDD.t195 211.112
R6273 VDD.t2423 VDD.t1820 211.112
R6274 VDD.n1080 VDD.t810 205.447
R6275 VDD.n1078 VDD.t1324 205.447
R6276 VDD.n999 VDD.t2032 205.447
R6277 VDD.n997 VDD.t4334 205.447
R6278 VDD.n951 VDD.t2210 205.447
R6279 VDD.n949 VDD.t1351 205.447
R6280 VDD.n870 VDD.t1647 205.447
R6281 VDD.n868 VDD.t1456 205.447
R6282 VDD.n822 VDD.t1726 205.447
R6283 VDD.n820 VDD.t3354 205.447
R6284 VDD.n741 VDD.t17 205.447
R6285 VDD.n739 VDD.t796 205.447
R6286 VDD.n693 VDD.t3574 205.447
R6287 VDD.n691 VDD.t4168 205.447
R6288 VDD.n590 VDD.t1367 205.447
R6289 VDD.n588 VDD.t3414 205.447
R6290 VDD.n542 VDD.t3957 205.447
R6291 VDD.n540 VDD.t233 205.447
R6292 VDD.n461 VDD.t1108 205.447
R6293 VDD.n459 VDD.t957 205.447
R6294 VDD.n413 VDD.t52 205.447
R6295 VDD.n411 VDD.t48 205.447
R6296 VDD.n332 VDD.t2491 205.447
R6297 VDD.n330 VDD.t167 205.447
R6298 VDD.n284 VDD.t2283 205.447
R6299 VDD.n282 VDD.t2570 205.447
R6300 VDD.n155 VDD.t416 205.447
R6301 VDD.n153 VDD.t2065 205.447
R6302 VDD.n203 VDD.t3339 205.447
R6303 VDD.n201 VDD.t863 205.447
R6304 VDD.n65 VDD.t99 205.447
R6305 VDD.n63 VDD.t3333 205.447
R6306 VDD.n2860 VDD.t1965 205.447
R6307 VDD.n2858 VDD.t1502 205.447
R6308 VDD.n3 VDD.t1945 205.447
R6309 VDD.n1 VDD.t1247 205.447
R6310 VDD.n1092 VDD.t3713 205.447
R6311 VDD.n963 VDD.t3853 205.447
R6312 VDD.n834 VDD.t3776 205.447
R6313 VDD.n705 VDD.t3701 205.447
R6314 VDD.n554 VDD.t3703 205.447
R6315 VDD.n425 VDD.t3828 205.447
R6316 VDD.n296 VDD.t3705 205.447
R6317 VDD.n167 VDD.t3833 205.447
R6318 VDD.n2872 VDD.t3781 205.447
R6319 VDD.n1023 VDD.t3181 205.421
R6320 VDD.n894 VDD.t2807 205.421
R6321 VDD.n765 VDD.t134 205.421
R6322 VDD.n614 VDD.t1379 205.421
R6323 VDD.n485 VDD.t3142 205.421
R6324 VDD.n356 VDD.t1512 205.421
R6325 VDD.n227 VDD.t430 205.421
R6326 VDD.n89 VDD.t1708 205.421
R6327 VDD.n27 VDD.t2888 205.421
R6328 VDD.t1460 VDD.t1462 205.405
R6329 VDD.n1112 VDD.t3747 205.349
R6330 VDD.n1085 VDD.t3711 205.349
R6331 VDD.n1111 VDD.t3696 205.349
R6332 VDD.n1100 VDD.t3835 205.349
R6333 VDD.n1086 VDD.t1061 205.349
R6334 VDD.n1099 VDD.t2383 205.349
R6335 VDD.n1123 VDD.t1600 205.349
R6336 VDD.n1032 VDD.t794 205.349
R6337 VDD.n1033 VDD.t3175 205.349
R6338 VDD.n1005 VDD.t951 205.349
R6339 VDD.n1004 VDD.t3179 205.349
R6340 VDD.n1044 VDD.t1533 205.349
R6341 VDD.n1045 VDD.t3171 205.349
R6342 VDD.n1056 VDD.t917 205.349
R6343 VDD.n983 VDD.t3719 205.349
R6344 VDD.n956 VDD.t3851 205.349
R6345 VDD.n982 VDD.t65 205.349
R6346 VDD.n971 VDD.t3784 205.349
R6347 VDD.n957 VDD.t626 205.349
R6348 VDD.n970 VDD.t1249 205.349
R6349 VDD.n994 VDD.t4296 205.349
R6350 VDD.n903 VDD.t436 205.349
R6351 VDD.n904 VDD.t2805 205.349
R6352 VDD.n876 VDD.t1491 205.349
R6353 VDD.n875 VDD.t2801 205.349
R6354 VDD.n915 VDD.t3 205.349
R6355 VDD.n916 VDD.t2811 205.349
R6356 VDD.n927 VDD.t2645 205.349
R6357 VDD.n854 VDD.t3717 205.349
R6358 VDD.n827 VDD.t3743 205.349
R6359 VDD.n853 VDD.t1210 205.349
R6360 VDD.n842 VDD.t3756 205.349
R6361 VDD.n828 VDD.t1139 205.349
R6362 VDD.n841 VDD.t3398 205.349
R6363 VDD.n865 VDD.t922 205.349
R6364 VDD.n774 VDD.t2793 205.349
R6365 VDD.n775 VDD.t132 205.349
R6366 VDD.n747 VDD.t410 205.349
R6367 VDD.n746 VDD.t128 205.349
R6368 VDD.n786 VDD.t240 205.349
R6369 VDD.n787 VDD.t122 205.349
R6370 VDD.n798 VDD.t2787 205.349
R6371 VDD.n725 VDD.t3849 205.349
R6372 VDD.n698 VDD.t3824 205.349
R6373 VDD.n724 VDD.t44 205.349
R6374 VDD.n713 VDD.t3867 205.349
R6375 VDD.n699 VDD.t1621 205.349
R6376 VDD.n712 VDD.t1865 205.349
R6377 VDD.n736 VDD.t4021 205.349
R6378 VDD.n636 VDD.t1383 205.349
R6379 VDD.n595 VDD.t1373 205.349
R6380 VDD.n635 VDD.t3348 205.349
R6381 VDD.n624 VDD.t1377 205.349
R6382 VDD.n596 VDD.t2042 205.349
R6383 VDD.n623 VDD.t873 205.349
R6384 VDD.n647 VDD.t1212 205.349
R6385 VDD.n574 VDD.t3857 205.349
R6386 VDD.n547 VDD.t3826 205.349
R6387 VDD.n573 VDD.t4131 205.349
R6388 VDD.n562 VDD.t3869 205.349
R6389 VDD.n548 VDD.t175 205.349
R6390 VDD.n561 VDD.t1487 205.349
R6391 VDD.n585 VDD.t1154 205.349
R6392 VDD.n494 VDD.t503 205.349
R6393 VDD.n495 VDD.t3140 205.349
R6394 VDD.n467 VDD.t149 205.349
R6395 VDD.n466 VDD.t3136 205.349
R6396 VDD.n506 VDD.t606 205.349
R6397 VDD.n507 VDD.t3130 205.349
R6398 VDD.n518 VDD.t511 205.349
R6399 VDD.n445 VDD.t3800 205.349
R6400 VDD.n418 VDD.t3773 205.349
R6401 VDD.n444 VDD.t1202 205.349
R6402 VDD.n433 VDD.t3806 205.349
R6403 VDD.n419 VDD.t2112 205.349
R6404 VDD.n432 VDD.t1568 205.349
R6405 VDD.n456 VDD.t2038 205.349
R6406 VDD.n365 VDD.t1233 205.349
R6407 VDD.n366 VDD.t1510 205.349
R6408 VDD.n338 VDD.t3144 205.349
R6409 VDD.n337 VDD.t1506 205.349
R6410 VDD.n377 VDD.t1498 205.349
R6411 VDD.n378 VDD.t1516 205.349
R6412 VDD.n389 VDD.t1471 205.349
R6413 VDD.n316 VDD.t3863 205.349
R6414 VDD.n289 VDD.t3830 205.349
R6415 VDD.n315 VDD.t3991 205.349
R6416 VDD.n304 VDD.t3875 205.349
R6417 VDD.n290 VDD.t1065 205.349
R6418 VDD.n303 VDD.t1861 205.349
R6419 VDD.n327 VDD.t2285 205.349
R6420 VDD.n187 VDD.t3749 205.349
R6421 VDD.n160 VDD.t3779 205.349
R6422 VDD.n186 VDD.t3266 205.349
R6423 VDD.n175 VDD.t3810 205.349
R6424 VDD.n161 VDD.t280 205.349
R6425 VDD.n174 VDD.t358 205.349
R6426 VDD.n198 VDD.t491 205.349
R6427 VDD.n236 VDD.t507 205.349
R6428 VDD.n237 VDD.t428 205.349
R6429 VDD.n209 VDD.t1223 205.349
R6430 VDD.n208 VDD.t424 205.349
R6431 VDD.n248 VDD.t3307 205.349
R6432 VDD.n249 VDD.t434 205.349
R6433 VDD.n260 VDD.t913 205.349
R6434 VDD.n98 VDD.t580 205.349
R6435 VDD.n99 VDD.t1718 205.349
R6436 VDD.n71 VDD.t881 205.349
R6437 VDD.n70 VDD.t1706 205.349
R6438 VDD.n110 VDD.t3358 205.349
R6439 VDD.n111 VDD.t1714 205.349
R6440 VDD.n122 VDD.t771 205.349
R6441 VDD.n2892 VDD.t3786 205.349
R6442 VDD.n2865 VDD.t3820 205.349
R6443 VDD.n2891 VDD.t1951 205.349
R6444 VDD.n2880 VDD.t3871 205.349
R6445 VDD.n2866 VDD.t2512 205.349
R6446 VDD.n2879 VDD.t1684 205.349
R6447 VDD.n2903 VDD.t1256 205.349
R6448 VDD.n36 VDD.t1915 205.349
R6449 VDD.n37 VDD.t2902 205.349
R6450 VDD.n9 VDD.t1921 205.349
R6451 VDD.n8 VDD.t2900 205.349
R6452 VDD.n48 VDD.t1581 205.349
R6453 VDD.n49 VDD.t2892 205.349
R6454 VDD.n60 VDD.t2206 205.349
R6455 VDD.t3974 VDD.t889 202.953
R6456 VDD.t1024 VDD.t1019 202.953
R6457 VDD.t2126 VDD.t2162 202.495
R6458 VDD.t2370 VDD.t2320 201.131
R6459 VDD.t485 VDD.t2592 196.715
R6460 VDD.n1955 VDD.n1954 195
R6461 VDD.n1957 VDD.n1956 195
R6462 VDD.n2331 VDD.n2330 195
R6463 VDD.n2333 VDD.n2332 195
R6464 VDD.n2321 VDD.n2320 195
R6465 VDD.n2323 VDD.n2322 195
R6466 VDD.n2311 VDD.n2310 195
R6467 VDD.n2313 VDD.n2312 195
R6468 VDD.n2300 VDD.n2299 195
R6469 VDD.n2302 VDD.n2301 195
R6470 VDD.n2290 VDD.n2289 195
R6471 VDD.n2292 VDD.n2291 195
R6472 VDD.n2280 VDD.n2279 195
R6473 VDD.n2282 VDD.n2281 195
R6474 VDD.n2270 VDD.n2269 195
R6475 VDD.n2272 VDD.n2271 195
R6476 VDD.n1068 VDD.n1067 195
R6477 VDD.n1066 VDD.n1065 195
R6478 VDD.n939 VDD.n938 195
R6479 VDD.n937 VDD.n936 195
R6480 VDD.n810 VDD.n809 195
R6481 VDD.n808 VDD.n807 195
R6482 VDD.n659 VDD.n658 195
R6483 VDD.n657 VDD.n656 195
R6484 VDD.n530 VDD.n529 195
R6485 VDD.n528 VDD.n527 195
R6486 VDD.n401 VDD.n400 195
R6487 VDD.n399 VDD.n398 195
R6488 VDD.n272 VDD.n271 195
R6489 VDD.n270 VDD.n269 195
R6490 VDD.n134 VDD.n133 195
R6491 VDD.n132 VDD.n131 195
R6492 VDD.n2918 VDD.n2917 195
R6493 VDD.n2916 VDD.n2915 195
R6494 VDD.t3613 VDD.t3592 190.044
R6495 VDD.t3500 VDD.t3498 190
R6496 VDD.t4192 VDD.t4190 187.655
R6497 VDD.t2583 VDD.t2601 187.655
R6498 VDD.t2601 VDD.t2607 187.655
R6499 VDD.t4093 VDD.t4113 187.655
R6500 VDD.t463 VDD.t473 187.655
R6501 VDD.t473 VDD.t476 187.655
R6502 VDD.t4223 VDD.t4192 187.655
R6503 VDD.t4081 VDD.t4093 187.655
R6504 VDD.n1114 VDD.n1113 185.16
R6505 VDD.n1082 VDD.n1081 185.16
R6506 VDD.n1080 VDD.n1079 185.16
R6507 VDD.n1084 VDD.n1083 185.16
R6508 VDD.n1108 VDD.n1107 185.16
R6509 VDD.n1110 VDD.n1109 185.16
R6510 VDD.n1102 VDD.n1101 185.16
R6511 VDD.n1090 VDD.n1089 185.16
R6512 VDD.n1088 VDD.n1087 185.16
R6513 VDD.n1092 VDD.n1091 185.16
R6514 VDD.n1096 VDD.n1095 185.16
R6515 VDD.n1098 VDD.n1097 185.16
R6516 VDD.n1078 VDD.n1077 185.16
R6517 VDD.n1120 VDD.n1119 185.16
R6518 VDD.n1122 VDD.n1121 185.16
R6519 VDD.n1025 VDD.n1024 185.16
R6520 VDD.n1029 VDD.n1028 185.16
R6521 VDD.n1031 VDD.n1030 185.16
R6522 VDD.n1035 VDD.n1034 185.16
R6523 VDD.n1009 VDD.n1008 185.16
R6524 VDD.n1007 VDD.n1006 185.16
R6525 VDD.n1003 VDD.n1002 185.16
R6526 VDD.n1041 VDD.n1040 185.16
R6527 VDD.n1043 VDD.n1042 185.16
R6528 VDD.n1047 VDD.n1046 185.16
R6529 VDD.n1001 VDD.n1000 185.16
R6530 VDD.n999 VDD.n998 185.16
R6531 VDD.n997 VDD.n996 185.16
R6532 VDD.n1053 VDD.n1052 185.16
R6533 VDD.n1055 VDD.n1054 185.16
R6534 VDD.n985 VDD.n984 185.16
R6535 VDD.n953 VDD.n952 185.16
R6536 VDD.n951 VDD.n950 185.16
R6537 VDD.n955 VDD.n954 185.16
R6538 VDD.n979 VDD.n978 185.16
R6539 VDD.n981 VDD.n980 185.16
R6540 VDD.n973 VDD.n972 185.16
R6541 VDD.n961 VDD.n960 185.16
R6542 VDD.n959 VDD.n958 185.16
R6543 VDD.n963 VDD.n962 185.16
R6544 VDD.n967 VDD.n966 185.16
R6545 VDD.n969 VDD.n968 185.16
R6546 VDD.n949 VDD.n948 185.16
R6547 VDD.n991 VDD.n990 185.16
R6548 VDD.n993 VDD.n992 185.16
R6549 VDD.n896 VDD.n895 185.16
R6550 VDD.n900 VDD.n899 185.16
R6551 VDD.n902 VDD.n901 185.16
R6552 VDD.n906 VDD.n905 185.16
R6553 VDD.n880 VDD.n879 185.16
R6554 VDD.n878 VDD.n877 185.16
R6555 VDD.n874 VDD.n873 185.16
R6556 VDD.n912 VDD.n911 185.16
R6557 VDD.n914 VDD.n913 185.16
R6558 VDD.n918 VDD.n917 185.16
R6559 VDD.n872 VDD.n871 185.16
R6560 VDD.n870 VDD.n869 185.16
R6561 VDD.n868 VDD.n867 185.16
R6562 VDD.n924 VDD.n923 185.16
R6563 VDD.n926 VDD.n925 185.16
R6564 VDD.n856 VDD.n855 185.16
R6565 VDD.n824 VDD.n823 185.16
R6566 VDD.n822 VDD.n821 185.16
R6567 VDD.n826 VDD.n825 185.16
R6568 VDD.n850 VDD.n849 185.16
R6569 VDD.n852 VDD.n851 185.16
R6570 VDD.n844 VDD.n843 185.16
R6571 VDD.n832 VDD.n831 185.16
R6572 VDD.n830 VDD.n829 185.16
R6573 VDD.n834 VDD.n833 185.16
R6574 VDD.n838 VDD.n837 185.16
R6575 VDD.n840 VDD.n839 185.16
R6576 VDD.n820 VDD.n819 185.16
R6577 VDD.n862 VDD.n861 185.16
R6578 VDD.n864 VDD.n863 185.16
R6579 VDD.n767 VDD.n766 185.16
R6580 VDD.n771 VDD.n770 185.16
R6581 VDD.n773 VDD.n772 185.16
R6582 VDD.n777 VDD.n776 185.16
R6583 VDD.n751 VDD.n750 185.16
R6584 VDD.n749 VDD.n748 185.16
R6585 VDD.n745 VDD.n744 185.16
R6586 VDD.n783 VDD.n782 185.16
R6587 VDD.n785 VDD.n784 185.16
R6588 VDD.n789 VDD.n788 185.16
R6589 VDD.n743 VDD.n742 185.16
R6590 VDD.n741 VDD.n740 185.16
R6591 VDD.n739 VDD.n738 185.16
R6592 VDD.n795 VDD.n794 185.16
R6593 VDD.n797 VDD.n796 185.16
R6594 VDD.n727 VDD.n726 185.16
R6595 VDD.n695 VDD.n694 185.16
R6596 VDD.n693 VDD.n692 185.16
R6597 VDD.n697 VDD.n696 185.16
R6598 VDD.n721 VDD.n720 185.16
R6599 VDD.n723 VDD.n722 185.16
R6600 VDD.n715 VDD.n714 185.16
R6601 VDD.n703 VDD.n702 185.16
R6602 VDD.n701 VDD.n700 185.16
R6603 VDD.n705 VDD.n704 185.16
R6604 VDD.n709 VDD.n708 185.16
R6605 VDD.n711 VDD.n710 185.16
R6606 VDD.n691 VDD.n690 185.16
R6607 VDD.n733 VDD.n732 185.16
R6608 VDD.n735 VDD.n734 185.16
R6609 VDD.n638 VDD.n637 185.16
R6610 VDD.n592 VDD.n591 185.16
R6611 VDD.n590 VDD.n589 185.16
R6612 VDD.n594 VDD.n593 185.16
R6613 VDD.n632 VDD.n631 185.16
R6614 VDD.n634 VDD.n633 185.16
R6615 VDD.n626 VDD.n625 185.16
R6616 VDD.n600 VDD.n599 185.16
R6617 VDD.n598 VDD.n597 185.16
R6618 VDD.n616 VDD.n615 185.16
R6619 VDD.n620 VDD.n619 185.16
R6620 VDD.n622 VDD.n621 185.16
R6621 VDD.n588 VDD.n587 185.16
R6622 VDD.n644 VDD.n643 185.16
R6623 VDD.n646 VDD.n645 185.16
R6624 VDD.n576 VDD.n575 185.16
R6625 VDD.n544 VDD.n543 185.16
R6626 VDD.n542 VDD.n541 185.16
R6627 VDD.n546 VDD.n545 185.16
R6628 VDD.n570 VDD.n569 185.16
R6629 VDD.n572 VDD.n571 185.16
R6630 VDD.n564 VDD.n563 185.16
R6631 VDD.n552 VDD.n551 185.16
R6632 VDD.n550 VDD.n549 185.16
R6633 VDD.n554 VDD.n553 185.16
R6634 VDD.n558 VDD.n557 185.16
R6635 VDD.n560 VDD.n559 185.16
R6636 VDD.n540 VDD.n539 185.16
R6637 VDD.n582 VDD.n581 185.16
R6638 VDD.n584 VDD.n583 185.16
R6639 VDD.n487 VDD.n486 185.16
R6640 VDD.n491 VDD.n490 185.16
R6641 VDD.n493 VDD.n492 185.16
R6642 VDD.n497 VDD.n496 185.16
R6643 VDD.n471 VDD.n470 185.16
R6644 VDD.n469 VDD.n468 185.16
R6645 VDD.n465 VDD.n464 185.16
R6646 VDD.n503 VDD.n502 185.16
R6647 VDD.n505 VDD.n504 185.16
R6648 VDD.n509 VDD.n508 185.16
R6649 VDD.n463 VDD.n462 185.16
R6650 VDD.n461 VDD.n460 185.16
R6651 VDD.n459 VDD.n458 185.16
R6652 VDD.n515 VDD.n514 185.16
R6653 VDD.n517 VDD.n516 185.16
R6654 VDD.n447 VDD.n446 185.16
R6655 VDD.n415 VDD.n414 185.16
R6656 VDD.n413 VDD.n412 185.16
R6657 VDD.n417 VDD.n416 185.16
R6658 VDD.n441 VDD.n440 185.16
R6659 VDD.n443 VDD.n442 185.16
R6660 VDD.n435 VDD.n434 185.16
R6661 VDD.n423 VDD.n422 185.16
R6662 VDD.n421 VDD.n420 185.16
R6663 VDD.n425 VDD.n424 185.16
R6664 VDD.n429 VDD.n428 185.16
R6665 VDD.n431 VDD.n430 185.16
R6666 VDD.n411 VDD.n410 185.16
R6667 VDD.n453 VDD.n452 185.16
R6668 VDD.n455 VDD.n454 185.16
R6669 VDD.n358 VDD.n357 185.16
R6670 VDD.n362 VDD.n361 185.16
R6671 VDD.n364 VDD.n363 185.16
R6672 VDD.n368 VDD.n367 185.16
R6673 VDD.n342 VDD.n341 185.16
R6674 VDD.n340 VDD.n339 185.16
R6675 VDD.n336 VDD.n335 185.16
R6676 VDD.n374 VDD.n373 185.16
R6677 VDD.n376 VDD.n375 185.16
R6678 VDD.n380 VDD.n379 185.16
R6679 VDD.n334 VDD.n333 185.16
R6680 VDD.n332 VDD.n331 185.16
R6681 VDD.n330 VDD.n329 185.16
R6682 VDD.n386 VDD.n385 185.16
R6683 VDD.n388 VDD.n387 185.16
R6684 VDD.n318 VDD.n317 185.16
R6685 VDD.n286 VDD.n285 185.16
R6686 VDD.n284 VDD.n283 185.16
R6687 VDD.n288 VDD.n287 185.16
R6688 VDD.n312 VDD.n311 185.16
R6689 VDD.n314 VDD.n313 185.16
R6690 VDD.n306 VDD.n305 185.16
R6691 VDD.n294 VDD.n293 185.16
R6692 VDD.n292 VDD.n291 185.16
R6693 VDD.n296 VDD.n295 185.16
R6694 VDD.n300 VDD.n299 185.16
R6695 VDD.n302 VDD.n301 185.16
R6696 VDD.n282 VDD.n281 185.16
R6697 VDD.n324 VDD.n323 185.16
R6698 VDD.n326 VDD.n325 185.16
R6699 VDD.n189 VDD.n188 185.16
R6700 VDD.n157 VDD.n156 185.16
R6701 VDD.n155 VDD.n154 185.16
R6702 VDD.n159 VDD.n158 185.16
R6703 VDD.n183 VDD.n182 185.16
R6704 VDD.n185 VDD.n184 185.16
R6705 VDD.n177 VDD.n176 185.16
R6706 VDD.n165 VDD.n164 185.16
R6707 VDD.n163 VDD.n162 185.16
R6708 VDD.n167 VDD.n166 185.16
R6709 VDD.n171 VDD.n170 185.16
R6710 VDD.n173 VDD.n172 185.16
R6711 VDD.n153 VDD.n152 185.16
R6712 VDD.n195 VDD.n194 185.16
R6713 VDD.n197 VDD.n196 185.16
R6714 VDD.n229 VDD.n228 185.16
R6715 VDD.n233 VDD.n232 185.16
R6716 VDD.n235 VDD.n234 185.16
R6717 VDD.n239 VDD.n238 185.16
R6718 VDD.n213 VDD.n212 185.16
R6719 VDD.n211 VDD.n210 185.16
R6720 VDD.n207 VDD.n206 185.16
R6721 VDD.n245 VDD.n244 185.16
R6722 VDD.n247 VDD.n246 185.16
R6723 VDD.n251 VDD.n250 185.16
R6724 VDD.n205 VDD.n204 185.16
R6725 VDD.n203 VDD.n202 185.16
R6726 VDD.n201 VDD.n200 185.16
R6727 VDD.n257 VDD.n256 185.16
R6728 VDD.n259 VDD.n258 185.16
R6729 VDD.n91 VDD.n90 185.16
R6730 VDD.n95 VDD.n94 185.16
R6731 VDD.n97 VDD.n96 185.16
R6732 VDD.n101 VDD.n100 185.16
R6733 VDD.n75 VDD.n74 185.16
R6734 VDD.n73 VDD.n72 185.16
R6735 VDD.n69 VDD.n68 185.16
R6736 VDD.n107 VDD.n106 185.16
R6737 VDD.n109 VDD.n108 185.16
R6738 VDD.n113 VDD.n112 185.16
R6739 VDD.n67 VDD.n66 185.16
R6740 VDD.n65 VDD.n64 185.16
R6741 VDD.n63 VDD.n62 185.16
R6742 VDD.n119 VDD.n118 185.16
R6743 VDD.n121 VDD.n120 185.16
R6744 VDD.n2894 VDD.n2893 185.16
R6745 VDD.n2862 VDD.n2861 185.16
R6746 VDD.n2860 VDD.n2859 185.16
R6747 VDD.n2864 VDD.n2863 185.16
R6748 VDD.n2888 VDD.n2887 185.16
R6749 VDD.n2890 VDD.n2889 185.16
R6750 VDD.n2882 VDD.n2881 185.16
R6751 VDD.n2870 VDD.n2869 185.16
R6752 VDD.n2868 VDD.n2867 185.16
R6753 VDD.n2872 VDD.n2871 185.16
R6754 VDD.n2876 VDD.n2875 185.16
R6755 VDD.n2878 VDD.n2877 185.16
R6756 VDD.n2858 VDD.n2857 185.16
R6757 VDD.n2900 VDD.n2899 185.16
R6758 VDD.n2902 VDD.n2901 185.16
R6759 VDD.n29 VDD.n28 185.16
R6760 VDD.n33 VDD.n32 185.16
R6761 VDD.n35 VDD.n34 185.16
R6762 VDD.n39 VDD.n38 185.16
R6763 VDD.n13 VDD.n12 185.16
R6764 VDD.n11 VDD.n10 185.16
R6765 VDD.n7 VDD.n6 185.16
R6766 VDD.n45 VDD.n44 185.16
R6767 VDD.n47 VDD.n46 185.16
R6768 VDD.n51 VDD.n50 185.16
R6769 VDD.n5 VDD.n4 185.16
R6770 VDD.n3 VDD.n2 185.16
R6771 VDD.n1 VDD.n0 185.16
R6772 VDD.n57 VDD.n56 185.16
R6773 VDD.n59 VDD.n58 185.16
R6774 VDD.t2116 VDD.n1063 182.756
R6775 VDD.t2615 VDD.n934 182.756
R6776 VDD.t962 VDD.n805 182.756
R6777 VDD.t690 VDD.n654 182.756
R6778 VDD.t3283 VDD.n525 182.756
R6779 VDD.t1110 VDD.n396 182.756
R6780 VDD.t696 VDD.n267 182.756
R6781 VDD.t1322 VDD.n129 182.756
R6782 VDD.t3124 VDD.n2913 182.756
R6783 VDD.t1356 VDD.t1352 182.4
R6784 VDD.n674 VDD.t1460 179.731
R6785 VDD.t2102 VDD.t2104 175.386
R6786 VDD.t2100 VDD.t2102 175.386
R6787 VDD.t866 VDD.t870 175.386
R6788 VDD.t870 VDD.t868 175.386
R6789 VDD.t1928 VDD.t1930 175.386
R6790 VDD.t1930 VDD.t1942 175.386
R6791 VDD.t3383 VDD.t3385 175.386
R6792 VDD.t3395 VDD.t3383 175.386
R6793 VDD.t3520 VDD.t3524 175.386
R6794 VDD.t3516 VDD.t3520 175.386
R6795 VDD.t1078 VDD.t1886 175.386
R6796 VDD.t1076 VDD.t1078 175.386
R6797 VDD.t4002 VDD.t4004 175.386
R6798 VDD.t4000 VDD.t4002 175.386
R6799 VDD.t3407 VDD.t3411 175.386
R6800 VDD.t3411 VDD.t3409 175.386
R6801 VDD.t2784 VDD.t2782 175.386
R6802 VDD.t2782 VDD.t2778 175.386
R6803 VDD.t2012 VDD.t2010 175.386
R6804 VDD.t2010 VDD.t2020 175.386
R6805 VDD.t4008 VDD.t4006 175.386
R6806 VDD.t4006 VDD.t4016 175.386
R6807 VDD.t1894 VDD.t1900 175.386
R6808 VDD.t1892 VDD.t1894 175.386
R6809 VDD.t1693 VDD.t1695 175.386
R6810 VDD.t1697 VDD.t1693 175.386
R6811 VDD.t1468 VDD.t1466 175.386
R6812 VDD.t1464 VDD.t1468 175.386
R6813 VDD.t834 VDD.t836 175.386
R6814 VDD.t842 VDD.t834 175.386
R6815 VDD.t1285 VDD.t1281 175.386
R6816 VDD.t1281 VDD.t1283 175.386
R6817 VDD.t2443 VDD.t2441 175.386
R6818 VDD.t2441 VDD.t2437 175.386
R6819 VDD.t158 VDD.t154 175.386
R6820 VDD.t152 VDD.t158 175.386
R6821 VDD.t2070 VDD.t2074 175.386
R6822 VDD.t2072 VDD.t2070 175.386
R6823 VDD.t969 VDD.t967 175.386
R6824 VDD.t967 VDD.t965 175.386
R6825 VDD.t944 VDD.t942 175.386
R6826 VDD.t942 VDD.t946 175.386
R6827 VDD.t3661 VDD.t3663 175.386
R6828 VDD.t3659 VDD.t3661 175.386
R6829 VDD.t3320 VDD.t3322 175.386
R6830 VDD.t3314 VDD.t3320 175.386
R6831 VDD.t4058 VDD.t4056 175.386
R6832 VDD.t4056 VDD.t4052 175.386
R6833 VDD.t2743 VDD.t2741 175.386
R6834 VDD.t2745 VDD.t2743 175.386
R6835 VDD.t2213 VDD.t2217 175.386
R6836 VDD.t2215 VDD.t2213 175.386
R6837 VDD.t1956 VDD.t1966 175.386
R6838 VDD.t1952 VDD.t1956 175.386
R6839 VDD.t601 VDD.t1588 175.386
R6840 VDD.t1588 VDD.t1592 175.386
R6841 VDD.t3192 VDD.t3194 175.386
R6842 VDD.t3194 VDD.t3186 175.386
R6843 VDD.t2497 VDD.t2499 175.386
R6844 VDD.t2499 VDD.t2503 175.386
R6845 VDD.t3681 VDD.t3683 175.386
R6846 VDD.t3683 VDD.t3685 175.386
R6847 VDD.t4265 VDD.t4267 175.386
R6848 VDD.t4267 VDD.t4269 175.386
R6849 VDD.t4291 VDD.t4279 175.386
R6850 VDD.t4279 VDD.t4285 175.386
R6851 VDD.t3887 VDD.t3889 175.386
R6852 VDD.t3889 VDD.t3895 175.386
R6853 VDD.t103 VDD.t105 175.386
R6854 VDD.t105 VDD.t107 175.386
R6855 VDD.t3269 VDD.t3273 175.386
R6856 VDD.t3273 VDD.t3279 175.386
R6857 VDD.t4040 VDD.t4038 175.386
R6858 VDD.t4038 VDD.t4042 175.386
R6859 VDD.t4044 VDD.t4046 175.386
R6860 VDD.t4046 VDD.t4048 175.386
R6861 VDD.t3669 VDD.t3673 175.386
R6862 VDD.t3673 VDD.t3677 175.386
R6863 VDD.t660 VDD.t662 175.386
R6864 VDD.t662 VDD.t668 175.386
R6865 VDD.t20 VDD.t24 175.386
R6866 VDD.t24 VDD.t30 175.386
R6867 VDD.t4026 VDD.t4024 175.386
R6868 VDD.t4024 VDD.t4030 175.386
R6869 VDD.t573 VDD.t571 175.386
R6870 VDD.t571 VDD.t575 175.386
R6871 VDD.t144 VDD.t146 175.386
R6872 VDD.t146 VDD.t142 175.386
R6873 VDD.t4148 VDD.t4154 175.386
R6874 VDD.t4154 VDD.t4152 175.386
R6875 VDD.t1048 VDD.t1050 175.386
R6876 VDD.t1050 VDD.t2250 175.386
R6877 VDD.t4243 VDD.t4249 175.386
R6878 VDD.t4249 VDD.t3936 175.386
R6879 VDD.t2724 VDD.t2712 175.386
R6880 VDD.t2712 VDD.t2716 175.386
R6881 VDD.t223 VDD.t221 175.386
R6882 VDD.t225 VDD.t223 175.386
R6883 VDD.t2425 VDD.t2248 175.386
R6884 VDD.t2246 VDD.t2425 175.386
R6885 VDD.t1980 VDD.t1910 175.386
R6886 VDD.t1978 VDD.t1980 175.386
R6887 VDD.t1603 VDD.t2052 175.386
R6888 VDD.t2052 VDD.t2056 175.386
R6889 VDD.t1293 VDD.t1295 175.386
R6890 VDD.t1295 VDD.t1299 175.386
R6891 VDD.t295 VDD.t293 175.386
R6892 VDD.t283 VDD.t295 175.386
R6893 VDD.t714 VDD.t712 175.386
R6894 VDD.t716 VDD.t714 175.386
R6895 VDD.t2517 VDD.t2515 175.386
R6896 VDD.t2519 VDD.t2517 175.386
R6897 VDD.t219 VDD.t217 175.386
R6898 VDD.t209 VDD.t219 175.386
R6899 VDD.t4173 VDD.t4175 175.386
R6900 VDD.t4175 VDD.t4181 175.386
R6901 VDD.t2314 VDD.t2302 175.386
R6902 VDD.t2302 VDD.t2304 175.386
R6903 VDD.t1330 VDD.t1334 175.386
R6904 VDD.t1334 VDD.t1336 175.386
R6905 VDD.t117 VDD.t1129 175.386
R6906 VDD.t1129 VDD.t1131 175.386
R6907 VDD.t1084 VDD.t563 175.386
R6908 VDD.t563 VDD.t1082 175.386
R6909 VDD.t700 VDD.t702 175.386
R6910 VDD.t702 VDD.t706 175.386
R6911 VDD.t461 VDD.t459 175.386
R6912 VDD.t449 VDD.t461 175.386
R6913 VDD.t247 VDD.t243 175.386
R6914 VDD.t253 VDD.t247 175.386
R6915 VDD.t2915 VDD.t2913 175.386
R6916 VDD.t2913 VDD.t2909 175.386
R6917 VDD.t722 VDD.t720 175.386
R6918 VDD.t720 VDD.t718 175.386
R6919 VDD.t4327 VDD.t4325 175.386
R6920 VDD.t4329 VDD.t4327 175.386
R6921 VDD.t2565 VDD.t2561 175.386
R6922 VDD.t2563 VDD.t2565 175.386
R6923 VDD.t2737 VDD.t2739 175.386
R6924 VDD.t2739 VDD.t496 175.386
R6925 VDD.t1609 VDD.t636 175.386
R6926 VDD.t636 VDD.t1605 175.386
R6927 VDD.t1932 VDD.t1926 175.386
R6928 VDD.t1926 VDD.t1972 175.386
R6929 VDD.t1826 VDD.t1824 175.386
R6930 VDD.t1822 VDD.t1826 175.386
R6931 VDD.t3405 VDD.t3403 175.386
R6932 VDD.t3401 VDD.t3405 175.386
R6933 VDD.t1769 VDD.t1775 175.386
R6934 VDD.t1761 VDD.t1769 175.386
R6935 VDD.t2254 VDD.t2252 175.386
R6936 VDD.t2252 VDD.t2256 175.386
R6937 VDD.t2223 VDD.t2221 175.386
R6938 VDD.t2221 VDD.t2219 175.386
R6939 VDD.t2090 VDD.t2092 175.386
R6940 VDD.t2084 VDD.t2090 175.386
R6941 VDD.t2539 VDD.t1327 175.386
R6942 VDD.t2537 VDD.t2539 175.386
R6943 VDD.t1360 VDD.t1362 175.386
R6944 VDD.t1358 VDD.t1360 175.386
R6945 VDD.t803 VDD.t805 175.386
R6946 VDD.t801 VDD.t803 175.386
R6947 VDD.t752 VDD.t750 175.386
R6948 VDD.t750 VDD.t748 175.386
R6949 VDD.t4206 VDD.t4204 175.386
R6950 VDD.t4204 VDD.t4202 175.386
R6951 VDD.t4134 VDD.t4136 175.386
R6952 VDD.t4138 VDD.t4134 175.386
R6953 VDD.t445 VDD.t447 175.386
R6954 VDD.t443 VDD.t445 175.386
R6955 VDD.t3326 VDD.t3328 175.386
R6956 VDD.t3324 VDD.t3326 175.386
R6957 VDD.t84 VDD.t94 175.386
R6958 VDD.t82 VDD.t84 175.386
R6959 VDD.t2470 VDD.t2468 175.386
R6960 VDD.t2468 VDD.t2466 175.386
R6961 VDD.t265 VDD.t545 175.386
R6962 VDD.t545 VDD.t541 175.386
R6963 VDD.t343 VDD.t341 175.386
R6964 VDD.t341 VDD.t337 175.386
R6965 VDD.t2189 VDD.t2187 175.386
R6966 VDD.t2187 VDD.t2185 175.386
R6967 VDD.t1856 VDD.t1854 175.386
R6968 VDD.t1854 VDD.t1858 175.386
R6969 VDD.t1733 VDD.t1737 175.386
R6970 VDD.t1737 VDD.t1735 175.386
R6971 VDD.t1558 VDD.t1560 175.386
R6972 VDD.t1560 VDD.t1562 175.386
R6973 VDD.t4105 VDD.t4109 175.386
R6974 VDD.t4109 VDD.t4096 175.386
R6975 VDD.t613 VDD.t615 175.386
R6976 VDD.t611 VDD.t613 175.386
R6977 VDD.t3464 VDD.t908 175.386
R6978 VDD.t3462 VDD.t3464 175.386
R6979 VDD.t3996 VDD.t3998 175.386
R6980 VDD.t3994 VDD.t3996 175.386
R6981 VDD.t3944 VDD.t3940 175.386
R6982 VDD.t3942 VDD.t3944 175.386
R6983 VDD.t297 VDD.t301 175.386
R6984 VDD.t301 VDD.t299 175.386
R6985 VDD.t1625 VDD.t1629 175.386
R6986 VDD.t1629 VDD.t1627 175.386
R6987 VDD.t1431 VDD.t1433 175.386
R6988 VDD.t1433 VDD.t1435 175.386
R6989 VDD.t2700 VDD.t2704 175.386
R6990 VDD.t2704 VDD.t2702 175.386
R6991 VDD.t1851 VDD.t1849 175.386
R6992 VDD.t1849 VDD.t1847 175.386
R6993 VDD.t2756 VDD.t2760 175.386
R6994 VDD.t2760 VDD.t2758 175.386
R6995 VDD.t3906 VDD.t3910 175.386
R6996 VDD.t3910 VDD.t3908 175.386
R6997 VDD.t403 VDD.t407 175.386
R6998 VDD.t407 VDD.t405 175.386
R6999 VDD.t2882 VDD.t2878 175.386
R7000 VDD.t2880 VDD.t2882 175.386
R7001 VDD.t2476 VDD.t2472 175.386
R7002 VDD.t2474 VDD.t2476 175.386
R7003 VDD.t1586 VDD.t1582 175.386
R7004 VDD.t1584 VDD.t1586 175.386
R7005 VDD.t1117 VDD.t1119 175.386
R7006 VDD.t1121 VDD.t1117 175.386
R7007 VDD.t2401 VDD.t2407 175.386
R7008 VDD.t2407 VDD.t2405 175.386
R7009 VDD.t2836 VDD.t2841 175.386
R7010 VDD.t2841 VDD.t2839 175.386
R7011 VDD.t3238 VDD.t3242 175.386
R7012 VDD.t3242 VDD.t3240 175.386
R7013 VDD.t1840 VDD.t1844 175.386
R7014 VDD.t1844 VDD.t1842 175.386
R7015 VDD.t2694 VDD.t2690 175.386
R7016 VDD.t2692 VDD.t2694 175.386
R7017 VDD.t1878 VDD.t170 175.386
R7018 VDD.t1880 VDD.t1878 175.386
R7019 VDD.t3473 VDD.t3479 175.386
R7020 VDD.t3479 VDD.t3475 175.386
R7021 VDD.t3432 VDD.t3430 175.386
R7022 VDD.t3430 VDD.t3436 175.386
R7023 VDD.t3643 VDD.t3649 175.386
R7024 VDD.t3649 VDD.t3647 175.386
R7025 VDD.t2234 VDD.t2240 172.727
R7026 VDD.t2240 VDD.t1665 172.727
R7027 VDD.t999 VDD.t991 172.727
R7028 VDD.t1021 VDD.t999 172.727
R7029 VDD.t4212 VDD.t4210 172.727
R7030 VDD.t4228 VDD.t4212 172.727
R7031 VDD.t1034 VDD.t583 172.727
R7032 VDD.t583 VDD.t989 172.727
R7033 VDD.t263 VDD.t553 172.727
R7034 VDD.t517 VDD.t263 172.727
R7035 VDD.t995 VDD.t1002 172.727
R7036 VDD.t1002 VDD.t1026 172.727
R7037 VDD.t4087 VDD.t4085 172.727
R7038 VDD.t4085 VDD.t4091 172.727
R7039 VDD.t593 VDD.t1015 172.727
R7040 VDD.t1015 VDD.t1017 172.727
R7041 VDD.t1393 VDD.t1167 169.833
R7042 VDD.t787 VDD.t789 169.833
R7043 VDD.t3486 VDD.t3488 169.833
R7044 VDD.t4186 VDD.t4219 168.267
R7045 VDD.t4219 VDD.t4241 168.267
R7046 VDD.t2138 VDD.t2178 168.267
R7047 VDD.t2178 VDD.t2172 168.267
R7048 VDD.t4111 VDD.t4107 168.267
R7049 VDD.t4107 VDD.t4079 168.267
R7050 VDD.t2145 VDD.t2141 168.267
R7051 VDD.t2141 VDD.t2124 168.267
R7052 VDD.t2136 VDD.t2176 168.267
R7053 VDD.t2176 VDD.t2134 168.267
R7054 VDD.t2236 VDD.t1681 168.267
R7055 VDD.t1681 VDD.t1674 168.267
R7056 VDD.t2174 VDD.t2170 168.267
R7057 VDD.t2170 VDD.t2143 168.267
R7058 VDD.t259 VDD.t555 168.267
R7059 VDD.t555 VDD.t533 168.267
R7060 VDD.t2598 VDD.t471 168.267
R7061 VDD.t471 VDD.t469 168.267
R7062 VDD.t2242 VDD.t1667 168.267
R7063 VDD.t1667 VDD.t1669 168.267
R7064 VDD.t2585 VDD.t2590 168.267
R7065 VDD.t2590 VDD.t2613 168.267
R7066 VDD.t535 VDD.t543 168.267
R7067 VDD.t543 VDD.t547 168.267
R7068 VDD.t4217 VDD.t4237 168.267
R7069 VDD.t4237 VDD.t4235 168.267
R7070 VDD.t2322 VDD.t2349 168.267
R7071 VDD.t2349 VDD.t2351 168.267
R7072 VDD.t4068 VDD.t4075 168.267
R7073 VDD.t4075 VDD.t4103 168.267
R7074 VDD.t2356 VDD.t2366 168.267
R7075 VDD.t2366 VDD.t2372 168.267
R7076 VDD.t2374 VDD.t2368 168.267
R7077 VDD.t2327 VDD.t2374 168.267
R7078 VDD.t514 VDD.t521 168.267
R7079 VDD.t521 VDD.t523 168.267
R7080 VDD.n1135 VDD.t3500 164.272
R7081 VDD.t2335 VDD.t2360 163.441
R7082 VDD.t2360 VDD.t2358 163.441
R7083 VDD.t2229 VDD.t1655 163.441
R7084 VDD.t1655 VDD.t1663 163.441
R7085 VDD.t1597 VDD.t1599 158.609
R7086 VDD.t632 VDD.t1597 158.609
R7087 VDD.t630 VDD.t632 158.609
R7088 VDD.t1308 VDD.t1306 158.609
R7089 VDD.t1306 VDD.t1325 158.609
R7090 VDD.t1325 VDD.t1323 158.609
R7091 VDD.t791 VDD.t793 158.609
R7092 VDD.t3220 VDD.t791 158.609
R7093 VDD.t3216 VDD.t3220 158.609
R7094 VDD.t4407 VDD.t4508 158.609
R7095 VDD.t4508 VDD.t3182 158.609
R7096 VDD.t3182 VDD.t3180 158.609
R7097 VDD.t914 VDD.t916 158.609
R7098 VDD.t2109 VDD.t914 158.609
R7099 VDD.t2107 VDD.t2109 158.609
R7100 VDD.t2397 VDD.t80 158.609
R7101 VDD.t80 VDD.t4331 158.609
R7102 VDD.t4331 VDD.t4333 158.609
R7103 VDD.t4293 VDD.t4295 158.609
R7104 VDD.t1540 VDD.t4293 158.609
R7105 VDD.t2848 VDD.t1540 158.609
R7106 VDD.t658 VDD.t656 158.609
R7107 VDD.t656 VDD.t1348 158.609
R7108 VDD.t1348 VDD.t1350 158.609
R7109 VDD.t437 VDD.t435 158.609
R7110 VDD.t2529 VDD.t437 158.609
R7111 VDD.t2531 VDD.t2529 158.609
R7112 VDD.t4474 VDD.t4367 158.609
R7113 VDD.t4367 VDD.t2798 158.609
R7114 VDD.t2798 VDD.t2806 158.609
R7115 VDD.t2642 VDD.t2644 158.609
R7116 VDD.t3115 VDD.t2642 158.609
R7117 VDD.t3117 VDD.t3115 158.609
R7118 VDD.t1191 VDD.t1193 158.609
R7119 VDD.t1193 VDD.t1457 158.609
R7120 VDD.t1457 VDD.t1455 158.609
R7121 VDD.t923 VDD.t921 158.609
R7122 VDD.t1218 VDD.t923 158.609
R7123 VDD.t1220 VDD.t1218 158.609
R7124 VDD.t2850 VDD.t2852 158.609
R7125 VDD.t2852 VDD.t3351 158.609
R7126 VDD.t3351 VDD.t3353 158.609
R7127 VDD.t2794 VDD.t2792 158.609
R7128 VDD.t3359 VDD.t2794 158.609
R7129 VDD.t3363 VDD.t3359 158.609
R7130 VDD.t4391 VDD.t4458 158.609
R7131 VDD.t4458 VDD.t125 158.609
R7132 VDD.t125 VDD.t133 158.609
R7133 VDD.t2788 VDD.t2786 158.609
R7134 VDD.t818 VDD.t2788 158.609
R7135 VDD.t820 VDD.t818 158.609
R7136 VDD.t1888 VDD.t1890 158.609
R7137 VDD.t1890 VDD.t2485 158.609
R7138 VDD.t2485 VDD.t795 158.609
R7139 VDD.t4022 VDD.t4020 158.609
R7140 VDD.t230 VDD.t4022 158.609
R7141 VDD.t228 VDD.t230 158.609
R7142 VDD.t1868 VDD.t1870 158.609
R7143 VDD.t1870 VDD.t4169 158.609
R7144 VDD.t4169 VDD.t4167 158.609
R7145 VDD.t1213 VDD.t1211 158.609
R7146 VDD.t1421 VDD.t1213 158.609
R7147 VDD.t1423 VDD.t1421 158.609
R7148 VDD.t3575 VDD.t3577 158.609
R7149 VDD.t3577 VDD.t3415 158.609
R7150 VDD.t3415 VDD.t3413 158.609
R7151 VDD.t1366 VDD.t1364 158.609
R7152 VDD.t1364 VDD.t3083 158.609
R7153 VDD.t3083 VDD.t3067 158.609
R7154 VDD.t3635 VDD.t3631 158.609
R7155 VDD.t1380 VDD.t3635 158.609
R7156 VDD.t1382 VDD.t1380 158.609
R7157 VDD.t3349 VDD.t3347 158.609
R7158 VDD.t1988 VDD.t3349 158.609
R7159 VDD.t1990 VDD.t1988 158.609
R7160 VDD.t3637 VDD.t3623 158.609
R7161 VDD.t3623 VDD.t1368 158.609
R7162 VDD.t1368 VDD.t1372 158.609
R7163 VDD.t2041 VDD.t2043 158.609
R7164 VDD.t2043 VDD.t2986 158.609
R7165 VDD.t2986 VDD.t3087 158.609
R7166 VDD.t4439 VDD.t4364 158.609
R7167 VDD.t1374 VDD.t4439 158.609
R7168 VDD.t1376 VDD.t1374 158.609
R7169 VDD.t874 VDD.t872 158.609
R7170 VDD.t1994 VDD.t874 158.609
R7171 VDD.t1721 VDD.t1994 158.609
R7172 VDD.t4510 VDD.t4417 158.609
R7173 VDD.t4417 VDD.t1370 158.609
R7174 VDD.t1370 VDD.t1378 158.609
R7175 VDD.t1155 VDD.t1153 158.609
R7176 VDD.t4247 VDD.t1155 158.609
R7177 VDD.t4245 VDD.t4247 158.609
R7178 VDD.t2696 VDD.t2698 158.609
R7179 VDD.t2698 VDD.t234 158.609
R7180 VDD.t234 VDD.t232 158.609
R7181 VDD.t504 VDD.t502 158.609
R7182 VDD.t2050 VDD.t504 158.609
R7183 VDD.t197 VDD.t2050 158.609
R7184 VDD.t4395 VDD.t4460 158.609
R7185 VDD.t4460 VDD.t3133 158.609
R7186 VDD.t3133 VDD.t3141 158.609
R7187 VDD.t512 VDD.t510 158.609
R7188 VDD.t4263 VDD.t512 158.609
R7189 VDD.t4261 VDD.t4263 158.609
R7190 VDD.t2547 VDD.t2549 158.609
R7191 VDD.t2549 VDD.t958 158.609
R7192 VDD.t958 VDD.t956 158.609
R7193 VDD.t2039 VDD.t2037 158.609
R7194 VDD.t2096 VDD.t2039 158.609
R7195 VDD.t2098 VDD.t2096 158.609
R7196 VDD.t2864 VDD.t2866 158.609
R7197 VDD.t2866 VDD.t49 158.609
R7198 VDD.t49 VDD.t47 158.609
R7199 VDD.t1234 VDD.t1232 158.609
R7200 VDD.t3159 VDD.t1234 158.609
R7201 VDD.t3161 VDD.t3159 158.609
R7202 VDD.t4467 VDD.t4351 158.609
R7203 VDD.t4351 VDD.t1503 158.609
R7204 VDD.t1503 VDD.t1511 158.609
R7205 VDD.t1472 VDD.t1470 158.609
R7206 VDD.t1160 VDD.t1472 158.609
R7207 VDD.t1162 VDD.t1160 158.609
R7208 VDD.t3334 VDD.t3336 158.609
R7209 VDD.t3336 VDD.t168 158.609
R7210 VDD.t168 VDD.t166 158.609
R7211 VDD.t2286 VDD.t2284 158.609
R7212 VDD.t355 VDD.t2286 158.609
R7213 VDD.t353 VDD.t355 158.609
R7214 VDD.t1442 VDD.t1444 158.609
R7215 VDD.t1444 VDD.t2571 158.609
R7216 VDD.t2571 VDD.t2569 158.609
R7217 VDD.t492 VDD.t490 158.609
R7218 VDD.t271 VDD.t492 158.609
R7219 VDD.t273 VDD.t271 158.609
R7220 VDD.t2025 VDD.t2027 158.609
R7221 VDD.t2027 VDD.t413 158.609
R7222 VDD.t413 VDD.t2064 158.609
R7223 VDD.t508 VDD.t506 158.609
R7224 VDD.t12 VDD.t508 158.609
R7225 VDD.t2453 VDD.t12 158.609
R7226 VDD.t4476 VDD.t4369 158.609
R7227 VDD.t4369 VDD.t421 158.609
R7228 VDD.t421 VDD.t429 158.609
R7229 VDD.t910 VDD.t912 158.609
R7230 VDD.t2765 VDD.t910 158.609
R7231 VDD.t2767 VDD.t2765 158.609
R7232 VDD.t1451 VDD.t1453 158.609
R7233 VDD.t1453 VDD.t864 158.609
R7234 VDD.t864 VDD.t862 158.609
R7235 VDD.t577 VDD.t579 158.609
R7236 VDD.t1269 VDD.t577 158.609
R7237 VDD.t1265 VDD.t1269 158.609
R7238 VDD.t4444 VDD.t4377 158.609
R7239 VDD.t4377 VDD.t1709 158.609
R7240 VDD.t1709 VDD.t1707 158.609
R7241 VDD.t768 VDD.t770 158.609
R7242 VDD.t4064 VDD.t768 158.609
R7243 VDD.t925 VDD.t4064 158.609
R7244 VDD.t932 VDD.t930 158.609
R7245 VDD.t930 VDD.t3330 158.609
R7246 VDD.t3330 VDD.t3332 158.609
R7247 VDD.t1257 VDD.t1255 158.609
R7248 VDD.t2066 VDD.t1257 158.609
R7249 VDD.t2068 VDD.t2066 158.609
R7250 VDD.t1070 VDD.t1068 158.609
R7251 VDD.t1068 VDD.t1499 158.609
R7252 VDD.t1499 VDD.t1501 158.609
R7253 VDD.t1968 VDD.t1914 158.609
R7254 VDD.t856 VDD.t1968 158.609
R7255 VDD.t858 VDD.t856 158.609
R7256 VDD.t4362 VDD.t4450 158.609
R7257 VDD.t4450 VDD.t2897 158.609
R7258 VDD.t2897 VDD.t2887 158.609
R7259 VDD.t2207 VDD.t2205 158.609
R7260 VDD.t1743 VDD.t2207 158.609
R7261 VDD.t1741 VDD.t1743 158.609
R7262 VDD.t372 VDD.t374 158.609
R7263 VDD.t374 VDD.t1244 158.609
R7264 VDD.t1244 VDD.t1246 158.609
R7265 VDD.t809 VDD.t807 158.333
R7266 VDD.t807 VDD.t3095 158.333
R7267 VDD.t3095 VDD.t2939 158.333
R7268 VDD.t76 VDD.t78 158.333
R7269 VDD.t3753 VDD.t76 158.333
R7270 VDD.t3746 VDD.t3753 158.333
R7271 VDD.t3693 VDD.t3695 158.333
R7272 VDD.t1263 VDD.t3693 158.333
R7273 VDD.t1259 VDD.t1263 158.333
R7274 VDD.t74 VDD.t70 158.333
R7275 VDD.t70 VDD.t3731 158.333
R7276 VDD.t3731 VDD.t3710 158.333
R7277 VDD.t1060 VDD.t1062 158.333
R7278 VDD.t1062 VDD.t2966 158.333
R7279 VDD.t2966 VDD.t3008 158.333
R7280 VDD.t4337 VDD.t4419 158.333
R7281 VDD.t3864 VDD.t4337 158.333
R7282 VDD.t3834 VDD.t3864 158.333
R7283 VDD.t2380 VDD.t2382 158.333
R7284 VDD.t1271 VDD.t2380 158.333
R7285 VDD.t1267 VDD.t1271 158.333
R7286 VDD.t4446 VDD.t4385 158.333
R7287 VDD.t4385 VDD.t3720 158.333
R7288 VDD.t3720 VDD.t3712 158.333
R7289 VDD.t2209 VDD.t2211 158.333
R7290 VDD.t2211 VDD.t2970 158.333
R7291 VDD.t2970 VDD.t2984 158.333
R7292 VDD.t3208 VDD.t3210 158.333
R7293 VDD.t3735 VDD.t3208 158.333
R7294 VDD.t3718 VDD.t3735 158.333
R7295 VDD.t62 VDD.t64 158.333
R7296 VDD.t3230 VDD.t62 158.333
R7297 VDD.t3226 VDD.t3230 158.333
R7298 VDD.t3206 VDD.t3202 158.333
R7299 VDD.t3202 VDD.t3877 158.333
R7300 VDD.t3877 VDD.t3850 158.333
R7301 VDD.t625 VDD.t623 158.333
R7302 VDD.t623 VDD.t2990 158.333
R7303 VDD.t2990 VDD.t3051 158.333
R7304 VDD.t4483 VDD.t4371 158.333
R7305 VDD.t3803 VDD.t4483 158.333
R7306 VDD.t3783 VDD.t3803 158.333
R7307 VDD.t1250 VDD.t1248 158.333
R7308 VDD.t3222 VDD.t1250 158.333
R7309 VDD.t3218 VDD.t3222 158.333
R7310 VDD.t4415 VDD.t4335 158.333
R7311 VDD.t4335 VDD.t3858 158.333
R7312 VDD.t3858 VDD.t3852 158.333
R7313 VDD.t1725 VDD.t1723 158.333
R7314 VDD.t1723 VDD.t3048 158.333
R7315 VDD.t3048 VDD.t3040 158.333
R7316 VDD.t2673 VDD.t2671 158.333
R7317 VDD.t3706 VDD.t2673 158.333
R7318 VDD.t3716 VDD.t3706 158.333
R7319 VDD.t1207 VDD.t1209 158.333
R7320 VDD.t2525 VDD.t1207 158.333
R7321 VDD.t2527 VDD.t2525 158.333
R7322 VDD.t2679 VDD.t2681 158.333
R7323 VDD.t2681 VDD.t3738 158.333
R7324 VDD.t3738 VDD.t3742 158.333
R7325 VDD.t1138 VDD.t1140 158.333
R7326 VDD.t1140 VDD.t3004 158.333
R7327 VDD.t3004 VDD.t2935 158.333
R7328 VDD.t4413 VDD.t4506 158.333
R7329 VDD.t3750 VDD.t4413 158.333
R7330 VDD.t3755 VDD.t3750 158.333
R7331 VDD.t3399 VDD.t3397 158.333
R7332 VDD.t2533 VDD.t3399 158.333
R7333 VDD.t2535 VDD.t2533 158.333
R7334 VDD.t4489 VDD.t4383 158.333
R7335 VDD.t4383 VDD.t3740 158.333
R7336 VDD.t3740 VDD.t3775 158.333
R7337 VDD.t3573 VDD.t3571 158.333
R7338 VDD.t3571 VDD.t3091 158.333
R7339 VDD.t3091 VDD.t3080 158.333
R7340 VDD.t3256 VDD.t3254 158.333
R7341 VDD.t3838 VDD.t3256 158.333
R7342 VDD.t3848 VDD.t3838 158.333
R7343 VDD.t45 VDD.t43 158.333
R7344 VDD.t3369 VDD.t45 158.333
R7345 VDD.t3373 VDD.t3369 158.333
R7346 VDD.t3248 VDD.t3252 158.333
R7347 VDD.t3252 VDD.t3807 158.333
R7348 VDD.t3807 VDD.t3823 158.333
R7349 VDD.t1620 VDD.t1622 158.333
R7350 VDD.t1622 VDD.t2925 158.333
R7351 VDD.t2925 VDD.t3030 158.333
R7352 VDD.t4491 VDD.t4427 158.333
R7353 VDD.t3846 VDD.t4491 158.333
R7354 VDD.t3866 VDD.t3846 158.333
R7355 VDD.t1866 VDD.t1864 158.333
R7356 VDD.t3361 VDD.t1866 158.333
R7357 VDD.t3365 VDD.t3361 158.333
R7358 VDD.t4399 VDD.t4463 158.333
R7359 VDD.t4463 VDD.t3813 158.333
R7360 VDD.t3813 VDD.t3700 158.333
R7361 VDD.t3956 VDD.t3954 158.333
R7362 VDD.t3954 VDD.t3089 158.333
R7363 VDD.t3089 VDD.t3074 158.333
R7364 VDD.t3633 VDD.t3629 158.333
R7365 VDD.t3842 VDD.t3633 158.333
R7366 VDD.t3856 VDD.t3842 158.333
R7367 VDD.t4132 VDD.t4130 158.333
R7368 VDD.t1992 VDD.t4132 158.333
R7369 VDD.t1996 VDD.t1992 158.333
R7370 VDD.t3625 VDD.t3627 158.333
R7371 VDD.t3627 VDD.t3811 158.333
R7372 VDD.t3811 VDD.t3825 158.333
R7373 VDD.t174 VDD.t176 158.333
R7374 VDD.t176 VDD.t3099 158.333
R7375 VDD.t3099 VDD.t3024 158.333
R7376 VDD.t4495 VDD.t4429 158.333
R7377 VDD.t3854 VDD.t4495 158.333
R7378 VDD.t3868 VDD.t3854 158.333
R7379 VDD.t1488 VDD.t1486 158.333
R7380 VDD.t1984 VDD.t1488 158.333
R7381 VDD.t1986 VDD.t1984 158.333
R7382 VDD.t4401 VDD.t4465 158.333
R7383 VDD.t4465 VDD.t3817 158.333
R7384 VDD.t3817 VDD.t3702 158.333
R7385 VDD.t51 VDD.t53 158.333
R7386 VDD.t53 VDD.t2961 158.333
R7387 VDD.t2961 VDD.t2947 158.333
R7388 VDD.t185 VDD.t183 158.333
R7389 VDD.t3787 VDD.t185 158.333
R7390 VDD.t3799 VDD.t3787 158.333
R7391 VDD.t1203 VDD.t1201 158.333
R7392 VDD.t199 VDD.t1203 158.333
R7393 VDD.t201 VDD.t199 158.333
R7394 VDD.t179 VDD.t181 158.333
R7395 VDD.t181 VDD.t3762 158.333
R7396 VDD.t3762 VDD.t3772 158.333
R7397 VDD.t2111 VDD.t844 158.333
R7398 VDD.t844 VDD.t2980 158.333
R7399 VDD.t2980 VDD.t3065 158.333
R7400 VDD.t4452 VDD.t4381 158.333
R7401 VDD.t3796 VDD.t4452 158.333
R7402 VDD.t3805 VDD.t3796 158.333
R7403 VDD.t2790 VDD.t1567 158.333
R7404 VDD.t207 VDD.t2790 158.333
R7405 VDD.t2048 VDD.t207 158.333
R7406 VDD.t4343 VDD.t4432 158.333
R7407 VDD.t4432 VDD.t3767 158.333
R7408 VDD.t3767 VDD.t3827 158.333
R7409 VDD.t2282 VDD.t2280 158.333
R7410 VDD.t2280 VDD.t3085 158.333
R7411 VDD.t3085 VDD.t3069 158.333
R7412 VDD.t2661 VDD.t2659 158.333
R7413 VDD.t3844 VDD.t2661 158.333
R7414 VDD.t3862 VDD.t3844 158.333
R7415 VDD.t3992 VDD.t3990 158.333
R7416 VDD.t3163 VDD.t3992 158.333
R7417 VDD.t3165 VDD.t3163 158.333
R7418 VDD.t2655 VDD.t2657 158.333
R7419 VDD.t2657 VDD.t3815 158.333
R7420 VDD.t3815 VDD.t3829 158.333
R7421 VDD.t1064 VDD.t1066 158.333
R7422 VDD.t1066 VDD.t3097 158.333
R7423 VDD.t3097 VDD.t3020 158.333
R7424 VDD.t4499 VDD.t4434 158.333
R7425 VDD.t3860 VDD.t4499 158.333
R7426 VDD.t3874 VDD.t3860 158.333
R7427 VDD.t1862 VDD.t1860 158.333
R7428 VDD.t3151 VDD.t1862 158.333
R7429 VDD.t3155 VDD.t3151 158.333
R7430 VDD.t4403 VDD.t4469 158.333
R7431 VDD.t4469 VDD.t3821 158.333
R7432 VDD.t3821 VDD.t3704 158.333
R7433 VDD.t415 VDD.t417 158.333
R7434 VDD.t417 VDD.t2997 158.333
R7435 VDD.t2997 VDD.t2992 158.333
R7436 VDD.t569 VDD.t567 158.333
R7437 VDD.t3744 VDD.t569 158.333
R7438 VDD.t3748 VDD.t3744 158.333
R7439 VDD.t3267 VDD.t3265 158.333
R7440 VDD.t10 VDD.t3267 158.333
R7441 VDD.t2451 VDD.t10 158.333
R7442 VDD.t323 VDD.t325 158.333
R7443 VDD.t325 VDD.t3764 158.333
R7444 VDD.t3764 VDD.t3778 158.333
R7445 VDD.t279 VDD.t281 158.333
R7446 VDD.t281 VDD.t2978 158.333
R7447 VDD.t2978 VDD.t3062 158.333
R7448 VDD.t4454 VDD.t4387 158.333
R7449 VDD.t3801 VDD.t4454 158.333
R7450 VDD.t3809 VDD.t3801 158.333
R7451 VDD.t359 VDD.t357 158.333
R7452 VDD.t2455 VDD.t359 158.333
R7453 VDD.t4 VDD.t2455 158.333
R7454 VDD.t4349 VDD.t4436 158.333
R7455 VDD.t4436 VDD.t3770 158.333
R7456 VDD.t3770 VDD.t3832 158.333
R7457 VDD.t1964 VDD.t1922 158.333
R7458 VDD.t1922 VDD.t2923 158.333
R7459 VDD.t2923 VDD.t3076 158.333
R7460 VDD.t650 VDD.t646 158.333
R7461 VDD.t3759 VDD.t650 158.333
R7462 VDD.t3785 VDD.t3759 158.333
R7463 VDD.t1908 VDD.t1950 158.333
R7464 VDD.t848 VDD.t1908 158.333
R7465 VDD.t850 VDD.t848 158.333
R7466 VDD.t652 VDD.t654 158.333
R7467 VDD.t654 VDD.t3793 158.333
R7468 VDD.t3793 VDD.t3819 158.333
R7469 VDD.t2511 VDD.t2513 158.333
R7470 VDD.t2513 VDD.t3046 158.333
R7471 VDD.t3046 VDD.t2931 158.333
R7472 VDD.t4472 VDD.t4341 158.333
R7473 VDD.t3840 VDD.t4472 158.333
R7474 VDD.t3870 VDD.t3840 158.333
R7475 VDD.t1685 VDD.t1683 158.333
R7476 VDD.t860 VDD.t1685 158.333
R7477 VDD.t846 VDD.t860 158.333
R7478 VDD.t4375 VDD.t4493 158.333
R7479 VDD.t4493 VDD.t3872 158.333
R7480 VDD.t3872 VDD.t3780 158.333
R7481 VDD.t1654 VDD.t1653 158.06
R7482 VDD.t1671 VDD.t1654 158.06
R7483 VDD.t1676 VDD.t1671 158.06
R7484 VDD.t2233 VDD.t1676 158.06
R7485 VDD.t587 VDD.t2233 158.06
R7486 VDD.t589 VDD.t587 158.06
R7487 VDD.t1006 VDD.t589 158.06
R7488 VDD.t1009 VDD.t1030 158.06
R7489 VDD.t4234 VDD.t4227 158.06
R7490 VDD.t4198 VDD.t4234 158.06
R7491 VDD.t4201 VDD.t4198 158.06
R7492 VDD.t4216 VDD.t4201 158.06
R7493 VDD.t2376 VDD.t4216 158.06
R7494 VDD.t2378 VDD.t2376 158.06
R7495 VDD.t2333 VDD.t2378 158.06
R7496 VDD.t2337 VDD.t2362 158.06
R7497 VDD.t528 VDD.t527 158.06
R7498 VDD.t551 VDD.t528 158.06
R7499 VDD.t552 VDD.t551 158.06
R7500 VDD.t516 VDD.t552 158.06
R7501 VDD.t2605 VDD.t516 158.06
R7502 VDD.t2611 VDD.t2605 158.06
R7503 VDD.t2575 VDD.t2611 158.06
R7504 VDD.t2577 VDD.t2596 158.06
R7505 VDD.t4098 VDD.t4095 158.06
R7506 VDD.t4115 VDD.t4098 158.06
R7507 VDD.t4118 VDD.t4115 158.06
R7508 VDD.t4072 VDD.t4118 158.06
R7509 VDD.t2160 VDD.t4072 158.06
R7510 VDD.t2166 VDD.t2160 158.06
R7511 VDD.t2122 VDD.t2166 158.06
R7512 VDD.t2128 VDD.t2147 158.06
R7513 VDD.t1643 VDD.t1642 158.06
R7514 VDD.t2203 VDD.t1643 158.06
R7515 VDD.t2204 VDD.t2203 158.06
R7516 VDD.t1637 VDD.t2204 158.06
R7517 VDD.t3606 VDD.t1637 158.06
R7518 VDD.t3608 VDD.t3606 158.06
R7519 VDD.t3586 VDD.t3608 158.06
R7520 VDD.t3590 VDD.t3598 158.06
R7521 VDD.t390 VDD.t389 158.06
R7522 VDD.t399 VDD.t390 158.06
R7523 VDD.t400 VDD.t399 158.06
R7524 VDD.t378 VDD.t400 158.06
R7525 VDD.t3961 VDD.t378 158.06
R7526 VDD.t3964 VDD.t3961 158.06
R7527 VDD.t3977 VDD.t3964 158.06
R7528 VDD.t3983 VDD.t895 158.06
R7529 VDD.t2816 VDD.t2838 158.06
R7530 VDD.t2821 VDD.t2816 158.06
R7531 VDD.t2822 VDD.t2821 158.06
R7532 VDD.t2829 VDD.t2822 158.06
R7533 VDD.t3535 VDD.t2829 158.06
R7534 VDD.t3541 VDD.t3535 158.06
R7535 VDD.t3550 VDD.t3541 158.06
R7536 VDD.t3552 VDD.t3566 158.06
R7537 VDD.t3449 VDD.t3446 158.06
R7538 VDD.t2298 VDD.t3449 158.06
R7539 VDD.t2299 VDD.t2298 158.06
R7540 VDD.t3429 VDD.t2299 158.06
R7541 VDD.t1170 VDD.t3429 158.06
R7542 VDD.t1172 VDD.t1170 158.06
R7543 VDD.t1398 VDD.t1172 158.06
R7544 VDD.t1400 VDD.t1416 158.06
R7545 VDD.t2031 VDD.t2029 158.06
R7546 VDD.t2029 VDD.t3078 158.06
R7547 VDD.t3078 VDD.t3101 158.06
R7548 VDD.t3212 VDD.t3214 158.06
R7549 VDD.t3172 VDD.t3212 158.06
R7550 VDD.t3170 VDD.t3172 158.06
R7551 VDD.t1534 VDD.t1532 158.06
R7552 VDD.t3228 VDD.t1534 158.06
R7553 VDD.t3224 VDD.t3228 158.06
R7554 VDD.t3204 VDD.t3200 158.06
R7555 VDD.t3200 VDD.t3184 158.06
R7556 VDD.t3184 VDD.t3178 158.06
R7557 VDD.t950 VDD.t948 158.06
R7558 VDD.t948 VDD.t2994 158.06
R7559 VDD.t2994 VDD.t3057 158.06
R7560 VDD.t4479 VDD.t4360 158.06
R7561 VDD.t3176 VDD.t4479 158.06
R7562 VDD.t3174 VDD.t3176 158.06
R7563 VDD.t2115 VDD.t2116 158.06
R7564 VDD.t2114 VDD.t2115 158.06
R7565 VDD.t2113 VDD.t2114 158.06
R7566 VDD.t2117 VDD.t2113 158.06
R7567 VDD.t40 VDD.t2117 158.06
R7568 VDD.t38 VDD.t40 158.06
R7569 VDD.t36 VDD.t38 158.06
R7570 VDD.t34 VDD.t32 158.06
R7571 VDD.t1646 VDD.t1648 158.06
R7572 VDD.t1648 VDD.t2959 158.06
R7573 VDD.t2959 VDD.t2945 158.06
R7574 VDD.t2669 VDD.t2667 158.06
R7575 VDD.t2808 VDD.t2669 158.06
R7576 VDD.t2810 VDD.t2808 158.06
R7577 VDD.t0 VDD.t2 158.06
R7578 VDD.t2521 VDD.t0 158.06
R7579 VDD.t2523 VDD.t2521 158.06
R7580 VDD.t2675 VDD.t2677 158.06
R7581 VDD.t2677 VDD.t2796 158.06
R7582 VDD.t2796 VDD.t2800 158.06
R7583 VDD.t1490 VDD.t1492 158.06
R7584 VDD.t1492 VDD.t3014 158.06
R7585 VDD.t3014 VDD.t2963 158.06
R7586 VDD.t4393 VDD.t4501 158.06
R7587 VDD.t2802 VDD.t4393 158.06
R7588 VDD.t2804 VDD.t2802 158.06
R7589 VDD.t2616 VDD.t2615 158.06
R7590 VDD.t2617 VDD.t2616 158.06
R7591 VDD.t2618 VDD.t2617 158.06
R7592 VDD.t2619 VDD.t2618 158.06
R7593 VDD.t3928 VDD.t2619 158.06
R7594 VDD.t3920 VDD.t3928 158.06
R7595 VDD.t3924 VDD.t3920 158.06
R7596 VDD.t3922 VDD.t3926 158.06
R7597 VDD.t16 VDD.t14 158.06
R7598 VDD.t14 VDD.t3034 158.06
R7599 VDD.t3034 VDD.t3018 158.06
R7600 VDD.t3260 VDD.t3258 158.06
R7601 VDD.t119 VDD.t3260 158.06
R7602 VDD.t121 VDD.t119 158.06
R7603 VDD.t241 VDD.t239 158.06
R7604 VDD.t3367 VDD.t241 158.06
R7605 VDD.t3371 VDD.t3367 158.06
R7606 VDD.t3246 VDD.t3250 158.06
R7607 VDD.t3250 VDD.t123 158.06
R7608 VDD.t123 VDD.t127 158.06
R7609 VDD.t409 VDD.t411 158.06
R7610 VDD.t411 VDD.t2929 158.06
R7611 VDD.t2929 VDD.t3036 158.06
R7612 VDD.t4485 VDD.t4422 158.06
R7613 VDD.t129 VDD.t4485 158.06
R7614 VDD.t131 VDD.t129 158.06
R7615 VDD.t963 VDD.t962 158.06
R7616 VDD.t964 VDD.t963 158.06
R7617 VDD.t960 VDD.t964 158.06
R7618 VDD.t961 VDD.t960 158.06
R7619 VDD.t1477 VDD.t961 158.06
R7620 VDD.t1479 VDD.t1477 158.06
R7621 VDD.t1226 VDD.t1479 158.06
R7622 VDD.t1481 VDD.t1228 158.06
R7623 VDD.t686 VDD.t690 158.06
R7624 VDD.t687 VDD.t686 158.06
R7625 VDD.t688 VDD.t687 158.06
R7626 VDD.t689 VDD.t688 158.06
R7627 VDD.t4305 VDD.t689 158.06
R7628 VDD.t4297 VDD.t4305 158.06
R7629 VDD.t4301 VDD.t4297 158.06
R7630 VDD.t4299 VDD.t4303 158.06
R7631 VDD.t1107 VDD.t1105 158.06
R7632 VDD.t1105 VDD.t3028 158.06
R7633 VDD.t3028 VDD.t3016 158.06
R7634 VDD.t193 VDD.t191 158.06
R7635 VDD.t3127 VDD.t193 158.06
R7636 VDD.t3129 VDD.t3127 158.06
R7637 VDD.t607 VDD.t605 158.06
R7638 VDD.t203 VDD.t607 158.06
R7639 VDD.t205 VDD.t203 158.06
R7640 VDD.t187 VDD.t189 158.06
R7641 VDD.t189 VDD.t3131 158.06
R7642 VDD.t3131 VDD.t3135 158.06
R7643 VDD.t148 VDD.t2646 158.06
R7644 VDD.t2646 VDD.t2927 158.06
R7645 VDD.t2927 VDD.t3032 158.06
R7646 VDD.t4487 VDD.t4424 158.06
R7647 VDD.t3137 VDD.t4487 158.06
R7648 VDD.t3139 VDD.t3137 158.06
R7649 VDD.t3284 VDD.t3283 158.06
R7650 VDD.t3285 VDD.t3284 158.06
R7651 VDD.t3281 VDD.t3285 158.06
R7652 VDD.t3282 VDD.t3281 158.06
R7653 VDD.t4251 VDD.t3282 158.06
R7654 VDD.t4253 VDD.t4251 158.06
R7655 VDD.t4257 VDD.t4253 158.06
R7656 VDD.t4255 VDD.t4259 158.06
R7657 VDD.t2490 VDD.t2492 158.06
R7658 VDD.t2492 VDD.t2974 158.06
R7659 VDD.t2974 VDD.t2955 158.06
R7660 VDD.t2653 VDD.t2651 158.06
R7661 VDD.t1513 VDD.t2653 158.06
R7662 VDD.t1515 VDD.t1513 158.06
R7663 VDD.t1495 VDD.t1497 158.06
R7664 VDD.t3153 VDD.t1495 158.06
R7665 VDD.t3157 VDD.t3153 158.06
R7666 VDD.t2663 VDD.t2665 158.06
R7667 VDD.t2665 VDD.t1133 158.06
R7668 VDD.t1133 VDD.t1505 158.06
R7669 VDD.t3143 VDD.t3145 158.06
R7670 VDD.t3145 VDD.t3022 158.06
R7671 VDD.t3022 VDD.t2976 158.06
R7672 VDD.t4389 VDD.t4497 158.06
R7673 VDD.t1507 VDD.t4389 158.06
R7674 VDD.t1509 VDD.t1507 158.06
R7675 VDD.t1111 VDD.t1110 158.06
R7676 VDD.t1112 VDD.t1111 158.06
R7677 VDD.t1113 VDD.t1112 158.06
R7678 VDD.t1114 VDD.t1113 158.06
R7679 VDD.t742 VDD.t1114 158.06
R7680 VDD.t734 VDD.t742 158.06
R7681 VDD.t738 VDD.t734 158.06
R7682 VDD.t736 VDD.t740 158.06
R7683 VDD.t3338 VDD.t3340 158.06
R7684 VDD.t3340 VDD.t2953 158.06
R7685 VDD.t2953 VDD.t2941 158.06
R7686 VDD.t329 VDD.t327 158.06
R7687 VDD.t431 VDD.t329 158.06
R7688 VDD.t433 VDD.t431 158.06
R7689 VDD.t3298 VDD.t3306 158.06
R7690 VDD.t6 VDD.t3298 158.06
R7691 VDD.t8 VDD.t6 158.06
R7692 VDD.t331 VDD.t565 158.06
R7693 VDD.t565 VDD.t419 158.06
R7694 VDD.t419 VDD.t423 158.06
R7695 VDD.t1222 VDD.t1224 158.06
R7696 VDD.t1224 VDD.t3010 158.06
R7697 VDD.t3010 VDD.t2957 158.06
R7698 VDD.t4397 VDD.t4503 158.06
R7699 VDD.t425 VDD.t4397 158.06
R7700 VDD.t427 VDD.t425 158.06
R7701 VDD.t697 VDD.t696 158.06
R7702 VDD.t698 VDD.t697 158.06
R7703 VDD.t694 VDD.t698 158.06
R7704 VDD.t695 VDD.t694 158.06
R7705 VDD.t982 VDD.t695 158.06
R7706 VDD.t984 VDD.t982 158.06
R7707 VDD.t2905 VDD.t984 158.06
R7708 VDD.t2903 VDD.t2907 158.06
R7709 VDD.t98 VDD.t96 158.06
R7710 VDD.t96 VDD.t3044 158.06
R7711 VDD.t3044 VDD.t3055 158.06
R7712 VDD.t1419 VDD.t66 158.06
R7713 VDD.t1715 VDD.t1419 158.06
R7714 VDD.t1713 VDD.t1715 158.06
R7715 VDD.t3355 VDD.t3357 158.06
R7716 VDD.t1261 VDD.t3355 158.06
R7717 VDD.t1273 VDD.t1261 158.06
R7718 VDD.t72 VDD.t68 158.06
R7719 VDD.t68 VDD.t1711 158.06
R7720 VDD.t1711 VDD.t1705 158.06
R7721 VDD.t880 VDD.t882 158.06
R7722 VDD.t882 VDD.t2972 158.06
R7723 VDD.t2972 VDD.t3012 158.06
R7724 VDD.t4512 VDD.t4411 158.06
R7725 VDD.t1719 VDD.t4512 158.06
R7726 VDD.t1717 VDD.t1719 158.06
R7727 VDD.t1321 VDD.t1322 158.06
R7728 VDD.t1320 VDD.t1321 158.06
R7729 VDD.t1319 VDD.t1320 158.06
R7730 VDD.t1318 VDD.t1319 158.06
R7731 VDD.t4314 VDD.t1318 158.06
R7732 VDD.t4322 VDD.t4314 158.06
R7733 VDD.t4320 VDD.t4322 158.06
R7734 VDD.t4318 VDD.t4316 158.06
R7735 VDD.t1944 VDD.t1918 158.06
R7736 VDD.t1918 VDD.t3072 158.06
R7737 VDD.t3072 VDD.t3038 158.06
R7738 VDD.t648 VDD.t644 158.06
R7739 VDD.t2889 VDD.t648 158.06
R7740 VDD.t2891 VDD.t2889 158.06
R7741 VDD.t1578 VDD.t1580 158.06
R7742 VDD.t852 VDD.t1578 158.06
R7743 VDD.t854 VDD.t852 158.06
R7744 VDD.t640 VDD.t642 158.06
R7745 VDD.t642 VDD.t2893 158.06
R7746 VDD.t2893 VDD.t2899 158.06
R7747 VDD.t1920 VDD.t1976 158.06
R7748 VDD.t1976 VDD.t3042 158.06
R7749 VDD.t3042 VDD.t2968 158.06
R7750 VDD.t4441 VDD.t4339 158.06
R7751 VDD.t2895 VDD.t4441 158.06
R7752 VDD.t2901 VDD.t2895 158.06
R7753 VDD.t3126 VDD.t3124 158.06
R7754 VDD.t3122 VDD.t3126 158.06
R7755 VDD.t3123 VDD.t3122 158.06
R7756 VDD.t3125 VDD.t3123 158.06
R7757 VDD.t3502 VDD.t3125 158.06
R7758 VDD.t3506 VDD.t3502 158.06
R7759 VDD.t3508 VDD.t3506 158.06
R7760 VDD.t3510 VDD.t3504 158.06
R7761 VDD.n670 VDD.t2422 148.181
R7762 VDD.n685 VDD.t2732 148.181
R7763 VDD.n1144 VDD.n1142 147.517
R7764 VDD.n1885 VDD.t826 145.268
R7765 VDD.n147 VDD.t1094 144.121
R7766 VDD.n670 VDD.n669 140.65
R7767 VDD.n685 VDD.n668 140.587
R7768 VDD.n2218 VDD.t3560 129.654
R7769 VDD.n2243 VDD.t317 129.654
R7770 VDD.n1884 VDD.t1569 129.654
R7771 VDD.n1885 VDD.t1356 117.8
R7772 VDD.t2273 VDD.n1134 116.552
R7773 VDD.t2819 VDD.n1919 116.552
R7774 VDD.n1909 VDD.t3434 116.552
R7775 VDD.t393 VDD.n1926 116.552
R7776 VDD.n1927 VDD.t2197 116.552
R7777 VDD.t4070 VDD.n1938 116.552
R7778 VDD.t531 VDD.n1945 116.552
R7779 VDD.n1946 VDD.t4208 116.552
R7780 VDD.n1899 VDD.t1661 116.552
R7781 VDD.n683 VDD.t2391 116.552
R7782 VDD.t1094 VDD.t1090 115.297
R7783 VDD.t1090 VDD.t1092 115.297
R7784 VDD.n2835 VDD.n2834 114.007
R7785 VDD.n2844 VDD.n2843 114.007
R7786 VDD.n2850 VDD.n2849 114.007
R7787 VDD.n2746 VDD.n2744 114.007
R7788 VDD.n2757 VDD.n2755 114.007
R7789 VDD.n2768 VDD.n2766 114.007
R7790 VDD.n2779 VDD.n2777 114.007
R7791 VDD.n2790 VDD.n2788 114.007
R7792 VDD.n2801 VDD.n2799 114.007
R7793 VDD.n2812 VDD.n2810 114.007
R7794 VDD.n2823 VDD.n2821 114.007
R7795 VDD.n2740 VDD.n2739 114.007
R7796 VDD.n2734 VDD.n2733 114.007
R7797 VDD.n2724 VDD.n2723 114.007
R7798 VDD.n1989 VDD.n1987 114.007
R7799 VDD.n2008 VDD.n2006 114.007
R7800 VDD.n2015 VDD.n2013 114.007
R7801 VDD.n1979 VDD.n1977 114.007
R7802 VDD.n2028 VDD.n2026 114.007
R7803 VDD.n2035 VDD.n2033 114.007
R7804 VDD.n1995 VDD.n1993 114.007
R7805 VDD.n1971 VDD.n1969 114.007
R7806 VDD.n2352 VDD.n2351 114.007
R7807 VDD.n2361 VDD.n2360 114.007
R7808 VDD.n1178 VDD.n1177 114.007
R7809 VDD.n1359 VDD.n1358 114.007
R7810 VDD.n1790 VDD.n1789 114.007
R7811 VDD.n1375 VDD.n1374 114.007
R7812 VDD.n1381 VDD.n1380 114.007
R7813 VDD.n1798 VDD.n1797 114.007
R7814 VDD.n1444 VDD.n1443 114.007
R7815 VDD.n1437 VDD.n1436 114.007
R7816 VDD.n1630 VDD.n1629 114.007
R7817 VDD.n1639 VDD.n1638 114.007
R7818 VDD.n1647 VDD.n1646 114.007
R7819 VDD.n1657 VDD.n1656 114.007
R7820 VDD.n1666 VDD.n1665 114.007
R7821 VDD.n1672 VDD.n1671 114.007
R7822 VDD.n1607 VDD.n1606 114.007
R7823 VDD.n1616 VDD.n1615 114.007
R7824 VDD.n1459 VDD.n1458 114.007
R7825 VDD.n1598 VDD.n1597 114.007
R7826 VDD.n1588 VDD.n1587 114.007
R7827 VDD.n1580 VDD.n1579 114.007
R7828 VDD.n1571 VDD.n1570 114.007
R7829 VDD.n1465 VDD.n1464 114.007
R7830 VDD.n2716 VDD.n2715 114.007
R7831 VDD.n2657 VDD.n2656 114.007
R7832 VDD.n2427 VDD.n2426 114.007
R7833 VDD.n2648 VDD.n2647 114.007
R7834 VDD.n2640 VDD.n2639 114.007
R7835 VDD.n2593 VDD.n2592 114.007
R7836 VDD.n2447 VDD.n2446 114.007
R7837 VDD.n2584 VDD.n2583 114.007
R7838 VDD.n2576 VDD.n2575 114.007
R7839 VDD.n2505 VDD.n2504 114.007
R7840 VDD.n2514 VDD.n2513 114.007
R7841 VDD.n2489 VDD.n2488 114.007
R7842 VDD.n2495 VDD.n2494 114.007
R7843 VDD.n2835 VDD.n2833 113.974
R7844 VDD.n2844 VDD.n2842 113.974
R7845 VDD.n2850 VDD.n2848 113.974
R7846 VDD.n2746 VDD.n2745 113.974
R7847 VDD.n2757 VDD.n2756 113.974
R7848 VDD.n2768 VDD.n2767 113.974
R7849 VDD.n2779 VDD.n2778 113.974
R7850 VDD.n2790 VDD.n2789 113.974
R7851 VDD.n2801 VDD.n2800 113.974
R7852 VDD.n2812 VDD.n2811 113.974
R7853 VDD.n2823 VDD.n2822 113.974
R7854 VDD.n2740 VDD.n2738 113.974
R7855 VDD.n2734 VDD.n2732 113.974
R7856 VDD.n2724 VDD.n2722 113.974
R7857 VDD.n1989 VDD.n1988 113.974
R7858 VDD.n2008 VDD.n2007 113.974
R7859 VDD.n2015 VDD.n2014 113.974
R7860 VDD.n1979 VDD.n1978 113.974
R7861 VDD.n2028 VDD.n2027 113.974
R7862 VDD.n2035 VDD.n2034 113.974
R7863 VDD.n1995 VDD.n1994 113.974
R7864 VDD.n1971 VDD.n1970 113.974
R7865 VDD.n2352 VDD.n2350 113.974
R7866 VDD.n2361 VDD.n2359 113.974
R7867 VDD.n1178 VDD.n1176 113.974
R7868 VDD.n1359 VDD.n1357 113.974
R7869 VDD.n1790 VDD.n1788 113.974
R7870 VDD.n1375 VDD.n1373 113.974
R7871 VDD.n1381 VDD.n1379 113.974
R7872 VDD.n1798 VDD.n1796 113.974
R7873 VDD.n1444 VDD.n1442 113.974
R7874 VDD.n1437 VDD.n1435 113.974
R7875 VDD.n1630 VDD.n1628 113.974
R7876 VDD.n1639 VDD.n1637 113.974
R7877 VDD.n1647 VDD.n1645 113.974
R7878 VDD.n1657 VDD.n1655 113.974
R7879 VDD.n1666 VDD.n1664 113.974
R7880 VDD.n1672 VDD.n1670 113.974
R7881 VDD.n1607 VDD.n1605 113.974
R7882 VDD.n1616 VDD.n1614 113.974
R7883 VDD.n1459 VDD.n1457 113.974
R7884 VDD.n1598 VDD.n1596 113.974
R7885 VDD.n1588 VDD.n1586 113.974
R7886 VDD.n1580 VDD.n1578 113.974
R7887 VDD.n1571 VDD.n1569 113.974
R7888 VDD.n1465 VDD.n1463 113.974
R7889 VDD.n2716 VDD.n2714 113.974
R7890 VDD.n2657 VDD.n2655 113.974
R7891 VDD.n2427 VDD.n2425 113.974
R7892 VDD.n2648 VDD.n2646 113.974
R7893 VDD.n2640 VDD.n2638 113.974
R7894 VDD.n2593 VDD.n2591 113.974
R7895 VDD.n2447 VDD.n2445 113.974
R7896 VDD.n2584 VDD.n2582 113.974
R7897 VDD.n2576 VDD.n2574 113.974
R7898 VDD.n2505 VDD.n2503 113.974
R7899 VDD.n2514 VDD.n2512 113.974
R7900 VDD.n2489 VDD.n2487 113.974
R7901 VDD.n2495 VDD.n2493 113.974
R7902 VDD.n1148 VDD.n1146 112.796
R7903 VDD.n2840 VDD.n2838 112.796
R7904 VDD.n2750 VDD.n2749 112.796
R7905 VDD.n2761 VDD.n2760 112.796
R7906 VDD.n2772 VDD.n2771 112.796
R7907 VDD.n2783 VDD.n2782 112.796
R7908 VDD.n2794 VDD.n2793 112.796
R7909 VDD.n2805 VDD.n2804 112.796
R7910 VDD.n2816 VDD.n2815 112.796
R7911 VDD.n2827 VDD.n2826 112.796
R7912 VDD.n1159 VDD.n1157 112.796
R7913 VDD.n2730 VDD.n2728 112.796
R7914 VDD.n2721 VDD.n2719 112.796
R7915 VDD.n1181 VDD.n1179 112.796
R7916 VDD.n2357 VDD.n2355 112.796
R7917 VDD.n1175 VDD.n1173 112.796
R7918 VDD.n1356 VDD.n1354 112.796
R7919 VDD.n1362 VDD.n1360 112.796
R7920 VDD.n1372 VDD.n1370 112.796
R7921 VDD.n1378 VDD.n1376 112.796
R7922 VDD.n1795 VDD.n1793 112.796
R7923 VDD.n1440 VDD.n1438 112.796
R7924 VDD.n1434 VDD.n1432 112.796
R7925 VDD.n1430 VDD.n1428 112.796
R7926 VDD.n1635 VDD.n1633 112.796
R7927 VDD.n1644 VDD.n1642 112.796
R7928 VDD.n1653 VDD.n1651 112.796
R7929 VDD.n1662 VDD.n1660 112.796
R7930 VDD.n1427 VDD.n1425 112.796
R7931 VDD.n1603 VDD.n1601 112.796
R7932 VDD.n1612 VDD.n1610 112.796
R7933 VDD.n1456 VDD.n1454 112.796
R7934 VDD.n1594 VDD.n1592 112.796
R7935 VDD.n1585 VDD.n1583 112.796
R7936 VDD.n1576 VDD.n1574 112.796
R7937 VDD.n1567 VDD.n1565 112.796
R7938 VDD.n1462 VDD.n1460 112.796
R7939 VDD.n1162 VDD.n1160 112.796
R7940 VDD.n2654 VDD.n2652 112.796
R7941 VDD.n2424 VDD.n2422 112.796
R7942 VDD.n2645 VDD.n2643 112.796
R7943 VDD.n2430 VDD.n2428 112.796
R7944 VDD.n2590 VDD.n2588 112.796
R7945 VDD.n2444 VDD.n2442 112.796
R7946 VDD.n2581 VDD.n2579 112.796
R7947 VDD.n2450 VDD.n2448 112.796
R7948 VDD.n2501 VDD.n2499 112.796
R7949 VDD.n2510 VDD.n2508 112.796
R7950 VDD.n2486 VDD.n2484 112.796
R7951 VDD.n2492 VDD.n2490 112.796
R7952 VDD.n1148 VDD.n1147 112.763
R7953 VDD.n2840 VDD.n2839 112.763
R7954 VDD.n2750 VDD.n2748 112.763
R7955 VDD.n2761 VDD.n2759 112.763
R7956 VDD.n2772 VDD.n2770 112.763
R7957 VDD.n2783 VDD.n2781 112.763
R7958 VDD.n2794 VDD.n2792 112.763
R7959 VDD.n2805 VDD.n2803 112.763
R7960 VDD.n2816 VDD.n2814 112.763
R7961 VDD.n2827 VDD.n2825 112.763
R7962 VDD.n1159 VDD.n1158 112.763
R7963 VDD.n2730 VDD.n2729 112.763
R7964 VDD.n2721 VDD.n2720 112.763
R7965 VDD.n1181 VDD.n1180 112.763
R7966 VDD.n2357 VDD.n2356 112.763
R7967 VDD.n1175 VDD.n1174 112.763
R7968 VDD.n1356 VDD.n1355 112.763
R7969 VDD.n1362 VDD.n1361 112.763
R7970 VDD.n1372 VDD.n1371 112.763
R7971 VDD.n1378 VDD.n1377 112.763
R7972 VDD.n1795 VDD.n1794 112.763
R7973 VDD.n1440 VDD.n1439 112.763
R7974 VDD.n1434 VDD.n1433 112.763
R7975 VDD.n1430 VDD.n1429 112.763
R7976 VDD.n1635 VDD.n1634 112.763
R7977 VDD.n1644 VDD.n1643 112.763
R7978 VDD.n1653 VDD.n1652 112.763
R7979 VDD.n1662 VDD.n1661 112.763
R7980 VDD.n1427 VDD.n1426 112.763
R7981 VDD.n1603 VDD.n1602 112.763
R7982 VDD.n1612 VDD.n1611 112.763
R7983 VDD.n1456 VDD.n1455 112.763
R7984 VDD.n1594 VDD.n1593 112.763
R7985 VDD.n1585 VDD.n1584 112.763
R7986 VDD.n1576 VDD.n1575 112.763
R7987 VDD.n1567 VDD.n1566 112.763
R7988 VDD.n1462 VDD.n1461 112.763
R7989 VDD.n1162 VDD.n1161 112.763
R7990 VDD.n2654 VDD.n2653 112.763
R7991 VDD.n2424 VDD.n2423 112.763
R7992 VDD.n2645 VDD.n2644 112.763
R7993 VDD.n2430 VDD.n2429 112.763
R7994 VDD.n2590 VDD.n2589 112.763
R7995 VDD.n2444 VDD.n2443 112.763
R7996 VDD.n2581 VDD.n2580 112.763
R7997 VDD.n2450 VDD.n2449 112.763
R7998 VDD.n2501 VDD.n2500 112.763
R7999 VDD.n2510 VDD.n2509 112.763
R8000 VDD.n2486 VDD.n2485 112.763
R8001 VDD.n2492 VDD.n2491 112.763
R8002 VDD.n1986 VDD.n1985 112.688
R8003 VDD.n2005 VDD.n2004 112.688
R8004 VDD.n1983 VDD.n1982 112.688
R8005 VDD.n1976 VDD.n1975 112.688
R8006 VDD.n2025 VDD.n2024 112.688
R8007 VDD.n1965 VDD.n1964 112.688
R8008 VDD.n1992 VDD.n1991 112.688
R8009 VDD.n1968 VDD.n1967 112.688
R8010 VDD.n1986 VDD.n1984 112.653
R8011 VDD.n2005 VDD.n2003 112.653
R8012 VDD.n1983 VDD.n1981 112.653
R8013 VDD.n1976 VDD.n1974 112.653
R8014 VDD.n2025 VDD.n2023 112.653
R8015 VDD.n1965 VDD.n1963 112.653
R8016 VDD.n1992 VDD.n1990 112.653
R8017 VDD.n1968 VDD.n1966 112.653
R8018 VDD.n1117 VDD.t630 109.043
R8019 VDD.n1026 VDD.t3216 109.043
R8020 VDD.n1050 VDD.t2107 109.043
R8021 VDD.n988 VDD.t2848 109.043
R8022 VDD.n897 VDD.t2531 109.043
R8023 VDD.n921 VDD.t3117 109.043
R8024 VDD.n859 VDD.t1220 109.043
R8025 VDD.n768 VDD.t3363 109.043
R8026 VDD.n792 VDD.t820 109.043
R8027 VDD.n730 VDD.t228 109.043
R8028 VDD.n641 VDD.t1423 109.043
R8029 VDD.t3067 VDD.n640 109.043
R8030 VDD.n629 VDD.t1990 109.043
R8031 VDD.t3087 VDD.n628 109.043
R8032 VDD.n617 VDD.t1721 109.043
R8033 VDD.n579 VDD.t4245 109.043
R8034 VDD.n488 VDD.t197 109.043
R8035 VDD.n512 VDD.t4261 109.043
R8036 VDD.n450 VDD.t2098 109.043
R8037 VDD.n359 VDD.t3161 109.043
R8038 VDD.n383 VDD.t1162 109.043
R8039 VDD.n321 VDD.t353 109.043
R8040 VDD.n192 VDD.t273 109.043
R8041 VDD.n230 VDD.t2453 109.043
R8042 VDD.n254 VDD.t2767 109.043
R8043 VDD.n92 VDD.t1265 109.043
R8044 VDD.n116 VDD.t925 109.043
R8045 VDD.n2897 VDD.t2068 109.043
R8046 VDD.n30 VDD.t858 109.043
R8047 VDD.n54 VDD.t1741 109.043
R8048 VDD.t2939 VDD.n1116 108.855
R8049 VDD.n1105 VDD.t1259 108.855
R8050 VDD.t3008 VDD.n1104 108.855
R8051 VDD.n1093 VDD.t1267 108.855
R8052 VDD.t2984 VDD.n987 108.855
R8053 VDD.n976 VDD.t3226 108.855
R8054 VDD.t3051 VDD.n975 108.855
R8055 VDD.n964 VDD.t3218 108.855
R8056 VDD.t3040 VDD.n858 108.855
R8057 VDD.n847 VDD.t2527 108.855
R8058 VDD.t2935 VDD.n846 108.855
R8059 VDD.n835 VDD.t2535 108.855
R8060 VDD.t3080 VDD.n729 108.855
R8061 VDD.n718 VDD.t3373 108.855
R8062 VDD.t3030 VDD.n717 108.855
R8063 VDD.n706 VDD.t3365 108.855
R8064 VDD.t3074 VDD.n578 108.855
R8065 VDD.n567 VDD.t1996 108.855
R8066 VDD.t3024 VDD.n566 108.855
R8067 VDD.n555 VDD.t1986 108.855
R8068 VDD.t2947 VDD.n449 108.855
R8069 VDD.n438 VDD.t201 108.855
R8070 VDD.t3065 VDD.n437 108.855
R8071 VDD.n426 VDD.t2048 108.855
R8072 VDD.t3069 VDD.n320 108.855
R8073 VDD.n309 VDD.t3165 108.855
R8074 VDD.t3020 VDD.n308 108.855
R8075 VDD.n297 VDD.t3155 108.855
R8076 VDD.t2992 VDD.n191 108.855
R8077 VDD.n180 VDD.t2451 108.855
R8078 VDD.t3062 VDD.n179 108.855
R8079 VDD.n168 VDD.t4 108.855
R8080 VDD.t3076 VDD.n2896 108.855
R8081 VDD.n2885 VDD.t850 108.855
R8082 VDD.t2931 VDD.n2884 108.855
R8083 VDD.n2873 VDD.t846 108.855
R8084 VDD.t3101 VDD.n1049 108.666
R8085 VDD.n1038 VDD.t3224 108.666
R8086 VDD.t3057 VDD.n1037 108.666
R8087 VDD.t2945 VDD.n920 108.666
R8088 VDD.n909 VDD.t2523 108.666
R8089 VDD.t2963 VDD.n908 108.666
R8090 VDD.t3018 VDD.n791 108.666
R8091 VDD.n780 VDD.t3371 108.666
R8092 VDD.t3036 VDD.n779 108.666
R8093 VDD.t3016 VDD.n511 108.666
R8094 VDD.n500 VDD.t205 108.666
R8095 VDD.t3032 VDD.n499 108.666
R8096 VDD.t2955 VDD.n382 108.666
R8097 VDD.n371 VDD.t3157 108.666
R8098 VDD.t2976 VDD.n370 108.666
R8099 VDD.t2941 VDD.n253 108.666
R8100 VDD.n242 VDD.t8 108.666
R8101 VDD.t2957 VDD.n241 108.666
R8102 VDD.t3055 VDD.n115 108.666
R8103 VDD.n104 VDD.t1273 108.666
R8104 VDD.t3012 VDD.n103 108.666
R8105 VDD.t3038 VDD.n53 108.666
R8106 VDD.n42 VDD.t854 108.666
R8107 VDD.t2968 VDD.n41 108.666
R8108 VDD.t4190 VDD.n1261 103.602
R8109 VDD.t4113 VDD.n1273 103.602
R8110 VDD.n1955 VDD.n1952 102.978
R8111 VDD.n2331 VDD.n2328 102.978
R8112 VDD.n2321 VDD.n2318 102.978
R8113 VDD.n2311 VDD.n2308 102.978
R8114 VDD.n2300 VDD.n2297 102.978
R8115 VDD.n2290 VDD.n2287 102.978
R8116 VDD.n2280 VDD.n2277 102.978
R8117 VDD.n2270 VDD.n2267 102.978
R8118 VDD.n1066 VDD.n1060 102.978
R8119 VDD.n937 VDD.n931 102.978
R8120 VDD.n808 VDD.n802 102.978
R8121 VDD.n657 VDD.n651 102.978
R8122 VDD.n528 VDD.n522 102.978
R8123 VDD.n399 VDD.n393 102.978
R8124 VDD.n270 VDD.n264 102.978
R8125 VDD.n132 VDD.n126 102.978
R8126 VDD.n2916 VDD.n2910 102.978
R8127 VDD.n1960 VDD.n1959 102.266
R8128 VDD.n2336 VDD.n2335 102.266
R8129 VDD.n2326 VDD.n2325 102.266
R8130 VDD.n2316 VDD.n2315 102.266
R8131 VDD.n2305 VDD.n2304 102.266
R8132 VDD.n2295 VDD.n2294 102.266
R8133 VDD.n2285 VDD.n2284 102.266
R8134 VDD.n2275 VDD.n2274 102.266
R8135 VDD.n1071 VDD.n1070 102.266
R8136 VDD.n942 VDD.n941 102.266
R8137 VDD.n813 VDD.n812 102.266
R8138 VDD.n662 VDD.n661 102.266
R8139 VDD.n533 VDD.n532 102.266
R8140 VDD.n404 VDD.n403 102.266
R8141 VDD.n275 VDD.n274 102.266
R8142 VDD.n137 VDD.n136 102.266
R8143 VDD.n2921 VDD.n2920 102.266
R8144 VDD.t1404 VDD.t1408 101.334
R8145 VDD.t1386 VDD.t1404 101.334
R8146 VDD.t2413 VDD.t1386 101.334
R8147 VDD.t2412 VDD.t2413 101.334
R8148 VDD.t2411 VDD.t2412 101.334
R8149 VDD.t3697 VDD.t3699 101.334
R8150 VDD.t3699 VDD.t3698 101.334
R8151 VDD.t3698 VDD.t1745 101.334
R8152 VDD.t1745 VDD.t1811 101.334
R8153 VDD.t1811 VDD.t1771 101.334
R8154 VDD.t3533 VDD.t3554 101.334
R8155 VDD.t3564 VDD.t3533 101.334
R8156 VDD.t2689 VDD.t3564 101.334
R8157 VDD.t2688 VDD.t2689 101.334
R8158 VDD.t2687 VDD.t2688 101.334
R8159 VDD.t4278 VDD.t4277 101.334
R8160 VDD.t4277 VDD.t4276 101.334
R8161 VDD.t4276 VDD.t766 101.334
R8162 VDD.t766 VDD.t1807 101.334
R8163 VDD.t1807 VDD.t1765 101.334
R8164 VDD.t891 VDD.t3966 101.334
R8165 VDD.t3981 VDD.t891 101.334
R8166 VDD.t2855 VDD.t3981 101.334
R8167 VDD.t2886 VDD.t2855 101.334
R8168 VDD.t2856 VDD.t2886 101.334
R8169 VDD.t1142 VDD.t1143 101.334
R8170 VDD.t1143 VDD.t2854 101.334
R8171 VDD.t2854 VDD.t1809 101.334
R8172 VDD.t1809 VDD.t1797 101.334
R8173 VDD.t1797 VDD.t1773 101.334
R8174 VDD.t3582 VDD.t3602 101.334
R8175 VDD.t3615 VDD.t3582 101.334
R8176 VDD.t2730 VDD.t3615 101.334
R8177 VDD.t2731 VDD.t2730 101.334
R8178 VDD.t2729 VDD.t2731 101.334
R8179 VDD.t1613 VDD.t1531 101.334
R8180 VDD.t1531 VDD.t1614 101.334
R8181 VDD.t1614 VDD.t1785 101.334
R8182 VDD.t1785 VDD.t1795 101.334
R8183 VDD.t1795 VDD.t1747 101.334
R8184 VDD.t2119 VDD.t2130 101.334
R8185 VDD.t2168 VDD.t2119 101.334
R8186 VDD.t684 VDD.t2168 101.334
R8187 VDD.t683 VDD.t684 101.334
R8188 VDD.t685 VDD.t683 101.334
R8189 VDD.t1447 VDD.t1446 101.334
R8190 VDD.t1446 VDD.t3381 101.334
R8191 VDD.t3381 VDD.t1779 101.334
R8192 VDD.t1779 VDD.t779 101.334
R8193 VDD.t779 VDD.t1805 101.334
R8194 VDD.t2594 VDD.t2603 101.334
R8195 VDD.t2579 VDD.t2594 101.334
R8196 VDD.t3986 VDD.t2579 101.334
R8197 VDD.t3985 VDD.t3986 101.334
R8198 VDD.t3987 VDD.t3985 101.334
R8199 VDD.t3958 VDD.t3960 101.334
R8200 VDD.t3960 VDD.t3959 101.334
R8201 VDD.t3959 VDD.t1755 101.334
R8202 VDD.t1755 VDD.t1803 101.334
R8203 VDD.t1803 VDD.t1783 101.334
R8204 VDD.t2341 VDD.t2353 101.334
R8205 VDD.t2324 VDD.t2341 101.334
R8206 VDD.t1199 VDD.t2324 101.334
R8207 VDD.t1198 VDD.t1199 101.334
R8208 VDD.t1200 VDD.t1198 101.334
R8209 VDD.t3953 VDD.t3952 101.334
R8210 VDD.t3952 VDD.t4185 101.334
R8211 VDD.t4185 VDD.t1749 101.334
R8212 VDD.t1749 VDD.t1799 101.334
R8213 VDD.t1799 VDD.t1777 101.334
R8214 VDD.t993 VDD.t1004 101.334
R8215 VDD.t1032 VDD.t993 101.334
R8216 VDD.t2081 VDD.t1032 101.334
R8217 VDD.t1645 VDD.t2081 101.334
R8218 VDD.t1644 VDD.t1645 101.334
R8219 VDD.t920 VDD.t919 101.334
R8220 VDD.t919 VDD.t918 101.334
R8221 VDD.t918 VDD.t764 101.334
R8222 VDD.t764 VDD.t1791 101.334
R8223 VDD.t1791 VDD.t1763 101.334
R8224 VDD.t2290 VDD.t3442 101.334
R8225 VDD.t2296 VDD.t2290 101.334
R8226 VDD.t1594 VDD.t2296 101.334
R8227 VDD.t1595 VDD.t1594 101.334
R8228 VDD.t1596 VDD.t1595 101.334
R8229 VDD.t971 VDD.t972 101.334
R8230 VDD.t972 VDD.t973 101.334
R8231 VDD.t973 VDD.t1412 101.334
R8232 VDD.t1412 VDD.t1176 101.334
R8233 VDD.t1176 VDD.t1396 101.334
R8234 VDD.t1659 VDD.t1657 101.334
R8235 VDD.t1679 VDD.t1659 101.334
R8236 VDD.t1149 VDD.t1679 101.334
R8237 VDD.t1150 VDD.t1149 101.334
R8238 VDD.t1148 VDD.t1150 101.334
R8239 VDD.t3692 VDD.t3690 101.334
R8240 VDD.t3687 VDD.t3692 101.334
R8241 VDD.t1037 VDD.t3687 101.334
R8242 VDD.t591 VDD.t1037 101.334
R8243 VDD.t987 VDD.t591 101.334
R8244 VDD.t980 VDD.t974 101.222
R8245 VDD.t974 VDD.t976 101.222
R8246 VDD.t976 VDD.t489 101.222
R8247 VDD.t489 VDD.t487 101.222
R8248 VDD.t487 VDD.t488 101.222
R8249 VDD.t1097 VDD.t1098 101.222
R8250 VDD.t1098 VDD.t1096 101.222
R8251 VDD.t1096 VDD.t1759 101.222
R8252 VDD.t1759 VDD.t1787 101.222
R8253 VDD.t1787 VDD.t783 101.222
R8254 VDD.t1406 VDD.t1410 101.222
R8255 VDD.t1410 VDD.t1384 101.222
R8256 VDD.t1384 VDD.t2769 101.222
R8257 VDD.t2769 VDD.t2770 101.222
R8258 VDD.t2770 VDD.t2771 101.222
R8259 VDD.t1474 VDD.t1846 101.222
R8260 VDD.t1846 VDD.t278 101.222
R8261 VDD.t278 VDD.t2292 101.222
R8262 VDD.t2292 VDD.t3417 101.222
R8263 VDD.t3417 VDD.t3425 101.222
R8264 VDD.t3308 VDD.t3304 101.222
R8265 VDD.t3302 VDD.t3308 101.222
R8266 VDD.t56 VDD.t3302 101.222
R8267 VDD.t4123 VDD.t56 101.222
R8268 VDD.t55 VDD.t4123 101.222
R8269 VDD.t2106 VDD.t1906 101.222
R8270 VDD.t1906 VDD.t1907 101.222
R8271 VDD.t1907 VDD.t2294 101.222
R8272 VDD.t2294 VDD.t3438 101.222
R8273 VDD.t3438 VDD.t3447 101.222
R8274 VDD.t2825 VDD.t2812 101.109
R8275 VDD.t2812 VDD.t2814 101.109
R8276 VDD.t2814 VDD.t2639 101.109
R8277 VDD.t2639 VDD.t2640 101.109
R8278 VDD.t2640 VDD.t2641 101.109
R8279 VDD.t1829 VDD.t1828 101.109
R8280 VDD.t1830 VDD.t1829 101.109
R8281 VDD.t3562 VDD.t1830 101.109
R8282 VDD.t3537 VDD.t3562 101.109
R8283 VDD.t3548 VDD.t3537 101.109
R8284 VDD.t401 VDD.t383 101.109
R8285 VDD.t383 VDD.t385 101.109
R8286 VDD.t385 VDD.t1817 101.109
R8287 VDD.t1817 VDD.t1818 101.109
R8288 VDD.t1818 VDD.t1819 101.109
R8289 VDD.t3291 VDD.t1459 101.109
R8290 VDD.t1459 VDD.t1835 101.109
R8291 VDD.t1835 VDD.t3979 101.109
R8292 VDD.t3979 VDD.t893 101.109
R8293 VDD.t893 VDD.t3968 101.109
R8294 VDD.t2195 VDD.t2193 101.109
R8295 VDD.t1631 VDD.t2195 101.109
R8296 VDD.t627 VDD.t1631 101.109
R8297 VDD.t628 VDD.t627 101.109
R8298 VDD.t629 VDD.t628 101.109
R8299 VDD.t4166 VDD.t4165 101.109
R8300 VDD.t4165 VDD.t3526 101.109
R8301 VDD.t3526 VDD.t3604 101.109
R8302 VDD.t3604 VDD.t3618 101.109
R8303 VDD.t3618 VDD.t3584 101.109
R8304 VDD.t4119 VDD.t4077 101.109
R8305 VDD.t4077 VDD.t4089 101.109
R8306 VDD.t4089 VDD.t2763 101.109
R8307 VDD.t2763 VDD.t2764 101.109
R8308 VDD.t2764 VDD.t2762 101.109
R8309 VDD.t42 VDD.t3452 101.109
R8310 VDD.t3490 VDD.t42 101.109
R8311 VDD.t2132 VDD.t3490 101.109
R8312 VDD.t2151 VDD.t2132 101.109
R8313 VDD.t2180 VDD.t2151 101.109
R8314 VDD.t525 VDD.t537 101.109
R8315 VDD.t537 VDD.t539 101.109
R8316 VDD.t539 VDD.t2414 101.109
R8317 VDD.t2414 VDD.t2415 101.109
R8318 VDD.t2415 VDD.t2416 101.109
R8319 VDD.t1236 VDD.t1237 101.109
R8320 VDD.t1237 VDD.t2871 101.109
R8321 VDD.t2871 VDD.t2588 101.109
R8322 VDD.t2588 VDD.t2609 101.109
R8323 VDD.t2609 VDD.t483 101.109
R8324 VDD.t4196 VDD.t4230 101.109
R8325 VDD.t4214 VDD.t4196 101.109
R8326 VDD.t1303 VDD.t4214 101.109
R8327 VDD.t1304 VDD.t1303 101.109
R8328 VDD.t1305 VDD.t1304 101.109
R8329 VDD.t2457 VDD.t2458 101.109
R8330 VDD.t2458 VDD.t2459 101.109
R8331 VDD.t2459 VDD.t1831 101.109
R8332 VDD.t1831 VDD.t2316 101.109
R8333 VDD.t2316 VDD.t2345 101.109
R8334 VDD.n2218 VDD.t1393 100.838
R8335 VDD.n2243 VDD.t787 100.838
R8336 VDD.n1884 VDD.t3486 100.838
R8337 VDD.t1974 VDD.t1982 100.111
R8338 VDD.t1962 VDD.t1974 100.111
R8339 VDD.t309 VDD.t1962 100.111
R8340 VDD.t310 VDD.t309 100.111
R8341 VDD.t308 VDD.t310 100.111
R8342 VDD.t368 VDD.t367 100.111
R8343 VDD.t1539 VDD.t368 100.111
R8344 VDD.t2058 VDD.t1539 100.111
R8345 VDD.t2060 VDD.t2058 100.111
R8346 VDD.t1601 VDD.t2060 100.111
R8347 VDD.t1301 VDD.t1297 100.111
R8348 VDD.t1291 VDD.t1301 100.111
R8349 VDD.t306 VDD.t1291 100.111
R8350 VDD.t307 VDD.t306 100.111
R8351 VDD.t305 VDD.t307 100.111
R8352 VDD.t2650 VDD.t2862 100.111
R8353 VDD.t2862 VDD.t2863 100.111
R8354 VDD.t2863 VDD.t289 100.111
R8355 VDD.t289 VDD.t285 100.111
R8356 VDD.t285 VDD.t287 100.111
R8357 VDD.t2417 VDD.t211 100.111
R8358 VDD.t211 VDD.t213 100.111
R8359 VDD.t213 VDD.t3286 100.111
R8360 VDD.t3286 VDD.t3287 100.111
R8361 VDD.t3287 VDD.t3342 100.111
R8362 VDD.t1151 VDD.t1152 100.111
R8363 VDD.t986 VDD.t1151 100.111
R8364 VDD.t4177 VDD.t986 100.111
R8365 VDD.t4183 VDD.t4177 100.111
R8366 VDD.t4171 VDD.t4183 100.111
R8367 VDD.t2308 VDD.t2310 100.111
R8368 VDD.t2312 VDD.t2308 100.111
R8369 VDD.t1525 VDD.t2312 100.111
R8370 VDD.t1526 VDD.t1525 100.111
R8371 VDD.t1527 VDD.t1526 100.111
R8372 VDD.t4163 VDD.t4164 100.111
R8373 VDD.t4164 VDD.t4162 100.111
R8374 VDD.t4162 VDD.t1332 100.111
R8375 VDD.t1332 VDD.t1340 100.111
R8376 VDD.t1340 VDD.t1338 100.111
R8377 VDD.t704 VDD.t708 100.111
R8378 VDD.t708 VDD.t710 100.111
R8379 VDD.t710 VDD.t928 100.111
R8380 VDD.t928 VDD.t927 100.111
R8381 VDD.t927 VDD.t929 100.111
R8382 VDD.t2270 VDD.t2269 100.111
R8383 VDD.t2269 VDD.t2268 100.111
R8384 VDD.t2268 VDD.t451 100.111
R8385 VDD.t451 VDD.t455 100.111
R8386 VDD.t455 VDD.t457 100.111
R8387 VDD.t245 VDD.t249 100.111
R8388 VDD.t249 VDD.t251 100.111
R8389 VDD.t251 VDD.t2394 100.111
R8390 VDD.t2394 VDD.t2395 100.111
R8391 VDD.t2395 VDD.t1853 100.111
R8392 VDD.t2427 VDD.t2428 100.111
R8393 VDD.t2428 VDD.t2429 100.111
R8394 VDD.t2429 VDD.t2917 100.111
R8395 VDD.t2917 VDD.t2919 100.111
R8396 VDD.t2919 VDD.t2921 100.111
R8397 VDD.t2567 VDD.t2555 100.111
R8398 VDD.t2555 VDD.t2557 100.111
R8399 VDD.t2557 VDD.t2845 100.111
R8400 VDD.t2845 VDD.t2846 100.111
R8401 VDD.t2846 VDD.t2847 100.111
R8402 VDD.t691 VDD.t692 100.111
R8403 VDD.t692 VDD.t693 100.111
R8404 VDD.t693 VDD.t498 100.111
R8405 VDD.t498 VDD.t500 100.111
R8406 VDD.t500 VDD.t2735 100.111
R8407 VDD.t1607 VDD.t1611 100.111
R8408 VDD.t1611 VDD.t634 100.111
R8409 VDD.t634 VDD.t2034 100.111
R8410 VDD.t2034 VDD.t2035 100.111
R8411 VDD.t2035 VDD.t2036 100.111
R8412 VDD.t744 VDD.t745 100.111
R8413 VDD.t745 VDD.t746 100.111
R8414 VDD.t746 VDD.t1940 100.111
R8415 VDD.t1940 VDD.t1936 100.111
R8416 VDD.t1936 VDD.t1912 100.111
R8417 VDD.t1954 VDD.t1946 100.111
R8418 VDD.t1958 VDD.t1954 100.111
R8419 VDD.t907 VDD.t1958 100.111
R8420 VDD.t906 VDD.t907 100.111
R8421 VDD.t905 VDD.t906 100.111
R8422 VDD.t2733 VDD.t2033 100.111
R8423 VDD.t2033 VDD.t2734 100.111
R8424 VDD.t2734 VDD.t3391 100.111
R8425 VDD.t3391 VDD.t3393 100.111
R8426 VDD.t3393 VDD.t3389 100.111
R8427 VDD.t3514 VDD.t3512 100.111
R8428 VDD.t3512 VDD.t3522 100.111
R8429 VDD.t3522 VDD.t2007 100.111
R8430 VDD.t2007 VDD.t2006 100.111
R8431 VDD.t2006 VDD.t2005 100.111
R8432 VDD.t1536 VDD.t1538 100.111
R8433 VDD.t1538 VDD.t1537 100.111
R8434 VDD.t1537 VDD.t1072 100.111
R8435 VDD.t1072 VDD.t1884 100.111
R8436 VDD.t1884 VDD.t1882 100.111
R8437 VDD.t2776 VDD.t2774 100.111
R8438 VDD.t2774 VDD.t2772 100.111
R8439 VDD.t2772 VDD.t4309 100.111
R8440 VDD.t4309 VDD.t4308 100.111
R8441 VDD.t4308 VDD.t4307 100.111
R8442 VDD.t1242 VDD.t1243 100.111
R8443 VDD.t1243 VDD.t1241 100.111
R8444 VDD.t1241 VDD.t2008 100.111
R8445 VDD.t2008 VDD.t2018 100.111
R8446 VDD.t2018 VDD.t2016 100.111
R8447 VDD.t4018 VDD.t4012 100.111
R8448 VDD.t4012 VDD.t4010 100.111
R8449 VDD.t4010 VDD.t1652 100.111
R8450 VDD.t1652 VDD.t1651 100.111
R8451 VDD.t1651 VDD.t1650 100.111
R8452 VDD.t2023 VDD.t2022 100.111
R8453 VDD.t2022 VDD.t2024 100.111
R8454 VDD.t2024 VDD.t1904 100.111
R8455 VDD.t1904 VDD.t1896 100.111
R8456 VDD.t1896 VDD.t1902 100.111
R8457 VDD.t830 VDD.t840 100.111
R8458 VDD.t840 VDD.t838 100.111
R8459 VDD.t838 VDD.t102 100.111
R8460 VDD.t102 VDD.t101 100.111
R8461 VDD.t101 VDD.t100 100.111
R8462 VDD.t1615 VDD.t1109 100.111
R8463 VDD.t1109 VDD.t1616 100.111
R8464 VDD.t1616 VDD.t1279 100.111
R8465 VDD.t1279 VDD.t1277 100.111
R8466 VDD.t1277 VDD.t1275 100.111
R8467 VDD.t2449 VDD.t2447 100.111
R8468 VDD.t2447 VDD.t2445 100.111
R8469 VDD.t2445 VDD.t2857 100.111
R8470 VDD.t2857 VDD.t2649 100.111
R8471 VDD.t2649 VDD.t2858 100.111
R8472 VDD.t1314 VDD.t1313 100.111
R8473 VDD.t1315 VDD.t1314 100.111
R8474 VDD.t1815 VDD.t1315 100.111
R8475 VDD.t160 VDD.t1815 100.111
R8476 VDD.t156 VDD.t160 100.111
R8477 VDD.t938 VDD.t936 100.111
R8478 VDD.t934 VDD.t938 100.111
R8479 VDD.t2728 VDD.t934 100.111
R8480 VDD.t2727 VDD.t2728 100.111
R8481 VDD.t2726 VDD.t2727 100.111
R8482 VDD.t1549 VDD.t1548 100.111
R8483 VDD.t1548 VDD.t2484 100.111
R8484 VDD.t2484 VDD.t3657 100.111
R8485 VDD.t3657 VDD.t3653 100.111
R8486 VDD.t3653 VDD.t3655 100.111
R8487 VDD.t3316 VDD.t3312 100.111
R8488 VDD.t3312 VDD.t3310 100.111
R8489 VDD.t3310 VDD.t2432 100.111
R8490 VDD.t2432 VDD.t2431 100.111
R8491 VDD.t2431 VDD.t2430 100.111
R8492 VDD.t3454 VDD.t3453 100.111
R8493 VDD.t3453 VDD.t3455 100.111
R8494 VDD.t3455 VDD.t4062 100.111
R8495 VDD.t4062 VDD.t4060 100.111
R8496 VDD.t4060 VDD.t4054 100.111
R8497 VDD.t1960 VDD.t1970 100.111
R8498 VDD.t1948 VDD.t1960 100.111
R8499 VDD.t1701 VDD.t1948 100.111
R8500 VDD.t1836 VDD.t1701 100.111
R8501 VDD.t1190 VDD.t1836 100.111
R8502 VDD.t1042 VDD.t1041 100.111
R8503 VDD.t1043 VDD.t1042 100.111
R8504 VDD.t1590 VDD.t1043 100.111
R8505 VDD.t597 VDD.t1590 100.111
R8506 VDD.t599 VDD.t597 100.111
R8507 VDD.t3198 VDD.t3196 100.111
R8508 VDD.t3190 VDD.t3198 100.111
R8509 VDD.t1080 VDD.t3190 100.111
R8510 VDD.t1081 VDD.t1080 100.111
R8511 VDD.t1347 VDD.t1081 100.111
R8512 VDD.t1699 VDD.t699 100.111
R8513 VDD.t1700 VDD.t1699 100.111
R8514 VDD.t2507 VDD.t1700 100.111
R8515 VDD.t2501 VDD.t2507 100.111
R8516 VDD.t2505 VDD.t2501 100.111
R8517 VDD.t4283 VDD.t4281 100.111
R8518 VDD.t4287 VDD.t4283 100.111
R8519 VDD.t2434 VDD.t4287 100.111
R8520 VDD.t3382 VDD.t2434 100.111
R8521 VDD.t2433 VDD.t3382 100.111
R8522 VDD.t1837 VDD.t1838 100.111
R8523 VDD.t1839 VDD.t1837 100.111
R8524 VDD.t3891 VDD.t1839 100.111
R8525 VDD.t3883 VDD.t3891 100.111
R8526 VDD.t3885 VDD.t3883 100.111
R8527 VDD.t111 VDD.t113 100.111
R8528 VDD.t115 VDD.t111 100.111
R8529 VDD.t3620 VDD.t115 100.111
R8530 VDD.t3621 VDD.t3620 100.111
R8531 VDD.t3622 VDD.t3621 100.111
R8532 VDD.t3689 VDD.t3691 100.111
R8533 VDD.t3688 VDD.t3689 100.111
R8534 VDD.t3271 VDD.t3688 100.111
R8535 VDD.t3277 VDD.t3271 100.111
R8536 VDD.t3275 VDD.t3277 100.111
R8537 VDD.t3675 VDD.t3671 100.111
R8538 VDD.t3679 VDD.t3675 100.111
R8539 VDD.t60 VDD.t3679 100.111
R8540 VDD.t59 VDD.t60 100.111
R8541 VDD.t61 VDD.t59 100.111
R8542 VDD.t1440 VDD.t1439 100.111
R8543 VDD.t2396 VDD.t1440 100.111
R8544 VDD.t664 VDD.t2396 100.111
R8545 VDD.t670 VDD.t664 100.111
R8546 VDD.t672 VDD.t670 100.111
R8547 VDD.t22 VDD.t18 100.111
R8548 VDD.t26 VDD.t22 100.111
R8549 VDD.t3290 VDD.t26 100.111
R8550 VDD.t3288 VDD.t3290 100.111
R8551 VDD.t3289 VDD.t3288 100.111
R8552 VDD.t732 VDD.t733 100.111
R8553 VDD.t733 VDD.t1040 100.111
R8554 VDD.t1040 VDD.t4034 100.111
R8555 VDD.t4034 VDD.t4036 100.111
R8556 VDD.t4036 VDD.t4028 100.111
R8557 VDD.t4150 VDD.t4156 100.111
R8558 VDD.t4156 VDD.t4158 100.111
R8559 VDD.t4158 VDD.t1345 100.111
R8560 VDD.t1345 VDD.t1346 100.111
R8561 VDD.t1346 VDD.t1344 100.111
R8562 VDD.t275 VDD.t276 100.111
R8563 VDD.t276 VDD.t277 100.111
R8564 VDD.t277 VDD.t1054 100.111
R8565 VDD.t1054 VDD.t1044 100.111
R8566 VDD.t1044 VDD.t1046 100.111
R8567 VDD.t4271 VDD.t3934 100.111
R8568 VDD.t3934 VDD.t4312 100.111
R8569 VDD.t4312 VDD.t2869 100.111
R8570 VDD.t2869 VDD.t2870 100.111
R8571 VDD.t2870 VDD.t2868 100.111
R8572 VDD.t2859 VDD.t2860 100.111
R8573 VDD.t2860 VDD.t2861 100.111
R8574 VDD.t2861 VDD.t2718 100.111
R8575 VDD.t2718 VDD.t2722 100.111
R8576 VDD.t2722 VDD.t2714 100.111
R8577 VDD.t1767 VDD.t1751 100.111
R8578 VDD.t1793 VDD.t1767 100.111
R8579 VDD.t2393 VDD.t1793 100.111
R8580 VDD.t1441 VDD.t2393 100.111
R8581 VDD.t3378 VDD.t1441 100.111
R8582 VDD.t3121 VDD.t3119 100.111
R8583 VDD.t3119 VDD.t3120 100.111
R8584 VDD.t3120 VDD.t2260 100.111
R8585 VDD.t2260 VDD.t2258 100.111
R8586 VDD.t2258 VDD.t2264 100.111
R8587 VDD.t1677 VDD.t2244 100.111
R8588 VDD.t2244 VDD.t2231 100.111
R8589 VDD.t2231 VDD.t1253 100.111
R8590 VDD.t1253 VDD.t1252 100.111
R8591 VDD.t1252 VDD.t1254 100.111
R8592 VDD.t581 VDD.t2554 100.111
R8593 VDD.t2554 VDD.t582 100.111
R8594 VDD.t582 VDD.t2088 100.111
R8595 VDD.t2088 VDD.t2082 100.111
R8596 VDD.t2082 VDD.t2094 100.111
R8597 VDD.t2624 VDD.t2630 100.111
R8598 VDD.t2630 VDD.t2628 100.111
R8599 VDD.t2628 VDD.t2266 100.111
R8600 VDD.t2266 VDD.t178 100.111
R8601 VDD.t178 VDD.t2267 100.111
R8602 VDD.t1543 VDD.t1624 100.111
R8603 VDD.t1624 VDD.t1542 100.111
R8604 VDD.t1542 VDD.t756 100.111
R8605 VDD.t756 VDD.t754 100.111
R8606 VDD.t754 VDD.t760 100.111
R8607 VDD.t4199 VDD.t4225 100.111
R8608 VDD.t4225 VDD.t4232 100.111
R8609 VDD.t4232 VDD.t1183 100.111
R8610 VDD.t1183 VDD.t1182 100.111
R8611 VDD.t1182 VDD.t3380 100.111
R8612 VDD.t799 VDD.t798 100.111
R8613 VDD.t798 VDD.t797 100.111
R8614 VDD.t797 VDD.t4142 100.111
R8615 VDD.t4142 VDD.t4140 100.111
R8616 VDD.t4140 VDD.t4144 100.111
R8617 VDD.t88 VDD.t86 100.111
R8618 VDD.t86 VDD.t90 100.111
R8619 VDD.t90 VDD.t885 100.111
R8620 VDD.t885 VDD.t886 100.111
R8621 VDD.t886 VDD.t884 100.111
R8622 VDD.t3379 VDD.t1231 100.111
R8623 VDD.t1230 VDD.t3379 100.111
R8624 VDD.t2462 VDD.t1230 100.111
R8625 VDD.t2460 VDD.t2462 100.111
R8626 VDD.t2435 VDD.t2460 100.111
R8627 VDD.t267 VDD.t529 100.111
R8628 VDD.t549 VDD.t267 100.111
R8629 VDD.t335 VDD.t549 100.111
R8630 VDD.t334 VDD.t335 100.111
R8631 VDD.t336 VDD.t334 100.111
R8632 VDD.t1517 VDD.t1518 100.111
R8633 VDD.t227 VDD.t1517 100.111
R8634 VDD.t345 VDD.t227 100.111
R8635 VDD.t339 VDD.t345 100.111
R8636 VDD.t878 VDD.t339 100.111
R8637 VDD.t1731 VDD.t1739 100.111
R8638 VDD.t1729 VDD.t1731 100.111
R8639 VDD.t2183 VDD.t1729 100.111
R8640 VDD.t333 VDD.t2183 100.111
R8641 VDD.t2184 VDD.t333 100.111
R8642 VDD.t1566 VDD.t1564 100.111
R8643 VDD.t1564 VDD.t1565 100.111
R8644 VDD.t1565 VDD.t1550 100.111
R8645 VDD.t1550 VDD.t1552 100.111
R8646 VDD.t1552 VDD.t1554 100.111
R8647 VDD.t4121 VDD.t4101 100.111
R8648 VDD.t4101 VDD.t4083 100.111
R8649 VDD.t4083 VDD.t955 100.111
R8650 VDD.t955 VDD.t954 100.111
R8651 VDD.t954 VDD.t953 100.111
R8652 VDD.t1575 VDD.t1577 100.111
R8653 VDD.t1577 VDD.t1576 100.111
R8654 VDD.t1576 VDD.t617 100.111
R8655 VDD.t617 VDD.t609 100.111
R8656 VDD.t609 VDD.t621 100.111
R8657 VDD.t3938 VDD.t3950 100.111
R8658 VDD.t3950 VDD.t3946 100.111
R8659 VDD.t3946 VDD.t772 100.111
R8660 VDD.t772 VDD.t774 100.111
R8661 VDD.t774 VDD.t773 100.111
R8662 VDD.t2076 VDD.t1164 100.111
R8663 VDD.t2747 VDD.t2076 100.111
R8664 VDD.t347 VDD.t2747 100.111
R8665 VDD.t303 VDD.t347 100.111
R8666 VDD.t351 VDD.t303 100.111
R8667 VDD.t2191 VDD.t2201 100.111
R8668 VDD.t1635 VDD.t2191 100.111
R8669 VDD.t557 VDD.t1635 100.111
R8670 VDD.t559 VDD.t557 100.111
R8671 VDD.t558 VDD.t559 100.111
R8672 VDD.t3377 VDD.t3375 100.111
R8673 VDD.t3376 VDD.t3377 100.111
R8674 VDD.t1427 VDD.t3376 100.111
R8675 VDD.t1429 VDD.t1427 100.111
R8676 VDD.t1437 VDD.t1429 100.111
R8677 VDD.t2754 VDD.t2748 100.111
R8678 VDD.t2750 VDD.t2754 100.111
R8679 VDD.t1483 VDD.t2750 100.111
R8680 VDD.t1485 VDD.t1483 100.111
R8681 VDD.t1484 VDD.t1485 100.111
R8682 VDD.t140 VDD.t139 100.111
R8683 VDD.t139 VDD.t141 100.111
R8684 VDD.t141 VDD.t3904 100.111
R8685 VDD.t3904 VDD.t3900 100.111
R8686 VDD.t3900 VDD.t3912 100.111
R8687 VDD.t387 VDD.t379 100.111
R8688 VDD.t379 VDD.t395 100.111
R8689 VDD.t395 VDD.t2046 100.111
R8690 VDD.t2046 VDD.t2045 100.111
R8691 VDD.t2045 VDD.t2047 100.111
R8692 VDD.t3899 VDD.t3898 100.111
R8693 VDD.t3898 VDD.t3897 100.111
R8694 VDD.t3897 VDD.t2876 100.111
R8695 VDD.t2876 VDD.t2872 100.111
R8696 VDD.t2872 VDD.t2874 100.111
R8697 VDD.t1144 VDD.t1123 100.111
R8698 VDD.t1123 VDD.t1146 100.111
R8699 VDD.t1146 VDD.t1449 100.111
R8700 VDD.t1449 VDD.t1448 100.111
R8701 VDD.t1448 VDD.t1450 100.111
R8702 VDD.t1544 VDD.t2648 100.111
R8703 VDD.t1494 VDD.t1544 100.111
R8704 VDD.t2399 VDD.t1494 100.111
R8705 VDD.t822 VDD.t2399 100.111
R8706 VDD.t2409 VDD.t822 100.111
R8707 VDD.t2834 VDD.t2817 100.111
R8708 VDD.t2827 VDD.t2834 100.111
R8709 VDD.t1216 VDD.t2827 100.111
R8710 VDD.t1215 VDD.t1216 100.111
R8711 VDD.t1217 VDD.t1215 100.111
R8712 VDD.t724 VDD.t1196 100.111
R8713 VDD.t1195 VDD.t724 100.111
R8714 VDD.t3232 VDD.t1195 100.111
R8715 VDD.t3236 VDD.t3232 100.111
R8716 VDD.t3234 VDD.t3236 100.111
R8717 VDD.t1872 VDD.t1874 100.111
R8718 VDD.t172 VDD.t1872 100.111
R8719 VDD.t1618 VDD.t172 100.111
R8720 VDD.t1617 VDD.t1618 100.111
R8721 VDD.t1619 VDD.t1617 100.111
R8722 VDD.t2487 VDD.t2488 100.111
R8723 VDD.t2489 VDD.t2487 100.111
R8724 VDD.t3477 VDD.t2489 100.111
R8725 VDD.t3469 VDD.t3477 100.111
R8726 VDD.t3471 VDD.t3469 100.111
R8727 VDD.t3421 VDD.t3427 100.111
R8728 VDD.t3444 VDD.t3421 100.111
R8729 VDD.t3882 VDD.t3444 100.111
R8730 VDD.t3881 VDD.t3882 100.111
R8731 VDD.t3880 VDD.t3881 100.111
R8732 VDD.t57 VDD.t3466 100.111
R8733 VDD.t3466 VDD.t58 100.111
R8734 VDD.t58 VDD.t3639 100.111
R8735 VDD.t3639 VDD.t3645 100.111
R8736 VDD.t3645 VDD.t3641 100.111
R8737 VDD.t1408 VDD.t1174 97.1116
R8738 VDD.t1771 VDD.t1789 97.1116
R8739 VDD.t3554 VDD.t3529 97.1116
R8740 VDD.t1765 VDD.t1753 97.1116
R8741 VDD.t3966 VDD.t3972 97.1116
R8742 VDD.t1773 VDD.t777 97.1116
R8743 VDD.t3602 VDD.t3596 97.1116
R8744 VDD.t1747 VDD.t1813 97.1116
R8745 VDD.t2130 VDD.t2155 97.1116
R8746 VDD.t1805 VDD.t1757 97.1116
R8747 VDD.t2603 VDD.t2573 97.1116
R8748 VDD.t1783 VDD.t762 97.1116
R8749 VDD.t2353 VDD.t1833 97.1116
R8750 VDD.t1777 VDD.t781 97.1116
R8751 VDD.t1004 VDD.t585 97.1116
R8752 VDD.t1763 VDD.t775 97.1116
R8753 VDD.t3442 VDD.t2288 97.1116
R8754 VDD.t1396 VDD.t1180 97.1116
R8755 VDD.t1657 VDD.t1672 97.1116
R8756 VDD.t595 VDD.t987 97.1116
R8757 VDD.t978 VDD.t980 97.0038
R8758 VDD.t783 VDD.t1781 97.0038
R8759 VDD.t1391 VDD.t1406 97.0038
R8760 VDD.t3425 VDD.t3450 97.0038
R8761 VDD.t3304 VDD.t3300 97.0038
R8762 VDD.t3447 VDD.t3423 97.0038
R8763 VDD.t2843 VDD.t2825 96.8963
R8764 VDD.t3539 VDD.t3548 96.8963
R8765 VDD.t376 VDD.t401 96.8963
R8766 VDD.t3968 VDD.t897 96.8963
R8767 VDD.t2193 VDD.t2199 96.8963
R8768 VDD.t3584 VDD.t3579 96.8963
R8769 VDD.t4073 VDD.t4119 96.8963
R8770 VDD.t2153 VDD.t2180 96.8963
R8771 VDD.t269 VDD.t525 96.8963
R8772 VDD.t483 VDD.t479 96.8963
R8773 VDD.t4230 VDD.t4194 96.8963
R8774 VDD.t2345 VDD.t2318 96.8963
R8775 VDD.n1422 VDD.t2100 96.8274
R8776 VDD.n1684 VDD.t1942 96.8274
R8777 VDD.n1691 VDD.t3516 96.8274
R8778 VDD.n1699 VDD.t4000 96.8274
R8779 VDD.t2778 VDD.n1698 96.8274
R8780 VDD.n1817 VDD.t4016 96.8274
R8781 VDD.n1824 VDD.t1697 96.8274
R8782 VDD.n1825 VDD.t842 96.8274
R8783 VDD.n1837 VDD.t2437 96.8274
R8784 VDD.n1838 VDD.t2072 96.8274
R8785 VDD.n1849 VDD.t946 96.8274
R8786 VDD.n1850 VDD.t3314 96.8274
R8787 VDD.n1474 VDD.t2745 96.8274
R8788 VDD.n1554 VDD.t1952 96.8274
R8789 VDD.t3186 VDD.n1553 96.8274
R8790 VDD.t3685 VDD.n1546 96.8274
R8791 VDD.t4285 VDD.n1539 96.8274
R8792 VDD.t107 VDD.n1529 96.8274
R8793 VDD.t4042 VDD.n1522 96.8274
R8794 VDD.t3677 VDD.n1515 96.8274
R8795 VDD.t30 VDD.n1505 96.8274
R8796 VDD.t575 VDD.n1498 96.8274
R8797 VDD.t4152 VDD.n1491 96.8274
R8798 VDD.t3936 VDD.n1481 96.8274
R8799 VDD.n1397 VDD.t225 96.8274
R8800 VDD.n1398 VDD.t1978 96.8274
R8801 VDD.n1713 VDD.t1299 96.8274
R8802 VDD.n1720 VDD.t716 96.8274
R8803 VDD.n1778 VDD.t209 96.8274
R8804 VDD.t2304 VDD.n1777 96.8274
R8805 VDD.t1131 VDD.n1770 96.8274
R8806 VDD.t706 VDD.n1763 96.8274
R8807 VDD.n1750 VDD.t253 96.8274
R8808 VDD.t718 VDD.n1749 96.8274
R8809 VDD.n1738 VDD.t2563 96.8274
R8810 VDD.t1605 VDD.n1737 96.8274
R8811 VDD.n2477 VDD.t1822 96.8274
R8812 VDD.n2478 VDD.t1761 96.8274
R8813 VDD.n2526 VDD.t2219 96.8274
R8814 VDD.n2530 VDD.t2537 96.8274
R8815 VDD.n2531 VDD.t801 96.8274
R8816 VDD.n2542 VDD.t4202 96.8274
R8817 VDD.n2546 VDD.t443 96.8274
R8818 VDD.n2565 VDD.t82 96.8274
R8819 VDD.t541 VDD.n2564 96.8274
R8820 VDD.t2185 VDD.n2560 96.8274
R8821 VDD.t1735 VDD.n2553 96.8274
R8822 VDD.n2606 VDD.t4096 96.8274
R8823 VDD.n2610 VDD.t3462 96.8274
R8824 VDD.n2629 VDD.t3942 96.8274
R8825 VDD.t1627 VDD.n2628 96.8274
R8826 VDD.t2702 VDD.n2624 96.8274
R8827 VDD.t2758 VDD.n2617 96.8274
R8828 VDD.n2670 VDD.t405 96.8274
R8829 VDD.n2674 VDD.t2474 96.8274
R8830 VDD.n2705 VDD.t1121 96.8274
R8831 VDD.t2839 VDD.n2704 96.8274
R8832 VDD.t1842 VDD.n2697 96.8274
R8833 VDD.n2687 VDD.t1880 96.8274
R8834 VDD.t3436 VDD.n2686 96.8274
R8835 VDD.t3558 VDD.n2218 96.6506
R8836 VDD.n2243 VDD.t321 96.6506
R8837 VDD.n1884 VDD.t1573 96.6506
R8838 VDD.t1982 VDD.t1924 95.939
R8839 VDD.t2054 VDD.t1601 95.939
R8840 VDD.t1297 VDD.t1289 95.939
R8841 VDD.t287 VDD.t291 95.939
R8842 VDD.t215 VDD.t2417 95.939
R8843 VDD.t4179 VDD.t4171 95.939
R8844 VDD.t2310 VDD.t2306 95.939
R8845 VDD.t1338 VDD.t1342 95.939
R8846 VDD.t3988 VDD.t704 95.939
R8847 VDD.t457 VDD.t453 95.939
R8848 VDD.t255 VDD.t245 95.939
R8849 VDD.t2921 VDD.t2911 95.939
R8850 VDD.t2559 VDD.t2567 95.939
R8851 VDD.t2735 VDD.t494 95.939
R8852 VDD.t638 VDD.t1607 95.939
R8853 VDD.t1912 VDD.t1938 95.939
R8854 VDD.t1946 VDD.t1934 95.939
R8855 VDD.t3389 VDD.t3387 95.939
R8856 VDD.t3518 VDD.t3514 95.939
R8857 VDD.t1882 VDD.t1074 95.939
R8858 VDD.t2780 VDD.t2776 95.939
R8859 VDD.t2016 VDD.t2014 95.939
R8860 VDD.t4014 VDD.t4018 95.939
R8861 VDD.t1902 VDD.t1898 95.939
R8862 VDD.t832 VDD.t830 95.939
R8863 VDD.t1275 VDD.t1287 95.939
R8864 VDD.t2439 VDD.t2449 95.939
R8865 VDD.t150 VDD.t156 95.939
R8866 VDD.t936 VDD.t940 95.939
R8867 VDD.t3655 VDD.t3665 95.939
R8868 VDD.t3318 VDD.t3316 95.939
R8869 VDD.t4054 VDD.t4050 95.939
R8870 VDD.t1970 VDD.t1916 95.939
R8871 VDD.t603 VDD.t599 95.939
R8872 VDD.t3196 VDD.t3188 95.939
R8873 VDD.t2509 VDD.t2505 95.939
R8874 VDD.t4281 VDD.t4289 95.939
R8875 VDD.t3893 VDD.t3885 95.939
R8876 VDD.t113 VDD.t109 95.939
R8877 VDD.t3494 VDD.t3275 95.939
R8878 VDD.t3671 VDD.t3667 95.939
R8879 VDD.t666 VDD.t672 95.939
R8880 VDD.t18 VDD.t28 95.939
R8881 VDD.t4028 VDD.t4032 95.939
R8882 VDD.t4160 VDD.t4150 95.939
R8883 VDD.t1046 VDD.t1052 95.939
R8884 VDD.t4310 VDD.t4271 95.939
R8885 VDD.t2714 VDD.t2720 95.939
R8886 VDD.t1751 VDD.t1801 95.939
R8887 VDD.t2264 VDD.t2262 95.939
R8888 VDD.t2227 VDD.t1677 95.939
R8889 VDD.t2094 VDD.t2086 95.939
R8890 VDD.t2626 VDD.t2624 95.939
R8891 VDD.t760 VDD.t758 95.939
R8892 VDD.t4221 VDD.t4199 95.939
R8893 VDD.t4144 VDD.t4146 95.939
R8894 VDD.t92 VDD.t88 95.939
R8895 VDD.t2464 VDD.t2435 95.939
R8896 VDD.t529 VDD.t261 95.939
R8897 VDD.t876 VDD.t878 95.939
R8898 VDD.t1739 VDD.t1727 95.939
R8899 VDD.t1554 VDD.t1556 95.939
R8900 VDD.t4099 VDD.t4121 95.939
R8901 VDD.t621 VDD.t619 95.939
R8902 VDD.t3948 VDD.t3938 95.939
R8903 VDD.t349 VDD.t351 95.939
R8904 VDD.t2201 VDD.t1638 95.939
R8905 VDD.t1425 VDD.t1437 95.939
R8906 VDD.t2748 VDD.t2752 95.939
R8907 VDD.t3912 VDD.t3902 95.939
R8908 VDD.t391 VDD.t387 95.939
R8909 VDD.t2874 VDD.t2884 95.939
R8910 VDD.t1115 VDD.t1144 95.939
R8911 VDD.t2403 VDD.t2409 95.939
R8912 VDD.t2817 VDD.t2823 95.939
R8913 VDD.t3244 VDD.t3234 95.939
R8914 VDD.t1874 VDD.t1876 95.939
R8915 VDD.t3467 VDD.t3471 95.939
R8916 VDD.t3427 VDD.t3440 95.939
R8917 VDD.t3641 VDD.t3651 95.939
R8918 VDD.n2378 VDD.t1665 95.3603
R8919 VDD.n2408 VDD.t4228 95.3603
R8920 VDD.n2401 VDD.t517 95.3603
R8921 VDD.t4091 VDD.n2396 95.3603
R8922 VDD.n1116 VDD.n1115 94.8255
R8923 VDD.n1106 VDD.n1105 94.8255
R8924 VDD.n1104 VDD.n1103 94.8255
R8925 VDD.n1094 VDD.n1093 94.8255
R8926 VDD.n1118 VDD.n1117 94.8255
R8927 VDD.n1027 VDD.n1026 94.8255
R8928 VDD.n1049 VDD.n1048 94.8255
R8929 VDD.n1039 VDD.n1038 94.8255
R8930 VDD.n1037 VDD.n1036 94.8255
R8931 VDD.n1051 VDD.n1050 94.8255
R8932 VDD.n987 VDD.n986 94.8255
R8933 VDD.n977 VDD.n976 94.8255
R8934 VDD.n975 VDD.n974 94.8255
R8935 VDD.n965 VDD.n964 94.8255
R8936 VDD.n989 VDD.n988 94.8255
R8937 VDD.n898 VDD.n897 94.8255
R8938 VDD.n920 VDD.n919 94.8255
R8939 VDD.n910 VDD.n909 94.8255
R8940 VDD.n908 VDD.n907 94.8255
R8941 VDD.n922 VDD.n921 94.8255
R8942 VDD.n858 VDD.n857 94.8255
R8943 VDD.n848 VDD.n847 94.8255
R8944 VDD.n846 VDD.n845 94.8255
R8945 VDD.n836 VDD.n835 94.8255
R8946 VDD.n860 VDD.n859 94.8255
R8947 VDD.n769 VDD.n768 94.8255
R8948 VDD.n791 VDD.n790 94.8255
R8949 VDD.n781 VDD.n780 94.8255
R8950 VDD.n779 VDD.n778 94.8255
R8951 VDD.n793 VDD.n792 94.8255
R8952 VDD.n729 VDD.n728 94.8255
R8953 VDD.n719 VDD.n718 94.8255
R8954 VDD.n717 VDD.n716 94.8255
R8955 VDD.n707 VDD.n706 94.8255
R8956 VDD.n731 VDD.n730 94.8255
R8957 VDD.n640 VDD.n639 94.8255
R8958 VDD.n630 VDD.n629 94.8255
R8959 VDD.n628 VDD.n627 94.8255
R8960 VDD.n618 VDD.n617 94.8255
R8961 VDD.n642 VDD.n641 94.8255
R8962 VDD.n578 VDD.n577 94.8255
R8963 VDD.n568 VDD.n567 94.8255
R8964 VDD.n566 VDD.n565 94.8255
R8965 VDD.n556 VDD.n555 94.8255
R8966 VDD.n580 VDD.n579 94.8255
R8967 VDD.n489 VDD.n488 94.8255
R8968 VDD.n511 VDD.n510 94.8255
R8969 VDD.n501 VDD.n500 94.8255
R8970 VDD.n499 VDD.n498 94.8255
R8971 VDD.n513 VDD.n512 94.8255
R8972 VDD.n449 VDD.n448 94.8255
R8973 VDD.n439 VDD.n438 94.8255
R8974 VDD.n437 VDD.n436 94.8255
R8975 VDD.n427 VDD.n426 94.8255
R8976 VDD.n451 VDD.n450 94.8255
R8977 VDD.n360 VDD.n359 94.8255
R8978 VDD.n382 VDD.n381 94.8255
R8979 VDD.n372 VDD.n371 94.8255
R8980 VDD.n370 VDD.n369 94.8255
R8981 VDD.n384 VDD.n383 94.8255
R8982 VDD.n320 VDD.n319 94.8255
R8983 VDD.n310 VDD.n309 94.8255
R8984 VDD.n308 VDD.n307 94.8255
R8985 VDD.n298 VDD.n297 94.8255
R8986 VDD.n322 VDD.n321 94.8255
R8987 VDD.n191 VDD.n190 94.8255
R8988 VDD.n181 VDD.n180 94.8255
R8989 VDD.n179 VDD.n178 94.8255
R8990 VDD.n169 VDD.n168 94.8255
R8991 VDD.n193 VDD.n192 94.8255
R8992 VDD.n231 VDD.n230 94.8255
R8993 VDD.n253 VDD.n252 94.8255
R8994 VDD.n243 VDD.n242 94.8255
R8995 VDD.n241 VDD.n240 94.8255
R8996 VDD.n255 VDD.n254 94.8255
R8997 VDD.n93 VDD.n92 94.8255
R8998 VDD.n115 VDD.n114 94.8255
R8999 VDD.n105 VDD.n104 94.8255
R9000 VDD.n103 VDD.n102 94.8255
R9001 VDD.n117 VDD.n116 94.8255
R9002 VDD.n2896 VDD.n2895 94.8255
R9003 VDD.n2886 VDD.n2885 94.8255
R9004 VDD.n2884 VDD.n2883 94.8255
R9005 VDD.n2874 VDD.n2873 94.8255
R9006 VDD.n2898 VDD.n2897 94.8255
R9007 VDD.n31 VDD.n30 94.8255
R9008 VDD.n53 VDD.n52 94.8255
R9009 VDD.n43 VDD.n42 94.8255
R9010 VDD.n41 VDD.n40 94.8255
R9011 VDD.n55 VDD.n54 94.8255
R9012 VDD.n1134 VDD.t4126 94.5607
R9013 VDD.n1919 VDD.t3543 94.5607
R9014 VDD.n1909 VDD.t1414 94.5607
R9015 VDD.n1926 VDD.t903 94.5607
R9016 VDD.n1927 VDD.t3600 94.5607
R9017 VDD.n1938 VDD.t2157 94.5607
R9018 VDD.n1945 VDD.t481 94.5607
R9019 VDD.n1946 VDD.t2364 94.5607
R9020 VDD.t997 VDD.n1899 94.5607
R9021 VDD.t195 VDD.n683 94.5607
R9022 VDD.t4241 VDD.n1309 92.8972
R9023 VDD.t4079 VDD.n1321 92.8972
R9024 VDD.t2134 VDD.n1285 92.8972
R9025 VDD.t2143 VDD.n1297 92.8972
R9026 VDD.t469 VDD.n1237 92.8972
R9027 VDD.t2613 VDD.n1249 92.8972
R9028 VDD.t4235 VDD.n1213 92.8972
R9029 VDD.t4103 VDD.n1225 92.8972
R9030 VDD.n1190 VDD.t2327 92.8972
R9031 VDD.t2358 VDD.n1200 90.2335
R9032 VDD.n1953 VDD.t1006 87.2622
R9033 VDD.n2329 VDD.t2333 87.2622
R9034 VDD.n2319 VDD.t2575 87.2622
R9035 VDD.n2309 VDD.t2122 87.2622
R9036 VDD.n2298 VDD.t3586 87.2622
R9037 VDD.n2288 VDD.t3977 87.2622
R9038 VDD.n2278 VDD.t3550 87.2622
R9039 VDD.n2268 VDD.t1398 87.2622
R9040 VDD.n1064 VDD.t36 87.2622
R9041 VDD.n935 VDD.t3924 87.2622
R9042 VDD.n806 VDD.t1226 87.2622
R9043 VDD.n655 VDD.t4301 87.2622
R9044 VDD.n526 VDD.t4257 87.2622
R9045 VDD.n397 VDD.t738 87.2622
R9046 VDD.n268 VDD.t2905 87.2622
R9047 VDD.n130 VDD.t4320 87.2622
R9048 VDD.n2914 VDD.t3508 87.2622
R9049 VDD.n1145 VDD.n1144 85.724
R9050 VDD.n1142 VDD.n1140 85.724
R9051 VDD.n1261 VDD.t2583 84.054
R9052 VDD.n1273 VDD.t463 84.054
R9053 VDD.n1422 VDD.t866 78.5582
R9054 VDD.t3385 VDD.n1684 78.5582
R9055 VDD.t1886 VDD.n1691 78.5582
R9056 VDD.n1699 VDD.t3407 78.5582
R9057 VDD.n1698 VDD.t2012 78.5582
R9058 VDD.t1900 VDD.n1817 78.5582
R9059 VDD.t1466 VDD.n1824 78.5582
R9060 VDD.n1825 VDD.t1285 78.5582
R9061 VDD.t154 VDD.n1837 78.5582
R9062 VDD.n1838 VDD.t969 78.5582
R9063 VDD.t3663 VDD.n1849 78.5582
R9064 VDD.n1850 VDD.t4058 78.5582
R9065 VDD.t2217 VDD.n1474 78.5582
R9066 VDD.n1554 VDD.t601 78.5582
R9067 VDD.n1553 VDD.t2497 78.5582
R9068 VDD.n1546 VDD.t4265 78.5582
R9069 VDD.n1539 VDD.t3887 78.5582
R9070 VDD.n1529 VDD.t3269 78.5582
R9071 VDD.n1522 VDD.t4044 78.5582
R9072 VDD.n1515 VDD.t660 78.5582
R9073 VDD.n1505 VDD.t4026 78.5582
R9074 VDD.n1498 VDD.t144 78.5582
R9075 VDD.n1491 VDD.t1048 78.5582
R9076 VDD.n1481 VDD.t2724 78.5582
R9077 VDD.t2248 VDD.n1397 78.5582
R9078 VDD.n1398 VDD.t1603 78.5582
R9079 VDD.t293 VDD.n1713 78.5582
R9080 VDD.t2515 VDD.n1720 78.5582
R9081 VDD.n1778 VDD.t4173 78.5582
R9082 VDD.n1777 VDD.t1330 78.5582
R9083 VDD.n1770 VDD.t1084 78.5582
R9084 VDD.n1763 VDD.t459 78.5582
R9085 VDD.n1750 VDD.t2915 78.5582
R9086 VDD.n1749 VDD.t4325 78.5582
R9087 VDD.n1738 VDD.t2737 78.5582
R9088 VDD.n1737 VDD.t1932 78.5582
R9089 VDD.t3403 VDD.n2477 78.5582
R9090 VDD.n2478 VDD.t2254 78.5582
R9091 VDD.t2092 VDD.n2526 78.5582
R9092 VDD.t1362 VDD.n2530 78.5582
R9093 VDD.n2531 VDD.t752 78.5582
R9094 VDD.t4136 VDD.n2542 78.5582
R9095 VDD.t3328 VDD.n2546 78.5582
R9096 VDD.n2565 VDD.t2470 78.5582
R9097 VDD.n2564 VDD.t343 78.5582
R9098 VDD.n2560 VDD.t1856 78.5582
R9099 VDD.n2553 VDD.t1558 78.5582
R9100 VDD.t615 VDD.n2606 78.5582
R9101 VDD.t3998 VDD.n2610 78.5582
R9102 VDD.n2629 VDD.t297 78.5582
R9103 VDD.n2628 VDD.t1431 78.5582
R9104 VDD.n2624 VDD.t1851 78.5582
R9105 VDD.n2617 VDD.t3906 78.5582
R9106 VDD.t2878 VDD.n2670 78.5582
R9107 VDD.t1582 VDD.n2674 78.5582
R9108 VDD.n2705 VDD.t2401 78.5582
R9109 VDD.n2704 VDD.t3238 78.5582
R9110 VDD.n2697 VDD.t2690 78.5582
R9111 VDD.n2687 VDD.t3473 78.5582
R9112 VDD.n2686 VDD.t3643 78.5582
R9113 VDD.t991 VDD.n2378 77.3679
R9114 VDD.n2408 VDD.t1034 77.3679
R9115 VDD.n2401 VDD.t995 77.3679
R9116 VDD.n2396 VDD.t593 77.3679
R9117 VDD.n1885 VDD.t824 76.0927
R9118 VDD.n1957 VDD.n1952 75.6711
R9119 VDD.n2333 VDD.n2328 75.6711
R9120 VDD.n2323 VDD.n2318 75.6711
R9121 VDD.n2313 VDD.n2308 75.6711
R9122 VDD.n2302 VDD.n2297 75.6711
R9123 VDD.n2292 VDD.n2287 75.6711
R9124 VDD.n2282 VDD.n2277 75.6711
R9125 VDD.n2272 VDD.n2267 75.6711
R9126 VDD.n1068 VDD.n1060 75.6711
R9127 VDD.n939 VDD.n931 75.6711
R9128 VDD.n810 VDD.n802 75.6711
R9129 VDD.n659 VDD.n651 75.6711
R9130 VDD.n530 VDD.n522 75.6711
R9131 VDD.n401 VDD.n393 75.6711
R9132 VDD.n272 VDD.n264 75.6711
R9133 VDD.n134 VDD.n126 75.6711
R9134 VDD.n2918 VDD.n2910 75.6711
R9135 VDD.n1309 VDD.t2138 75.3695
R9136 VDD.n1321 VDD.t2145 75.3695
R9137 VDD.n1285 VDD.t2236 75.3695
R9138 VDD.n1297 VDD.t259 75.3695
R9139 VDD.n1237 VDD.t2242 75.3695
R9140 VDD.n1249 VDD.t535 75.3695
R9141 VDD.n1213 VDD.t2322 75.3695
R9142 VDD.n1225 VDD.t2356 75.3695
R9143 VDD.n1190 VDD.t514 75.3695
R9144 VDD.n685 VDD.n684 74.2572
R9145 VDD.n684 VDD.n671 74.2572
R9146 VDD.n1960 VDD.n1953 74.0005
R9147 VDD.n2336 VDD.n2329 74.0005
R9148 VDD.n2326 VDD.n2319 74.0005
R9149 VDD.n2316 VDD.n2309 74.0005
R9150 VDD.n2305 VDD.n2298 74.0005
R9151 VDD.n2295 VDD.n2288 74.0005
R9152 VDD.n2285 VDD.n2278 74.0005
R9153 VDD.n2275 VDD.n2268 74.0005
R9154 VDD.n1071 VDD.n1064 74.0005
R9155 VDD.n942 VDD.n935 74.0005
R9156 VDD.n813 VDD.n806 74.0005
R9157 VDD.n662 VDD.n655 74.0005
R9158 VDD.n533 VDD.n526 74.0005
R9159 VDD.n404 VDD.n397 74.0005
R9160 VDD.n275 VDD.n268 74.0005
R9161 VDD.n137 VDD.n130 74.0005
R9162 VDD.n2921 VDD.n2914 74.0005
R9163 VDD.n1200 VDD.t2229 73.2084
R9164 VDD.n1144 VDD.n1143 73.1255
R9165 VDD.n1142 VDD.n1141 73.1255
R9166 VDD.n1953 VDD.t1009 70.7977
R9167 VDD.n2329 VDD.t2337 70.7977
R9168 VDD.n2319 VDD.t2577 70.7977
R9169 VDD.n2309 VDD.t2128 70.7977
R9170 VDD.n2298 VDD.t3590 70.7977
R9171 VDD.n2288 VDD.t3983 70.7977
R9172 VDD.n2278 VDD.t3552 70.7977
R9173 VDD.n2268 VDD.t1400 70.7977
R9174 VDD.n1064 VDD.t34 70.7977
R9175 VDD.n935 VDD.t3922 70.7977
R9176 VDD.n806 VDD.t1481 70.7977
R9177 VDD.n655 VDD.t4299 70.7977
R9178 VDD.n526 VDD.t4255 70.7977
R9179 VDD.n397 VDD.t736 70.7977
R9180 VDD.n268 VDD.t2903 70.7977
R9181 VDD.n130 VDD.t4318 70.7977
R9182 VDD.n2914 VDD.t3510 70.7977
R9183 VDD.n2218 VDD.t1165 68.9949
R9184 VDD.n2243 VDD.t785 68.9949
R9185 VDD.n1884 VDD.t3484 68.9949
R9186 VDD.t1354 VDD.n1885 64.6005
R9187 VDD.n1876 VDD.t674 59.3755
R9188 VDD.n684 VDD.t2421 59.2645
R9189 VDD.n2189 VDD.n2188 53.374
R9190 VDD.n2081 VDD.n2080 53.374
R9191 VDD.n2747 VDD.t2411 52.7783
R9192 VDD.n2758 VDD.t2687 52.7783
R9193 VDD.n2769 VDD.t2856 52.7783
R9194 VDD.n2780 VDD.t2729 52.7783
R9195 VDD.n2791 VDD.t685 52.7783
R9196 VDD.n2802 VDD.t3987 52.7783
R9197 VDD.n2813 VDD.t1200 52.7783
R9198 VDD.n2824 VDD.t1644 52.7783
R9199 VDD.n1996 VDD.t971 52.7783
R9200 VDD.t3690 VDD.n1973 52.7783
R9201 VDD.n2846 VDD.t1097 52.7197
R9202 VDD.n2837 VDD.t1474 52.7197
R9203 VDD.n2847 VDD.t2106 52.7197
R9204 VDD.n2002 VDD.t1828 52.6613
R9205 VDD.n2011 VDD.t3291 52.6613
R9206 VDD.n2012 VDD.t4166 52.6613
R9207 VDD.n2022 VDD.t3452 52.6613
R9208 VDD.n2031 VDD.t1236 52.6613
R9209 VDD.n2032 VDD.t2457 52.6613
R9210 VDD.t367 VDD.n1383 52.141
R9211 VDD.n1384 VDD.t2650 52.141
R9212 VDD.t1152 VDD.n1792 52.141
R9213 VDD.n1802 VDD.t4163 52.141
R9214 VDD.n1801 VDD.t2270 52.141
R9215 VDD.n2364 VDD.t2427 52.141
R9216 VDD.n2363 VDD.t691 52.141
R9217 VDD.n2354 VDD.t744 52.141
R9218 VDD.n1669 VDD.t2733 52.141
R9219 VDD.n1668 VDD.t1536 52.141
R9220 VDD.n1659 VDD.t1242 52.141
R9221 VDD.n1650 VDD.t2023 52.141
R9222 VDD.n1641 VDD.t1615 52.141
R9223 VDD.n1632 VDD.t1313 52.141
R9224 VDD.n1447 VDD.t1549 52.141
R9225 VDD.n1446 VDD.t3454 52.141
R9226 VDD.t1041 VDD.n1564 52.141
R9227 VDD.t699 VDD.n1573 52.141
R9228 VDD.t1838 VDD.n1582 52.141
R9229 VDD.t3691 VDD.n1591 52.141
R9230 VDD.t1439 VDD.n1600 52.141
R9231 VDD.n1619 VDD.t732 52.141
R9232 VDD.n1618 VDD.t275 52.141
R9233 VDD.n1609 VDD.t2859 52.141
R9234 VDD.n2517 VDD.t3121 52.141
R9235 VDD.n2516 VDD.t581 52.141
R9236 VDD.n2507 VDD.t1543 52.141
R9237 VDD.n2498 VDD.t799 52.141
R9238 VDD.t1231 VDD.n2578 52.141
R9239 VDD.t1518 VDD.n2587 52.141
R9240 VDD.n2597 VDD.t1566 52.141
R9241 VDD.n2596 VDD.t1575 52.141
R9242 VDD.t1164 VDD.n2642 52.141
R9243 VDD.t3375 VDD.n2651 52.141
R9244 VDD.n2661 VDD.t140 52.141
R9245 VDD.n2660 VDD.t3899 52.141
R9246 VDD.t2648 VDD.n2718 52.141
R9247 VDD.t1196 VDD.n2727 52.141
R9248 VDD.t2488 VDD.n2736 52.141
R9249 VDD.n2737 VDD.t57 52.141
R9250 VDD.n2747 VDD.t3697 48.5561
R9251 VDD.n2758 VDD.t4278 48.5561
R9252 VDD.n2769 VDD.t1142 48.5561
R9253 VDD.n2780 VDD.t1613 48.5561
R9254 VDD.n2791 VDD.t1447 48.5561
R9255 VDD.n2802 VDD.t3958 48.5561
R9256 VDD.n2813 VDD.t3953 48.5561
R9257 VDD.n2824 VDD.t920 48.5561
R9258 VDD.n1996 VDD.t1596 48.5561
R9259 VDD.n1973 VDD.t1148 48.5561
R9260 VDD.t488 VDD.n2846 48.5022
R9261 VDD.t2771 VDD.n2837 48.5022
R9262 VDD.n2847 VDD.t55 48.5022
R9263 VDD.t2641 VDD.n2002 48.4484
R9264 VDD.t1819 VDD.n2011 48.4484
R9265 VDD.n2012 VDD.t629 48.4484
R9266 VDD.t2762 VDD.n2022 48.4484
R9267 VDD.t2416 VDD.n2031 48.4484
R9268 VDD.n2032 VDD.t1305 48.4484
R9269 VDD.n1383 VDD.t308 47.9698
R9270 VDD.n1384 VDD.t305 47.9698
R9271 VDD.n1792 VDD.t3342 47.9698
R9272 VDD.n1802 VDD.t1527 47.9698
R9273 VDD.t929 VDD.n1801 47.9698
R9274 VDD.n2364 VDD.t1853 47.9698
R9275 VDD.t2847 VDD.n2363 47.9698
R9276 VDD.t2036 VDD.n2354 47.9698
R9277 VDD.n1669 VDD.t905 47.9698
R9278 VDD.t2005 VDD.n1668 47.9698
R9279 VDD.t4307 VDD.n1659 47.9698
R9280 VDD.t1650 VDD.n1650 47.9698
R9281 VDD.t100 VDD.n1641 47.9698
R9282 VDD.t2858 VDD.n1632 47.9698
R9283 VDD.n1447 VDD.t2726 47.9698
R9284 VDD.t2430 VDD.n1446 47.9698
R9285 VDD.n1564 VDD.t1190 47.9698
R9286 VDD.n1573 VDD.t1347 47.9698
R9287 VDD.n1582 VDD.t2433 47.9698
R9288 VDD.n1591 VDD.t3622 47.9698
R9289 VDD.n1600 VDD.t61 47.9698
R9290 VDD.n1619 VDD.t3289 47.9698
R9291 VDD.t1344 VDD.n1618 47.9698
R9292 VDD.t2868 VDD.n1609 47.9698
R9293 VDD.n2517 VDD.t3378 47.9698
R9294 VDD.t1254 VDD.n2516 47.9698
R9295 VDD.t2267 VDD.n2507 47.9698
R9296 VDD.t3380 VDD.n2498 47.9698
R9297 VDD.n2578 VDD.t884 47.9698
R9298 VDD.n2587 VDD.t336 47.9698
R9299 VDD.n2597 VDD.t2184 47.9698
R9300 VDD.t953 VDD.n2596 47.9698
R9301 VDD.n2642 VDD.t773 47.9698
R9302 VDD.n2651 VDD.t558 47.9698
R9303 VDD.n2661 VDD.t1484 47.9698
R9304 VDD.t2047 VDD.n2660 47.9698
R9305 VDD.n2718 VDD.t1450 47.9698
R9306 VDD.n2727 VDD.t1217 47.9698
R9307 VDD.n2736 VDD.t1619 47.9698
R9308 VDD.n2737 VDD.t3880 47.9698
R9309 VDD.t676 VDD.t678 47.5005
R9310 VDD.n1134 VDD.n1133 47.413
R9311 VDD.n2396 VDD.n2395 47.413
R9312 VDD.n2402 VDD.n2401 47.413
R9313 VDD.n2409 VDD.n2408 47.413
R9314 VDD.n2378 VDD.n2377 47.413
R9315 VDD.n1947 VDD.n1946 47.413
R9316 VDD.n1945 VDD.n1944 47.413
R9317 VDD.n1938 VDD.n1937 47.413
R9318 VDD.n1928 VDD.n1927 47.413
R9319 VDD.n1926 VDD.n1925 47.413
R9320 VDD.n1919 VDD.n1918 47.413
R9321 VDD.n1910 VDD.n1909 47.413
R9322 VDD.n1899 VDD.n1898 47.413
R9323 VDD.n1309 VDD.n1308 47.413
R9324 VDD.n1321 VDD.n1320 47.413
R9325 VDD.n1285 VDD.n1284 47.413
R9326 VDD.n1297 VDD.n1296 47.413
R9327 VDD.n1261 VDD.n1260 47.413
R9328 VDD.n1273 VDD.n1272 47.413
R9329 VDD.n1237 VDD.n1236 47.413
R9330 VDD.n1249 VDD.n1248 47.413
R9331 VDD.n1213 VDD.n1212 47.413
R9332 VDD.n1225 VDD.n1224 47.413
R9333 VDD.n1200 VDD.n1199 47.413
R9334 VDD.n1191 VDD.n1190 47.413
R9335 VDD.n1739 VDD.n1738 47.413
R9336 VDD.n1749 VDD.n1748 47.413
R9337 VDD.n1849 VDD.n1848 47.413
R9338 VDD.n1839 VDD.n1838 47.413
R9339 VDD.n1824 VDD.n1823 47.413
R9340 VDD.n1423 VDD.n1422 47.413
R9341 VDD.n1684 VDD.n1683 47.413
R9342 VDD.n1691 VDD.n1690 47.413
R9343 VDD.n1700 VDD.n1699 47.413
R9344 VDD.n1698 VDD.n1697 47.413
R9345 VDD.n1817 VDD.n1816 47.413
R9346 VDD.n1826 VDD.n1825 47.413
R9347 VDD.n1837 VDD.n1836 47.413
R9348 VDD.n1851 VDD.n1850 47.413
R9349 VDD.n1491 VDD.n1490 47.413
R9350 VDD.n1498 VDD.n1497 47.413
R9351 VDD.n1522 VDD.n1521 47.413
R9352 VDD.n1474 VDD.n1473 47.413
R9353 VDD.n1555 VDD.n1554 47.413
R9354 VDD.n1553 VDD.n1552 47.413
R9355 VDD.n1546 VDD.n1545 47.413
R9356 VDD.n1539 VDD.n1538 47.413
R9357 VDD.n1529 VDD.n1528 47.413
R9358 VDD.n1515 VDD.n1514 47.413
R9359 VDD.n1505 VDD.n1504 47.413
R9360 VDD.n1481 VDD.n1480 47.413
R9361 VDD.n1397 VDD.n1396 47.413
R9362 VDD.n1399 VDD.n1398 47.413
R9363 VDD.n1713 VDD.n1712 47.413
R9364 VDD.n1720 VDD.n1719 47.413
R9365 VDD.n1779 VDD.n1778 47.413
R9366 VDD.n1777 VDD.n1776 47.413
R9367 VDD.n1770 VDD.n1769 47.413
R9368 VDD.n1763 VDD.n1762 47.413
R9369 VDD.n1751 VDD.n1750 47.413
R9370 VDD.n1737 VDD.n1736 47.413
R9371 VDD.n2530 VDD.n2529 47.413
R9372 VDD.n2479 VDD.n2478 47.413
R9373 VDD.n2477 VDD.n2476 47.413
R9374 VDD.n2532 VDD.n2531 47.413
R9375 VDD.n2542 VDD.n2541 47.413
R9376 VDD.n2546 VDD.n2545 47.413
R9377 VDD.n2566 VDD.n2565 47.413
R9378 VDD.n2564 VDD.n2563 47.413
R9379 VDD.n2560 VDD.n2559 47.413
R9380 VDD.n2553 VDD.n2552 47.413
R9381 VDD.n2606 VDD.n2605 47.413
R9382 VDD.n2610 VDD.n2609 47.413
R9383 VDD.n2630 VDD.n2629 47.413
R9384 VDD.n2628 VDD.n2627 47.413
R9385 VDD.n2624 VDD.n2623 47.413
R9386 VDD.n2617 VDD.n2616 47.413
R9387 VDD.n2670 VDD.n2669 47.413
R9388 VDD.n2674 VDD.n2673 47.413
R9389 VDD.n2706 VDD.n2705 47.413
R9390 VDD.n2704 VDD.n2703 47.413
R9391 VDD.n2697 VDD.n2696 47.413
R9392 VDD.n2688 VDD.n2687 47.413
R9393 VDD.n2686 VDD.n2685 47.413
R9394 VDD.n2526 VDD.n2525 47.413
R9395 VDD.n683 VDD.n682 47.413
R9396 VDD.t561 VDD.t560 46.7697
R9397 VDD.t562 VDD.t561 46.7697
R9398 VDD.t3167 VDD.t562 46.7697
R9399 VDD.t3168 VDD.t3167 46.7697
R9400 VDD.t3169 VDD.t3168 46.7697
R9401 VDD.t1529 VDD.t3169 46.7697
R9402 VDD.t1530 VDD.t1529 46.7697
R9403 VDD.t1528 VDD.t1530 46.7697
R9404 VDD.t2003 VDD.t1528 46.7697
R9405 VDD.t2001 VDD.t2003 46.7697
R9406 VDD.t2421 VDD.t2001 46.7697
R9407 VDD.n2229 VDD.t1011 39.9193
R9408 VDD.n2244 VDD.t311 39.9193
R9409 VDD.n1958 VDD.n1955 36.2404
R9410 VDD.n1959 VDD.n1958 36.2404
R9411 VDD.n2334 VDD.n2331 36.2404
R9412 VDD.n2335 VDD.n2334 36.2404
R9413 VDD.n2324 VDD.n2321 36.2404
R9414 VDD.n2325 VDD.n2324 36.2404
R9415 VDD.n2314 VDD.n2311 36.2404
R9416 VDD.n2315 VDD.n2314 36.2404
R9417 VDD.n2303 VDD.n2300 36.2404
R9418 VDD.n2304 VDD.n2303 36.2404
R9419 VDD.n2293 VDD.n2290 36.2404
R9420 VDD.n2294 VDD.n2293 36.2404
R9421 VDD.n2283 VDD.n2280 36.2404
R9422 VDD.n2284 VDD.n2283 36.2404
R9423 VDD.n2273 VDD.n2270 36.2404
R9424 VDD.n2274 VDD.n2273 36.2404
R9425 VDD.n1070 VDD.n1069 36.2404
R9426 VDD.n1069 VDD.n1066 36.2404
R9427 VDD.n941 VDD.n940 36.2404
R9428 VDD.n940 VDD.n937 36.2404
R9429 VDD.n812 VDD.n811 36.2404
R9430 VDD.n811 VDD.n808 36.2404
R9431 VDD.n661 VDD.n660 36.2404
R9432 VDD.n660 VDD.n657 36.2404
R9433 VDD.n532 VDD.n531 36.2404
R9434 VDD.n531 VDD.n528 36.2404
R9435 VDD.n403 VDD.n402 36.2404
R9436 VDD.n402 VDD.n399 36.2404
R9437 VDD.n274 VDD.n273 36.2404
R9438 VDD.n273 VDD.n270 36.2404
R9439 VDD.n136 VDD.n135 36.2404
R9440 VDD.n135 VDD.n132 36.2404
R9441 VDD.n2920 VDD.n2919 36.2404
R9442 VDD.n2919 VDD.n2916 36.2404
R9443 VDD.n1958 VDD.n1957 36.0299
R9444 VDD.n2334 VDD.n2333 36.0299
R9445 VDD.n2324 VDD.n2323 36.0299
R9446 VDD.n2314 VDD.n2313 36.0299
R9447 VDD.n2303 VDD.n2302 36.0299
R9448 VDD.n2293 VDD.n2292 36.0299
R9449 VDD.n2283 VDD.n2282 36.0299
R9450 VDD.n2273 VDD.n2272 36.0299
R9451 VDD.n1069 VDD.n1068 36.0299
R9452 VDD.n940 VDD.n939 36.0299
R9453 VDD.n811 VDD.n810 36.0299
R9454 VDD.n660 VDD.n659 36.0299
R9455 VDD.n531 VDD.n530 36.0299
R9456 VDD.n402 VDD.n401 36.0299
R9457 VDD.n273 VDD.n272 36.0299
R9458 VDD.n135 VDD.n134 36.0299
R9459 VDD.n2919 VDD.n2918 36.0299
R9460 VDD.t2347 VDD.t1013 31.8684
R9461 VDD.t2480 VDD.t315 31.8684
R9462 VDD.n1117 VDD 31.3918
R9463 VDD.n1026 VDD 31.3918
R9464 VDD.n1050 VDD 31.3918
R9465 VDD.n988 VDD 31.3918
R9466 VDD.n897 VDD 31.3918
R9467 VDD.n921 VDD 31.3918
R9468 VDD.n859 VDD 31.3918
R9469 VDD.n768 VDD 31.3918
R9470 VDD.n792 VDD 31.3918
R9471 VDD.n730 VDD 31.3918
R9472 VDD.n641 VDD 31.3918
R9473 VDD.n640 VDD 31.3918
R9474 VDD.n629 VDD 31.3918
R9475 VDD.n628 VDD 31.3918
R9476 VDD.n617 VDD 31.3918
R9477 VDD.n579 VDD 31.3918
R9478 VDD.n488 VDD 31.3918
R9479 VDD.n512 VDD 31.3918
R9480 VDD.n450 VDD 31.3918
R9481 VDD.n359 VDD 31.3918
R9482 VDD.n383 VDD 31.3918
R9483 VDD.n321 VDD 31.3918
R9484 VDD.n192 VDD 31.3918
R9485 VDD.n230 VDD 31.3918
R9486 VDD.n254 VDD 31.3918
R9487 VDD.n92 VDD 31.3918
R9488 VDD.n116 VDD 31.3918
R9489 VDD.n2897 VDD 31.3918
R9490 VDD.n30 VDD 31.3918
R9491 VDD.n54 VDD 31.3918
R9492 VDD.n1116 VDD 31.3373
R9493 VDD.n1105 VDD 31.3373
R9494 VDD.n1104 VDD 31.3373
R9495 VDD.n1093 VDD 31.3373
R9496 VDD.n987 VDD 31.3373
R9497 VDD.n976 VDD 31.3373
R9498 VDD.n975 VDD 31.3373
R9499 VDD.n964 VDD 31.3373
R9500 VDD.n858 VDD 31.3373
R9501 VDD.n847 VDD 31.3373
R9502 VDD.n846 VDD 31.3373
R9503 VDD.n835 VDD 31.3373
R9504 VDD.n729 VDD 31.3373
R9505 VDD.n718 VDD 31.3373
R9506 VDD.n717 VDD 31.3373
R9507 VDD.n706 VDD 31.3373
R9508 VDD.n578 VDD 31.3373
R9509 VDD.n567 VDD 31.3373
R9510 VDD.n566 VDD 31.3373
R9511 VDD.n555 VDD 31.3373
R9512 VDD.n449 VDD 31.3373
R9513 VDD.n438 VDD 31.3373
R9514 VDD.n437 VDD 31.3373
R9515 VDD.n426 VDD 31.3373
R9516 VDD.n320 VDD 31.3373
R9517 VDD.n309 VDD 31.3373
R9518 VDD.n308 VDD 31.3373
R9519 VDD.n297 VDD 31.3373
R9520 VDD.n191 VDD 31.3373
R9521 VDD.n180 VDD 31.3373
R9522 VDD.n179 VDD 31.3373
R9523 VDD.n168 VDD 31.3373
R9524 VDD.n2896 VDD 31.3373
R9525 VDD.n2885 VDD 31.3373
R9526 VDD.n2884 VDD 31.3373
R9527 VDD.n2873 VDD 31.3373
R9528 VDD.n1049 VDD 31.283
R9529 VDD.n1038 VDD 31.283
R9530 VDD.n1037 VDD 31.283
R9531 VDD.n920 VDD 31.283
R9532 VDD.n909 VDD 31.283
R9533 VDD.n908 VDD 31.283
R9534 VDD.n791 VDD 31.283
R9535 VDD.n780 VDD 31.283
R9536 VDD.n779 VDD 31.283
R9537 VDD.n511 VDD 31.283
R9538 VDD.n500 VDD 31.283
R9539 VDD.n499 VDD 31.283
R9540 VDD.n382 VDD 31.283
R9541 VDD.n371 VDD 31.283
R9542 VDD.n370 VDD 31.283
R9543 VDD.n253 VDD 31.283
R9544 VDD.n242 VDD 31.283
R9545 VDD.n241 VDD 31.283
R9546 VDD.n115 VDD 31.283
R9547 VDD.n104 VDD 31.283
R9548 VDD.n103 VDD 31.283
R9549 VDD.n53 VDD 31.283
R9550 VDD.n42 VDD 31.283
R9551 VDD.n41 VDD 31.283
R9552 VDD.n1885 VDD.t676 30.6776
R9553 VDD.n1131 VDD.t4127 30.379
R9554 VDD.n1131 VDD.t4129 30.379
R9555 VDD.n1127 VDD.t2272 30.379
R9556 VDD.n1127 VDD.t2274 30.379
R9557 VDD.n1129 VDD.t3501 30.379
R9558 VDD.n1129 VDD.t3499 30.379
R9559 VDD.n2527 VDD.t1363 30.379
R9560 VDD.n2527 VDD.t1361 30.379
R9561 VDD.n2462 VDD.t2540 30.379
R9562 VDD.n2462 VDD.t2538 30.379
R9563 VDD.n2533 VDD.t804 30.379
R9564 VDD.n2533 VDD.t802 30.379
R9565 VDD.n2465 VDD.t753 30.379
R9566 VDD.n2465 VDD.t751 30.379
R9567 VDD.n2539 VDD.t4137 30.379
R9568 VDD.n2539 VDD.t4135 30.379
R9569 VDD.n2459 VDD.t4205 30.379
R9570 VDD.n2459 VDD.t4203 30.379
R9571 VDD.n2689 VDD.t1879 30.379
R9572 VDD.n2689 VDD.t1881 30.379
R9573 VDD.n2678 VDD.t3474 30.379
R9574 VDD.n2678 VDD.t3480 30.379
R9575 VDD.n2694 VDD.t2691 30.379
R9576 VDD.n2694 VDD.t2695 30.379
R9577 VDD.n2675 VDD.t1845 30.379
R9578 VDD.n2675 VDD.t1843 30.379
R9579 VDD.n2683 VDD.t3644 30.379
R9580 VDD.n2683 VDD.t3650 30.379
R9581 VDD.n2680 VDD.t3431 30.379
R9582 VDD.n2680 VDD.t3437 30.379
R9583 VDD.n2707 VDD.t1118 30.379
R9584 VDD.n2707 VDD.t1122 30.379
R9585 VDD.n2417 VDD.t2402 30.379
R9586 VDD.n2417 VDD.t2408 30.379
R9587 VDD.n2671 VDD.t1583 30.379
R9588 VDD.n2671 VDD.t1587 30.379
R9589 VDD.n2414 VDD.t2477 30.379
R9590 VDD.n2414 VDD.t2475 30.379
R9591 VDD.n2701 VDD.t3239 30.379
R9592 VDD.n2701 VDD.t3243 30.379
R9593 VDD.n2698 VDD.t2842 30.379
R9594 VDD.n2698 VDD.t2840 30.379
R9595 VDD.n2397 VDD.t1205 30.379
R9596 VDD.n2397 VDD.t1158 30.379
R9597 VDD.n2393 VDD.t594 30.379
R9598 VDD.n2393 VDD.t1016 30.379
R9599 VDD.n2390 VDD.t4086 30.379
R9600 VDD.n2390 VDD.t4092 30.379
R9601 VDD.n2383 VDD.t237 30.379
R9602 VDD.n2383 VDD.t238 30.379
R9603 VDD.n2388 VDD.t996 30.379
R9604 VDD.n2388 VDD.t1003 30.379
R9605 VDD.n2386 VDD.t264 30.379
R9606 VDD.n2386 VDD.t518 30.379
R9607 VDD.n2379 VDD.t1058 30.379
R9608 VDD.n2379 VDD.t1059 30.379
R9609 VDD.n1167 VDD.t1035 30.379
R9610 VDD.n1167 VDD.t584 30.379
R9611 VDD.n1165 VDD.t4213 30.379
R9612 VDD.n1165 VDD.t4229 30.379
R9613 VDD.n2369 VDD.t164 30.379
R9614 VDD.n2369 VDD.t165 30.379
R9615 VDD.n2375 VDD.t992 30.379
R9616 VDD.n2375 VDD.t1000 30.379
R9617 VDD.n1169 VDD.t2241 30.379
R9618 VDD.n1169 VDD.t1666 30.379
R9619 VDD.n2200 VDD.t2344 30.379
R9620 VDD.n2200 VDD.t2348 30.379
R9621 VDD.n2202 VDD.t2582 30.379
R9622 VDD.n2202 VDD.t2600 30.379
R9623 VDD.n2211 VDD.t2121 30.379
R9624 VDD.n2211 VDD.t2140 30.379
R9625 VDD.n2205 VDD.t3611 30.379
R9626 VDD.n2205 VDD.t3594 30.379
R9627 VDD.n2208 VDD.t3971 30.379
R9628 VDD.n2208 VDD.t888 30.379
R9629 VDD.n2215 VDD.t1168 30.379
R9630 VDD.n2215 VDD.t1394 30.379
R9631 VDD.n2213 VDD.t3546 30.379
R9632 VDD.n2213 VDD.t3561 30.379
R9633 VDD.n2225 VDD.t1014 30.379
R9634 VDD.n2225 VDD.t1039 30.379
R9635 VDD.n2122 VDD.t1036 30.379
R9636 VDD.n2122 VDD.t1008 30.379
R9637 VDD.n2120 VDD.t1238 30.379
R9638 VDD.n2120 VDD.t1240 30.379
R9639 VDD.n2125 VDD.t2355 30.379
R9640 VDD.n2125 VDD.t2330 30.379
R9641 VDD.n2181 VDD.t3264 30.379
R9642 VDD.n2181 VDD.t3263 30.379
R9643 VDD.n2128 VDD.t2587 30.379
R9644 VDD.n2128 VDD.t468 30.379
R9645 VDD.n2151 VDD.t1184 30.379
R9646 VDD.n2151 VDD.t1186 30.379
R9647 VDD.n2131 VDD.t2182 30.379
R9648 VDD.n2131 VDD.t2150 30.379
R9649 VDD.n2172 VDD.t2553 30.379
R9650 VDD.n2172 VDD.t2552 30.379
R9651 VDD.n2134 VDD.t3595 30.379
R9652 VDD.n2134 VDD.t3617 30.379
R9653 VDD.n2167 VDD.t1197 30.379
R9654 VDD.n2167 VDD.t2063 30.379
R9655 VDD.n2137 VDD.t3976 30.379
R9656 VDD.n2137 VDD.t901 30.379
R9657 VDD.n2162 VDD.t817 30.379
R9658 VDD.n2162 VDD.t816 30.379
R9659 VDD.n2140 VDD.t3547 30.379
R9660 VDD.n2140 VDD.t3528 30.379
R9661 VDD.n2157 VDD.t1312 30.379
R9662 VDD.n2157 VDD.t1311 30.379
R9663 VDD.n2143 VDD.t1395 30.379
R9664 VDD.n2143 VDD.t1169 30.379
R9665 VDD.n2153 VDD.t136 30.379
R9666 VDD.n2153 VDD.t1206 30.379
R9667 VDD.n2186 VDD.t3112 30.379
R9668 VDD.n2186 VDD.t3114 30.379
R9669 VDD.n2042 VDD.t1704 30.379
R9670 VDD.n2042 VDD.t1702 30.379
R9671 VDD.n2040 VDD.t1029 30.379
R9672 VDD.n2040 VDD.t1023 30.379
R9673 VDD.n2047 VDD.t366 30.379
R9674 VDD.n2047 VDD.t362 30.379
R9675 VDD.n2051 VDD.t2332 30.379
R9676 VDD.n2051 VDD.t2329 30.379
R9677 VDD.n2082 VDD.t2000 30.379
R9678 VDD.n2082 VDD.t1998 30.379
R9679 VDD.n2055 VDD.t478 30.379
R9680 VDD.n2055 VDD.t466 30.379
R9681 VDD.n2087 VDD.t2496 30.379
R9682 VDD.n2087 VDD.t2494 30.379
R9683 VDD.n2059 VDD.t2165 30.379
R9684 VDD.n2059 VDD.t2159 30.379
R9685 VDD.n2092 VDD.t747 30.379
R9686 VDD.n2092 VDD.t800 30.379
R9687 VDD.n2063 VDD.t3589 30.379
R9688 VDD.n2063 VDD.t3581 30.379
R9689 VDD.n2097 VDD.t682 30.379
R9690 VDD.n2097 VDD.t680 30.379
R9691 VDD.n2067 VDD.t3963 30.379
R9692 VDD.n2067 VDD.t900 30.379
R9693 VDD.n2102 VDD.t3493 30.379
R9694 VDD.n2102 VDD.t3491 30.379
R9695 VDD.n2071 VDD.t3532 30.379
R9696 VDD.n2071 VDD.t3527 30.379
R9697 VDD.n2107 VDD.t1189 30.379
R9698 VDD.n2107 VDD.t1187 30.379
R9699 VDD.n2075 VDD.t1390 30.379
R9700 VDD.n2075 VDD.t1388 30.379
R9701 VDD.n2078 VDD.t3106 30.379
R9702 VDD.n2078 VDD.t3110 30.379
R9703 VDD.n2245 VDD.t316 30.379
R9704 VDD.n2245 VDD.t314 30.379
R9705 VDD.n2253 VDD.t2483 30.379
R9706 VDD.n2253 VDD.t2481 30.379
R9707 VDD.n2248 VDD.t1547 30.379
R9708 VDD.n2248 VDD.t1546 30.379
R9709 VDD.n2251 VDD.t729 30.379
R9710 VDD.n2251 VDD.t731 30.379
R9711 VDD.n2235 VDD.t2279 30.379
R9712 VDD.n2235 VDD.t2278 30.379
R9713 VDD.n2237 VDD.t790 30.379
R9714 VDD.n2237 VDD.t788 30.379
R9715 VDD.n2240 VDD.t320 30.379
R9716 VDD.n2240 VDD.t318 30.379
R9717 VDD.n2260 VDD.t371 30.379
R9718 VDD.n2260 VDD.t370 30.379
R9719 VDD.n1892 VDD.t4189 30.379
R9720 VDD.n1892 VDD.t4209 30.379
R9721 VDD.n1894 VDD.t2365 30.379
R9722 VDD.n1894 VDD.t2371 30.379
R9723 VDD.n1939 VDD.t520 30.379
R9724 VDD.n1939 VDD.t532 30.379
R9725 VDD.n1941 VDD.t482 30.379
R9726 VDD.n1941 VDD.t486 30.379
R9727 VDD.n1900 VDD.t4067 30.379
R9728 VDD.n1900 VDD.t4071 30.379
R9729 VDD.n1934 VDD.t2158 30.379
R9730 VDD.n1934 VDD.t2163 30.379
R9731 VDD.n1903 VDD.t1641 30.379
R9732 VDD.n1903 VDD.t2198 30.379
R9733 VDD.n1929 VDD.t3601 30.379
R9734 VDD.n1929 VDD.t3614 30.379
R9735 VDD.n1920 VDD.t382 30.379
R9736 VDD.n1920 VDD.t394 30.379
R9737 VDD.n1922 VDD.t904 30.379
R9738 VDD.n1922 VDD.t3975 30.379
R9739 VDD.n1905 VDD.t2833 30.379
R9740 VDD.n1905 VDD.t2820 30.379
R9741 VDD.n1915 VDD.t3544 30.379
R9742 VDD.n1915 VDD.t3557 30.379
R9743 VDD.n1907 VDD.t3420 30.379
R9744 VDD.n1907 VDD.t3435 30.379
R9745 VDD.n1911 VDD.t1415 30.379
R9746 VDD.n1911 VDD.t1179 30.379
R9747 VDD.n1896 VDD.t2239 30.379
R9748 VDD.n1896 VDD.t1662 30.379
R9749 VDD.n1888 VDD.t998 30.379
R9750 VDD.n1888 VDD.t1020 30.379
R9751 VDD.n1871 VDD.t3483 30.379
R9752 VDD.n1871 VDD.t3482 30.379
R9753 VDD.n1865 VDD.t2384 30.379
R9754 VDD.n1865 VDD.t2386 30.379
R9755 VDD.n1868 VDD.t679 30.379
R9756 VDD.n1868 VDD.t677 30.379
R9757 VDD.n1863 VDD.t2638 30.379
R9758 VDD.n1863 VDD.t2637 30.379
R9759 VDD.n1855 VDD.t1353 30.379
R9760 VDD.n1855 VDD.t1357 30.379
R9761 VDD.n1857 VDD.t829 30.379
R9762 VDD.n1857 VDD.t827 30.379
R9763 VDD.n1879 VDD.t1572 30.379
R9764 VDD.n1879 VDD.t1570 30.379
R9765 VDD.n1860 VDD.t3489 30.379
R9766 VDD.n1860 VDD.t3487 30.379
R9767 VDD.n1310 VDD.t3932 30.379
R9768 VDD.n1310 VDD.t3933 30.379
R9769 VDD.n1306 VDD.t2139 30.379
R9770 VDD.n1306 VDD.t2179 30.379
R9771 VDD.n1303 VDD.t4220 30.379
R9772 VDD.n1303 VDD.t4242 30.379
R9773 VDD.n1322 VDD.t2685 30.379
R9774 VDD.n1322 VDD.t2686 30.379
R9775 VDD.n1318 VDD.t2146 30.379
R9776 VDD.n1318 VDD.t2142 30.379
R9777 VDD.n1315 VDD.t4108 30.379
R9778 VDD.n1315 VDD.t4080 30.379
R9779 VDD.n1286 VDD.t727 30.379
R9780 VDD.n1286 VDD.t728 30.379
R9781 VDD.n1282 VDD.t2237 30.379
R9782 VDD.n1282 VDD.t1682 30.379
R9783 VDD.n1279 VDD.t2177 30.379
R9784 VDD.n1279 VDD.t2135 30.379
R9785 VDD.n1298 VDD.t2635 30.379
R9786 VDD.n1298 VDD.t2633 30.379
R9787 VDD.n1294 VDD.t260 30.379
R9788 VDD.n1294 VDD.t556 30.379
R9789 VDD.n1291 VDD.t2171 30.379
R9790 VDD.n1291 VDD.t2144 30.379
R9791 VDD.n1262 VDD.t2078 30.379
R9792 VDD.n1262 VDD.t2079 30.379
R9793 VDD.n1258 VDD.t2584 30.379
R9794 VDD.n1258 VDD.t2602 30.379
R9795 VDD.n1255 VDD.t4193 30.379
R9796 VDD.n1255 VDD.t4191 30.379
R9797 VDD.n1274 VDD.t4324 30.379
R9798 VDD.n1274 VDD.t4274 30.379
R9799 VDD.n1270 VDD.t464 30.379
R9800 VDD.n1270 VDD.t474 30.379
R9801 VDD.n1267 VDD.t4094 30.379
R9802 VDD.n1267 VDD.t4114 30.379
R9803 VDD.n1238 VDD.t1088 30.379
R9804 VDD.n1238 VDD.t1089 30.379
R9805 VDD.n1234 VDD.t2243 30.379
R9806 VDD.n1234 VDD.t1668 30.379
R9807 VDD.n1231 VDD.t472 30.379
R9808 VDD.n1231 VDD.t470 30.379
R9809 VDD.n1250 VDD.t813 30.379
R9810 VDD.n1250 VDD.t814 30.379
R9811 VDD.n1246 VDD.t536 30.379
R9812 VDD.n1246 VDD.t544 30.379
R9813 VDD.n1243 VDD.t2591 30.379
R9814 VDD.n1243 VDD.t2614 30.379
R9815 VDD.n1214 VDD.t3148 30.379
R9816 VDD.n1214 VDD.t3149 30.379
R9817 VDD.n1210 VDD.t2323 30.379
R9818 VDD.n1210 VDD.t2350 30.379
R9819 VDD.n1207 VDD.t4238 30.379
R9820 VDD.n1207 VDD.t4236 30.379
R9821 VDD.n1226 VDD.t2623 30.379
R9822 VDD.n1226 VDD.t2621 30.379
R9823 VDD.n1222 VDD.t2357 30.379
R9824 VDD.n1222 VDD.t2367 30.379
R9825 VDD.n1219 VDD.t4076 30.379
R9826 VDD.n1219 VDD.t4104 30.379
R9827 VDD.n1201 VDD.t1127 30.379
R9828 VDD.n1201 VDD.t1128 30.379
R9829 VDD.n1197 VDD.t2230 30.379
R9830 VDD.n1197 VDD.t1656 30.379
R9831 VDD.n1194 VDD.t2361 30.379
R9832 VDD.n1194 VDD.t2359 30.379
R9833 VDD.n1183 VDD.t441 30.379
R9834 VDD.n1183 VDD.t442 30.379
R9835 VDD.n1188 VDD.t515 30.379
R9836 VDD.n1188 VDD.t522 30.379
R9837 VDD.n1186 VDD.t2375 30.379
R9838 VDD.n1186 VDD.t2328 30.379
R9839 VDD.n1729 VDD.t2738 30.379
R9840 VDD.n1729 VDD.t2740 30.379
R9841 VDD.n1740 VDD.t2566 30.379
R9842 VDD.n1740 VDD.t2564 30.379
R9843 VDD.n1746 VDD.t4326 30.379
R9844 VDD.n1746 VDD.t4328 30.379
R9845 VDD.n1725 VDD.t721 30.379
R9846 VDD.n1725 VDD.t719 30.379
R9847 VDD.n1394 VDD.t2249 30.379
R9848 VDD.n1394 VDD.t2426 30.379
R9849 VDD.n1389 VDD.t224 30.379
R9850 VDD.n1389 VDD.t226 30.379
R9851 VDD.n1400 VDD.t1981 30.379
R9852 VDD.n1400 VDD.t1979 30.379
R9853 VDD.n1392 VDD.t1604 30.379
R9854 VDD.n1392 VDD.t2053 30.379
R9855 VDD.n1710 VDD.t294 30.379
R9856 VDD.n1710 VDD.t296 30.379
R9857 VDD.n1367 VDD.t1296 30.379
R9858 VDD.n1367 VDD.t1300 30.379
R9859 VDD.n1780 VDD.t220 30.379
R9860 VDD.n1780 VDD.t210 30.379
R9861 VDD.n1365 VDD.t4174 30.379
R9862 VDD.n1365 VDD.t4176 30.379
R9863 VDD.n1717 VDD.t2516 30.379
R9864 VDD.n1717 VDD.t2518 30.379
R9865 VDD.n1714 VDD.t715 30.379
R9866 VDD.n1714 VDD.t717 30.379
R9867 VDD.n1774 VDD.t1331 30.379
R9868 VDD.n1774 VDD.t1335 30.379
R9869 VDD.n1771 VDD.t2303 30.379
R9870 VDD.n1771 VDD.t2305 30.379
R9871 VDD.n1758 VDD.t703 30.379
R9872 VDD.n1758 VDD.t707 30.379
R9873 VDD.n1760 VDD.t460 30.379
R9874 VDD.n1760 VDD.t462 30.379
R9875 VDD.n1767 VDD.t1085 30.379
R9876 VDD.n1767 VDD.t564 30.379
R9877 VDD.n1764 VDD.t1130 30.379
R9878 VDD.n1764 VDD.t1132 30.379
R9879 VDD.n1723 VDD.t2916 30.379
R9880 VDD.n1723 VDD.t2914 30.379
R9881 VDD.n1721 VDD.t248 30.379
R9882 VDD.n1721 VDD.t254 30.379
R9883 VDD.n1846 VDD.t3664 30.379
R9884 VDD.n1846 VDD.t3662 30.379
R9885 VDD.n1844 VDD.t943 30.379
R9886 VDD.n1844 VDD.t947 30.379
R9887 VDD.n1334 VDD.t970 30.379
R9888 VDD.n1334 VDD.t968 30.379
R9889 VDD.n1332 VDD.t2071 30.379
R9890 VDD.n1332 VDD.t2073 30.379
R9891 VDD.n1821 VDD.t1467 30.379
R9892 VDD.n1821 VDD.t1469 30.379
R9893 VDD.n1818 VDD.t1694 30.379
R9894 VDD.n1818 VDD.t1698 30.379
R9895 VDD.n1827 VDD.t835 30.379
R9896 VDD.n1827 VDD.t843 30.379
R9897 VDD.n1340 VDD.t1286 30.379
R9898 VDD.n1340 VDD.t1282 30.379
R9899 VDD.n1834 VDD.t155 30.379
R9900 VDD.n1834 VDD.t159 30.379
R9901 VDD.n1336 VDD.t2442 30.379
R9902 VDD.n1336 VDD.t2438 30.379
R9903 VDD.n1420 VDD.t867 30.379
R9904 VDD.n1420 VDD.t871 30.379
R9905 VDD.n1418 VDD.t2103 30.379
R9906 VDD.n1418 VDD.t2101 30.379
R9907 VDD.n1679 VDD.t1931 30.379
R9908 VDD.n1679 VDD.t1943 30.379
R9909 VDD.n1681 VDD.t3386 30.379
R9910 VDD.n1681 VDD.t3384 30.379
R9911 VDD.n1688 VDD.t1887 30.379
R9912 VDD.n1688 VDD.t1079 30.379
R9913 VDD.n1685 VDD.t3521 30.379
R9914 VDD.n1685 VDD.t3517 30.379
R9915 VDD.n1693 VDD.t2783 30.379
R9916 VDD.n1693 VDD.t2779 30.379
R9917 VDD.n1695 VDD.t2013 30.379
R9918 VDD.n1695 VDD.t2011 30.379
R9919 VDD.n1416 VDD.t3408 30.379
R9920 VDD.n1416 VDD.t3412 30.379
R9921 VDD.n1414 VDD.t4003 30.379
R9922 VDD.n1414 VDD.t4001 30.379
R9923 VDD.n1814 VDD.t1901 30.379
R9924 VDD.n1814 VDD.t1895 30.379
R9925 VDD.n1342 VDD.t4007 30.379
R9926 VDD.n1342 VDD.t4017 30.379
R9927 VDD.n1329 VDD.t4059 30.379
R9928 VDD.n1329 VDD.t4057 30.379
R9929 VDD.n1327 VDD.t3321 30.379
R9930 VDD.n1327 VDD.t3315 30.379
R9931 VDD.n1488 VDD.t1049 30.379
R9932 VDD.n1488 VDD.t1051 30.379
R9933 VDD.n1486 VDD.t4155 30.379
R9934 VDD.n1486 VDD.t4153 30.379
R9935 VDD.n1495 VDD.t145 30.379
R9936 VDD.n1495 VDD.t147 30.379
R9937 VDD.n1492 VDD.t572 30.379
R9938 VDD.n1492 VDD.t576 30.379
R9939 VDD.n1519 VDD.t4045 30.379
R9940 VDD.n1519 VDD.t4047 30.379
R9941 VDD.n1516 VDD.t4039 30.379
R9942 VDD.n1516 VDD.t4043 30.379
R9943 VDD.n1510 VDD.t3674 30.379
R9944 VDD.n1510 VDD.t3678 30.379
R9945 VDD.n1512 VDD.t661 30.379
R9946 VDD.n1512 VDD.t663 30.379
R9947 VDD.n1502 VDD.t4027 30.379
R9948 VDD.n1502 VDD.t4025 30.379
R9949 VDD.n1499 VDD.t25 30.379
R9950 VDD.n1499 VDD.t31 30.379
R9951 VDD.n1471 VDD.t2218 30.379
R9952 VDD.n1471 VDD.t2214 30.379
R9953 VDD.n1466 VDD.t2744 30.379
R9954 VDD.n1466 VDD.t2746 30.379
R9955 VDD.n1556 VDD.t1957 30.379
R9956 VDD.n1556 VDD.t1953 30.379
R9957 VDD.n1469 VDD.t602 30.379
R9958 VDD.n1469 VDD.t1589 30.379
R9959 VDD.n1550 VDD.t2498 30.379
R9960 VDD.n1550 VDD.t2500 30.379
R9961 VDD.n1547 VDD.t3195 30.379
R9962 VDD.n1547 VDD.t3187 30.379
R9963 VDD.n1534 VDD.t4280 30.379
R9964 VDD.n1534 VDD.t4286 30.379
R9965 VDD.n1536 VDD.t3888 30.379
R9966 VDD.n1536 VDD.t3890 30.379
R9967 VDD.n1543 VDD.t4266 30.379
R9968 VDD.n1543 VDD.t4268 30.379
R9969 VDD.n1540 VDD.t3684 30.379
R9970 VDD.n1540 VDD.t3686 30.379
R9971 VDD.n1526 VDD.t3270 30.379
R9972 VDD.n1526 VDD.t3274 30.379
R9973 VDD.n1523 VDD.t106 30.379
R9974 VDD.n1523 VDD.t108 30.379
R9975 VDD.n1478 VDD.t2725 30.379
R9976 VDD.n1478 VDD.t2713 30.379
R9977 VDD.n1475 VDD.t4250 30.379
R9978 VDD.n1475 VDD.t3937 30.379
R9979 VDD.n1734 VDD.t1933 30.379
R9980 VDD.n1734 VDD.t1927 30.379
R9981 VDD.n1731 VDD.t637 30.379
R9982 VDD.n1731 VDD.t1606 30.379
R9983 VDD.n2612 VDD.t2761 30.379
R9984 VDD.n2612 VDD.t2759 30.379
R9985 VDD.n2614 VDD.t3907 30.379
R9986 VDD.n2614 VDD.t3911 30.379
R9987 VDD.n2621 VDD.t1852 30.379
R9988 VDD.n2621 VDD.t1850 30.379
R9989 VDD.n2618 VDD.t2705 30.379
R9990 VDD.n2618 VDD.t2703 30.379
R9991 VDD.n2667 VDD.t2879 30.379
R9992 VDD.n2667 VDD.t2883 30.379
R9993 VDD.n2419 VDD.t408 30.379
R9994 VDD.n2419 VDD.t406 30.379
R9995 VDD.n2631 VDD.t3945 30.379
R9996 VDD.n2631 VDD.t3943 30.379
R9997 VDD.n2437 VDD.t298 30.379
R9998 VDD.n2437 VDD.t302 30.379
R9999 VDD.n2607 VDD.t3999 30.379
R10000 VDD.n2607 VDD.t3997 30.379
R10001 VDD.n2434 VDD.t3465 30.379
R10002 VDD.n2434 VDD.t3463 30.379
R10003 VDD.n2625 VDD.t1432 30.379
R10004 VDD.n2625 VDD.t1434 30.379
R10005 VDD.n2431 VDD.t1630 30.379
R10006 VDD.n2431 VDD.t1628 30.379
R10007 VDD.n2548 VDD.t1738 30.379
R10008 VDD.n2548 VDD.t1736 30.379
R10009 VDD.n2550 VDD.t1559 30.379
R10010 VDD.n2550 VDD.t1561 30.379
R10011 VDD.n2557 VDD.t1857 30.379
R10012 VDD.n2557 VDD.t1855 30.379
R10013 VDD.n2554 VDD.t2188 30.379
R10014 VDD.n2554 VDD.t2186 30.379
R10015 VDD.n2603 VDD.t616 30.379
R10016 VDD.n2603 VDD.t614 30.379
R10017 VDD.n2439 VDD.t4110 30.379
R10018 VDD.n2439 VDD.t4097 30.379
R10019 VDD.n2567 VDD.t85 30.379
R10020 VDD.n2567 VDD.t83 30.379
R10021 VDD.n2457 VDD.t2471 30.379
R10022 VDD.n2457 VDD.t2469 30.379
R10023 VDD.n2543 VDD.t3329 30.379
R10024 VDD.n2543 VDD.t3327 30.379
R10025 VDD.n2454 VDD.t446 30.379
R10026 VDD.n2454 VDD.t444 30.379
R10027 VDD.n2561 VDD.t344 30.379
R10028 VDD.n2561 VDD.t342 30.379
R10029 VDD.n2451 VDD.t546 30.379
R10030 VDD.n2451 VDD.t542 30.379
R10031 VDD.n2472 VDD.t2255 30.379
R10032 VDD.n2472 VDD.t2253 30.379
R10033 VDD.n2480 VDD.t1770 30.379
R10034 VDD.n2480 VDD.t1762 30.379
R10035 VDD.n2474 VDD.t3404 30.379
R10036 VDD.n2474 VDD.t3406 30.379
R10037 VDD.n2469 VDD.t1827 30.379
R10038 VDD.n2469 VDD.t1823 30.379
R10039 VDD.n2523 VDD.t2093 30.379
R10040 VDD.n2523 VDD.t2091 30.379
R10041 VDD.n2467 VDD.t2222 30.379
R10042 VDD.n2467 VDD.t2220 30.379
R10043 VDD.n1015 VDD.t3777 30.379
R10044 VDD.n1015 VDD.t3782 30.379
R10045 VDD.n1013 VDD.t4354 30.379
R10046 VDD.n1013 VDD.t4366 30.379
R10047 VDD.n1010 VDD.t3082 30.379
R10048 VDD.n1010 VDD.t3071 30.379
R10049 VDD.n1057 VDD.t1524 30.379
R10050 VDD.n1057 VDD.t1520 30.379
R10051 VDD.n886 VDD.t3795 30.379
R10052 VDD.n886 VDD.t3879 30.379
R10053 VDD.n884 VDD.t4380 30.379
R10054 VDD.n884 VDD.t4443 30.379
R10055 VDD.n881 VDD.t3060 30.379
R10056 VDD.n881 VDD.t3002 30.379
R10057 VDD.n928 VDD.t3917 30.379
R10058 VDD.n928 VDD.t3919 30.379
R10059 VDD.n757 VDD.t3798 30.379
R10060 VDD.n757 VDD.t3876 30.379
R10061 VDD.n755 VDD.t4456 30.379
R10062 VDD.n755 VDD.t4505 30.379
R10063 VDD.n752 VDD.t3093 30.379
R10064 VDD.n752 VDD.t3027 30.379
R10065 VDD.n799 VDD.t3461 30.379
R10066 VDD.n799 VDD.t3457 30.379
R10067 VDD.n606 VDD.t3723 30.379
R10068 VDD.n606 VDD.t3769 30.379
R10069 VDD.n604 VDD.t4356 30.379
R10070 VDD.n604 VDD.t4438 30.379
R10071 VDD.n601 VDD.t3003 30.379
R10072 VDD.n601 VDD.t2938 30.379
R10073 VDD.n648 VDD.t3346 30.379
R10074 VDD.n648 VDD.t1317 30.379
R10075 VDD.n477 VDD.t3752 30.379
R10076 VDD.n477 VDD.t3757 30.379
R10077 VDD.n475 VDD.t4421 30.379
R10078 VDD.n475 VDD.t4426 30.379
R10079 VDD.n472 VDD.t2965 30.379
R10080 VDD.n472 VDD.t2952 30.379
R10081 VDD.n519 VDD.t2544 30.379
R10082 VDD.n519 VDD.t2546 30.379
R10083 VDD.n348 VDD.t3725 30.379
R10084 VDD.n348 VDD.t3737 30.379
R10085 VDD.n346 VDD.t4358 30.379
R10086 VDD.n346 VDD.t4379 30.379
R10087 VDD.n343 VDD.t3000 30.379
R10088 VDD.n343 VDD.t2989 30.379
R10089 VDD.n390 VDD.t2711 30.379
R10090 VDD.n390 VDD.t2707 30.379
R10091 VDD.n219 VDD.t3726 30.379
R10092 VDD.n219 VDD.t3758 30.379
R10093 VDD.n217 VDD.t4359 30.379
R10094 VDD.n217 VDD.t4431 30.379
R10095 VDD.n214 VDD.t2999 30.379
R10096 VDD.n214 VDD.t2950 30.379
R10097 VDD.n261 VDD.t1690 30.379
R10098 VDD.n261 VDD.t1692 30.379
R10099 VDD.n145 VDD.t1135 30.379
R10100 VDD.n145 VDD.t1136 30.379
R10101 VDD.n142 VDD.t1091 30.379
R10102 VDD.n142 VDD.t1093 30.379
R10103 VDD.n679 VDD.t196 30.379
R10104 VDD.n679 VDD.t1821 30.379
R10105 VDD.n677 VDD.t2390 30.379
R10106 VDD.n677 VDD.t2392 30.379
R10107 VDD.n672 VDD.t1461 30.379
R10108 VDD.n672 VDD.t1463 30.379
R10109 VDD.n81 VDD.t3766 30.379
R10110 VDD.n81 VDD.t3774 30.379
R10111 VDD.n79 VDD.t4462 30.379
R10112 VDD.n79 VDD.t4471 30.379
R10113 VDD.n76 VDD.t3053 30.379
R10114 VDD.n76 VDD.t3050 30.379
R10115 VDD.n123 VDD.t1100 30.379
R10116 VDD.n123 VDD.t1102 30.379
R10117 VDD.n19 VDD.t3728 30.379
R10118 VDD.n19 VDD.t3837 30.379
R10119 VDD.n17 VDD.t4406 30.379
R10120 VDD.n17 VDD.t4514 30.379
R10121 VDD.n14 VDD.t2944 30.379
R10122 VDD.n14 VDD.t2996 30.379
R10123 VDD.n2907 VDD.t3295 30.379
R10124 VDD.n2907 VDD.t3293 30.379
R10125 VDD.t3496 VDD.n1135 25.7302
R10126 VDD.t1475 VDD.n674 25.6762
R10127 VDD.n1954 VDD.t588 25.395
R10128 VDD.n1954 VDD.t590 25.395
R10129 VDD.n1956 VDD.t1007 25.395
R10130 VDD.n1956 VDD.t1010 25.395
R10131 VDD.n2330 VDD.t2377 25.395
R10132 VDD.n2330 VDD.t2379 25.395
R10133 VDD.n2332 VDD.t2334 25.395
R10134 VDD.n2332 VDD.t2338 25.395
R10135 VDD.n2320 VDD.t2606 25.395
R10136 VDD.n2320 VDD.t2612 25.395
R10137 VDD.n2322 VDD.t2576 25.395
R10138 VDD.n2322 VDD.t2578 25.395
R10139 VDD.n2310 VDD.t2161 25.395
R10140 VDD.n2310 VDD.t2167 25.395
R10141 VDD.n2312 VDD.t2123 25.395
R10142 VDD.n2312 VDD.t2129 25.395
R10143 VDD.n2299 VDD.t3607 25.395
R10144 VDD.n2299 VDD.t3609 25.395
R10145 VDD.n2301 VDD.t3587 25.395
R10146 VDD.n2301 VDD.t3591 25.395
R10147 VDD.n2289 VDD.t3962 25.395
R10148 VDD.n2289 VDD.t3965 25.395
R10149 VDD.n2291 VDD.t3978 25.395
R10150 VDD.n2291 VDD.t3984 25.395
R10151 VDD.n2279 VDD.t3536 25.395
R10152 VDD.n2279 VDD.t3542 25.395
R10153 VDD.n2281 VDD.t3551 25.395
R10154 VDD.n2281 VDD.t3553 25.395
R10155 VDD.n2269 VDD.t1171 25.395
R10156 VDD.n2269 VDD.t1173 25.395
R10157 VDD.n2271 VDD.t1399 25.395
R10158 VDD.n2271 VDD.t1401 25.395
R10159 VDD.n1065 VDD.t41 25.395
R10160 VDD.n1065 VDD.t39 25.395
R10161 VDD.n1067 VDD.t37 25.395
R10162 VDD.n1067 VDD.t35 25.395
R10163 VDD.n936 VDD.t3929 25.395
R10164 VDD.n936 VDD.t3921 25.395
R10165 VDD.n938 VDD.t3925 25.395
R10166 VDD.n938 VDD.t3923 25.395
R10167 VDD.n807 VDD.t1478 25.395
R10168 VDD.n807 VDD.t1480 25.395
R10169 VDD.n809 VDD.t1227 25.395
R10170 VDD.n809 VDD.t1482 25.395
R10171 VDD.n656 VDD.t4306 25.395
R10172 VDD.n656 VDD.t4298 25.395
R10173 VDD.n658 VDD.t4302 25.395
R10174 VDD.n658 VDD.t4300 25.395
R10175 VDD.n527 VDD.t4252 25.395
R10176 VDD.n527 VDD.t4254 25.395
R10177 VDD.n529 VDD.t4258 25.395
R10178 VDD.n529 VDD.t4256 25.395
R10179 VDD.n398 VDD.t743 25.395
R10180 VDD.n398 VDD.t735 25.395
R10181 VDD.n400 VDD.t739 25.395
R10182 VDD.n400 VDD.t737 25.395
R10183 VDD.n269 VDD.t983 25.395
R10184 VDD.n269 VDD.t985 25.395
R10185 VDD.n271 VDD.t2906 25.395
R10186 VDD.n271 VDD.t2904 25.395
R10187 VDD.n131 VDD.t4315 25.395
R10188 VDD.n131 VDD.t4323 25.395
R10189 VDD.n133 VDD.t4321 25.395
R10190 VDD.n133 VDD.t4319 25.395
R10191 VDD.n2915 VDD.t3503 25.395
R10192 VDD.n2915 VDD.t3507 25.395
R10193 VDD.n2917 VDD.t3509 25.395
R10194 VDD.n2917 VDD.t3511 25.395
R10195 VDD.n2001 VDD.n1986 23.447
R10196 VDD.n2010 VDD.n2005 23.447
R10197 VDD.n2016 VDD.n1983 23.447
R10198 VDD.n2021 VDD.n1976 23.447
R10199 VDD.n2030 VDD.n2025 23.447
R10200 VDD.n2036 VDD.n1965 23.447
R10201 VDD.n1997 VDD.n1992 23.447
R10202 VDD.n1972 VDD.n1968 23.447
R10203 VDD.n2836 VDD.n1148 23.3925
R10204 VDD.n2845 VDD.n2840 23.3925
R10205 VDD.n2751 VDD.n2750 23.3925
R10206 VDD.n2762 VDD.n2761 23.3925
R10207 VDD.n2773 VDD.n2772 23.3925
R10208 VDD.n2784 VDD.n2783 23.3925
R10209 VDD.n2795 VDD.n2794 23.3925
R10210 VDD.n2806 VDD.n2805 23.3925
R10211 VDD.n2817 VDD.n2816 23.3925
R10212 VDD.n2828 VDD.n2827 23.3925
R10213 VDD.n2741 VDD.n1159 23.3925
R10214 VDD.n2735 VDD.n2730 23.3925
R10215 VDD.n2726 VDD.n2721 23.3925
R10216 VDD.n2353 VDD.n1181 23.3925
R10217 VDD.n2362 VDD.n2357 23.3925
R10218 VDD.n2365 VDD.n1175 23.3925
R10219 VDD.n1803 VDD.n1356 23.3925
R10220 VDD.n1791 VDD.n1362 23.3925
R10221 VDD.n1385 VDD.n1372 23.3925
R10222 VDD.n1382 VDD.n1378 23.3925
R10223 VDD.n1800 VDD.n1795 23.3925
R10224 VDD.n1445 VDD.n1440 23.3925
R10225 VDD.n1448 VDD.n1434 23.3925
R10226 VDD.n1631 VDD.n1430 23.3925
R10227 VDD.n1640 VDD.n1635 23.3925
R10228 VDD.n1649 VDD.n1644 23.3925
R10229 VDD.n1658 VDD.n1653 23.3925
R10230 VDD.n1667 VDD.n1662 23.3925
R10231 VDD.n1673 VDD.n1427 23.3925
R10232 VDD.n1608 VDD.n1603 23.3925
R10233 VDD.n1617 VDD.n1612 23.3925
R10234 VDD.n1620 VDD.n1456 23.3925
R10235 VDD.n1599 VDD.n1594 23.3925
R10236 VDD.n1590 VDD.n1585 23.3925
R10237 VDD.n1581 VDD.n1576 23.3925
R10238 VDD.n1572 VDD.n1567 23.3925
R10239 VDD.n1563 VDD.n1462 23.3925
R10240 VDD.n2717 VDD.n1162 23.3925
R10241 VDD.n2659 VDD.n2654 23.3925
R10242 VDD.n2662 VDD.n2424 23.3925
R10243 VDD.n2650 VDD.n2645 23.3925
R10244 VDD.n2641 VDD.n2430 23.3925
R10245 VDD.n2595 VDD.n2590 23.3925
R10246 VDD.n2598 VDD.n2444 23.3925
R10247 VDD.n2586 VDD.n2581 23.3925
R10248 VDD.n2577 VDD.n2450 23.3925
R10249 VDD.n2506 VDD.n2501 23.3925
R10250 VDD.n2515 VDD.n2510 23.3925
R10251 VDD.n2518 VDD.n2486 23.3925
R10252 VDD.n2497 VDD.n2492 23.3925
R10253 VDD.n2836 VDD.n2835 23.3556
R10254 VDD.n2845 VDD.n2844 23.3556
R10255 VDD.n2851 VDD.n2850 23.3556
R10256 VDD.n2751 VDD.n2746 23.3556
R10257 VDD.n2762 VDD.n2757 23.3556
R10258 VDD.n2773 VDD.n2768 23.3556
R10259 VDD.n2784 VDD.n2779 23.3556
R10260 VDD.n2795 VDD.n2790 23.3556
R10261 VDD.n2806 VDD.n2801 23.3556
R10262 VDD.n2817 VDD.n2812 23.3556
R10263 VDD.n2828 VDD.n2823 23.3556
R10264 VDD.n2741 VDD.n2740 23.3556
R10265 VDD.n2735 VDD.n2734 23.3556
R10266 VDD.n2726 VDD.n2724 23.3556
R10267 VDD.n2001 VDD.n1989 23.3556
R10268 VDD.n2010 VDD.n2008 23.3556
R10269 VDD.n2016 VDD.n2015 23.3556
R10270 VDD.n2021 VDD.n1979 23.3556
R10271 VDD.n2030 VDD.n2028 23.3556
R10272 VDD.n2036 VDD.n2035 23.3556
R10273 VDD.n1997 VDD.n1995 23.3556
R10274 VDD.n1972 VDD.n1971 23.3556
R10275 VDD.n2353 VDD.n2352 23.3556
R10276 VDD.n2362 VDD.n2361 23.3556
R10277 VDD.n2365 VDD.n1178 23.3556
R10278 VDD.n1803 VDD.n1359 23.3556
R10279 VDD.n1791 VDD.n1790 23.3556
R10280 VDD.n1385 VDD.n1375 23.3556
R10281 VDD.n1382 VDD.n1381 23.3556
R10282 VDD.n1800 VDD.n1798 23.3556
R10283 VDD.n1445 VDD.n1444 23.3556
R10284 VDD.n1448 VDD.n1437 23.3556
R10285 VDD.n1631 VDD.n1630 23.3556
R10286 VDD.n1640 VDD.n1639 23.3556
R10287 VDD.n1649 VDD.n1647 23.3556
R10288 VDD.n1658 VDD.n1657 23.3556
R10289 VDD.n1667 VDD.n1666 23.3556
R10290 VDD.n1673 VDD.n1672 23.3556
R10291 VDD.n1608 VDD.n1607 23.3556
R10292 VDD.n1617 VDD.n1616 23.3556
R10293 VDD.n1620 VDD.n1459 23.3556
R10294 VDD.n1599 VDD.n1598 23.3556
R10295 VDD.n1590 VDD.n1588 23.3556
R10296 VDD.n1581 VDD.n1580 23.3556
R10297 VDD.n1572 VDD.n1571 23.3556
R10298 VDD.n1563 VDD.n1465 23.3556
R10299 VDD.n2717 VDD.n2716 23.3556
R10300 VDD.n2659 VDD.n2657 23.3556
R10301 VDD.n2662 VDD.n2427 23.3556
R10302 VDD.n2650 VDD.n2648 23.3556
R10303 VDD.n2641 VDD.n2640 23.3556
R10304 VDD.n2595 VDD.n2593 23.3556
R10305 VDD.n2598 VDD.n2447 23.3556
R10306 VDD.n2586 VDD.n2584 23.3556
R10307 VDD.n2577 VDD.n2576 23.3556
R10308 VDD.n2506 VDD.n2505 23.3556
R10309 VDD.n2515 VDD.n2514 23.3556
R10310 VDD.n2518 VDD.n2489 23.3556
R10311 VDD.n2497 VDD.n2495 23.3556
R10312 VDD.n2218 VDD.t887 23.1467
R10313 VDD.n2243 VDD.t313 23.1467
R10314 VDD.n2837 VDD.n2836 22.3465
R10315 VDD.n2846 VDD.n2845 22.3465
R10316 VDD.n2851 VDD.n2847 22.3465
R10317 VDD.n2751 VDD.n2747 22.3465
R10318 VDD.n2762 VDD.n2758 22.3465
R10319 VDD.n2773 VDD.n2769 22.3465
R10320 VDD.n2784 VDD.n2780 22.3465
R10321 VDD.n2795 VDD.n2791 22.3465
R10322 VDD.n2806 VDD.n2802 22.3465
R10323 VDD.n2817 VDD.n2813 22.3465
R10324 VDD.n2828 VDD.n2824 22.3465
R10325 VDD.n2736 VDD.n2735 22.3465
R10326 VDD.n1997 VDD.n1996 22.3465
R10327 VDD.n2002 VDD.n2001 22.3465
R10328 VDD.n2011 VDD.n2010 22.3465
R10329 VDD.n2016 VDD.n2012 22.3465
R10330 VDD.n2022 VDD.n2021 22.3465
R10331 VDD.n2031 VDD.n2030 22.3465
R10332 VDD.n2036 VDD.n2032 22.3465
R10333 VDD.n1973 VDD.n1972 22.3465
R10334 VDD.n2354 VDD.n2353 22.3465
R10335 VDD.n2363 VDD.n2362 22.3465
R10336 VDD.n2365 VDD.n2364 22.3465
R10337 VDD.n1803 VDD.n1802 22.3465
R10338 VDD.n1792 VDD.n1791 22.3465
R10339 VDD.n1385 VDD.n1384 22.3465
R10340 VDD.n1383 VDD.n1382 22.3465
R10341 VDD.n1801 VDD.n1800 22.3465
R10342 VDD.n1446 VDD.n1445 22.3465
R10343 VDD.n1448 VDD.n1447 22.3465
R10344 VDD.n1632 VDD.n1631 22.3465
R10345 VDD.n1641 VDD.n1640 22.3465
R10346 VDD.n1659 VDD.n1658 22.3465
R10347 VDD.n1668 VDD.n1667 22.3465
R10348 VDD.n1650 VDD.n1649 22.3465
R10349 VDD.n1673 VDD.n1669 22.3465
R10350 VDD.n1609 VDD.n1608 22.3465
R10351 VDD.n1618 VDD.n1617 22.3465
R10352 VDD.n1620 VDD.n1619 22.3465
R10353 VDD.n1600 VDD.n1599 22.3465
R10354 VDD.n1582 VDD.n1581 22.3465
R10355 VDD.n1573 VDD.n1572 22.3465
R10356 VDD.n1591 VDD.n1590 22.3465
R10357 VDD.n1564 VDD.n1563 22.3465
R10358 VDD.n2718 VDD.n2717 22.3465
R10359 VDD.n2662 VDD.n2661 22.3465
R10360 VDD.n2642 VDD.n2641 22.3465
R10361 VDD.n2598 VDD.n2597 22.3465
R10362 VDD.n2578 VDD.n2577 22.3465
R10363 VDD.n2507 VDD.n2506 22.3465
R10364 VDD.n2516 VDD.n2515 22.3465
R10365 VDD.n2518 VDD.n2517 22.3465
R10366 VDD.n2587 VDD.n2586 22.3465
R10367 VDD.n2596 VDD.n2595 22.3465
R10368 VDD.n2651 VDD.n2650 22.3465
R10369 VDD.n2660 VDD.n2659 22.3465
R10370 VDD.n2727 VDD.n2726 22.3465
R10371 VDD.n2741 VDD.n2737 22.3465
R10372 VDD.n2498 VDD.n2497 22.3465
R10373 VDD.n1113 VDD.t77 20.1899
R10374 VDD.n1113 VDD.t3754 20.1899
R10375 VDD.n1081 VDD.t2940 20.1899
R10376 VDD.n1081 VDD.t79 20.1899
R10377 VDD.n1079 VDD.t808 20.1899
R10378 VDD.n1079 VDD.t3096 20.1899
R10379 VDD.n1083 VDD.t71 20.1899
R10380 VDD.n1083 VDD.t3732 20.1899
R10381 VDD.n1107 VDD.t1260 20.1899
R10382 VDD.n1107 VDD.t75 20.1899
R10383 VDD.n1109 VDD.t3694 20.1899
R10384 VDD.n1109 VDD.t1264 20.1899
R10385 VDD.n1101 VDD.t4338 20.1899
R10386 VDD.n1101 VDD.t3865 20.1899
R10387 VDD.n1089 VDD.t3009 20.1899
R10388 VDD.n1089 VDD.t4420 20.1899
R10389 VDD.n1087 VDD.t1063 20.1899
R10390 VDD.n1087 VDD.t2967 20.1899
R10391 VDD.n1091 VDD.t4386 20.1899
R10392 VDD.n1091 VDD.t3721 20.1899
R10393 VDD.n1095 VDD.t1268 20.1899
R10394 VDD.n1095 VDD.t4447 20.1899
R10395 VDD.n1097 VDD.t2381 20.1899
R10396 VDD.n1097 VDD.t1272 20.1899
R10397 VDD.n1077 VDD.t1307 20.1899
R10398 VDD.n1077 VDD.t1326 20.1899
R10399 VDD.n1119 VDD.t631 20.1899
R10400 VDD.n1119 VDD.t1309 20.1899
R10401 VDD.n1121 VDD.t1598 20.1899
R10402 VDD.n1121 VDD.t633 20.1899
R10403 VDD.n1024 VDD.t4509 20.1899
R10404 VDD.n1024 VDD.t3183 20.1899
R10405 VDD.n1028 VDD.t3217 20.1899
R10406 VDD.n1028 VDD.t4408 20.1899
R10407 VDD.n1030 VDD.t792 20.1899
R10408 VDD.n1030 VDD.t3221 20.1899
R10409 VDD.n1034 VDD.t4480 20.1899
R10410 VDD.n1034 VDD.t3177 20.1899
R10411 VDD.n1008 VDD.t3058 20.1899
R10412 VDD.n1008 VDD.t4361 20.1899
R10413 VDD.n1006 VDD.t949 20.1899
R10414 VDD.n1006 VDD.t2995 20.1899
R10415 VDD.n1002 VDD.t3201 20.1899
R10416 VDD.n1002 VDD.t3185 20.1899
R10417 VDD.n1040 VDD.t3225 20.1899
R10418 VDD.n1040 VDD.t3205 20.1899
R10419 VDD.n1042 VDD.t1535 20.1899
R10420 VDD.n1042 VDD.t3229 20.1899
R10421 VDD.n1046 VDD.t3213 20.1899
R10422 VDD.n1046 VDD.t3173 20.1899
R10423 VDD.n1000 VDD.t3102 20.1899
R10424 VDD.n1000 VDD.t3215 20.1899
R10425 VDD.n998 VDD.t2030 20.1899
R10426 VDD.n998 VDD.t3079 20.1899
R10427 VDD.n996 VDD.t81 20.1899
R10428 VDD.n996 VDD.t4332 20.1899
R10429 VDD.n1052 VDD.t2108 20.1899
R10430 VDD.n1052 VDD.t2398 20.1899
R10431 VDD.n1054 VDD.t915 20.1899
R10432 VDD.n1054 VDD.t2110 20.1899
R10433 VDD.n984 VDD.t3209 20.1899
R10434 VDD.n984 VDD.t3736 20.1899
R10435 VDD.n952 VDD.t2985 20.1899
R10436 VDD.n952 VDD.t3211 20.1899
R10437 VDD.n950 VDD.t2212 20.1899
R10438 VDD.n950 VDD.t2971 20.1899
R10439 VDD.n954 VDD.t3203 20.1899
R10440 VDD.n954 VDD.t3878 20.1899
R10441 VDD.n978 VDD.t3227 20.1899
R10442 VDD.n978 VDD.t3207 20.1899
R10443 VDD.n980 VDD.t63 20.1899
R10444 VDD.n980 VDD.t3231 20.1899
R10445 VDD.n972 VDD.t4484 20.1899
R10446 VDD.n972 VDD.t3804 20.1899
R10447 VDD.n960 VDD.t3052 20.1899
R10448 VDD.n960 VDD.t4372 20.1899
R10449 VDD.n958 VDD.t624 20.1899
R10450 VDD.n958 VDD.t2991 20.1899
R10451 VDD.n962 VDD.t4336 20.1899
R10452 VDD.n962 VDD.t3859 20.1899
R10453 VDD.n966 VDD.t3219 20.1899
R10454 VDD.n966 VDD.t4416 20.1899
R10455 VDD.n968 VDD.t1251 20.1899
R10456 VDD.n968 VDD.t3223 20.1899
R10457 VDD.n948 VDD.t657 20.1899
R10458 VDD.n948 VDD.t1349 20.1899
R10459 VDD.n990 VDD.t2849 20.1899
R10460 VDD.n990 VDD.t659 20.1899
R10461 VDD.n992 VDD.t4294 20.1899
R10462 VDD.n992 VDD.t1541 20.1899
R10463 VDD.n895 VDD.t4368 20.1899
R10464 VDD.n895 VDD.t2799 20.1899
R10465 VDD.n899 VDD.t2532 20.1899
R10466 VDD.n899 VDD.t4475 20.1899
R10467 VDD.n901 VDD.t438 20.1899
R10468 VDD.n901 VDD.t2530 20.1899
R10469 VDD.n905 VDD.t4394 20.1899
R10470 VDD.n905 VDD.t2803 20.1899
R10471 VDD.n879 VDD.t2964 20.1899
R10472 VDD.n879 VDD.t4502 20.1899
R10473 VDD.n877 VDD.t1493 20.1899
R10474 VDD.n877 VDD.t3015 20.1899
R10475 VDD.n873 VDD.t2678 20.1899
R10476 VDD.n873 VDD.t2797 20.1899
R10477 VDD.n911 VDD.t2524 20.1899
R10478 VDD.n911 VDD.t2676 20.1899
R10479 VDD.n913 VDD.t1 20.1899
R10480 VDD.n913 VDD.t2522 20.1899
R10481 VDD.n917 VDD.t2670 20.1899
R10482 VDD.n917 VDD.t2809 20.1899
R10483 VDD.n871 VDD.t2946 20.1899
R10484 VDD.n871 VDD.t2668 20.1899
R10485 VDD.n869 VDD.t1649 20.1899
R10486 VDD.n869 VDD.t2960 20.1899
R10487 VDD.n867 VDD.t1194 20.1899
R10488 VDD.n867 VDD.t1458 20.1899
R10489 VDD.n923 VDD.t3118 20.1899
R10490 VDD.n923 VDD.t1192 20.1899
R10491 VDD.n925 VDD.t2643 20.1899
R10492 VDD.n925 VDD.t3116 20.1899
R10493 VDD.n855 VDD.t2674 20.1899
R10494 VDD.n855 VDD.t3707 20.1899
R10495 VDD.n823 VDD.t3041 20.1899
R10496 VDD.n823 VDD.t2672 20.1899
R10497 VDD.n821 VDD.t1724 20.1899
R10498 VDD.n821 VDD.t3049 20.1899
R10499 VDD.n825 VDD.t2682 20.1899
R10500 VDD.n825 VDD.t3739 20.1899
R10501 VDD.n849 VDD.t2528 20.1899
R10502 VDD.n849 VDD.t2680 20.1899
R10503 VDD.n851 VDD.t1208 20.1899
R10504 VDD.n851 VDD.t2526 20.1899
R10505 VDD.n843 VDD.t4414 20.1899
R10506 VDD.n843 VDD.t3751 20.1899
R10507 VDD.n831 VDD.t2936 20.1899
R10508 VDD.n831 VDD.t4507 20.1899
R10509 VDD.n829 VDD.t1141 20.1899
R10510 VDD.n829 VDD.t3005 20.1899
R10511 VDD.n833 VDD.t4384 20.1899
R10512 VDD.n833 VDD.t3741 20.1899
R10513 VDD.n837 VDD.t2536 20.1899
R10514 VDD.n837 VDD.t4490 20.1899
R10515 VDD.n839 VDD.t3400 20.1899
R10516 VDD.n839 VDD.t2534 20.1899
R10517 VDD.n819 VDD.t2853 20.1899
R10518 VDD.n819 VDD.t3352 20.1899
R10519 VDD.n861 VDD.t1221 20.1899
R10520 VDD.n861 VDD.t2851 20.1899
R10521 VDD.n863 VDD.t924 20.1899
R10522 VDD.n863 VDD.t1219 20.1899
R10523 VDD.n766 VDD.t4459 20.1899
R10524 VDD.n766 VDD.t126 20.1899
R10525 VDD.n770 VDD.t3364 20.1899
R10526 VDD.n770 VDD.t4392 20.1899
R10527 VDD.n772 VDD.t2795 20.1899
R10528 VDD.n772 VDD.t3360 20.1899
R10529 VDD.n776 VDD.t4486 20.1899
R10530 VDD.n776 VDD.t130 20.1899
R10531 VDD.n750 VDD.t3037 20.1899
R10532 VDD.n750 VDD.t4423 20.1899
R10533 VDD.n748 VDD.t412 20.1899
R10534 VDD.n748 VDD.t2930 20.1899
R10535 VDD.n744 VDD.t3251 20.1899
R10536 VDD.n744 VDD.t124 20.1899
R10537 VDD.n782 VDD.t3372 20.1899
R10538 VDD.n782 VDD.t3247 20.1899
R10539 VDD.n784 VDD.t242 20.1899
R10540 VDD.n784 VDD.t3368 20.1899
R10541 VDD.n788 VDD.t3261 20.1899
R10542 VDD.n788 VDD.t120 20.1899
R10543 VDD.n742 VDD.t3019 20.1899
R10544 VDD.n742 VDD.t3259 20.1899
R10545 VDD.n740 VDD.t15 20.1899
R10546 VDD.n740 VDD.t3035 20.1899
R10547 VDD.n738 VDD.t1891 20.1899
R10548 VDD.n738 VDD.t2486 20.1899
R10549 VDD.n794 VDD.t821 20.1899
R10550 VDD.n794 VDD.t1889 20.1899
R10551 VDD.n796 VDD.t2789 20.1899
R10552 VDD.n796 VDD.t819 20.1899
R10553 VDD.n726 VDD.t3257 20.1899
R10554 VDD.n726 VDD.t3839 20.1899
R10555 VDD.n694 VDD.t3081 20.1899
R10556 VDD.n694 VDD.t3255 20.1899
R10557 VDD.n692 VDD.t3572 20.1899
R10558 VDD.n692 VDD.t3092 20.1899
R10559 VDD.n696 VDD.t3253 20.1899
R10560 VDD.n696 VDD.t3808 20.1899
R10561 VDD.n720 VDD.t3374 20.1899
R10562 VDD.n720 VDD.t3249 20.1899
R10563 VDD.n722 VDD.t46 20.1899
R10564 VDD.n722 VDD.t3370 20.1899
R10565 VDD.n714 VDD.t4492 20.1899
R10566 VDD.n714 VDD.t3847 20.1899
R10567 VDD.n702 VDD.t3031 20.1899
R10568 VDD.n702 VDD.t4428 20.1899
R10569 VDD.n700 VDD.t1623 20.1899
R10570 VDD.n700 VDD.t2926 20.1899
R10571 VDD.n704 VDD.t4464 20.1899
R10572 VDD.n704 VDD.t3814 20.1899
R10573 VDD.n708 VDD.t3366 20.1899
R10574 VDD.n708 VDD.t4400 20.1899
R10575 VDD.n710 VDD.t1867 20.1899
R10576 VDD.n710 VDD.t3362 20.1899
R10577 VDD.n690 VDD.t1871 20.1899
R10578 VDD.n690 VDD.t4170 20.1899
R10579 VDD.n732 VDD.t229 20.1899
R10580 VDD.n732 VDD.t1869 20.1899
R10581 VDD.n734 VDD.t4023 20.1899
R10582 VDD.n734 VDD.t231 20.1899
R10583 VDD.n637 VDD.t3636 20.1899
R10584 VDD.n637 VDD.t1381 20.1899
R10585 VDD.n591 VDD.t3068 20.1899
R10586 VDD.n591 VDD.t3632 20.1899
R10587 VDD.n589 VDD.t1365 20.1899
R10588 VDD.n589 VDD.t3084 20.1899
R10589 VDD.n593 VDD.t3624 20.1899
R10590 VDD.n593 VDD.t1369 20.1899
R10591 VDD.n631 VDD.t1991 20.1899
R10592 VDD.n631 VDD.t3638 20.1899
R10593 VDD.n633 VDD.t3350 20.1899
R10594 VDD.n633 VDD.t1989 20.1899
R10595 VDD.n625 VDD.t4440 20.1899
R10596 VDD.n625 VDD.t1375 20.1899
R10597 VDD.n599 VDD.t3088 20.1899
R10598 VDD.n599 VDD.t4365 20.1899
R10599 VDD.n597 VDD.t2044 20.1899
R10600 VDD.n597 VDD.t2987 20.1899
R10601 VDD.n615 VDD.t4418 20.1899
R10602 VDD.n615 VDD.t1371 20.1899
R10603 VDD.n619 VDD.t1722 20.1899
R10604 VDD.n619 VDD.t4511 20.1899
R10605 VDD.n621 VDD.t875 20.1899
R10606 VDD.n621 VDD.t1995 20.1899
R10607 VDD.n587 VDD.t3578 20.1899
R10608 VDD.n587 VDD.t3416 20.1899
R10609 VDD.n643 VDD.t1424 20.1899
R10610 VDD.n643 VDD.t3576 20.1899
R10611 VDD.n645 VDD.t1214 20.1899
R10612 VDD.n645 VDD.t1422 20.1899
R10613 VDD.n575 VDD.t3634 20.1899
R10614 VDD.n575 VDD.t3843 20.1899
R10615 VDD.n543 VDD.t3075 20.1899
R10616 VDD.n543 VDD.t3630 20.1899
R10617 VDD.n541 VDD.t3955 20.1899
R10618 VDD.n541 VDD.t3090 20.1899
R10619 VDD.n545 VDD.t3628 20.1899
R10620 VDD.n545 VDD.t3812 20.1899
R10621 VDD.n569 VDD.t1997 20.1899
R10622 VDD.n569 VDD.t3626 20.1899
R10623 VDD.n571 VDD.t4133 20.1899
R10624 VDD.n571 VDD.t1993 20.1899
R10625 VDD.n563 VDD.t4496 20.1899
R10626 VDD.n563 VDD.t3855 20.1899
R10627 VDD.n551 VDD.t3025 20.1899
R10628 VDD.n551 VDD.t4430 20.1899
R10629 VDD.n549 VDD.t177 20.1899
R10630 VDD.n549 VDD.t3100 20.1899
R10631 VDD.n553 VDD.t4466 20.1899
R10632 VDD.n553 VDD.t3818 20.1899
R10633 VDD.n557 VDD.t1987 20.1899
R10634 VDD.n557 VDD.t4402 20.1899
R10635 VDD.n559 VDD.t1489 20.1899
R10636 VDD.n559 VDD.t1985 20.1899
R10637 VDD.n539 VDD.t2699 20.1899
R10638 VDD.n539 VDD.t235 20.1899
R10639 VDD.n581 VDD.t4246 20.1899
R10640 VDD.n581 VDD.t2697 20.1899
R10641 VDD.n583 VDD.t1156 20.1899
R10642 VDD.n583 VDD.t4248 20.1899
R10643 VDD.n486 VDD.t4461 20.1899
R10644 VDD.n486 VDD.t3134 20.1899
R10645 VDD.n490 VDD.t198 20.1899
R10646 VDD.n490 VDD.t4396 20.1899
R10647 VDD.n492 VDD.t505 20.1899
R10648 VDD.n492 VDD.t2051 20.1899
R10649 VDD.n496 VDD.t4488 20.1899
R10650 VDD.n496 VDD.t3138 20.1899
R10651 VDD.n470 VDD.t3033 20.1899
R10652 VDD.n470 VDD.t4425 20.1899
R10653 VDD.n468 VDD.t2647 20.1899
R10654 VDD.n468 VDD.t2928 20.1899
R10655 VDD.n464 VDD.t190 20.1899
R10656 VDD.n464 VDD.t3132 20.1899
R10657 VDD.n502 VDD.t206 20.1899
R10658 VDD.n502 VDD.t188 20.1899
R10659 VDD.n504 VDD.t608 20.1899
R10660 VDD.n504 VDD.t204 20.1899
R10661 VDD.n508 VDD.t194 20.1899
R10662 VDD.n508 VDD.t3128 20.1899
R10663 VDD.n462 VDD.t3017 20.1899
R10664 VDD.n462 VDD.t192 20.1899
R10665 VDD.n460 VDD.t1106 20.1899
R10666 VDD.n460 VDD.t3029 20.1899
R10667 VDD.n458 VDD.t2550 20.1899
R10668 VDD.n458 VDD.t959 20.1899
R10669 VDD.n514 VDD.t4262 20.1899
R10670 VDD.n514 VDD.t2548 20.1899
R10671 VDD.n516 VDD.t513 20.1899
R10672 VDD.n516 VDD.t4264 20.1899
R10673 VDD.n446 VDD.t186 20.1899
R10674 VDD.n446 VDD.t3788 20.1899
R10675 VDD.n414 VDD.t2948 20.1899
R10676 VDD.n414 VDD.t184 20.1899
R10677 VDD.n412 VDD.t54 20.1899
R10678 VDD.n412 VDD.t2962 20.1899
R10679 VDD.n416 VDD.t182 20.1899
R10680 VDD.n416 VDD.t3763 20.1899
R10681 VDD.n440 VDD.t202 20.1899
R10682 VDD.n440 VDD.t180 20.1899
R10683 VDD.n442 VDD.t1204 20.1899
R10684 VDD.n442 VDD.t200 20.1899
R10685 VDD.n434 VDD.t4453 20.1899
R10686 VDD.n434 VDD.t3797 20.1899
R10687 VDD.n422 VDD.t3066 20.1899
R10688 VDD.n422 VDD.t4382 20.1899
R10689 VDD.n420 VDD.t845 20.1899
R10690 VDD.n420 VDD.t2981 20.1899
R10691 VDD.n424 VDD.t4433 20.1899
R10692 VDD.n424 VDD.t3768 20.1899
R10693 VDD.n428 VDD.t2049 20.1899
R10694 VDD.n428 VDD.t4344 20.1899
R10695 VDD.n430 VDD.t2791 20.1899
R10696 VDD.n430 VDD.t208 20.1899
R10697 VDD.n410 VDD.t2867 20.1899
R10698 VDD.n410 VDD.t50 20.1899
R10699 VDD.n452 VDD.t2099 20.1899
R10700 VDD.n452 VDD.t2865 20.1899
R10701 VDD.n454 VDD.t2040 20.1899
R10702 VDD.n454 VDD.t2097 20.1899
R10703 VDD.n357 VDD.t4352 20.1899
R10704 VDD.n357 VDD.t1504 20.1899
R10705 VDD.n361 VDD.t3162 20.1899
R10706 VDD.n361 VDD.t4468 20.1899
R10707 VDD.n363 VDD.t1235 20.1899
R10708 VDD.n363 VDD.t3160 20.1899
R10709 VDD.n367 VDD.t4390 20.1899
R10710 VDD.n367 VDD.t1508 20.1899
R10711 VDD.n341 VDD.t2977 20.1899
R10712 VDD.n341 VDD.t4498 20.1899
R10713 VDD.n339 VDD.t3146 20.1899
R10714 VDD.n339 VDD.t3023 20.1899
R10715 VDD.n335 VDD.t2666 20.1899
R10716 VDD.n335 VDD.t1134 20.1899
R10717 VDD.n373 VDD.t3158 20.1899
R10718 VDD.n373 VDD.t2664 20.1899
R10719 VDD.n375 VDD.t1496 20.1899
R10720 VDD.n375 VDD.t3154 20.1899
R10721 VDD.n379 VDD.t2654 20.1899
R10722 VDD.n379 VDD.t1514 20.1899
R10723 VDD.n333 VDD.t2956 20.1899
R10724 VDD.n333 VDD.t2652 20.1899
R10725 VDD.n331 VDD.t2493 20.1899
R10726 VDD.n331 VDD.t2975 20.1899
R10727 VDD.n329 VDD.t3337 20.1899
R10728 VDD.n329 VDD.t169 20.1899
R10729 VDD.n385 VDD.t1163 20.1899
R10730 VDD.n385 VDD.t3335 20.1899
R10731 VDD.n387 VDD.t1473 20.1899
R10732 VDD.n387 VDD.t1161 20.1899
R10733 VDD.n317 VDD.t2662 20.1899
R10734 VDD.n317 VDD.t3845 20.1899
R10735 VDD.n285 VDD.t3070 20.1899
R10736 VDD.n285 VDD.t2660 20.1899
R10737 VDD.n283 VDD.t2281 20.1899
R10738 VDD.n283 VDD.t3086 20.1899
R10739 VDD.n287 VDD.t2658 20.1899
R10740 VDD.n287 VDD.t3816 20.1899
R10741 VDD.n311 VDD.t3166 20.1899
R10742 VDD.n311 VDD.t2656 20.1899
R10743 VDD.n313 VDD.t3993 20.1899
R10744 VDD.n313 VDD.t3164 20.1899
R10745 VDD.n305 VDD.t4500 20.1899
R10746 VDD.n305 VDD.t3861 20.1899
R10747 VDD.n293 VDD.t3021 20.1899
R10748 VDD.n293 VDD.t4435 20.1899
R10749 VDD.n291 VDD.t1067 20.1899
R10750 VDD.n291 VDD.t3098 20.1899
R10751 VDD.n295 VDD.t4470 20.1899
R10752 VDD.n295 VDD.t3822 20.1899
R10753 VDD.n299 VDD.t3156 20.1899
R10754 VDD.n299 VDD.t4404 20.1899
R10755 VDD.n301 VDD.t1863 20.1899
R10756 VDD.n301 VDD.t3152 20.1899
R10757 VDD.n281 VDD.t1445 20.1899
R10758 VDD.n281 VDD.t2572 20.1899
R10759 VDD.n323 VDD.t354 20.1899
R10760 VDD.n323 VDD.t1443 20.1899
R10761 VDD.n325 VDD.t2287 20.1899
R10762 VDD.n325 VDD.t356 20.1899
R10763 VDD.n188 VDD.t570 20.1899
R10764 VDD.n188 VDD.t3745 20.1899
R10765 VDD.n156 VDD.t2993 20.1899
R10766 VDD.n156 VDD.t568 20.1899
R10767 VDD.n154 VDD.t418 20.1899
R10768 VDD.n154 VDD.t2998 20.1899
R10769 VDD.n158 VDD.t326 20.1899
R10770 VDD.n158 VDD.t3765 20.1899
R10771 VDD.n182 VDD.t2452 20.1899
R10772 VDD.n182 VDD.t324 20.1899
R10773 VDD.n184 VDD.t3268 20.1899
R10774 VDD.n184 VDD.t11 20.1899
R10775 VDD.n176 VDD.t4455 20.1899
R10776 VDD.n176 VDD.t3802 20.1899
R10777 VDD.n164 VDD.t3063 20.1899
R10778 VDD.n164 VDD.t4388 20.1899
R10779 VDD.n162 VDD.t282 20.1899
R10780 VDD.n162 VDD.t2979 20.1899
R10781 VDD.n166 VDD.t4437 20.1899
R10782 VDD.n166 VDD.t3771 20.1899
R10783 VDD.n170 VDD.t5 20.1899
R10784 VDD.n170 VDD.t4350 20.1899
R10785 VDD.n172 VDD.t360 20.1899
R10786 VDD.n172 VDD.t2456 20.1899
R10787 VDD.n152 VDD.t2028 20.1899
R10788 VDD.n152 VDD.t414 20.1899
R10789 VDD.n194 VDD.t274 20.1899
R10790 VDD.n194 VDD.t2026 20.1899
R10791 VDD.n196 VDD.t493 20.1899
R10792 VDD.n196 VDD.t272 20.1899
R10793 VDD.n228 VDD.t4370 20.1899
R10794 VDD.n228 VDD.t422 20.1899
R10795 VDD.n232 VDD.t2454 20.1899
R10796 VDD.n232 VDD.t4477 20.1899
R10797 VDD.n234 VDD.t509 20.1899
R10798 VDD.n234 VDD.t13 20.1899
R10799 VDD.n238 VDD.t4398 20.1899
R10800 VDD.n238 VDD.t426 20.1899
R10801 VDD.n212 VDD.t2958 20.1899
R10802 VDD.n212 VDD.t4504 20.1899
R10803 VDD.n210 VDD.t1225 20.1899
R10804 VDD.n210 VDD.t3011 20.1899
R10805 VDD.n206 VDD.t566 20.1899
R10806 VDD.n206 VDD.t420 20.1899
R10807 VDD.n244 VDD.t9 20.1899
R10808 VDD.n244 VDD.t332 20.1899
R10809 VDD.n246 VDD.t3299 20.1899
R10810 VDD.n246 VDD.t7 20.1899
R10811 VDD.n250 VDD.t330 20.1899
R10812 VDD.n250 VDD.t432 20.1899
R10813 VDD.n204 VDD.t2942 20.1899
R10814 VDD.n204 VDD.t328 20.1899
R10815 VDD.n202 VDD.t3341 20.1899
R10816 VDD.n202 VDD.t2954 20.1899
R10817 VDD.n200 VDD.t1454 20.1899
R10818 VDD.n200 VDD.t865 20.1899
R10819 VDD.n256 VDD.t2768 20.1899
R10820 VDD.n256 VDD.t1452 20.1899
R10821 VDD.n258 VDD.t911 20.1899
R10822 VDD.n258 VDD.t2766 20.1899
R10823 VDD.n90 VDD.t4378 20.1899
R10824 VDD.n90 VDD.t1710 20.1899
R10825 VDD.n94 VDD.t1266 20.1899
R10826 VDD.n94 VDD.t4445 20.1899
R10827 VDD.n96 VDD.t578 20.1899
R10828 VDD.n96 VDD.t1270 20.1899
R10829 VDD.n100 VDD.t4513 20.1899
R10830 VDD.n100 VDD.t1720 20.1899
R10831 VDD.n74 VDD.t3013 20.1899
R10832 VDD.n74 VDD.t4412 20.1899
R10833 VDD.n72 VDD.t883 20.1899
R10834 VDD.n72 VDD.t2973 20.1899
R10835 VDD.n68 VDD.t69 20.1899
R10836 VDD.n68 VDD.t1712 20.1899
R10837 VDD.n106 VDD.t1274 20.1899
R10838 VDD.n106 VDD.t73 20.1899
R10839 VDD.n108 VDD.t3356 20.1899
R10840 VDD.n108 VDD.t1262 20.1899
R10841 VDD.n112 VDD.t1420 20.1899
R10842 VDD.n112 VDD.t1716 20.1899
R10843 VDD.n66 VDD.t3056 20.1899
R10844 VDD.n66 VDD.t67 20.1899
R10845 VDD.n64 VDD.t97 20.1899
R10846 VDD.n64 VDD.t3045 20.1899
R10847 VDD.n62 VDD.t931 20.1899
R10848 VDD.n62 VDD.t3331 20.1899
R10849 VDD.n118 VDD.t926 20.1899
R10850 VDD.n118 VDD.t933 20.1899
R10851 VDD.n120 VDD.t769 20.1899
R10852 VDD.n120 VDD.t4065 20.1899
R10853 VDD.n2893 VDD.t651 20.1899
R10854 VDD.n2893 VDD.t3760 20.1899
R10855 VDD.n2861 VDD.t3077 20.1899
R10856 VDD.n2861 VDD.t647 20.1899
R10857 VDD.n2859 VDD.t1923 20.1899
R10858 VDD.n2859 VDD.t2924 20.1899
R10859 VDD.n2863 VDD.t655 20.1899
R10860 VDD.n2863 VDD.t3794 20.1899
R10861 VDD.n2887 VDD.t851 20.1899
R10862 VDD.n2887 VDD.t653 20.1899
R10863 VDD.n2889 VDD.t1909 20.1899
R10864 VDD.n2889 VDD.t849 20.1899
R10865 VDD.n2881 VDD.t4473 20.1899
R10866 VDD.n2881 VDD.t3841 20.1899
R10867 VDD.n2869 VDD.t2932 20.1899
R10868 VDD.n2869 VDD.t4342 20.1899
R10869 VDD.n2867 VDD.t2514 20.1899
R10870 VDD.n2867 VDD.t3047 20.1899
R10871 VDD.n2871 VDD.t4494 20.1899
R10872 VDD.n2871 VDD.t3873 20.1899
R10873 VDD.n2875 VDD.t847 20.1899
R10874 VDD.n2875 VDD.t4376 20.1899
R10875 VDD.n2877 VDD.t1686 20.1899
R10876 VDD.n2877 VDD.t861 20.1899
R10877 VDD.n2857 VDD.t1069 20.1899
R10878 VDD.n2857 VDD.t1500 20.1899
R10879 VDD.n2899 VDD.t2069 20.1899
R10880 VDD.n2899 VDD.t1071 20.1899
R10881 VDD.n2901 VDD.t1258 20.1899
R10882 VDD.n2901 VDD.t2067 20.1899
R10883 VDD.n28 VDD.t4451 20.1899
R10884 VDD.n28 VDD.t2898 20.1899
R10885 VDD.n32 VDD.t859 20.1899
R10886 VDD.n32 VDD.t4363 20.1899
R10887 VDD.n34 VDD.t1969 20.1899
R10888 VDD.n34 VDD.t857 20.1899
R10889 VDD.n38 VDD.t4442 20.1899
R10890 VDD.n38 VDD.t2896 20.1899
R10891 VDD.n12 VDD.t2969 20.1899
R10892 VDD.n12 VDD.t4340 20.1899
R10893 VDD.n10 VDD.t1977 20.1899
R10894 VDD.n10 VDD.t3043 20.1899
R10895 VDD.n6 VDD.t643 20.1899
R10896 VDD.n6 VDD.t2894 20.1899
R10897 VDD.n44 VDD.t855 20.1899
R10898 VDD.n44 VDD.t641 20.1899
R10899 VDD.n46 VDD.t1579 20.1899
R10900 VDD.n46 VDD.t853 20.1899
R10901 VDD.n50 VDD.t649 20.1899
R10902 VDD.n50 VDD.t2890 20.1899
R10903 VDD.n4 VDD.t3039 20.1899
R10904 VDD.n4 VDD.t645 20.1899
R10905 VDD.n2 VDD.t1919 20.1899
R10906 VDD.n2 VDD.t3073 20.1899
R10907 VDD.n0 VDD.t375 20.1899
R10908 VDD.n0 VDD.t1245 20.1899
R10909 VDD.n56 VDD.t1742 20.1899
R10910 VDD.n56 VDD.t373 20.1899
R10911 VDD.n58 VDD.t2208 20.1899
R10912 VDD.n58 VDD.t1744 20.1899
R10913 VDD VDD.t1308 18.1744
R10914 VDD VDD.t4407 18.1744
R10915 VDD VDD.t2397 18.1744
R10916 VDD VDD.t658 18.1744
R10917 VDD VDD.t4474 18.1744
R10918 VDD VDD.t1191 18.1744
R10919 VDD VDD.t2850 18.1744
R10920 VDD VDD.t4391 18.1744
R10921 VDD VDD.t1888 18.1744
R10922 VDD VDD.t1868 18.1744
R10923 VDD VDD.t3575 18.1744
R10924 VDD.t3631 VDD 18.1744
R10925 VDD VDD.t3637 18.1744
R10926 VDD.t4364 VDD 18.1744
R10927 VDD VDD.t4510 18.1744
R10928 VDD VDD.t2696 18.1744
R10929 VDD VDD.t4395 18.1744
R10930 VDD VDD.t2547 18.1744
R10931 VDD VDD.t2864 18.1744
R10932 VDD VDD.t4467 18.1744
R10933 VDD VDD.t3334 18.1744
R10934 VDD VDD.t1442 18.1744
R10935 VDD VDD.t2025 18.1744
R10936 VDD VDD.t4476 18.1744
R10937 VDD VDD.t1451 18.1744
R10938 VDD VDD.t4444 18.1744
R10939 VDD VDD.t932 18.1744
R10940 VDD VDD.t1070 18.1744
R10941 VDD VDD.t4362 18.1744
R10942 VDD VDD.t372 18.1744
R10943 VDD.t78 VDD 18.1429
R10944 VDD VDD.t74 18.1429
R10945 VDD.t4419 VDD 18.1429
R10946 VDD VDD.t4446 18.1429
R10947 VDD.t3210 VDD 18.1429
R10948 VDD VDD.t3206 18.1429
R10949 VDD.t4371 VDD 18.1429
R10950 VDD VDD.t4415 18.1429
R10951 VDD.t2671 VDD 18.1429
R10952 VDD VDD.t2679 18.1429
R10953 VDD.t4506 VDD 18.1429
R10954 VDD VDD.t4489 18.1429
R10955 VDD.t3254 VDD 18.1429
R10956 VDD VDD.t3248 18.1429
R10957 VDD.t4427 VDD 18.1429
R10958 VDD VDD.t4399 18.1429
R10959 VDD.t3629 VDD 18.1429
R10960 VDD VDD.t3625 18.1429
R10961 VDD.t4429 VDD 18.1429
R10962 VDD VDD.t4401 18.1429
R10963 VDD.t183 VDD 18.1429
R10964 VDD VDD.t179 18.1429
R10965 VDD.t4381 VDD 18.1429
R10966 VDD VDD.t4343 18.1429
R10967 VDD.t2659 VDD 18.1429
R10968 VDD VDD.t2655 18.1429
R10969 VDD.t4434 VDD 18.1429
R10970 VDD VDD.t4403 18.1429
R10971 VDD.t567 VDD 18.1429
R10972 VDD VDD.t323 18.1429
R10973 VDD.t4387 VDD 18.1429
R10974 VDD VDD.t4349 18.1429
R10975 VDD.t646 VDD 18.1429
R10976 VDD VDD.t652 18.1429
R10977 VDD.t4341 VDD 18.1429
R10978 VDD VDD.t4375 18.1429
R10979 VDD.t3214 VDD 18.1114
R10980 VDD VDD.t3204 18.1114
R10981 VDD.t4360 VDD 18.1114
R10982 VDD.t2667 VDD 18.1114
R10983 VDD VDD.t2675 18.1114
R10984 VDD.t4501 VDD 18.1114
R10985 VDD.t3258 VDD 18.1114
R10986 VDD VDD.t3246 18.1114
R10987 VDD.t4422 VDD 18.1114
R10988 VDD.t191 VDD 18.1114
R10989 VDD VDD.t187 18.1114
R10990 VDD.t4424 VDD 18.1114
R10991 VDD.t2651 VDD 18.1114
R10992 VDD VDD.t2663 18.1114
R10993 VDD.t4497 VDD 18.1114
R10994 VDD.t327 VDD 18.1114
R10995 VDD VDD.t331 18.1114
R10996 VDD.t4503 VDD 18.1114
R10997 VDD.t66 VDD 18.1114
R10998 VDD VDD.t72 18.1114
R10999 VDD.t4411 VDD 18.1114
R11000 VDD.t644 VDD 18.1114
R11001 VDD VDD.t640 18.1114
R11002 VDD.t4339 VDD 18.1114
R11003 VDD.n2256 VDD 16.4024
R11004 VDD.n1914 VDD.n1913 16.3773
R11005 VDD.n2192 VDD.t137 16.3704
R11006 VDD.n2114 VDD.t363 16.3704
R11007 VDD.n2220 VDD 16.3534
R11008 VDD VDD.n2234 16.3534
R11009 VDD VDD.n1882 16.2755
R11010 VDD.n2231 VDD 16.2729
R11011 VDD.n2256 VDD 16.2724
R11012 VDD VDD.n1854 16.2724
R11013 VDD VDD.n2199 16.27
R11014 VDD VDD.n2223 16.27
R11015 VDD.n2257 VDD 16.27
R11016 VDD VDD.n2258 16.27
R11017 VDD VDD.n1874 16.27
R11018 VDD.n1873 VDD 16.27
R11019 VDD.n2222 VDD 16.2628
R11020 VDD VDD.n2233 16.2628
R11021 VDD VDD.n1862 16.2628
R11022 VDD.n2221 VDD 16.258
R11023 VDD.n2265 VDD 16.258
R11024 VDD.n1878 VDD 16.258
R11025 VDD VDD.n2198 16.2556
R11026 VDD.n1887 VDD 16.2556
R11027 VDD.n2220 VDD 16.2195
R11028 VDD VDD.n2234 16.2195
R11029 VDD.n1882 VDD 16.2195
R11030 VDD.n2339 VDD 16.21
R11031 VDD.n2306 VDD 16.1803
R11032 VDD.n2286 VDD 16.1803
R11033 VDD.n2161 VDD.n2156 16.1788
R11034 VDD.n2327 VDD 16.1769
R11035 VDD.n2296 VDD 16.1769
R11036 VDD.n1950 VDD.n1890 16.1752
R11037 VDD.n2317 VDD 16.1735
R11038 VDD.n2337 VDD 16.1702
R11039 VDD.n2276 VDD 16.1702
R11040 VDD.n1924 VDD.n1902 16.1382
R11041 VDD.n1917 VDD.n1914 16.1214
R11042 VDD.n1932 VDD.n1931 16.0978
R11043 VDD.n1949 VDD.n1948 16.0952
R11044 VDD.n1936 VDD.n1933 16.0952
R11045 VDD.n1943 VDD.n1891 16.0939
R11046 VDD.n151 VDD.n150 15.8946
R11047 VDD.n2196 VDD.n2195 15.847
R11048 VDD.n2183 VDD.n2119 15.847
R11049 VDD.n2178 VDD.n2177 15.847
R11050 VDD.n2176 VDD.n2175 15.847
R11051 VDD.n2171 VDD.n2170 15.847
R11052 VDD.n2166 VDD.n2165 15.847
R11053 VDD.n2161 VDD.n2160 15.847
R11054 VDD.n2117 VDD.n2116 15.847
R11055 VDD.n2050 VDD.n2039 15.847
R11056 VDD.n2086 VDD.n2085 15.847
R11057 VDD.n2091 VDD.n2090 15.847
R11058 VDD.n2096 VDD.n2095 15.847
R11059 VDD.n2101 VDD.n2100 15.847
R11060 VDD.n2106 VDD.n2105 15.847
R11061 VDD.n2111 VDD.n2110 15.847
R11062 VDD.n1884 VDD.t674 13.3599
R11063 VDD.t467 VDD.t135 13.0964
R11064 VDD.t137 VDD.t467 13.0964
R11065 VDD.t361 VDD.t365 13.0964
R11066 VDD.t363 VDD.t361 13.0964
R11067 VDD.n2833 VDD.t2293 11.8205
R11068 VDD.n2833 VDD.t3418 11.8205
R11069 VDD.n2834 VDD.t3426 11.8205
R11070 VDD.n1146 VDD.t1407 11.8205
R11071 VDD.n1147 VDD.t1411 11.8205
R11072 VDD.n1147 VDD.t1385 11.8205
R11073 VDD.n2842 VDD.t1760 11.8205
R11074 VDD.n2842 VDD.t1788 11.8205
R11075 VDD.n2843 VDD.t784 11.8205
R11076 VDD.n2838 VDD.t981 11.8205
R11077 VDD.n2839 VDD.t975 11.8205
R11078 VDD.n2839 VDD.t977 11.8205
R11079 VDD.n2848 VDD.t2295 11.8205
R11080 VDD.n2848 VDD.t3439 11.8205
R11081 VDD.n2849 VDD.t3448 11.8205
R11082 VDD.n1141 VDD.t3305 11.8205
R11083 VDD.n1143 VDD.t3309 11.8205
R11084 VDD.n1143 VDD.t3303 11.8205
R11085 VDD.n2748 VDD.t1746 11.8205
R11086 VDD.n2748 VDD.t1812 11.8205
R11087 VDD.n2749 VDD.t1772 11.8205
R11088 VDD.n2744 VDD.t1409 11.8205
R11089 VDD.n2745 VDD.t1405 11.8205
R11090 VDD.n2745 VDD.t1387 11.8205
R11091 VDD.n2759 VDD.t767 11.8205
R11092 VDD.n2759 VDD.t1808 11.8205
R11093 VDD.n2760 VDD.t1766 11.8205
R11094 VDD.n2755 VDD.t3555 11.8205
R11095 VDD.n2756 VDD.t3534 11.8205
R11096 VDD.n2756 VDD.t3565 11.8205
R11097 VDD.n2770 VDD.t1810 11.8205
R11098 VDD.n2770 VDD.t1798 11.8205
R11099 VDD.n2771 VDD.t1774 11.8205
R11100 VDD.n2766 VDD.t3967 11.8205
R11101 VDD.n2767 VDD.t892 11.8205
R11102 VDD.n2767 VDD.t3982 11.8205
R11103 VDD.n2781 VDD.t1786 11.8205
R11104 VDD.n2781 VDD.t1796 11.8205
R11105 VDD.n2782 VDD.t1748 11.8205
R11106 VDD.n2777 VDD.t3603 11.8205
R11107 VDD.n2778 VDD.t3583 11.8205
R11108 VDD.n2778 VDD.t3616 11.8205
R11109 VDD.n2792 VDD.t1780 11.8205
R11110 VDD.n2792 VDD.t780 11.8205
R11111 VDD.n2793 VDD.t1806 11.8205
R11112 VDD.n2788 VDD.t2131 11.8205
R11113 VDD.n2789 VDD.t2120 11.8205
R11114 VDD.n2789 VDD.t2169 11.8205
R11115 VDD.n2803 VDD.t1756 11.8205
R11116 VDD.n2803 VDD.t1804 11.8205
R11117 VDD.n2804 VDD.t1784 11.8205
R11118 VDD.n2799 VDD.t2604 11.8205
R11119 VDD.n2800 VDD.t2595 11.8205
R11120 VDD.n2800 VDD.t2580 11.8205
R11121 VDD.n2814 VDD.t1750 11.8205
R11122 VDD.n2814 VDD.t1800 11.8205
R11123 VDD.n2815 VDD.t1778 11.8205
R11124 VDD.n2810 VDD.t2354 11.8205
R11125 VDD.n2811 VDD.t2342 11.8205
R11126 VDD.n2811 VDD.t2325 11.8205
R11127 VDD.n2825 VDD.t765 11.8205
R11128 VDD.n2825 VDD.t1792 11.8205
R11129 VDD.n2826 VDD.t1764 11.8205
R11130 VDD.n2821 VDD.t1005 11.8205
R11131 VDD.n2822 VDD.t994 11.8205
R11132 VDD.n2822 VDD.t1033 11.8205
R11133 VDD.n2738 VDD.t3640 11.8205
R11134 VDD.n2738 VDD.t3646 11.8205
R11135 VDD.n2739 VDD.t3642 11.8205
R11136 VDD.n1157 VDD.t3428 11.8205
R11137 VDD.n1158 VDD.t3422 11.8205
R11138 VDD.n1158 VDD.t3445 11.8205
R11139 VDD.n2732 VDD.t3478 11.8205
R11140 VDD.n2732 VDD.t3470 11.8205
R11141 VDD.n2733 VDD.t3472 11.8205
R11142 VDD.n2728 VDD.t1875 11.8205
R11143 VDD.n2729 VDD.t1873 11.8205
R11144 VDD.n2729 VDD.t173 11.8205
R11145 VDD.n2722 VDD.t3233 11.8205
R11146 VDD.n2722 VDD.t3237 11.8205
R11147 VDD.n2723 VDD.t3235 11.8205
R11148 VDD.n2719 VDD.t2818 11.8205
R11149 VDD.n2720 VDD.t2835 11.8205
R11150 VDD.n2720 VDD.t2828 11.8205
R11151 VDD.n1984 VDD.t2813 11.8205
R11152 VDD.n1984 VDD.t2815 11.8205
R11153 VDD.n1985 VDD.t2826 11.8205
R11154 VDD.n1987 VDD.t3549 11.8205
R11155 VDD.n1988 VDD.t3563 11.8205
R11156 VDD.n1988 VDD.t3538 11.8205
R11157 VDD.n2003 VDD.t384 11.8205
R11158 VDD.n2003 VDD.t386 11.8205
R11159 VDD.n2004 VDD.t402 11.8205
R11160 VDD.n2006 VDD.t3969 11.8205
R11161 VDD.n2007 VDD.t3980 11.8205
R11162 VDD.n2007 VDD.t894 11.8205
R11163 VDD.n1981 VDD.t2196 11.8205
R11164 VDD.n1981 VDD.t1632 11.8205
R11165 VDD.n1982 VDD.t2194 11.8205
R11166 VDD.n2013 VDD.t3585 11.8205
R11167 VDD.n2014 VDD.t3605 11.8205
R11168 VDD.n2014 VDD.t3619 11.8205
R11169 VDD.n1974 VDD.t4078 11.8205
R11170 VDD.n1974 VDD.t4090 11.8205
R11171 VDD.n1975 VDD.t4120 11.8205
R11172 VDD.n1977 VDD.t2181 11.8205
R11173 VDD.n1978 VDD.t2133 11.8205
R11174 VDD.n1978 VDD.t2152 11.8205
R11175 VDD.n2023 VDD.t538 11.8205
R11176 VDD.n2023 VDD.t540 11.8205
R11177 VDD.n2024 VDD.t526 11.8205
R11178 VDD.n2026 VDD.t484 11.8205
R11179 VDD.n2027 VDD.t2589 11.8205
R11180 VDD.n2027 VDD.t2610 11.8205
R11181 VDD.n1963 VDD.t4197 11.8205
R11182 VDD.n1963 VDD.t4215 11.8205
R11183 VDD.n1964 VDD.t4231 11.8205
R11184 VDD.n2033 VDD.t2346 11.8205
R11185 VDD.n2034 VDD.t1832 11.8205
R11186 VDD.n2034 VDD.t2317 11.8205
R11187 VDD.n1990 VDD.t2291 11.8205
R11188 VDD.n1990 VDD.t2297 11.8205
R11189 VDD.n1991 VDD.t3443 11.8205
R11190 VDD.n1993 VDD.t1397 11.8205
R11191 VDD.n1994 VDD.t1413 11.8205
R11192 VDD.n1994 VDD.t1177 11.8205
R11193 VDD.n1966 VDD.t1660 11.8205
R11194 VDD.n1966 VDD.t1680 11.8205
R11195 VDD.n1967 VDD.t1658 11.8205
R11196 VDD.n1969 VDD.t988 11.8205
R11197 VDD.n1970 VDD.t1038 11.8205
R11198 VDD.n1970 VDD.t592 11.8205
R11199 VDD.n2350 VDD.t1941 11.8205
R11200 VDD.n2350 VDD.t1937 11.8205
R11201 VDD.n2351 VDD.t1913 11.8205
R11202 VDD.n1179 VDD.t1608 11.8205
R11203 VDD.n1180 VDD.t1612 11.8205
R11204 VDD.n1180 VDD.t635 11.8205
R11205 VDD.n2359 VDD.t499 11.8205
R11206 VDD.n2359 VDD.t501 11.8205
R11207 VDD.n2360 VDD.t2736 11.8205
R11208 VDD.n2355 VDD.t2568 11.8205
R11209 VDD.n2356 VDD.t2556 11.8205
R11210 VDD.n2356 VDD.t2558 11.8205
R11211 VDD.n1176 VDD.t2918 11.8205
R11212 VDD.n1176 VDD.t2920 11.8205
R11213 VDD.n1177 VDD.t2922 11.8205
R11214 VDD.n1173 VDD.t246 11.8205
R11215 VDD.n1174 VDD.t250 11.8205
R11216 VDD.n1174 VDD.t252 11.8205
R11217 VDD.n1357 VDD.t1333 11.8205
R11218 VDD.n1357 VDD.t1341 11.8205
R11219 VDD.n1358 VDD.t1339 11.8205
R11220 VDD.n1354 VDD.t2311 11.8205
R11221 VDD.n1355 VDD.t2309 11.8205
R11222 VDD.n1355 VDD.t2313 11.8205
R11223 VDD.n1788 VDD.t4178 11.8205
R11224 VDD.n1788 VDD.t4184 11.8205
R11225 VDD.n1789 VDD.t4172 11.8205
R11226 VDD.n1360 VDD.t2418 11.8205
R11227 VDD.n1361 VDD.t212 11.8205
R11228 VDD.n1361 VDD.t214 11.8205
R11229 VDD.n1373 VDD.t290 11.8205
R11230 VDD.n1373 VDD.t286 11.8205
R11231 VDD.n1374 VDD.t288 11.8205
R11232 VDD.n1370 VDD.t1298 11.8205
R11233 VDD.n1371 VDD.t1302 11.8205
R11234 VDD.n1371 VDD.t1292 11.8205
R11235 VDD.n1379 VDD.t2059 11.8205
R11236 VDD.n1379 VDD.t2061 11.8205
R11237 VDD.n1380 VDD.t1602 11.8205
R11238 VDD.n1376 VDD.t1983 11.8205
R11239 VDD.n1377 VDD.t1975 11.8205
R11240 VDD.n1377 VDD.t1963 11.8205
R11241 VDD.n1796 VDD.t452 11.8205
R11242 VDD.n1796 VDD.t456 11.8205
R11243 VDD.n1797 VDD.t458 11.8205
R11244 VDD.n1793 VDD.t705 11.8205
R11245 VDD.n1794 VDD.t709 11.8205
R11246 VDD.n1794 VDD.t711 11.8205
R11247 VDD.n1442 VDD.t4063 11.8205
R11248 VDD.n1442 VDD.t4061 11.8205
R11249 VDD.n1443 VDD.t4055 11.8205
R11250 VDD.n1438 VDD.t3317 11.8205
R11251 VDD.n1439 VDD.t3313 11.8205
R11252 VDD.n1439 VDD.t3311 11.8205
R11253 VDD.n1435 VDD.t3658 11.8205
R11254 VDD.n1435 VDD.t3654 11.8205
R11255 VDD.n1436 VDD.t3656 11.8205
R11256 VDD.n1432 VDD.t937 11.8205
R11257 VDD.n1433 VDD.t939 11.8205
R11258 VDD.n1433 VDD.t935 11.8205
R11259 VDD.n1628 VDD.t1816 11.8205
R11260 VDD.n1628 VDD.t161 11.8205
R11261 VDD.n1629 VDD.t157 11.8205
R11262 VDD.n1428 VDD.t2450 11.8205
R11263 VDD.n1429 VDD.t2448 11.8205
R11264 VDD.n1429 VDD.t2446 11.8205
R11265 VDD.n1637 VDD.t1280 11.8205
R11266 VDD.n1637 VDD.t1278 11.8205
R11267 VDD.n1638 VDD.t1276 11.8205
R11268 VDD.n1633 VDD.t831 11.8205
R11269 VDD.n1634 VDD.t841 11.8205
R11270 VDD.n1634 VDD.t839 11.8205
R11271 VDD.n1645 VDD.t1905 11.8205
R11272 VDD.n1645 VDD.t1897 11.8205
R11273 VDD.n1646 VDD.t1903 11.8205
R11274 VDD.n1642 VDD.t4019 11.8205
R11275 VDD.n1643 VDD.t4013 11.8205
R11276 VDD.n1643 VDD.t4011 11.8205
R11277 VDD.n1655 VDD.t2009 11.8205
R11278 VDD.n1655 VDD.t2019 11.8205
R11279 VDD.n1656 VDD.t2017 11.8205
R11280 VDD.n1651 VDD.t2777 11.8205
R11281 VDD.n1652 VDD.t2775 11.8205
R11282 VDD.n1652 VDD.t2773 11.8205
R11283 VDD.n1664 VDD.t1073 11.8205
R11284 VDD.n1664 VDD.t1885 11.8205
R11285 VDD.n1665 VDD.t1883 11.8205
R11286 VDD.n1660 VDD.t3515 11.8205
R11287 VDD.n1661 VDD.t3513 11.8205
R11288 VDD.n1661 VDD.t3523 11.8205
R11289 VDD.n1670 VDD.t3392 11.8205
R11290 VDD.n1670 VDD.t3394 11.8205
R11291 VDD.n1671 VDD.t3390 11.8205
R11292 VDD.n1425 VDD.t1947 11.8205
R11293 VDD.n1426 VDD.t1955 11.8205
R11294 VDD.n1426 VDD.t1959 11.8205
R11295 VDD.n1605 VDD.t2719 11.8205
R11296 VDD.n1605 VDD.t2723 11.8205
R11297 VDD.n1606 VDD.t2715 11.8205
R11298 VDD.n1601 VDD.t4272 11.8205
R11299 VDD.n1602 VDD.t3935 11.8205
R11300 VDD.n1602 VDD.t4313 11.8205
R11301 VDD.n1614 VDD.t1055 11.8205
R11302 VDD.n1614 VDD.t1045 11.8205
R11303 VDD.n1615 VDD.t1047 11.8205
R11304 VDD.n1610 VDD.t4151 11.8205
R11305 VDD.n1611 VDD.t4157 11.8205
R11306 VDD.n1611 VDD.t4159 11.8205
R11307 VDD.n1457 VDD.t4035 11.8205
R11308 VDD.n1457 VDD.t4037 11.8205
R11309 VDD.n1458 VDD.t4029 11.8205
R11310 VDD.n1454 VDD.t19 11.8205
R11311 VDD.n1455 VDD.t23 11.8205
R11312 VDD.n1455 VDD.t27 11.8205
R11313 VDD.n1596 VDD.t665 11.8205
R11314 VDD.n1596 VDD.t671 11.8205
R11315 VDD.n1597 VDD.t673 11.8205
R11316 VDD.n1592 VDD.t3672 11.8205
R11317 VDD.n1593 VDD.t3676 11.8205
R11318 VDD.n1593 VDD.t3680 11.8205
R11319 VDD.n1586 VDD.t3272 11.8205
R11320 VDD.n1586 VDD.t3278 11.8205
R11321 VDD.n1587 VDD.t3276 11.8205
R11322 VDD.n1583 VDD.t114 11.8205
R11323 VDD.n1584 VDD.t112 11.8205
R11324 VDD.n1584 VDD.t116 11.8205
R11325 VDD.n1578 VDD.t3892 11.8205
R11326 VDD.n1578 VDD.t3884 11.8205
R11327 VDD.n1579 VDD.t3886 11.8205
R11328 VDD.n1574 VDD.t4282 11.8205
R11329 VDD.n1575 VDD.t4284 11.8205
R11330 VDD.n1575 VDD.t4288 11.8205
R11331 VDD.n1569 VDD.t2508 11.8205
R11332 VDD.n1569 VDD.t2502 11.8205
R11333 VDD.n1570 VDD.t2506 11.8205
R11334 VDD.n1565 VDD.t3197 11.8205
R11335 VDD.n1566 VDD.t3199 11.8205
R11336 VDD.n1566 VDD.t3191 11.8205
R11337 VDD.n1463 VDD.t1591 11.8205
R11338 VDD.n1463 VDD.t598 11.8205
R11339 VDD.n1464 VDD.t600 11.8205
R11340 VDD.n1460 VDD.t1971 11.8205
R11341 VDD.n1461 VDD.t1961 11.8205
R11342 VDD.n1461 VDD.t1949 11.8205
R11343 VDD.n2714 VDD.t2400 11.8205
R11344 VDD.n2714 VDD.t823 11.8205
R11345 VDD.n2715 VDD.t2410 11.8205
R11346 VDD.n1160 VDD.t1145 11.8205
R11347 VDD.n1161 VDD.t1124 11.8205
R11348 VDD.n1161 VDD.t1147 11.8205
R11349 VDD.n2655 VDD.t2877 11.8205
R11350 VDD.n2655 VDD.t2873 11.8205
R11351 VDD.n2656 VDD.t2875 11.8205
R11352 VDD.n2652 VDD.t388 11.8205
R11353 VDD.n2653 VDD.t380 11.8205
R11354 VDD.n2653 VDD.t396 11.8205
R11355 VDD.n2425 VDD.t3905 11.8205
R11356 VDD.n2425 VDD.t3901 11.8205
R11357 VDD.n2426 VDD.t3913 11.8205
R11358 VDD.n2422 VDD.t2749 11.8205
R11359 VDD.n2423 VDD.t2755 11.8205
R11360 VDD.n2423 VDD.t2751 11.8205
R11361 VDD.n2646 VDD.t1428 11.8205
R11362 VDD.n2646 VDD.t1430 11.8205
R11363 VDD.n2647 VDD.t1438 11.8205
R11364 VDD.n2643 VDD.t2202 11.8205
R11365 VDD.n2644 VDD.t2192 11.8205
R11366 VDD.n2644 VDD.t1636 11.8205
R11367 VDD.n2638 VDD.t348 11.8205
R11368 VDD.n2638 VDD.t304 11.8205
R11369 VDD.n2639 VDD.t352 11.8205
R11370 VDD.n2428 VDD.t3939 11.8205
R11371 VDD.n2429 VDD.t3951 11.8205
R11372 VDD.n2429 VDD.t3947 11.8205
R11373 VDD.n2591 VDD.t618 11.8205
R11374 VDD.n2591 VDD.t610 11.8205
R11375 VDD.n2592 VDD.t622 11.8205
R11376 VDD.n2588 VDD.t4122 11.8205
R11377 VDD.n2589 VDD.t4102 11.8205
R11378 VDD.n2589 VDD.t4084 11.8205
R11379 VDD.n2445 VDD.t1551 11.8205
R11380 VDD.n2445 VDD.t1553 11.8205
R11381 VDD.n2446 VDD.t1555 11.8205
R11382 VDD.n2442 VDD.t1740 11.8205
R11383 VDD.n2443 VDD.t1732 11.8205
R11384 VDD.n2443 VDD.t1730 11.8205
R11385 VDD.n2582 VDD.t346 11.8205
R11386 VDD.n2582 VDD.t340 11.8205
R11387 VDD.n2583 VDD.t879 11.8205
R11388 VDD.n2579 VDD.t530 11.8205
R11389 VDD.n2580 VDD.t268 11.8205
R11390 VDD.n2580 VDD.t550 11.8205
R11391 VDD.n2574 VDD.t2463 11.8205
R11392 VDD.n2574 VDD.t2461 11.8205
R11393 VDD.n2575 VDD.t2436 11.8205
R11394 VDD.n2448 VDD.t89 11.8205
R11395 VDD.n2449 VDD.t87 11.8205
R11396 VDD.n2449 VDD.t91 11.8205
R11397 VDD.n2503 VDD.t757 11.8205
R11398 VDD.n2503 VDD.t755 11.8205
R11399 VDD.n2504 VDD.t761 11.8205
R11400 VDD.n2499 VDD.t2625 11.8205
R11401 VDD.n2500 VDD.t2631 11.8205
R11402 VDD.n2500 VDD.t2629 11.8205
R11403 VDD.n2512 VDD.t2089 11.8205
R11404 VDD.n2512 VDD.t2083 11.8205
R11405 VDD.n2513 VDD.t2095 11.8205
R11406 VDD.n2508 VDD.t1678 11.8205
R11407 VDD.n2509 VDD.t2245 11.8205
R11408 VDD.n2509 VDD.t2232 11.8205
R11409 VDD.n2487 VDD.t2261 11.8205
R11410 VDD.n2487 VDD.t2259 11.8205
R11411 VDD.n2488 VDD.t2265 11.8205
R11412 VDD.n2484 VDD.t1752 11.8205
R11413 VDD.n2485 VDD.t1768 11.8205
R11414 VDD.n2485 VDD.t1794 11.8205
R11415 VDD.n2493 VDD.t4143 11.8205
R11416 VDD.n2493 VDD.t4141 11.8205
R11417 VDD.n2494 VDD.t4145 11.8205
R11418 VDD.n2490 VDD.t4200 11.8205
R11419 VDD.n2491 VDD.t4226 11.8205
R11420 VDD.n2491 VDD.t4233 11.8205
R11421 VDD.n2834 VDD.t3451 10.3878
R11422 VDD.n1146 VDD.t1392 10.3878
R11423 VDD.n2843 VDD.t1782 10.3878
R11424 VDD.n2838 VDD.t979 10.3878
R11425 VDD.n2849 VDD.t3424 10.3878
R11426 VDD.n1141 VDD.t3301 10.3878
R11427 VDD.n2749 VDD.t1790 10.3878
R11428 VDD.n2744 VDD.t1175 10.3878
R11429 VDD.n2760 VDD.t1754 10.3878
R11430 VDD.n2755 VDD.t3530 10.3878
R11431 VDD.n2771 VDD.t778 10.3878
R11432 VDD.n2766 VDD.t3973 10.3878
R11433 VDD.n2782 VDD.t1814 10.3878
R11434 VDD.n2777 VDD.t3597 10.3878
R11435 VDD.n2793 VDD.t1758 10.3878
R11436 VDD.n2788 VDD.t2156 10.3878
R11437 VDD.n2804 VDD.t763 10.3878
R11438 VDD.n2799 VDD.t2574 10.3878
R11439 VDD.n2815 VDD.t782 10.3878
R11440 VDD.n2810 VDD.t1834 10.3878
R11441 VDD.n2826 VDD.t776 10.3878
R11442 VDD.n2821 VDD.t586 10.3878
R11443 VDD.n2739 VDD.t3652 10.3878
R11444 VDD.n1157 VDD.t3441 10.3878
R11445 VDD.n2733 VDD.t3468 10.3878
R11446 VDD.n2728 VDD.t1877 10.3878
R11447 VDD.n2723 VDD.t3245 10.3878
R11448 VDD.n2719 VDD.t2824 10.3878
R11449 VDD.n1985 VDD.t2844 10.3878
R11450 VDD.n1987 VDD.t3540 10.3878
R11451 VDD.n2004 VDD.t377 10.3878
R11452 VDD.n2006 VDD.t898 10.3878
R11453 VDD.n1982 VDD.t2200 10.3878
R11454 VDD.n2013 VDD.t3580 10.3878
R11455 VDD.n1975 VDD.t4074 10.3878
R11456 VDD.n1977 VDD.t2154 10.3878
R11457 VDD.n2024 VDD.t270 10.3878
R11458 VDD.n2026 VDD.t480 10.3878
R11459 VDD.n1964 VDD.t4195 10.3878
R11460 VDD.n2033 VDD.t2319 10.3878
R11461 VDD.n1991 VDD.t2289 10.3878
R11462 VDD.n1993 VDD.t1181 10.3878
R11463 VDD.n1967 VDD.t1673 10.3878
R11464 VDD.n1969 VDD.t596 10.3878
R11465 VDD.n2351 VDD.t1939 10.3878
R11466 VDD.n1179 VDD.t639 10.3878
R11467 VDD.n2360 VDD.t495 10.3878
R11468 VDD.n2355 VDD.t2560 10.3878
R11469 VDD.n1177 VDD.t2912 10.3878
R11470 VDD.n1173 VDD.t256 10.3878
R11471 VDD.n1358 VDD.t1343 10.3878
R11472 VDD.n1354 VDD.t2307 10.3878
R11473 VDD.n1789 VDD.t4180 10.3878
R11474 VDD.n1360 VDD.t216 10.3878
R11475 VDD.n1374 VDD.t292 10.3878
R11476 VDD.n1370 VDD.t1290 10.3878
R11477 VDD.n1380 VDD.t2055 10.3878
R11478 VDD.n1376 VDD.t1925 10.3878
R11479 VDD.n1797 VDD.t454 10.3878
R11480 VDD.n1793 VDD.t3989 10.3878
R11481 VDD.n1443 VDD.t4051 10.3878
R11482 VDD.n1438 VDD.t3319 10.3878
R11483 VDD.n1436 VDD.t3666 10.3878
R11484 VDD.n1432 VDD.t941 10.3878
R11485 VDD.n1629 VDD.t151 10.3878
R11486 VDD.n1428 VDD.t2440 10.3878
R11487 VDD.n1638 VDD.t1288 10.3878
R11488 VDD.n1633 VDD.t833 10.3878
R11489 VDD.n1646 VDD.t1899 10.3878
R11490 VDD.n1642 VDD.t4015 10.3878
R11491 VDD.n1656 VDD.t2015 10.3878
R11492 VDD.n1651 VDD.t2781 10.3878
R11493 VDD.n1665 VDD.t1075 10.3878
R11494 VDD.n1660 VDD.t3519 10.3878
R11495 VDD.n1671 VDD.t3388 10.3878
R11496 VDD.n1425 VDD.t1935 10.3878
R11497 VDD.n1606 VDD.t2721 10.3878
R11498 VDD.n1601 VDD.t4311 10.3878
R11499 VDD.n1615 VDD.t1053 10.3878
R11500 VDD.n1610 VDD.t4161 10.3878
R11501 VDD.n1458 VDD.t4033 10.3878
R11502 VDD.n1454 VDD.t29 10.3878
R11503 VDD.n1597 VDD.t667 10.3878
R11504 VDD.n1592 VDD.t3668 10.3878
R11505 VDD.n1587 VDD.t3495 10.3878
R11506 VDD.n1583 VDD.t110 10.3878
R11507 VDD.n1579 VDD.t3894 10.3878
R11508 VDD.n1574 VDD.t4290 10.3878
R11509 VDD.n1570 VDD.t2510 10.3878
R11510 VDD.n1565 VDD.t3189 10.3878
R11511 VDD.n1464 VDD.t604 10.3878
R11512 VDD.n1460 VDD.t1917 10.3878
R11513 VDD.n2715 VDD.t2404 10.3878
R11514 VDD.n1160 VDD.t1116 10.3878
R11515 VDD.n2656 VDD.t2885 10.3878
R11516 VDD.n2652 VDD.t392 10.3878
R11517 VDD.n2426 VDD.t3903 10.3878
R11518 VDD.n2422 VDD.t2753 10.3878
R11519 VDD.n2647 VDD.t1426 10.3878
R11520 VDD.n2643 VDD.t1639 10.3878
R11521 VDD.n2639 VDD.t350 10.3878
R11522 VDD.n2428 VDD.t3949 10.3878
R11523 VDD.n2592 VDD.t620 10.3878
R11524 VDD.n2588 VDD.t4100 10.3878
R11525 VDD.n2446 VDD.t1557 10.3878
R11526 VDD.n2442 VDD.t1728 10.3878
R11527 VDD.n2583 VDD.t877 10.3878
R11528 VDD.n2579 VDD.t262 10.3878
R11529 VDD.n2575 VDD.t2465 10.3878
R11530 VDD.n2448 VDD.t93 10.3878
R11531 VDD.n2504 VDD.t759 10.3878
R11532 VDD.n2499 VDD.t2627 10.3878
R11533 VDD.n2513 VDD.t2087 10.3878
R11534 VDD.n2508 VDD.t2228 10.3878
R11535 VDD.n2488 VDD.t2263 10.3878
R11536 VDD.n2484 VDD.t1802 10.3878
R11537 VDD.n2494 VDD.t4147 10.3878
R11538 VDD.n2490 VDD.t4222 10.3878
R11539 VDD.n681 VDD 9.42895
R11540 VDD VDD.n2111 9.3597
R11541 VDD VDD.n2118 9.10566
R11542 VDD.n2218 VDD.t2339 8.72225
R11543 VDD.t2478 VDD.n2243 8.72225
R11544 VDD.n1193 VDD.n1185 7.98309
R11545 VDD.n1325 VDD.n1324 7.9105
R11546 VDD.n1313 VDD.n1312 7.9105
R11547 VDD.n1301 VDD.n1300 7.9105
R11548 VDD.n1289 VDD.n1288 7.9105
R11549 VDD.n1277 VDD.n1276 7.9105
R11550 VDD.n1265 VDD.n1264 7.9105
R11551 VDD.n1253 VDD.n1252 7.9105
R11552 VDD.n1241 VDD.n1240 7.9105
R11553 VDD.n1229 VDD.n1228 7.9105
R11554 VDD.n1217 VDD.n1216 7.9105
R11555 VDD.n1204 VDD.n1203 7.9105
R11556 VDD.n2372 VDD.n2371 7.9105
R11557 VDD.n2381 VDD.n1163 7.9105
R11558 VDD.n2406 VDD.n2405 7.9105
R11559 VDD.n2399 VDD.n2385 7.9105
R11560 VDD.n669 VDD.t2420 7.59513
R11561 VDD.n669 VDD.t2419 7.59513
R11562 VDD.n668 VDD.t2004 7.59513
R11563 VDD.n668 VDD.t2002 7.59513
R11564 VDD.n1062 VDD.t1521 6.98579
R11565 VDD.n933 VDD.t3914 6.98579
R11566 VDD.n804 VDD.t3458 6.98579
R11567 VDD.n653 VDD.t3343 6.98579
R11568 VDD.n524 VDD.t2541 6.98579
R11569 VDD.n395 VDD.t2708 6.98579
R11570 VDD.n266 VDD.t1687 6.98579
R11571 VDD.n128 VDD.t1103 6.98579
R11572 VDD.n2912 VDD.t3296 6.98579
R11573 VDD.n2538 VDD.n2537 4.98339
R11574 VDD.n2682 VDD.n2677 4.98339
R11575 VDD.n2666 VDD.n2665 4.98339
R11576 VDD.n2635 VDD.n2433 4.98339
R11577 VDD.n2602 VDD.n2601 4.98339
R11578 VDD.n2571 VDD.n2453 4.98339
R11579 VDD.n2522 VDD.n2521 4.98339
R11580 VDD.n2693 VDD.n2692 4.89827
R11581 VDD.n2710 VDD.n2416 4.89827
R11582 VDD.n2620 VDD.n2421 4.89827
R11583 VDD.n2634 VDD.n2436 4.89827
R11584 VDD.n2556 VDD.n2441 4.89827
R11585 VDD.n2570 VDD.n2456 4.89827
R11586 VDD.n2536 VDD.n2464 4.89827
R11587 VDD.n2483 VDD.n2471 4.89827
R11588 VDD.n2700 VDD.n2413 4.87738
R11589 VDD.n1677 VDD.n1424 4.75
R11590 VDD.n1559 VDD.n1468 4.75
R11591 VDD.n1403 VDD.n1391 4.75
R11592 VDD.n2536 VDD.n2535 4.52383
R11593 VDD.n2692 VDD.n2691 4.52383
R11594 VDD.n2710 VDD.n2709 4.52383
R11595 VDD.n1403 VDD.n1402 4.52383
R11596 VDD.n1709 VDD.n1708 4.52383
R11597 VDD.n1783 VDD.n1782 4.52383
R11598 VDD.n1716 VDD.n1364 4.52383
R11599 VDD.n1773 VDD.n1352 4.52383
R11600 VDD.n1757 VDD.n1756 4.52383
R11601 VDD.n1766 VDD.n1351 4.52383
R11602 VDD.n1753 VDD.n1752 4.52383
R11603 VDD.n1830 VDD.n1829 4.52383
R11604 VDD.n1833 VDD.n1832 4.52383
R11605 VDD.n1820 VDD.n1339 4.52383
R11606 VDD.n1678 VDD.n1677 4.52383
R11607 VDD.n1687 VDD.n1412 4.52383
R11608 VDD.n1692 VDD.n1413 4.52383
R11609 VDD.n1702 VDD.n1701 4.52383
R11610 VDD.n1813 VDD.n1812 4.52383
R11611 VDD.n1853 VDD.n1852 4.52383
R11612 VDD.n1841 VDD.n1840 4.52383
R11613 VDD.n1843 VDD.n1842 4.52383
R11614 VDD.n1509 VDD.n1508 4.52383
R11615 VDD.n1501 VDD.n1451 4.52383
R11616 VDD.n1518 VDD.n1347 4.52383
R11617 VDD.n1559 VDD.n1558 4.52383
R11618 VDD.n1549 VDD.n1407 4.52383
R11619 VDD.n1533 VDD.n1532 4.52383
R11620 VDD.n1542 VDD.n1408 4.52383
R11621 VDD.n1525 VDD.n1348 4.52383
R11622 VDD.n1477 VDD.n1278 4.52383
R11623 VDD.n1494 VDD.n1452 4.52383
R11624 VDD.n1485 VDD.n1484 4.52383
R11625 VDD.n1733 VDD.n1230 4.52383
R11626 VDD.n1745 VDD.n1744 4.52383
R11627 VDD.n1743 VDD.n1742 4.52383
R11628 VDD.n2611 VDD.n2421 4.52383
R11629 VDD.n2634 VDD.n2633 4.52383
R11630 VDD.n2547 VDD.n2441 4.52383
R11631 VDD.n2570 VDD.n2569 4.52383
R11632 VDD.n2483 VDD.n2482 4.52383
R11633 VDD.n687 VDD.n686 3.9555
R11634 VDD.n1885 VDD.n1884 3.46404
R11635 VDD.n1063 VDD.n1062 3.29339
R11636 VDD.n934 VDD.n933 3.29339
R11637 VDD.n805 VDD.n804 3.29339
R11638 VDD.n654 VDD.n653 3.29339
R11639 VDD.n525 VDD.n524 3.29339
R11640 VDD.n396 VDD.n395 3.29339
R11641 VDD.n267 VDD.n266 3.29339
R11642 VDD.n129 VDD.n128 3.29339
R11643 VDD.n2913 VDD.n2912 3.29339
R11644 VDD.n1021 VDD.t4353 1.95523
R11645 VDD.n1017 VDD.t3733 1.95523
R11646 VDD.n892 VDD.t4373 1.95523
R11647 VDD.n888 VDD.t3789 1.95523
R11648 VDD.n763 VDD.t4448 1.95523
R11649 VDD.n759 VDD.t3791 1.95523
R11650 VDD.n612 VDD.t4355 1.95523
R11651 VDD.n608 VDD.t3722 1.95523
R11652 VDD.n483 VDD.t4345 1.95523
R11653 VDD.n479 VDD.t3708 1.95523
R11654 VDD.n354 VDD.t4357 1.95523
R11655 VDD.n350 VDD.t3724 1.95523
R11656 VDD.n225 VDD.t4347 1.95523
R11657 VDD.n221 VDD.t3714 1.95523
R11658 VDD.n87 VDD.t4409 1.95523
R11659 VDD.n83 VDD.t3729 1.95523
R11660 VDD.n25 VDD.t4405 1.95523
R11661 VDD.n21 VDD.t3727 1.95523
R11662 VDD.n1124 VDD.n1123 1.92718
R11663 VDD.n995 VDD.n994 1.92718
R11664 VDD.n866 VDD.n865 1.92718
R11665 VDD.n737 VDD.n736 1.92718
R11666 VDD.n586 VDD.n585 1.92718
R11667 VDD.n457 VDD.n456 1.92718
R11668 VDD.n328 VDD.n327 1.92718
R11669 VDD.n199 VDD.n198 1.92718
R11670 VDD.n2904 VDD.n2903 1.92718
R11671 VDD.n1072 VDD.n1071 1.92682
R11672 VDD.n943 VDD.n942 1.92682
R11673 VDD.n814 VDD.n813 1.92682
R11674 VDD.n663 VDD.n662 1.92682
R11675 VDD.n534 VDD.n533 1.92682
R11676 VDD.n405 VDD.n404 1.92682
R11677 VDD.n276 VDD.n275 1.92682
R11678 VDD.n138 VDD.n137 1.92682
R11679 VDD.n2922 VDD.n2921 1.92682
R11680 VDD VDD.n1960 1.91624
R11681 VDD VDD.n2336 1.91624
R11682 VDD VDD.n2326 1.91624
R11683 VDD VDD.n2316 1.91624
R11684 VDD VDD.n2305 1.91624
R11685 VDD VDD.n2295 1.91624
R11686 VDD VDD.n2285 1.91624
R11687 VDD VDD.n2275 1.91624
R11688 VDD.n2854 VDD 1.82215
R11689 VDD.t1056 VDD.n2382 1.79974
R11690 VDD.n2407 VDD.t236 1.79974
R11691 VDD.n2400 VDD.t1157 1.79974
R11692 VDD.n140 VDD.n139 1.76513
R11693 VDD.n1074 VDD.n1073 1.7634
R11694 VDD.n945 VDD.n944 1.7634
R11695 VDD.n816 VDD.n815 1.7634
R11696 VDD.n665 VDD.n664 1.7634
R11697 VDD.n536 VDD.n535 1.7634
R11698 VDD.n407 VDD.n406 1.7634
R11699 VDD.n278 VDD.n277 1.7634
R11700 VDD.n2906 VDD.n2905 1.7634
R11701 VDD.n2118 VDD.n2117 1.68666
R11702 VDD.n2413 VDD.n2412 1.57187
R11703 VDD.n1023 VDD.n1022 1.50655
R11704 VDD.n894 VDD.n893 1.50655
R11705 VDD.n765 VDD.n764 1.50655
R11706 VDD.n614 VDD.n613 1.50655
R11707 VDD.n485 VDD.n484 1.50655
R11708 VDD.n356 VDD.n355 1.50655
R11709 VDD.n227 VDD.n226 1.50655
R11710 VDD.n89 VDD.n88 1.50655
R11711 VDD.n27 VDD.n26 1.50655
R11712 VDD.n1999 VDD.n1998 1.46141
R11713 VDD.n1313 VDD.n1305 1.36656
R11714 VDD.n1217 VDD.n1209 1.36638
R11715 VDD.n1265 VDD.n1257 1.36637
R11716 VDD.n1204 VDD.n1196 1.36607
R11717 VDD.n2392 VDD.n2385 1.36269
R11718 VDD.n1289 VDD.n1281 1.34299
R11719 VDD.n1241 VDD.n1233 1.34283
R11720 VDD.n2411 VDD.n2410 1.29371
R11721 VDD.n2404 VDD.n2403 1.29371
R11722 VDD.n2374 VDD.n2373 1.29371
R11723 VDD.n1317 VDD.n1314 1.29371
R11724 VDD.n1293 VDD.n1290 1.29371
R11725 VDD.n1269 VDD.n1266 1.29371
R11726 VDD.n1245 VDD.n1242 1.29371
R11727 VDD.n1221 VDD.n1218 1.29371
R11728 VDD.n1193 VDD.n1192 1.29371
R11729 VDD.n2198 VDD.n2197 1.17983
R11730 VDD.n2038 VDD.n1962 1.09646
R11731 VDD.n2019 VDD.n2018 1.02596
R11732 VDD.n2018 VDD.n1980 0.975598
R11733 VDD.n1999 VDD.n1980 0.966646
R11734 VDD.n2019 VDD.n1962 0.955456
R11735 VDD.n2338 VDD.n2232 0.94433
R11736 VDD.n2232 VDD.n1961 0.890873
R11737 VDD.n2190 VDD.n2189 0.808212
R11738 VDD.n2112 VDD.n2081 0.808212
R11739 VDD.n2731 VDD.n1156 0.717237
R11740 VDD.n2713 VDD.n2712 0.717237
R11741 VDD.n2664 VDD.n2663 0.717237
R11742 VDD.n2637 VDD.n2636 0.717237
R11743 VDD.n2600 VDD.n2599 0.717237
R11744 VDD.n2573 VDD.n2572 0.717237
R11745 VDD.n2502 VDD.n2461 0.717237
R11746 VDD.n2520 VDD.n2519 0.717237
R11747 VDD.n1960 VDD.n1952 0.711611
R11748 VDD.n2336 VDD.n2328 0.711611
R11749 VDD.n2326 VDD.n2318 0.711611
R11750 VDD.n2316 VDD.n2308 0.711611
R11751 VDD.n2305 VDD.n2297 0.711611
R11752 VDD.n2295 VDD.n2287 0.711611
R11753 VDD.n2285 VDD.n2277 0.711611
R11754 VDD.n2275 VDD.n2267 0.711611
R11755 VDD.n1071 VDD.n1060 0.711611
R11756 VDD.n942 VDD.n931 0.711611
R11757 VDD.n813 VDD.n802 0.711611
R11758 VDD.n662 VDD.n651 0.711611
R11759 VDD.n533 VDD.n522 0.711611
R11760 VDD.n404 VDD.n393 0.711611
R11761 VDD.n275 VDD.n264 0.711611
R11762 VDD.n137 VDD.n126 0.711611
R11763 VDD.n2921 VDD.n2910 0.711611
R11764 VDD VDD.n2743 0.69574
R11765 VDD.n2232 VDD.n2231 0.690704
R11766 VDD.n1388 VDD.n1369 0.651821
R11767 VDD.n2905 VDD.n2904 0.629987
R11768 VDD.n2831 VDD.n2830 0.628071
R11769 VDD.n1675 VDD.n1674 0.627546
R11770 VDD.n1562 VDD.n1561 0.627546
R11771 VDD.n2754 VDD.n1155 0.612134
R11772 VDD.n2765 VDD.n1154 0.612134
R11773 VDD.n2776 VDD.n1153 0.612134
R11774 VDD.n2787 VDD.n1152 0.612134
R11775 VDD.n2798 VDD.n1151 0.612134
R11776 VDD.n2809 VDD.n1150 0.612134
R11777 VDD.n2820 VDD.n1149 0.612134
R11778 VDD.n2232 VDD.n2038 0.543454
R11779 VDD.n2905 VDD.n61 0.533877
R11780 VDD.n1951 VDD.n1950 0.530556
R11781 VDD.n2836 VDD.n2832 0.529912
R11782 VDD.n2845 VDD.n2841 0.529912
R11783 VDD.n2852 VDD.n2851 0.529912
R11784 VDD.n2752 VDD.n2751 0.529912
R11785 VDD.n2763 VDD.n2762 0.529912
R11786 VDD.n2774 VDD.n2773 0.529912
R11787 VDD.n2785 VDD.n2784 0.529912
R11788 VDD.n2796 VDD.n2795 0.529912
R11789 VDD.n2807 VDD.n2806 0.529912
R11790 VDD.n2818 VDD.n2817 0.529912
R11791 VDD.n2829 VDD.n2828 0.529912
R11792 VDD.n2742 VDD.n2741 0.529912
R11793 VDD.n2735 VDD.n2731 0.529912
R11794 VDD.n2726 VDD.n2725 0.529912
R11795 VDD.n2001 VDD.n2000 0.529912
R11796 VDD.n2010 VDD.n2009 0.529912
R11797 VDD.n2017 VDD.n2016 0.529912
R11798 VDD.n2021 VDD.n2020 0.529912
R11799 VDD.n2030 VDD.n2029 0.529912
R11800 VDD.n2037 VDD.n2036 0.529912
R11801 VDD.n1998 VDD.n1997 0.529912
R11802 VDD.n1972 VDD.n1961 0.529912
R11803 VDD.n2353 VDD.n2349 0.529912
R11804 VDD.n2362 VDD.n2358 0.529912
R11805 VDD.n2366 VDD.n2365 0.529912
R11806 VDD.n1804 VDD.n1803 0.529912
R11807 VDD.n1791 VDD.n1787 0.529912
R11808 VDD.n1386 VDD.n1385 0.529912
R11809 VDD.n1382 VDD.n1369 0.529912
R11810 VDD.n1800 VDD.n1799 0.529912
R11811 VDD.n1445 VDD.n1441 0.529912
R11812 VDD.n1449 VDD.n1448 0.529912
R11813 VDD.n1631 VDD.n1627 0.529912
R11814 VDD.n1640 VDD.n1636 0.529912
R11815 VDD.n1649 VDD.n1648 0.529912
R11816 VDD.n1658 VDD.n1654 0.529912
R11817 VDD.n1667 VDD.n1663 0.529912
R11818 VDD.n1674 VDD.n1673 0.529912
R11819 VDD.n1608 VDD.n1604 0.529912
R11820 VDD.n1617 VDD.n1613 0.529912
R11821 VDD.n1621 VDD.n1620 0.529912
R11822 VDD.n1599 VDD.n1595 0.529912
R11823 VDD.n1590 VDD.n1589 0.529912
R11824 VDD.n1581 VDD.n1577 0.529912
R11825 VDD.n1572 VDD.n1568 0.529912
R11826 VDD.n1563 VDD.n1562 0.529912
R11827 VDD.n2717 VDD.n2713 0.529912
R11828 VDD.n2659 VDD.n2658 0.529912
R11829 VDD.n2663 VDD.n2662 0.529912
R11830 VDD.n2650 VDD.n2649 0.529912
R11831 VDD.n2641 VDD.n2637 0.529912
R11832 VDD.n2595 VDD.n2594 0.529912
R11833 VDD.n2599 VDD.n2598 0.529912
R11834 VDD.n2586 VDD.n2585 0.529912
R11835 VDD.n2577 VDD.n2573 0.529912
R11836 VDD.n2506 VDD.n2502 0.529912
R11837 VDD.n2515 VDD.n2511 0.529912
R11838 VDD.n2519 VDD.n2518 0.529912
R11839 VDD.n2497 VDD.n2496 0.529912
R11840 VDD.n2341 VDD.n2340 0.5175
R11841 VDD.n278 VDD.n199 0.516382
R11842 VDD.n1206 VDD.n1182 0.50246
R11843 VDD.n686 VDD.n685 0.49871
R11844 VDD.n2853 VDD.n2852 0.487643
R11845 VDD.n2753 VDD.n2752 0.487643
R11846 VDD.n2764 VDD.n2763 0.487643
R11847 VDD.n2775 VDD.n2774 0.487643
R11848 VDD.n2786 VDD.n2785 0.487643
R11849 VDD.n2797 VDD.n2796 0.487643
R11850 VDD.n2808 VDD.n2807 0.487643
R11851 VDD.n2819 VDD.n2818 0.487643
R11852 VDD.n2830 VDD.n2829 0.487643
R11853 VDD.n2743 VDD.n2742 0.487643
R11854 VDD.n2725 VDD.n1155 0.487643
R11855 VDD.n2000 VDD.n1999 0.487643
R11856 VDD.n2009 VDD.n1980 0.487643
R11857 VDD.n2018 VDD.n2017 0.487643
R11858 VDD.n2020 VDD.n2019 0.487643
R11859 VDD.n2029 VDD.n1962 0.487643
R11860 VDD.n2038 VDD.n2037 0.487643
R11861 VDD.n1799 VDD.n1353 0.487643
R11862 VDD.n1648 VDD.n1345 0.487643
R11863 VDD.n1654 VDD.n1410 0.487643
R11864 VDD.n1663 VDD.n1411 0.487643
R11865 VDD.n1450 VDD.n1449 0.487643
R11866 VDD.n1441 VDD.n1302 0.487643
R11867 VDD.n1636 VDD.n1346 0.487643
R11868 VDD.n1627 VDD.n1626 0.487643
R11869 VDD.n1589 VDD.n1349 0.487643
R11870 VDD.n1577 VDD.n1405 0.487643
R11871 VDD.n1568 VDD.n1406 0.487643
R11872 VDD.n1613 VDD.n1453 0.487643
R11873 VDD.n1604 VDD.n1254 0.487643
R11874 VDD.n1595 VDD.n1350 0.487643
R11875 VDD.n1622 VDD.n1621 0.487643
R11876 VDD.n2367 VDD.n2366 0.487643
R11877 VDD.n1787 VDD.n1786 0.487643
R11878 VDD.n1805 VDD.n1804 0.487643
R11879 VDD.n1387 VDD.n1386 0.487643
R11880 VDD.n2358 VDD.n1171 0.487643
R11881 VDD.n2349 VDD.n2348 0.487643
R11882 VDD.n2658 VDD.n1154 0.487643
R11883 VDD.n2649 VDD.n1153 0.487643
R11884 VDD.n2594 VDD.n1152 0.487643
R11885 VDD.n2585 VDD.n1151 0.487643
R11886 VDD.n2496 VDD.n1150 0.487643
R11887 VDD.n2511 VDD.n1149 0.487643
R11888 VDD.n2841 VDD.n1125 0.487643
R11889 VDD.n2832 VDD.n2831 0.487643
R11890 VDD.n1019 VDD.n1018 0.471681
R11891 VDD.n1020 VDD.n1012 0.471681
R11892 VDD.n890 VDD.n889 0.471681
R11893 VDD.n891 VDD.n883 0.471681
R11894 VDD.n761 VDD.n760 0.471681
R11895 VDD.n762 VDD.n754 0.471681
R11896 VDD.n610 VDD.n609 0.471681
R11897 VDD.n611 VDD.n603 0.471681
R11898 VDD.n481 VDD.n480 0.471681
R11899 VDD.n482 VDD.n474 0.471681
R11900 VDD.n352 VDD.n351 0.471681
R11901 VDD.n353 VDD.n345 0.471681
R11902 VDD.n223 VDD.n222 0.471681
R11903 VDD.n224 VDD.n216 0.471681
R11904 VDD.n85 VDD.n84 0.471681
R11905 VDD.n86 VDD.n78 0.471681
R11906 VDD.n23 VDD.n22 0.471681
R11907 VDD.n24 VDD.n16 0.471681
R11908 VDD.n1074 VDD.n995 0.46479
R11909 VDD.n2677 VDD.n1156 0.461787
R11910 VDD.n2712 VDD.n2711 0.461787
R11911 VDD.n2665 VDD.n2664 0.461787
R11912 VDD.n2636 VDD.n2635 0.461787
R11913 VDD.n2601 VDD.n2600 0.461787
R11914 VDD.n2572 VDD.n2571 0.461787
R11915 VDD.n2537 VDD.n2461 0.461787
R11916 VDD.n2521 VDD.n2520 0.461787
R11917 VDD.n407 VDD.n328 0.461646
R11918 VDD.n665 VDD.n586 0.454935
R11919 VDD.n816 VDD.n737 0.448963
R11920 VDD.n1755 VDD.n1754 0.44832
R11921 VDD.n1785 VDD.n1784 0.44832
R11922 VDD.n1404 VDD.n1388 0.44832
R11923 VDD.n1728 VDD.n1727 0.44832
R11924 VDD.n945 VDD.n866 0.445564
R11925 VDD.n686 VDD.n667 0.438133
R11926 VDD.n2340 VDD.n2339 0.438122
R11927 VDD.n536 VDD.n457 0.437262
R11928 VDD.n1507 VDD.n1506 0.430365
R11929 VDD.n1531 VDD.n1530 0.430365
R11930 VDD.n1561 VDD.n1560 0.430365
R11931 VDD.n1483 VDD.n1482 0.430365
R11932 VDD.n1831 VDD.n1338 0.428253
R11933 VDD.n1409 VDD.n1344 0.428253
R11934 VDD.n1676 VDD.n1675 0.428253
R11935 VDD.n1431 VDD.n1326 0.428253
R11936 VDD.n1136 VDD.n1130 0.409094
R11937 VDD.n1206 VDD.n1205 0.396608
R11938 VDD.n2820 VDD.n2819 0.387346
R11939 VDD.n2809 VDD.n2808 0.387346
R11940 VDD.n2787 VDD.n2786 0.387346
R11941 VDD.n2765 VDD.n2764 0.387346
R11942 VDD.n2754 VDD.n2753 0.387346
R11943 VDD.n2798 VDD.n2797 0.387196
R11944 VDD.n1951 VDD.n1887 0.378552
R11945 VDD.n279 VDD.n151 0.368946
R11946 VDD.n817 VDD.n689 0.368387
R11947 VDD VDD.n2853 0.361938
R11948 VDD.n2854 VDD.n1124 0.355568
R11949 VDD.n408 VDD.n280 0.344607
R11950 VDD.n666 VDD.n538 0.343488
R11951 VDD.n2851 VDD.n1145 0.338713
R11952 VDD.n1075 VDD.n947 0.338173
R11953 VDD.n946 VDD.n818 0.337054
R11954 VDD.t1013 VDD.t2343 0.335952
R11955 VDD.t887 VDD.t2347 0.335952
R11956 VDD.t2339 VDD.t1011 0.335952
R11957 VDD.n2229 VDD.n2228 0.335952
R11958 VDD.t315 VDD.t2482 0.335952
R11959 VDD.t313 VDD.t2480 0.335952
R11960 VDD.t311 VDD.t2478 0.335952
R11961 VDD.n2263 VDD.n2244 0.335952
R11962 VDD.n2086 VDD.n2039 0.332336
R11963 VDD.n2091 VDD.n2086 0.332336
R11964 VDD.n2101 VDD.n2096 0.332336
R11965 VDD.n2106 VDD.n2101 0.332336
R11966 VDD.n2111 VDD.n2106 0.332336
R11967 VDD.n2196 VDD.n2119 0.332336
R11968 VDD.n2177 VDD.n2119 0.332336
R11969 VDD.n2177 VDD.n2176 0.332336
R11970 VDD.n2171 VDD.n2166 0.332336
R11971 VDD.n2166 VDD.n2161 0.332336
R11972 VDD.n199 VDD.n151 0.32198
R11973 VDD.n1140 VDD.n1139 0.317305
R11974 VDD.n1076 VDD.n141 0.316911
R11975 VDD.n537 VDD.n409 0.314393
R11976 VDD.n141 VDD.n140 0.305233
R11977 VDD.n2117 VDD.n2039 0.287639
R11978 VDD.n1755 VDD.n1753 0.278084
R11979 VDD.n1832 VDD.n1831 0.278084
R11980 VDD.n1676 VDD.n1412 0.278084
R11981 VDD.n1812 VDD.n1344 0.278084
R11982 VDD.n1853 VDD.n1326 0.278084
R11983 VDD.n1507 VDD.n1451 0.278084
R11984 VDD.n1560 VDD.n1407 0.278084
R11985 VDD.n1531 VDD.n1348 0.278084
R11986 VDD.n1483 VDD.n1278 0.278084
R11987 VDD.n1784 VDD.n1352 0.278084
R11988 VDD.n1708 VDD.n1404 0.278084
R11989 VDD.n1728 VDD.n1230 0.278084
R11990 VDD.n676 VDD.n675 0.276668
R11991 VDD.n737 VDD.n689 0.271625
R11992 VDD.n688 VDD.n687 0.263336
R11993 VDD.n2307 VDD.n2266 0.258832
R11994 VDD.n2853 VDD.n1125 0.257192
R11995 VDD.n2368 VDD.n1172 0.25526
R11996 VDD.n1707 VDD.n1363 0.25526
R11997 VDD.n2346 VDD.n2345 0.253566
R11998 VDD.n1624 VDD.n1623 0.248344
R11999 VDD.n1809 VDD.n1808 0.248344
R12000 VDD.n1706 VDD.n1705 0.248344
R12001 VDD.n2344 VDD.n2343 0.248344
R12002 VDD.n1625 VDD.n1331 0.247215
R12003 VDD.n1811 VDD.n1810 0.247215
R12004 VDD.n1704 VDD.n1703 0.247215
R12005 VDD.n2342 VDD.n2341 0.247215
R12006 VDD VDD.n2775 0.24258
R12007 VDD.n1807 VDD 0.242557
R12008 VDD.n2856 VDD.n2855 0.241224
R12009 VDD.n2743 VDD.n1156 0.240983
R12010 VDD.n2712 VDD.n1155 0.240983
R12011 VDD.n2664 VDD.n1154 0.240983
R12012 VDD.n2636 VDD.n1153 0.240983
R12013 VDD.n2600 VDD.n1152 0.240983
R12014 VDD.n2572 VDD.n1151 0.240983
R12015 VDD.n2461 VDD.n1150 0.240983
R12016 VDD.n2520 VDD.n1149 0.240983
R12017 VDD.n995 VDD.n947 0.240454
R12018 VDD.n1124 VDD.n1076 0.240164
R12019 VDD.n866 VDD.n818 0.239745
R12020 VDD.n328 VDD.n280 0.238136
R12021 VDD.n457 VDD.n409 0.237663
R12022 VDD.n2372 VDD.n2368 0.236898
R12023 VDD.n586 VDD.n538 0.236282
R12024 VDD.n1914 VDD.n1902 0.228189
R12025 VDD.n1830 VDD.n1339 0.226668
R12026 VDD.n1702 VDD.n1413 0.226668
R12027 VDD.n1842 VDD.n1841 0.226668
R12028 VDD.n1508 VDD.n1347 0.226668
R12029 VDD.n1532 VDD.n1408 0.226668
R12030 VDD.n1484 VDD.n1452 0.226668
R12031 VDD.n1756 VDD.n1351 0.226668
R12032 VDD.n1783 VDD.n1364 0.226668
R12033 VDD.n1744 VDD.n1743 0.226668
R12034 VDD.n141 VDD.n61 0.224589
R12035 VDD.n409 VDD.n408 0.217875
R12036 VDD.n1949 VDD.n1891 0.214959
R12037 VDD.n1625 VDD.n1624 0.214047
R12038 VDD.n1810 VDD.n1809 0.214047
R12039 VDD.n1705 VDD.n1704 0.214047
R12040 VDD.n2343 VDD.n2342 0.214047
R12041 VDD.n1623 VDD.n1172 0.213905
R12042 VDD.n1808 VDD.n1807 0.213905
R12043 VDD.n1707 VDD.n1706 0.213905
R12044 VDD.n2345 VDD.n2344 0.213905
R12045 VDD.n947 VDD.n946 0.210042
R12046 VDD.n2856 VDD.n61 0.208923
R12047 VDD.n1932 VDD.n1902 0.208693
R12048 VDD.n1933 VDD.n1932 0.208344
R12049 VDD.n818 VDD.n817 0.208083
R12050 VDD.n2832 VDD 0.204865
R12051 VDD.n2841 VDD 0.204865
R12052 VDD.n2852 VDD 0.204865
R12053 VDD.n2742 VDD 0.204865
R12054 VDD.n2731 VDD 0.204865
R12055 VDD.n2725 VDD 0.204865
R12056 VDD.n2000 VDD 0.204865
R12057 VDD.n2009 VDD 0.204865
R12058 VDD.n2017 VDD 0.204865
R12059 VDD.n2020 VDD 0.204865
R12060 VDD.n2029 VDD 0.204865
R12061 VDD.n2037 VDD 0.204865
R12062 VDD.n1998 VDD 0.204865
R12063 VDD.n1961 VDD 0.204865
R12064 VDD.n2349 VDD 0.204865
R12065 VDD.n2358 VDD 0.204865
R12066 VDD.n2366 VDD 0.204865
R12067 VDD.n1804 VDD 0.204865
R12068 VDD.n1787 VDD 0.204865
R12069 VDD.n1386 VDD 0.204865
R12070 VDD.n1369 VDD 0.204865
R12071 VDD.n1799 VDD 0.204865
R12072 VDD.n1441 VDD 0.204865
R12073 VDD.n1449 VDD 0.204865
R12074 VDD.n1627 VDD 0.204865
R12075 VDD.n1636 VDD 0.204865
R12076 VDD.n1648 VDD 0.204865
R12077 VDD.n1654 VDD 0.204865
R12078 VDD.n1663 VDD 0.204865
R12079 VDD.n1674 VDD 0.204865
R12080 VDD.n1604 VDD 0.204865
R12081 VDD.n1613 VDD 0.204865
R12082 VDD.n1621 VDD 0.204865
R12083 VDD.n1595 VDD 0.204865
R12084 VDD.n1589 VDD 0.204865
R12085 VDD.n1577 VDD 0.204865
R12086 VDD.n1568 VDD 0.204865
R12087 VDD.n1562 VDD 0.204865
R12088 VDD.n2713 VDD 0.204865
R12089 VDD.n2658 VDD 0.204865
R12090 VDD.n2663 VDD 0.204865
R12091 VDD.n2649 VDD 0.204865
R12092 VDD.n2637 VDD 0.204865
R12093 VDD.n2594 VDD 0.204865
R12094 VDD.n2599 VDD 0.204865
R12095 VDD.n2585 VDD 0.204865
R12096 VDD.n2573 VDD 0.204865
R12097 VDD.n2502 VDD 0.204865
R12098 VDD.n2511 VDD 0.204865
R12099 VDD.n2519 VDD 0.204865
R12100 VDD.n2496 VDD 0.204865
R12101 VDD.n408 VDD.n407 0.197247
R12102 VDD.n1075 VDD.n1074 0.196954
R12103 VDD.n280 VDD.n279 0.196613
R12104 VDD.n538 VDD.n537 0.196054
R12105 VDD.n946 VDD.n945 0.195517
R12106 VDD.n279 VDD.n278 0.194526
R12107 VDD.n537 VDD.n536 0.194526
R12108 VDD.n666 VDD.n665 0.194526
R12109 VDD.n817 VDD.n816 0.194526
R12110 VDD.n1933 VDD.n1891 0.194419
R12111 VDD.n149 VDD.n144 0.19425
R12112 VDD.n2195 VDD 0.193208
R12113 VDD.n2183 VDD 0.193208
R12114 VDD.n2178 VDD 0.193208
R12115 VDD.n2175 VDD 0.193208
R12116 VDD.n2170 VDD 0.193208
R12117 VDD.n2165 VDD 0.193208
R12118 VDD.n2160 VDD 0.193208
R12119 VDD.n2156 VDD 0.193208
R12120 VDD.n2116 VDD 0.193208
R12121 VDD VDD.n2050 0.193208
R12122 VDD.n2085 VDD 0.193208
R12123 VDD.n2090 VDD 0.193208
R12124 VDD.n2095 VDD 0.193208
R12125 VDD.n2100 VDD 0.193208
R12126 VDD.n2105 VDD 0.193208
R12127 VDD.n2110 VDD 0.193208
R12128 VDD.n1076 VDD.n1075 0.187381
R12129 VDD.n2345 VDD.n1229 0.184287
R12130 VDD.n2341 VDD.n1325 0.183322
R12131 VDD.n2343 VDD.n1277 0.182523
R12132 VDD.n2341 VDD.n1853 0.172413
R12133 VDD.n2343 VDD.n1278 0.172413
R12134 VDD.n2345 VDD.n1230 0.172413
R12135 VDD.n1182 VDD.n1164 0.171845
R12136 VDD.n2327 VDD.n2317 0.170814
R12137 VDD.n2368 VDD.n1171 0.170687
R12138 VDD.n2306 VDD.n2296 0.170572
R12139 VDD.n2296 VDD.n2286 0.17033
R12140 VDD.n1786 VDD.n1363 0.16897
R12141 VDD.n2337 VDD.n2327 0.168392
R12142 VDD.n2176 VDD 0.167836
R12143 VDD.n2286 VDD.n2276 0.167665
R12144 VDD VDD.n2091 0.166621
R12145 VDD.n2096 VDD 0.166216
R12146 VDD.n1806 VDD.n1353 0.165966
R12147 VDD VDD.n2171 0.165
R12148 VDD.n1841 VDD.n1331 0.164842
R12149 VDD.n1624 VDD.n1452 0.164842
R12150 VDD.n1744 VDD.n1172 0.164842
R12151 VDD.n1786 VDD.n1785 0.164678
R12152 VDD.n1727 VDD.n1171 0.164678
R12153 VDD.n1703 VDD.n1702 0.162319
R12154 VDD.n1705 VDD.n1408 0.162319
R12155 VDD.n1707 VDD.n1364 0.162319
R12156 VDD.n2404 VDD.n2385 0.161112
R12157 VDD.n2197 VDD.n2118 0.160543
R12158 VDD.n1811 VDD.n1339 0.157903
R12159 VDD.n1809 VDD.n1347 0.157903
R12160 VDD.n1807 VDD.n1351 0.157903
R12161 VDD.n2348 VDD.n2347 0.155021
R12162 VDD.n1625 VDD.n1450 0.145523
R12163 VDD.n1623 VDD.n1453 0.145523
R12164 VDD.n2776 VDD 0.145266
R12165 VDD.n1704 VDD.n1410 0.14406
R12166 VDD.n1706 VDD.n1405 0.14406
R12167 VDD VDD.n1125 0.143458
R12168 VDD.n1812 VDD.n1811 0.143393
R12169 VDD.n1809 VDD.n1348 0.143393
R12170 VDD.n1807 VDD.n1352 0.143393
R12171 VDD.n1810 VDD.n1346 0.1415
R12172 VDD.n1808 VDD.n1350 0.1415
R12173 VDD.n1410 VDD.n1409 0.140403
R12174 VDD.n1450 VDD.n1431 0.140403
R12175 VDD.n1530 VDD.n1405 0.140403
R12176 VDD.n1482 VDD.n1453 0.140403
R12177 VDD.n2257 VDD.n2256 0.13977
R12178 VDD.n1703 VDD.n1412 0.138977
R12179 VDD.n1705 VDD.n1407 0.138977
R12180 VDD.n1708 VDD.n1707 0.138977
R12181 VDD.n2367 VDD 0.138281
R12182 VDD.n1805 VDD 0.138281
R12183 VDD VDD.n1387 0.138281
R12184 VDD.n2348 VDD 0.138281
R12185 VDD.n1218 VDD.n1217 0.137041
R12186 VDD.n1753 VDD.n1172 0.136453
R12187 VDD.n1832 VDD.n1331 0.136453
R12188 VDD.n1624 VDD.n1451 0.136453
R12189 VDD.n1314 VDD.n1313 0.136451
R12190 VDD.n1266 VDD.n1265 0.135985
R12191 VDD.n149 VDD.n148 0.135917
R12192 VDD.n2223 VDD.n2222 0.135733
R12193 VDD.n2258 VDD.n2233 0.135733
R12194 VDD.n1806 VDD.n1805 0.135276
R12195 VDD.n2221 VDD.n2220 0.13458
R12196 VDD.n2265 VDD.n2234 0.13458
R12197 VDD.n2222 VDD.n2221 0.132273
R12198 VDD.n1387 VDD.n1363 0.132272
R12199 VDD.n2342 VDD.n1302 0.132173
R12200 VDD.n2344 VDD.n1254 0.132173
R12201 VDD.n688 VDD.n666 0.131988
R12202 VDD.n2373 VDD.n1163 0.130567
R12203 VDD.n2368 VDD.n2367 0.130555
R12204 VDD.n1754 VDD 0.122829
R12205 VDD.n2692 VDD.n2677 0.121133
R12206 VDD.n2711 VDD.n2710 0.121133
R12207 VDD.n2665 VDD.n2421 0.121133
R12208 VDD.n2635 VDD.n2634 0.121133
R12209 VDD.n2601 VDD.n2441 0.121133
R12210 VDD.n2571 VDD.n2570 0.121133
R12211 VDD.n2537 VDD.n2536 0.121133
R12212 VDD.n2521 VDD.n2483 0.121133
R12213 VDD.n2231 VDD.n2198 0.118721
R12214 VDD VDD.n1345 0.117909
R12215 VDD VDD.n1411 0.117909
R12216 VDD VDD.n1302 0.117909
R12217 VDD.n1626 VDD 0.117909
R12218 VDD VDD.n1349 0.117909
R12219 VDD VDD.n1406 0.117909
R12220 VDD VDD.n1254 0.117909
R12221 VDD.n1622 VDD 0.117909
R12222 VDD.n2340 VDD.n1951 0.115563
R12223 VDD.n1810 VDD.n1345 0.115348
R12224 VDD.n1808 VDD.n1349 0.115348
R12225 VDD.n1704 VDD.n1411 0.112788
R12226 VDD.n1706 VDD.n1406 0.112788
R12227 VDD VDD.n2199 0.112666
R12228 VDD VDD.n2257 0.112666
R12229 VDD.n2752 VDD 0.111611
R12230 VDD.n2763 VDD 0.111611
R12231 VDD.n2774 VDD 0.111611
R12232 VDD.n2785 VDD 0.111611
R12233 VDD.n2796 VDD 0.111611
R12234 VDD.n2807 VDD 0.111611
R12235 VDD.n2818 VDD 0.111611
R12236 VDD.n2829 VDD 0.111611
R12237 VDD.n1626 VDD.n1625 0.111325
R12238 VDD.n1623 VDD.n1622 0.111325
R12239 VDD.n678 VDD.n676 0.109591
R12240 VDD.n2344 VDD.n1253 0.107732
R12241 VDD.n2342 VDD.n1301 0.107427
R12242 VDD.n2711 VDD.n2413 0.106511
R12243 VDD VDD.n1056 0.106084
R12244 VDD VDD.n927 0.106084
R12245 VDD VDD.n798 0.106084
R12246 VDD VDD.n647 0.106084
R12247 VDD VDD.n518 0.106084
R12248 VDD VDD.n389 0.106084
R12249 VDD VDD.n260 0.106084
R12250 VDD VDD.n122 0.106084
R12251 VDD VDD.n60 0.106084
R12252 VDD VDD.n1338 0.104741
R12253 VDD.n1506 VDD 0.104741
R12254 VDD.n1138 VDD.n1137 0.100535
R12255 VDD.n1082 VDD.n1080 0.0996736
R12256 VDD.n1114 VDD.n1112 0.0996736
R12257 VDD.n1123 VDD.n1122 0.0996736
R12258 VDD.n1122 VDD.n1120 0.0996736
R12259 VDD.n1001 VDD.n999 0.0996736
R12260 VDD.n1047 VDD.n1045 0.0996736
R12261 VDD.n1044 VDD.n1043 0.0996736
R12262 VDD.n1043 VDD.n1041 0.0996736
R12263 VDD.n1004 VDD.n1003 0.0996736
R12264 VDD.n1007 VDD.n1005 0.0996736
R12265 VDD.n1009 VDD.n1007 0.0996736
R12266 VDD.n1035 VDD.n1033 0.0996736
R12267 VDD.n1032 VDD.n1031 0.0996736
R12268 VDD.n1031 VDD.n1029 0.0996736
R12269 VDD.n1056 VDD.n1055 0.0996736
R12270 VDD.n1055 VDD.n1053 0.0996736
R12271 VDD.n953 VDD.n951 0.0996736
R12272 VDD.n985 VDD.n983 0.0996736
R12273 VDD.n994 VDD.n993 0.0996736
R12274 VDD.n993 VDD.n991 0.0996736
R12275 VDD.n872 VDD.n870 0.0996736
R12276 VDD.n918 VDD.n916 0.0996736
R12277 VDD.n915 VDD.n914 0.0996736
R12278 VDD.n914 VDD.n912 0.0996736
R12279 VDD.n875 VDD.n874 0.0996736
R12280 VDD.n878 VDD.n876 0.0996736
R12281 VDD.n880 VDD.n878 0.0996736
R12282 VDD.n906 VDD.n904 0.0996736
R12283 VDD.n903 VDD.n902 0.0996736
R12284 VDD.n902 VDD.n900 0.0996736
R12285 VDD.n927 VDD.n926 0.0996736
R12286 VDD.n926 VDD.n924 0.0996736
R12287 VDD.n824 VDD.n822 0.0996736
R12288 VDD.n856 VDD.n854 0.0996736
R12289 VDD.n865 VDD.n864 0.0996736
R12290 VDD.n864 VDD.n862 0.0996736
R12291 VDD.n743 VDD.n741 0.0996736
R12292 VDD.n789 VDD.n787 0.0996736
R12293 VDD.n786 VDD.n785 0.0996736
R12294 VDD.n785 VDD.n783 0.0996736
R12295 VDD.n746 VDD.n745 0.0996736
R12296 VDD.n749 VDD.n747 0.0996736
R12297 VDD.n751 VDD.n749 0.0996736
R12298 VDD.n777 VDD.n775 0.0996736
R12299 VDD.n774 VDD.n773 0.0996736
R12300 VDD.n773 VDD.n771 0.0996736
R12301 VDD.n798 VDD.n797 0.0996736
R12302 VDD.n797 VDD.n795 0.0996736
R12303 VDD.n695 VDD.n693 0.0996736
R12304 VDD.n727 VDD.n725 0.0996736
R12305 VDD.n736 VDD.n735 0.0996736
R12306 VDD.n735 VDD.n733 0.0996736
R12307 VDD.n623 VDD.n622 0.0996736
R12308 VDD.n622 VDD.n620 0.0996736
R12309 VDD.n598 VDD.n596 0.0996736
R12310 VDD.n600 VDD.n598 0.0996736
R12311 VDD.n626 VDD.n624 0.0996736
R12312 VDD.n635 VDD.n634 0.0996736
R12313 VDD.n634 VDD.n632 0.0996736
R12314 VDD.n595 VDD.n594 0.0996736
R12315 VDD.n592 VDD.n590 0.0996736
R12316 VDD.n638 VDD.n636 0.0996736
R12317 VDD.n647 VDD.n646 0.0996736
R12318 VDD.n646 VDD.n644 0.0996736
R12319 VDD.n544 VDD.n542 0.0996736
R12320 VDD.n576 VDD.n574 0.0996736
R12321 VDD.n585 VDD.n584 0.0996736
R12322 VDD.n584 VDD.n582 0.0996736
R12323 VDD.n463 VDD.n461 0.0996736
R12324 VDD.n509 VDD.n507 0.0996736
R12325 VDD.n506 VDD.n505 0.0996736
R12326 VDD.n505 VDD.n503 0.0996736
R12327 VDD.n466 VDD.n465 0.0996736
R12328 VDD.n469 VDD.n467 0.0996736
R12329 VDD.n471 VDD.n469 0.0996736
R12330 VDD.n497 VDD.n495 0.0996736
R12331 VDD.n494 VDD.n493 0.0996736
R12332 VDD.n493 VDD.n491 0.0996736
R12333 VDD.n518 VDD.n517 0.0996736
R12334 VDD.n517 VDD.n515 0.0996736
R12335 VDD.n415 VDD.n413 0.0996736
R12336 VDD.n447 VDD.n445 0.0996736
R12337 VDD.n456 VDD.n455 0.0996736
R12338 VDD.n455 VDD.n453 0.0996736
R12339 VDD.n334 VDD.n332 0.0996736
R12340 VDD.n380 VDD.n378 0.0996736
R12341 VDD.n377 VDD.n376 0.0996736
R12342 VDD.n376 VDD.n374 0.0996736
R12343 VDD.n337 VDD.n336 0.0996736
R12344 VDD.n340 VDD.n338 0.0996736
R12345 VDD.n342 VDD.n340 0.0996736
R12346 VDD.n368 VDD.n366 0.0996736
R12347 VDD.n365 VDD.n364 0.0996736
R12348 VDD.n364 VDD.n362 0.0996736
R12349 VDD.n389 VDD.n388 0.0996736
R12350 VDD.n388 VDD.n386 0.0996736
R12351 VDD.n286 VDD.n284 0.0996736
R12352 VDD.n318 VDD.n316 0.0996736
R12353 VDD.n327 VDD.n326 0.0996736
R12354 VDD.n326 VDD.n324 0.0996736
R12355 VDD.n157 VDD.n155 0.0996736
R12356 VDD.n189 VDD.n187 0.0996736
R12357 VDD.n198 VDD.n197 0.0996736
R12358 VDD.n197 VDD.n195 0.0996736
R12359 VDD.n205 VDD.n203 0.0996736
R12360 VDD.n251 VDD.n249 0.0996736
R12361 VDD.n248 VDD.n247 0.0996736
R12362 VDD.n247 VDD.n245 0.0996736
R12363 VDD.n208 VDD.n207 0.0996736
R12364 VDD.n211 VDD.n209 0.0996736
R12365 VDD.n213 VDD.n211 0.0996736
R12366 VDD.n239 VDD.n237 0.0996736
R12367 VDD.n236 VDD.n235 0.0996736
R12368 VDD.n235 VDD.n233 0.0996736
R12369 VDD.n260 VDD.n259 0.0996736
R12370 VDD.n259 VDD.n257 0.0996736
R12371 VDD.n67 VDD.n65 0.0996736
R12372 VDD.n113 VDD.n111 0.0996736
R12373 VDD.n110 VDD.n109 0.0996736
R12374 VDD.n109 VDD.n107 0.0996736
R12375 VDD.n70 VDD.n69 0.0996736
R12376 VDD.n73 VDD.n71 0.0996736
R12377 VDD.n75 VDD.n73 0.0996736
R12378 VDD.n101 VDD.n99 0.0996736
R12379 VDD.n98 VDD.n97 0.0996736
R12380 VDD.n97 VDD.n95 0.0996736
R12381 VDD.n122 VDD.n121 0.0996736
R12382 VDD.n121 VDD.n119 0.0996736
R12383 VDD.n2862 VDD.n2860 0.0996736
R12384 VDD.n2894 VDD.n2892 0.0996736
R12385 VDD.n2903 VDD.n2902 0.0996736
R12386 VDD.n2902 VDD.n2900 0.0996736
R12387 VDD.n5 VDD.n3 0.0996736
R12388 VDD.n51 VDD.n49 0.0996736
R12389 VDD.n48 VDD.n47 0.0996736
R12390 VDD.n47 VDD.n45 0.0996736
R12391 VDD.n8 VDD.n7 0.0996736
R12392 VDD.n11 VDD.n9 0.0996736
R12393 VDD.n13 VDD.n11 0.0996736
R12394 VDD.n39 VDD.n37 0.0996736
R12395 VDD.n36 VDD.n35 0.0996736
R12396 VDD.n35 VDD.n33 0.0996736
R12397 VDD.n60 VDD.n59 0.0996736
R12398 VDD.n59 VDD.n57 0.0996736
R12399 VDD.n2831 VDD 0.0994712
R12400 VDD.n1099 VDD.n1098 0.0992654
R12401 VDD.n1098 VDD.n1096 0.0992654
R12402 VDD.n1088 VDD.n1086 0.0992654
R12403 VDD.n1090 VDD.n1088 0.0992654
R12404 VDD.n1102 VDD.n1100 0.0992654
R12405 VDD.n1111 VDD.n1110 0.0992654
R12406 VDD.n1110 VDD.n1108 0.0992654
R12407 VDD.n1085 VDD.n1084 0.0992654
R12408 VDD.n970 VDD.n969 0.0992654
R12409 VDD.n969 VDD.n967 0.0992654
R12410 VDD.n959 VDD.n957 0.0992654
R12411 VDD.n961 VDD.n959 0.0992654
R12412 VDD.n973 VDD.n971 0.0992654
R12413 VDD.n982 VDD.n981 0.0992654
R12414 VDD.n981 VDD.n979 0.0992654
R12415 VDD.n956 VDD.n955 0.0992654
R12416 VDD.n841 VDD.n840 0.0992654
R12417 VDD.n840 VDD.n838 0.0992654
R12418 VDD.n830 VDD.n828 0.0992654
R12419 VDD.n832 VDD.n830 0.0992654
R12420 VDD.n844 VDD.n842 0.0992654
R12421 VDD.n853 VDD.n852 0.0992654
R12422 VDD.n852 VDD.n850 0.0992654
R12423 VDD.n827 VDD.n826 0.0992654
R12424 VDD.n712 VDD.n711 0.0992654
R12425 VDD.n711 VDD.n709 0.0992654
R12426 VDD.n701 VDD.n699 0.0992654
R12427 VDD.n703 VDD.n701 0.0992654
R12428 VDD.n715 VDD.n713 0.0992654
R12429 VDD.n724 VDD.n723 0.0992654
R12430 VDD.n723 VDD.n721 0.0992654
R12431 VDD.n698 VDD.n697 0.0992654
R12432 VDD.n561 VDD.n560 0.0992654
R12433 VDD.n560 VDD.n558 0.0992654
R12434 VDD.n550 VDD.n548 0.0992654
R12435 VDD.n552 VDD.n550 0.0992654
R12436 VDD.n564 VDD.n562 0.0992654
R12437 VDD.n573 VDD.n572 0.0992654
R12438 VDD.n572 VDD.n570 0.0992654
R12439 VDD.n547 VDD.n546 0.0992654
R12440 VDD.n432 VDD.n431 0.0992654
R12441 VDD.n431 VDD.n429 0.0992654
R12442 VDD.n421 VDD.n419 0.0992654
R12443 VDD.n423 VDD.n421 0.0992654
R12444 VDD.n435 VDD.n433 0.0992654
R12445 VDD.n444 VDD.n443 0.0992654
R12446 VDD.n443 VDD.n441 0.0992654
R12447 VDD.n418 VDD.n417 0.0992654
R12448 VDD.n303 VDD.n302 0.0992654
R12449 VDD.n302 VDD.n300 0.0992654
R12450 VDD.n292 VDD.n290 0.0992654
R12451 VDD.n294 VDD.n292 0.0992654
R12452 VDD.n306 VDD.n304 0.0992654
R12453 VDD.n315 VDD.n314 0.0992654
R12454 VDD.n314 VDD.n312 0.0992654
R12455 VDD.n289 VDD.n288 0.0992654
R12456 VDD.n174 VDD.n173 0.0992654
R12457 VDD.n173 VDD.n171 0.0992654
R12458 VDD.n163 VDD.n161 0.0992654
R12459 VDD.n165 VDD.n163 0.0992654
R12460 VDD.n177 VDD.n175 0.0992654
R12461 VDD.n186 VDD.n185 0.0992654
R12462 VDD.n185 VDD.n183 0.0992654
R12463 VDD.n160 VDD.n159 0.0992654
R12464 VDD.n2879 VDD.n2878 0.0992654
R12465 VDD.n2878 VDD.n2876 0.0992654
R12466 VDD.n2868 VDD.n2866 0.0992654
R12467 VDD.n2870 VDD.n2868 0.0992654
R12468 VDD.n2882 VDD.n2880 0.0992654
R12469 VDD.n2891 VDD.n2890 0.0992654
R12470 VDD.n2890 VDD.n2888 0.0992654
R12471 VDD.n2865 VDD.n2864 0.0992654
R12472 VDD.n2317 VDD.n2307 0.0953479
R12473 VDD.n624 VDD.n623 0.0937345
R12474 VDD.n1033 VDD.n1032 0.0937345
R12475 VDD.n904 VDD.n903 0.0937345
R12476 VDD.n775 VDD.n774 0.0937345
R12477 VDD.n495 VDD.n494 0.0937345
R12478 VDD.n366 VDD.n365 0.0937345
R12479 VDD.n237 VDD.n236 0.0937345
R12480 VDD.n99 VDD.n98 0.0937345
R12481 VDD.n37 VDD.n36 0.0937345
R12482 VDD.n1100 VDD.n1099 0.0936091
R12483 VDD.n971 VDD.n970 0.0936091
R12484 VDD.n842 VDD.n841 0.0936091
R12485 VDD.n713 VDD.n712 0.0936091
R12486 VDD.n562 VDD.n561 0.0936091
R12487 VDD.n433 VDD.n432 0.0936091
R12488 VDD.n304 VDD.n303 0.0936091
R12489 VDD.n175 VDD.n174 0.0936091
R12490 VDD.n2880 VDD.n2879 0.0936091
R12491 VDD.n1242 VDD.n1241 0.0926298
R12492 VDD.n1290 VDD.n1289 0.0924671
R12493 VDD.n2231 VDD.n2199 0.0904632
R12494 VDD.n1115 VDD.n1114 0.090376
R12495 VDD.n1118 VDD.n1078 0.090376
R12496 VDD.n1048 VDD.n1047 0.090376
R12497 VDD.n1039 VDD.n1003 0.090376
R12498 VDD.n1036 VDD.n1035 0.090376
R12499 VDD.n1027 VDD.n1025 0.090376
R12500 VDD.n1051 VDD.n997 0.090376
R12501 VDD.n986 VDD.n985 0.090376
R12502 VDD.n989 VDD.n949 0.090376
R12503 VDD.n919 VDD.n918 0.090376
R12504 VDD.n910 VDD.n874 0.090376
R12505 VDD.n907 VDD.n906 0.090376
R12506 VDD.n898 VDD.n896 0.090376
R12507 VDD.n922 VDD.n868 0.090376
R12508 VDD.n857 VDD.n856 0.090376
R12509 VDD.n860 VDD.n820 0.090376
R12510 VDD.n790 VDD.n789 0.090376
R12511 VDD.n781 VDD.n745 0.090376
R12512 VDD.n778 VDD.n777 0.090376
R12513 VDD.n769 VDD.n767 0.090376
R12514 VDD.n793 VDD.n739 0.090376
R12515 VDD.n728 VDD.n727 0.090376
R12516 VDD.n731 VDD.n691 0.090376
R12517 VDD.n618 VDD.n616 0.090376
R12518 VDD.n627 VDD.n626 0.090376
R12519 VDD.n630 VDD.n594 0.090376
R12520 VDD.n639 VDD.n638 0.090376
R12521 VDD.n642 VDD.n588 0.090376
R12522 VDD.n577 VDD.n576 0.090376
R12523 VDD.n580 VDD.n540 0.090376
R12524 VDD.n510 VDD.n509 0.090376
R12525 VDD.n501 VDD.n465 0.090376
R12526 VDD.n498 VDD.n497 0.090376
R12527 VDD.n489 VDD.n487 0.090376
R12528 VDD.n513 VDD.n459 0.090376
R12529 VDD.n448 VDD.n447 0.090376
R12530 VDD.n451 VDD.n411 0.090376
R12531 VDD.n381 VDD.n380 0.090376
R12532 VDD.n372 VDD.n336 0.090376
R12533 VDD.n369 VDD.n368 0.090376
R12534 VDD.n360 VDD.n358 0.090376
R12535 VDD.n384 VDD.n330 0.090376
R12536 VDD.n319 VDD.n318 0.090376
R12537 VDD.n322 VDD.n282 0.090376
R12538 VDD.n190 VDD.n189 0.090376
R12539 VDD.n193 VDD.n153 0.090376
R12540 VDD.n252 VDD.n251 0.090376
R12541 VDD.n243 VDD.n207 0.090376
R12542 VDD.n240 VDD.n239 0.090376
R12543 VDD.n231 VDD.n229 0.090376
R12544 VDD.n255 VDD.n201 0.090376
R12545 VDD.n114 VDD.n113 0.090376
R12546 VDD.n105 VDD.n69 0.090376
R12547 VDD.n102 VDD.n101 0.090376
R12548 VDD.n93 VDD.n91 0.090376
R12549 VDD.n117 VDD.n63 0.090376
R12550 VDD.n2895 VDD.n2894 0.090376
R12551 VDD.n2898 VDD.n2858 0.090376
R12552 VDD.n52 VDD.n51 0.090376
R12553 VDD.n43 VDD.n7 0.090376
R12554 VDD.n40 VDD.n39 0.090376
R12555 VDD.n31 VDD.n29 0.090376
R12556 VDD.n55 VDD.n1 0.090376
R12557 VDD.n1094 VDD.n1092 0.0900062
R12558 VDD.n1103 VDD.n1102 0.0900062
R12559 VDD.n1106 VDD.n1084 0.0900062
R12560 VDD.n965 VDD.n963 0.0900062
R12561 VDD.n974 VDD.n973 0.0900062
R12562 VDD.n977 VDD.n955 0.0900062
R12563 VDD.n836 VDD.n834 0.0900062
R12564 VDD.n845 VDD.n844 0.0900062
R12565 VDD.n848 VDD.n826 0.0900062
R12566 VDD.n707 VDD.n705 0.0900062
R12567 VDD.n716 VDD.n715 0.0900062
R12568 VDD.n719 VDD.n697 0.0900062
R12569 VDD.n556 VDD.n554 0.0900062
R12570 VDD.n565 VDD.n564 0.0900062
R12571 VDD.n568 VDD.n546 0.0900062
R12572 VDD.n427 VDD.n425 0.0900062
R12573 VDD.n436 VDD.n435 0.0900062
R12574 VDD.n439 VDD.n417 0.0900062
R12575 VDD.n298 VDD.n296 0.0900062
R12576 VDD.n307 VDD.n306 0.0900062
R12577 VDD.n310 VDD.n288 0.0900062
R12578 VDD.n169 VDD.n167 0.0900062
R12579 VDD.n178 VDD.n177 0.0900062
R12580 VDD.n181 VDD.n159 0.0900062
R12581 VDD.n2874 VDD.n2872 0.0900062
R12582 VDD.n2883 VDD.n2882 0.0900062
R12583 VDD.n2886 VDD.n2864 0.0900062
R12584 VDD.n1072 VDD.n1059 0.0880141
R12585 VDD.n943 VDD.n930 0.0880141
R12586 VDD.n814 VDD.n801 0.0880141
R12587 VDD.n663 VDD.n650 0.0880141
R12588 VDD.n534 VDD.n521 0.0880141
R12589 VDD.n405 VDD.n392 0.0880141
R12590 VDD.n276 VDD.n263 0.0880141
R12591 VDD.n138 VDD.n125 0.0880141
R12592 VDD.n2922 VDD.n2909 0.0880141
R12593 VDD.n2338 VDD.n2337 0.0877165
R12594 VDD.n1005 VDD.n1004 0.0875105
R12595 VDD.n876 VDD.n875 0.0875105
R12596 VDD.n747 VDD.n746 0.0875105
R12597 VDD.n596 VDD.n595 0.0875105
R12598 VDD.n467 VDD.n466 0.0875105
R12599 VDD.n338 VDD.n337 0.0875105
R12600 VDD.n209 VDD.n208 0.0875105
R12601 VDD.n71 VDD.n70 0.0875105
R12602 VDD.n9 VDD.n8 0.0875105
R12603 VDD.n1086 VDD.n1085 0.0873851
R12604 VDD.n957 VDD.n956 0.0873851
R12605 VDD.n828 VDD.n827 0.0873851
R12606 VDD.n699 VDD.n698 0.0873851
R12607 VDD.n548 VDD.n547 0.0873851
R12608 VDD.n419 VDD.n418 0.0873851
R12609 VDD.n290 VDD.n289 0.0873851
R12610 VDD.n161 VDD.n160 0.0873851
R12611 VDD.n2866 VDD.n2865 0.0873851
R12612 VDD.n1045 VDD.n1044 0.0849171
R12613 VDD.n916 VDD.n915 0.0849171
R12614 VDD.n787 VDD.n786 0.0849171
R12615 VDD.n636 VDD.n635 0.0849171
R12616 VDD.n507 VDD.n506 0.0849171
R12617 VDD.n378 VDD.n377 0.0849171
R12618 VDD.n249 VDD.n248 0.0849171
R12619 VDD.n111 VDD.n110 0.0849171
R12620 VDD.n49 VDD.n48 0.0849171
R12621 VDD.n1112 VDD.n1111 0.0848555
R12622 VDD.n983 VDD.n982 0.0848555
R12623 VDD.n854 VDD.n853 0.0848555
R12624 VDD.n725 VDD.n724 0.0848555
R12625 VDD.n574 VDD.n573 0.0848555
R12626 VDD.n445 VDD.n444 0.0848555
R12627 VDD.n316 VDD.n315 0.0848555
R12628 VDD.n187 VDD.n186 0.0848555
R12629 VDD.n2892 VDD.n2891 0.0848555
R12630 VDD VDD.n2820 0.0841058
R12631 VDD VDD.n2809 0.0841058
R12632 VDD VDD.n2798 0.0841058
R12633 VDD VDD.n2787 0.0841058
R12634 VDD VDD.n2776 0.0841058
R12635 VDD VDD.n2765 0.0841058
R12636 VDD VDD.n2754 0.0841058
R12637 VDD.n2124 VDD.n2123 0.0839821
R12638 VDD.n2127 VDD.n2126 0.0839821
R12639 VDD.n2130 VDD.n2129 0.0839821
R12640 VDD.n2133 VDD.n2132 0.0839821
R12641 VDD.n2136 VDD.n2135 0.0839821
R12642 VDD.n2139 VDD.n2138 0.0839821
R12643 VDD.n2142 VDD.n2141 0.0839821
R12644 VDD.n2145 VDD.n2144 0.0839821
R12645 VDD.n2115 VDD.n2041 0.0839821
R12646 VDD.n2053 VDD.n2052 0.0839821
R12647 VDD.n2057 VDD.n2056 0.0839821
R12648 VDD.n2061 VDD.n2060 0.0839821
R12649 VDD.n2065 VDD.n2064 0.0839821
R12650 VDD.n2069 VDD.n2068 0.0839821
R12651 VDD.n2073 VDD.n2072 0.0839821
R12652 VDD.n2077 VDD.n2076 0.0839821
R12653 VDD.n1018 VDD.n1016 0.0839821
R12654 VDD.n889 VDD.n887 0.0839821
R12655 VDD.n760 VDD.n758 0.0839821
R12656 VDD.n609 VDD.n607 0.0839821
R12657 VDD.n480 VDD.n478 0.0839821
R12658 VDD.n351 VDD.n349 0.0839821
R12659 VDD.n222 VDD.n220 0.0839821
R12660 VDD.n144 VDD.n143 0.0839821
R12661 VDD.n84 VDD.n82 0.0839821
R12662 VDD.n22 VDD.n20 0.0839821
R12663 VDD.n2399 VDD.n2398 0.0829405
R12664 VDD.n2406 VDD.n2384 0.0829405
R12665 VDD.n2381 VDD.n2380 0.0829405
R12666 VDD.n2371 VDD.n2370 0.0829405
R12667 VDD.n1312 VDD.n1311 0.0829405
R12668 VDD.n1324 VDD.n1323 0.0829405
R12669 VDD.n1288 VDD.n1287 0.0829405
R12670 VDD.n1300 VDD.n1299 0.0829405
R12671 VDD.n1264 VDD.n1263 0.0829405
R12672 VDD.n1276 VDD.n1275 0.0829405
R12673 VDD.n1252 VDD.n1251 0.0829405
R12674 VDD.n1216 VDD.n1215 0.0829405
R12675 VDD.n1228 VDD.n1227 0.0829405
R12676 VDD.n1203 VDD.n1202 0.0829405
R12677 VDD.n1185 VDD.n1184 0.0829405
R12678 VDD.n1139 VDD.n1126 0.0822901
R12679 VDD.n1240 VDD.n1239 0.0818988
R12680 VDD.n1950 VDD.n1949 0.0817926
R12681 VDD.n1205 VDD.n1193 0.078355
R12682 VDD VDD.n2194 0.0775833
R12683 VDD.n2184 VDD 0.0775833
R12684 VDD.n2179 VDD 0.0775833
R12685 VDD VDD.n2174 0.0775833
R12686 VDD VDD.n2169 0.0775833
R12687 VDD VDD.n2164 0.0775833
R12688 VDD VDD.n2159 0.0775833
R12689 VDD VDD.n2155 0.0775833
R12690 VDD.n2044 VDD 0.0765417
R12691 VDD VDD.n2049 0.0765417
R12692 VDD VDD.n2084 0.0765417
R12693 VDD VDD.n2089 0.0765417
R12694 VDD VDD.n2094 0.0765417
R12695 VDD VDD.n2099 0.0765417
R12696 VDD VDD.n2104 0.0765417
R12697 VDD VDD.n2109 0.0765417
R12698 VDD.n2307 VDD.n2306 0.0745129
R12699 VDD.n1145 VDD.n1140 0.0741196
R12700 VDD.n1831 VDD.n1830 0.0733658
R12701 VDD.n1413 VDD.n1344 0.0733658
R12702 VDD.n1677 VDD.n1676 0.0733658
R12703 VDD.n1842 VDD.n1326 0.0733658
R12704 VDD.n1508 VDD.n1507 0.0733658
R12705 VDD.n1532 VDD.n1531 0.0733658
R12706 VDD.n1560 VDD.n1559 0.0733658
R12707 VDD.n1484 VDD.n1483 0.0733658
R12708 VDD.n1756 VDD.n1755 0.0733658
R12709 VDD.n1784 VDD.n1783 0.0733658
R12710 VDD.n1404 VDD.n1403 0.0733658
R12711 VDD.n1743 VDD.n1728 0.0733658
R12712 VDD.n1277 VDD.n1266 0.0732781
R12713 VDD.n1229 VDD.n1218 0.0729282
R12714 VDD.n1325 VDD.n1314 0.0723824
R12715 VDD.n2373 VDD.n2372 0.0709436
R12716 VDD.n2405 VDD.n2404 0.0675623
R12717 VDD.n2194 VDD.n2193 0.066125
R12718 VDD.n2185 VDD.n2184 0.066125
R12719 VDD.n2180 VDD.n2179 0.066125
R12720 VDD.n2174 VDD.n2150 0.066125
R12721 VDD.n2169 VDD.n2149 0.066125
R12722 VDD.n2164 VDD.n2148 0.066125
R12723 VDD.n2159 VDD.n2147 0.066125
R12724 VDD.n2155 VDD.n2146 0.066125
R12725 VDD.n2045 VDD.n2044 0.066125
R12726 VDD.n2049 VDD.n2046 0.066125
R12727 VDD.n2084 VDD.n2054 0.066125
R12728 VDD.n2089 VDD.n2058 0.066125
R12729 VDD.n2094 VDD.n2062 0.066125
R12730 VDD.n2099 VDD.n2066 0.066125
R12731 VDD.n2104 VDD.n2070 0.066125
R12732 VDD.n2109 VDD.n2074 0.066125
R12733 VDD.n1020 VDD.n1019 0.066125
R12734 VDD.n1022 VDD.n1012 0.066125
R12735 VDD.n891 VDD.n890 0.066125
R12736 VDD.n893 VDD.n883 0.066125
R12737 VDD.n762 VDD.n761 0.066125
R12738 VDD.n764 VDD.n754 0.066125
R12739 VDD.n611 VDD.n610 0.066125
R12740 VDD.n613 VDD.n603 0.066125
R12741 VDD.n482 VDD.n481 0.066125
R12742 VDD.n484 VDD.n474 0.066125
R12743 VDD.n353 VDD.n352 0.066125
R12744 VDD.n355 VDD.n345 0.066125
R12745 VDD.n224 VDD.n223 0.066125
R12746 VDD.n226 VDD.n216 0.066125
R12747 VDD.n86 VDD.n85 0.066125
R12748 VDD.n88 VDD.n78 0.066125
R12749 VDD.n24 VDD.n23 0.066125
R12750 VDD.n26 VDD.n16 0.066125
R12751 VDD.n2346 VDD.n1206 0.0651856
R12752 VDD.n2405 VDD.n1164 0.06497
R12753 VDD.n1887 VDD.n1854 0.0648091
R12754 VDD.n2411 VDD.n1164 0.0639556
R12755 VDD.n2412 VDD.n1163 0.0631667
R12756 VDD.n1874 VDD.n1854 0.0615242
R12757 VDD.n1059 VDD.n1058 0.0614987
R12758 VDD.n930 VDD.n929 0.0614987
R12759 VDD.n801 VDD.n800 0.0614987
R12760 VDD.n650 VDD.n649 0.0614987
R12761 VDD.n521 VDD.n520 0.0614987
R12762 VDD.n392 VDD.n391 0.0614987
R12763 VDD.n263 VDD.n262 0.0614987
R12764 VDD.n125 VDD.n124 0.0614987
R12765 VDD.n2909 VDD.n2908 0.0614987
R12766 VDD.n1073 VDD 0.0612752
R12767 VDD.n944 VDD 0.0612752
R12768 VDD.n815 VDD 0.0612752
R12769 VDD.n664 VDD 0.0612752
R12770 VDD.n535 VDD 0.0612752
R12771 VDD.n406 VDD 0.0612752
R12772 VDD.n277 VDD 0.0612752
R12773 VDD.n139 VDD 0.0612752
R12774 VDD VDD.n2906 0.0612752
R12775 VDD.n150 VDD 0.0597672
R12776 VDD.n1873 VDD.n1862 0.0597554
R12777 VDD.n1882 VDD.n1878 0.05925
R12778 VDD.n2195 VDD 0.0588333
R12779 VDD VDD.n2183 0.0588333
R12780 VDD VDD.n2178 0.0588333
R12781 VDD.n2175 VDD 0.0588333
R12782 VDD.n2170 VDD 0.0588333
R12783 VDD.n2165 VDD 0.0588333
R12784 VDD.n2160 VDD 0.0588333
R12785 VDD.n2156 VDD 0.0588333
R12786 VDD.n2116 VDD 0.0588333
R12787 VDD.n2050 VDD 0.0588333
R12788 VDD.n2085 VDD 0.0588333
R12789 VDD.n2090 VDD 0.0588333
R12790 VDD.n2095 VDD 0.0588333
R12791 VDD.n2100 VDD 0.0588333
R12792 VDD.n2105 VDD 0.0588333
R12793 VDD.n2110 VDD 0.0588333
R12794 VDD.n1133 VDD.n1132 0.0585357
R12795 VDD.n1878 VDD.n1862 0.0582392
R12796 VDD.n1205 VDD.n1204 0.0579046
R12797 VDD VDD.n2391 0.056838
R12798 VDD VDD.n2387 0.056838
R12799 VDD VDD.n1166 0.056838
R12800 VDD VDD.n1170 0.056838
R12801 VDD VDD.n1940 0.056838
R12802 VDD VDD.n1901 0.056838
R12803 VDD VDD.n1904 0.056838
R12804 VDD VDD.n1921 0.056838
R12805 VDD VDD.n1906 0.056838
R12806 VDD VDD.n1908 0.056838
R12807 VDD VDD.n1897 0.056838
R12808 VDD VDD.n1304 0.056838
R12809 VDD VDD.n1316 0.056838
R12810 VDD VDD.n1280 0.056838
R12811 VDD VDD.n1292 0.056838
R12812 VDD VDD.n1256 0.056838
R12813 VDD VDD.n1268 0.056838
R12814 VDD VDD.n1232 0.056838
R12815 VDD VDD.n1244 0.056838
R12816 VDD VDD.n1208 0.056838
R12817 VDD VDD.n1220 0.056838
R12818 VDD VDD.n1195 0.056838
R12819 VDD VDD.n1187 0.056838
R12820 VDD.n1948 VDD.n1893 0.0556643
R12821 VDD VDD.n678 0.0550455
R12822 VDD.n2534 VDD 0.0546373
R12823 VDD.n2690 VDD 0.0546373
R12824 VDD.n2708 VDD 0.0546373
R12825 VDD.n1741 VDD 0.0546373
R12826 VDD.n1401 VDD 0.0546373
R12827 VDD.n1781 VDD 0.0546373
R12828 VDD VDD.n1759 0.0546373
R12829 VDD VDD.n1845 0.0546373
R12830 VDD.n1828 VDD 0.0546373
R12831 VDD VDD.n1680 0.0546373
R12832 VDD VDD.n1694 0.0546373
R12833 VDD VDD.n1487 0.0546373
R12834 VDD VDD.n1511 0.0546373
R12835 VDD.n1557 VDD 0.0546373
R12836 VDD VDD.n1535 0.0546373
R12837 VDD VDD.n2613 0.0546373
R12838 VDD.n2632 VDD 0.0546373
R12839 VDD VDD.n2549 0.0546373
R12840 VDD.n2568 VDD 0.0546373
R12841 VDD.n2481 VDD 0.0546373
R12842 VDD.n2532 VDD.n2466 0.0539038
R12843 VDD.n2688 VDD.n2679 0.0539038
R12844 VDD.n2706 VDD.n2418 0.0539038
R12845 VDD.n2395 VDD.n2394 0.0539038
R12846 VDD.n2402 VDD.n2389 0.0539038
R12847 VDD.n2409 VDD.n1168 0.0539038
R12848 VDD.n2377 VDD.n2376 0.0539038
R12849 VDD.n1947 VDD.n1895 0.0539038
R12850 VDD.n1308 VDD.n1307 0.0539038
R12851 VDD.n1320 VDD.n1319 0.0539038
R12852 VDD.n1284 VDD.n1283 0.0539038
R12853 VDD.n1296 VDD.n1295 0.0539038
R12854 VDD.n1260 VDD.n1259 0.0539038
R12855 VDD.n1272 VDD.n1271 0.0539038
R12856 VDD.n1236 VDD.n1235 0.0539038
R12857 VDD.n1248 VDD.n1247 0.0539038
R12858 VDD.n1212 VDD.n1211 0.0539038
R12859 VDD.n1224 VDD.n1223 0.0539038
R12860 VDD.n1199 VDD.n1198 0.0539038
R12861 VDD.n1191 VDD.n1189 0.0539038
R12862 VDD.n1739 VDD.n1730 0.0539038
R12863 VDD.n1399 VDD.n1393 0.0539038
R12864 VDD.n1779 VDD.n1366 0.0539038
R12865 VDD.n1762 VDD.n1761 0.0539038
R12866 VDD.n1848 VDD.n1847 0.0539038
R12867 VDD.n1826 VDD.n1341 0.0539038
R12868 VDD.n1683 VDD.n1682 0.0539038
R12869 VDD.n1697 VDD.n1696 0.0539038
R12870 VDD.n1490 VDD.n1489 0.0539038
R12871 VDD.n1514 VDD.n1513 0.0539038
R12872 VDD.n1555 VDD.n1470 0.0539038
R12873 VDD.n1538 VDD.n1537 0.0539038
R12874 VDD.n2616 VDD.n2615 0.0539038
R12875 VDD.n2630 VDD.n2438 0.0539038
R12876 VDD.n2552 VDD.n2551 0.0539038
R12877 VDD.n2566 VDD.n2458 0.0539038
R12878 VDD.n2479 VDD.n2473 0.0539038
R12879 VDD VDD.n2460 0.0531316
R12880 VDD VDD.n2681 0.0531316
R12881 VDD VDD.n2699 0.0531316
R12882 VDD VDD.n1368 0.0531316
R12883 VDD VDD.n1772 0.0531316
R12884 VDD VDD.n1722 0.0531316
R12885 VDD VDD.n1337 0.0531316
R12886 VDD VDD.n1686 0.0531316
R12887 VDD VDD.n1343 0.0531316
R12888 VDD VDD.n1328 0.0531316
R12889 VDD VDD.n1500 0.0531316
R12890 VDD VDD.n1548 0.0531316
R12891 VDD VDD.n1524 0.0531316
R12892 VDD VDD.n1476 0.0531316
R12893 VDD VDD.n1732 0.0531316
R12894 VDD VDD.n2420 0.0531316
R12895 VDD VDD.n2432 0.0531316
R12896 VDD VDD.n2440 0.0531316
R12897 VDD VDD.n2452 0.0531316
R12898 VDD VDD.n2468 0.0531316
R12899 VDD.n2855 VDD.n2854 0.0531298
R12900 VDD.n2230 VDD.n2201 0.0528198
R12901 VDD.n2204 VDD.n2203 0.0528198
R12902 VDD.n2224 VDD.n2212 0.0528198
R12903 VDD.n2207 VDD.n2206 0.0528198
R12904 VDD.n2210 VDD.n2209 0.0528198
R12905 VDD.n2217 VDD.n2216 0.0528198
R12906 VDD.n2219 VDD.n2214 0.0528198
R12907 VDD.n2227 VDD.n2226 0.0528198
R12908 VDD.n2191 VDD.n2187 0.0528198
R12909 VDD.n2113 VDD.n2079 0.0528198
R12910 VDD.n2247 VDD.n2246 0.0528198
R12911 VDD.n2255 VDD.n2254 0.0528198
R12912 VDD.n2250 VDD.n2249 0.0528198
R12913 VDD.n2259 VDD.n2252 0.0528198
R12914 VDD.n2264 VDD.n2236 0.0528198
R12915 VDD.n2239 VDD.n2238 0.0528198
R12916 VDD.n2242 VDD.n2241 0.0528198
R12917 VDD.n2262 VDD.n2261 0.0528198
R12918 VDD.n1875 VDD.n1872 0.0528198
R12919 VDD.n1867 VDD.n1866 0.0528198
R12920 VDD.n1870 VDD.n1869 0.0528198
R12921 VDD.n1877 VDD.n1864 0.0528198
R12922 VDD.n1886 VDD.n1856 0.0528198
R12923 VDD.n1859 VDD.n1858 0.0528198
R12924 VDD.n1881 VDD.n1880 0.0528198
R12925 VDD.n1883 VDD.n1861 0.0528198
R12926 VDD.n1924 VDD.n1923 0.0521432
R12927 VDD.n1890 VDD.n1889 0.0515563
R12928 VDD.n1138 VDD 0.0515204
R12929 VDD.n1913 VDD.n1912 0.0509695
R12930 VDD.n2541 VDD.n2540 0.0503904
R12931 VDD.n2696 VDD.n2695 0.0503904
R12932 VDD.n2685 VDD.n2684 0.0503904
R12933 VDD.n2673 VDD.n2672 0.0503904
R12934 VDD.n2703 VDD.n2702 0.0503904
R12935 VDD.n1748 VDD.n1747 0.0503904
R12936 VDD.n1712 VDD.n1711 0.0503904
R12937 VDD.n1719 VDD.n1718 0.0503904
R12938 VDD.n1776 VDD.n1775 0.0503904
R12939 VDD.n1769 VDD.n1768 0.0503904
R12940 VDD.n1751 VDD.n1724 0.0503904
R12941 VDD.n1839 VDD.n1335 0.0503904
R12942 VDD.n1836 VDD.n1835 0.0503904
R12943 VDD.n1823 VDD.n1822 0.0503904
R12944 VDD.n1690 VDD.n1689 0.0503904
R12945 VDD.n1700 VDD.n1417 0.0503904
R12946 VDD.n1816 VDD.n1815 0.0503904
R12947 VDD.n1423 VDD.n1421 0.0503904
R12948 VDD.n1851 VDD.n1330 0.0503904
R12949 VDD.n1497 VDD.n1496 0.0503904
R12950 VDD.n1504 VDD.n1503 0.0503904
R12951 VDD.n1521 VDD.n1520 0.0503904
R12952 VDD.n1552 VDD.n1551 0.0503904
R12953 VDD.n1545 VDD.n1544 0.0503904
R12954 VDD.n1528 VDD.n1527 0.0503904
R12955 VDD.n1473 VDD.n1472 0.0503904
R12956 VDD.n1480 VDD.n1479 0.0503904
R12957 VDD.n1396 VDD.n1395 0.0503904
R12958 VDD.n1736 VDD.n1735 0.0503904
R12959 VDD.n2623 VDD.n2622 0.0503904
R12960 VDD.n2669 VDD.n2668 0.0503904
R12961 VDD.n2609 VDD.n2608 0.0503904
R12962 VDD.n2627 VDD.n2626 0.0503904
R12963 VDD.n2559 VDD.n2558 0.0503904
R12964 VDD.n2605 VDD.n2604 0.0503904
R12965 VDD.n2545 VDD.n2544 0.0503904
R12966 VDD.n2563 VDD.n2562 0.0503904
R12967 VDD.n2529 VDD.n2528 0.0503904
R12968 VDD.n2476 VDD.n2475 0.0503904
R12969 VDD.n2525 VDD.n2524 0.0503904
R12970 VDD.n1936 VDD.n1935 0.0497958
R12971 VDD.n1931 VDD.n1930 0.0497958
R12972 VDD.n1874 VDD 0.0496479
R12973 VDD.n1301 VDD.n1290 0.0494516
R12974 VDD.n1253 VDD.n1242 0.0494516
R12975 VDD.n1917 VDD.n1916 0.0486221
R12976 VDD.n2693 VDD.n2676 0.0471009
R12977 VDD.n2416 VDD.n2415 0.0471009
R12978 VDD.n1745 VDD.n1726 0.0471009
R12979 VDD.n1716 VDD.n1715 0.0471009
R12980 VDD.n1766 VDD.n1765 0.0471009
R12981 VDD.n1840 VDD.n1333 0.0471009
R12982 VDD.n1820 VDD.n1819 0.0471009
R12983 VDD.n1701 VDD.n1415 0.0471009
R12984 VDD.n1424 VDD.n1419 0.0471009
R12985 VDD.n1494 VDD.n1493 0.0471009
R12986 VDD.n1518 VDD.n1517 0.0471009
R12987 VDD.n1542 VDD.n1541 0.0471009
R12988 VDD.n1468 VDD.n1467 0.0471009
R12989 VDD.n1391 VDD.n1390 0.0471009
R12990 VDD.n2620 VDD.n2619 0.0471009
R12991 VDD.n2436 VDD.n2435 0.0471009
R12992 VDD.n2556 VDD.n2555 0.0471009
R12993 VDD.n2456 VDD.n2455 0.0471009
R12994 VDD.n2464 VDD.n2463 0.0471009
R12995 VDD.n2471 VDD.n2470 0.0471009
R12996 VDD.n1943 VDD.n1942 0.0468615
R12997 VDD.n2266 VDD.n2233 0.0460583
R12998 VDD.n681 VDD.n680 0.0448182
R12999 VDD.n2535 VDD.n2534 0.0443596
R13000 VDD.n2691 VDD.n2690 0.0443596
R13001 VDD.n2709 VDD.n2708 0.0443596
R13002 VDD.n1742 VDD.n1741 0.0443596
R13003 VDD.n1402 VDD.n1401 0.0443596
R13004 VDD.n1782 VDD.n1781 0.0443596
R13005 VDD.n1759 VDD.n1757 0.0443596
R13006 VDD.n1845 VDD.n1843 0.0443596
R13007 VDD.n1829 VDD.n1828 0.0443596
R13008 VDD.n1680 VDD.n1678 0.0443596
R13009 VDD.n1694 VDD.n1692 0.0443596
R13010 VDD.n1487 VDD.n1485 0.0443596
R13011 VDD.n1511 VDD.n1509 0.0443596
R13012 VDD.n1558 VDD.n1557 0.0443596
R13013 VDD.n1535 VDD.n1533 0.0443596
R13014 VDD.n2613 VDD.n2611 0.0443596
R13015 VDD.n2633 VDD.n2632 0.0443596
R13016 VDD.n2549 VDD.n2547 0.0443596
R13017 VDD.n2569 VDD.n2568 0.0443596
R13018 VDD.n2482 VDD.n2481 0.0443596
R13019 VDD VDD.n1353 0.0423493
R13020 VDD.n1139 VDD.n1138 0.0414154
R13021 VDD.n2223 VDD 0.0388497
R13022 VDD.n2258 VDD 0.0388497
R13023 VDD.n1132 VDD.n1126 0.0387653
R13024 VDD.n1346 VDD 0.0361615
R13025 VDD VDD.n1350 0.0361615
R13026 VDD VDD.n2230 0.0361308
R13027 VDD.n2204 VDD 0.0361308
R13028 VDD.n2224 VDD 0.0361308
R13029 VDD VDD.n2207 0.0361308
R13030 VDD VDD.n2210 0.0361308
R13031 VDD.n2217 VDD 0.0361308
R13032 VDD VDD.n2219 0.0361308
R13033 VDD.n2227 VDD 0.0361308
R13034 VDD VDD.n2247 0.0361308
R13035 VDD VDD.n2255 0.0361308
R13036 VDD VDD.n2250 0.0361308
R13037 VDD.n2259 VDD 0.0361308
R13038 VDD VDD.n2264 0.0361308
R13039 VDD.n2239 VDD 0.0361308
R13040 VDD.n2242 VDD 0.0361308
R13041 VDD.n2262 VDD 0.0361308
R13042 VDD.n1875 VDD 0.0361308
R13043 VDD VDD.n1867 0.0361308
R13044 VDD.n1870 VDD 0.0361308
R13045 VDD VDD.n1877 0.0361308
R13046 VDD VDD.n1886 0.0361308
R13047 VDD.n1859 VDD 0.0361308
R13048 VDD VDD.n1881 0.0361308
R13049 VDD.n1883 VDD 0.0361308
R13050 VDD.n1073 VDD 0.0347938
R13051 VDD.n944 VDD 0.0347938
R13052 VDD.n815 VDD 0.0347938
R13053 VDD.n664 VDD 0.0347938
R13054 VDD.n535 VDD 0.0347938
R13055 VDD.n406 VDD 0.0347938
R13056 VDD.n277 VDD 0.0347938
R13057 VDD.n139 VDD 0.0347938
R13058 VDD.n2906 VDD 0.0347938
R13059 VDD.n2904 VDD.n2856 0.0339315
R13060 VDD.n1754 VDD 0.033121
R13061 VDD.n1785 VDD 0.033121
R13062 VDD.n1388 VDD 0.033121
R13063 VDD.n1727 VDD 0.033121
R13064 VDD.n2197 VDD.n2196 0.0284569
R13065 VDD.n1025 VDD.n1023 0.0283926
R13066 VDD.n896 VDD.n894 0.0283926
R13067 VDD.n767 VDD.n765 0.0283926
R13068 VDD.n616 VDD.n614 0.0283926
R13069 VDD.n487 VDD.n485 0.0283926
R13070 VDD.n358 VDD.n356 0.0283926
R13071 VDD.n229 VDD.n227 0.0283926
R13072 VDD.n91 VDD.n89 0.0283926
R13073 VDD.n29 VDD.n27 0.0283926
R13074 VDD.n1409 VDD 0.0282977
R13075 VDD.n1675 VDD 0.0282977
R13076 VDD.n1431 VDD 0.0282977
R13077 VDD VDD.n1338 0.0282977
R13078 VDD.n1530 VDD 0.0282977
R13079 VDD.n1561 VDD 0.0282977
R13080 VDD.n1482 VDD 0.0282977
R13081 VDD.n1506 VDD 0.0282977
R13082 VDD.n2830 VDD 0.0258077
R13083 VDD.n2819 VDD 0.0258077
R13084 VDD.n2808 VDD 0.0258077
R13085 VDD.n2797 VDD 0.0258077
R13086 VDD.n2786 VDD 0.0258077
R13087 VDD.n2775 VDD 0.0258077
R13088 VDD.n2764 VDD 0.0258077
R13089 VDD.n2753 VDD 0.0258077
R13090 VDD.n671 VDD.n670 0.0243095
R13091 VDD.n2339 VDD.n2338 0.0230309
R13092 VDD.n1061 VDD 0.0206477
R13093 VDD.n932 VDD 0.0206477
R13094 VDD.n803 VDD 0.0206477
R13095 VDD.n652 VDD 0.0206477
R13096 VDD.n523 VDD 0.0206477
R13097 VDD.n394 VDD 0.0206477
R13098 VDD.n265 VDD 0.0206477
R13099 VDD.n127 VDD 0.0206477
R13100 VDD.n2911 VDD 0.0206477
R13101 VDD.n2190 VDD 0.0186075
R13102 VDD.n2112 VDD 0.0186075
R13103 VDD.n2194 VDD.n2121 0.0183571
R13104 VDD.n2184 VDD.n2182 0.0183571
R13105 VDD.n2179 VDD.n2152 0.0183571
R13106 VDD.n2174 VDD.n2173 0.0183571
R13107 VDD.n2169 VDD.n2168 0.0183571
R13108 VDD.n2164 VDD.n2163 0.0183571
R13109 VDD.n2159 VDD.n2158 0.0183571
R13110 VDD.n2155 VDD.n2154 0.0183571
R13111 VDD.n2044 VDD.n2043 0.0183571
R13112 VDD.n2049 VDD.n2048 0.0183571
R13113 VDD.n2084 VDD.n2083 0.0183571
R13114 VDD.n2089 VDD.n2088 0.0183571
R13115 VDD.n2094 VDD.n2093 0.0183571
R13116 VDD.n2099 VDD.n2098 0.0183571
R13117 VDD.n2104 VDD.n2103 0.0183571
R13118 VDD.n2109 VDD.n2108 0.0183571
R13119 VDD.n1019 VDD.n1014 0.0183571
R13120 VDD.n1012 VDD.n1011 0.0183571
R13121 VDD.n890 VDD.n885 0.0183571
R13122 VDD.n883 VDD.n882 0.0183571
R13123 VDD.n761 VDD.n756 0.0183571
R13124 VDD.n754 VDD.n753 0.0183571
R13125 VDD.n610 VDD.n605 0.0183571
R13126 VDD.n603 VDD.n602 0.0183571
R13127 VDD.n481 VDD.n476 0.0183571
R13128 VDD.n474 VDD.n473 0.0183571
R13129 VDD.n352 VDD.n347 0.0183571
R13130 VDD.n345 VDD.n344 0.0183571
R13131 VDD.n223 VDD.n218 0.0183571
R13132 VDD.n216 VDD.n215 0.0183571
R13133 VDD.n148 VDD.n146 0.0183571
R13134 VDD.n675 VDD.n673 0.0183571
R13135 VDD.n85 VDD.n80 0.0183571
R13136 VDD.n78 VDD.n77 0.0183571
R13137 VDD.n23 VDD.n18 0.0183571
R13138 VDD.n16 VDD.n15 0.0183571
R13139 VDD.n2191 VDD.n2190 0.0180234
R13140 VDD.n2113 VDD.n2112 0.0180234
R13141 VDD.n1137 VDD.n1136 0.0176233
R13142 VDD VDD.n1873 0.0173038
R13143 VDD.n2347 VDD.n1182 0.0141907
R13144 VDD VDD.n1806 0.0132027
R13145 VDD.n1138 VDD.n1128 0.0107041
R13146 VDD.n671 VDD.n667 0.0104206
R13147 VDD.n1115 VDD.n1082 0.00979752
R13148 VDD.n1120 VDD.n1118 0.00979752
R13149 VDD.n1048 VDD.n1001 0.00979752
R13150 VDD.n1041 VDD.n1039 0.00979752
R13151 VDD.n1036 VDD.n1009 0.00979752
R13152 VDD.n1029 VDD.n1027 0.00979752
R13153 VDD.n1053 VDD.n1051 0.00979752
R13154 VDD.n986 VDD.n953 0.00979752
R13155 VDD.n991 VDD.n989 0.00979752
R13156 VDD.n919 VDD.n872 0.00979752
R13157 VDD.n912 VDD.n910 0.00979752
R13158 VDD.n907 VDD.n880 0.00979752
R13159 VDD.n900 VDD.n898 0.00979752
R13160 VDD.n924 VDD.n922 0.00979752
R13161 VDD.n857 VDD.n824 0.00979752
R13162 VDD.n862 VDD.n860 0.00979752
R13163 VDD.n790 VDD.n743 0.00979752
R13164 VDD.n783 VDD.n781 0.00979752
R13165 VDD.n778 VDD.n751 0.00979752
R13166 VDD.n771 VDD.n769 0.00979752
R13167 VDD.n795 VDD.n793 0.00979752
R13168 VDD.n728 VDD.n695 0.00979752
R13169 VDD.n733 VDD.n731 0.00979752
R13170 VDD.n620 VDD.n618 0.00979752
R13171 VDD.n627 VDD.n600 0.00979752
R13172 VDD.n632 VDD.n630 0.00979752
R13173 VDD.n639 VDD.n592 0.00979752
R13174 VDD.n644 VDD.n642 0.00979752
R13175 VDD.n577 VDD.n544 0.00979752
R13176 VDD.n582 VDD.n580 0.00979752
R13177 VDD.n510 VDD.n463 0.00979752
R13178 VDD.n503 VDD.n501 0.00979752
R13179 VDD.n498 VDD.n471 0.00979752
R13180 VDD.n491 VDD.n489 0.00979752
R13181 VDD.n515 VDD.n513 0.00979752
R13182 VDD.n448 VDD.n415 0.00979752
R13183 VDD.n453 VDD.n451 0.00979752
R13184 VDD.n381 VDD.n334 0.00979752
R13185 VDD.n374 VDD.n372 0.00979752
R13186 VDD.n369 VDD.n342 0.00979752
R13187 VDD.n362 VDD.n360 0.00979752
R13188 VDD.n386 VDD.n384 0.00979752
R13189 VDD.n319 VDD.n286 0.00979752
R13190 VDD.n324 VDD.n322 0.00979752
R13191 VDD.n190 VDD.n157 0.00979752
R13192 VDD.n195 VDD.n193 0.00979752
R13193 VDD.n252 VDD.n205 0.00979752
R13194 VDD.n245 VDD.n243 0.00979752
R13195 VDD.n240 VDD.n213 0.00979752
R13196 VDD.n233 VDD.n231 0.00979752
R13197 VDD.n257 VDD.n255 0.00979752
R13198 VDD.n114 VDD.n67 0.00979752
R13199 VDD.n107 VDD.n105 0.00979752
R13200 VDD.n102 VDD.n75 0.00979752
R13201 VDD.n95 VDD.n93 0.00979752
R13202 VDD.n119 VDD.n117 0.00979752
R13203 VDD.n2895 VDD.n2862 0.00979752
R13204 VDD.n2900 VDD.n2898 0.00979752
R13205 VDD.n52 VDD.n5 0.00979752
R13206 VDD.n45 VDD.n43 0.00979752
R13207 VDD.n40 VDD.n13 0.00979752
R13208 VDD.n33 VDD.n31 0.00979752
R13209 VDD.n57 VDD.n55 0.00979752
R13210 VDD.n1096 VDD.n1094 0.00975926
R13211 VDD.n1103 VDD.n1090 0.00975926
R13212 VDD.n1108 VDD.n1106 0.00975926
R13213 VDD.n967 VDD.n965 0.00975926
R13214 VDD.n974 VDD.n961 0.00975926
R13215 VDD.n979 VDD.n977 0.00975926
R13216 VDD.n838 VDD.n836 0.00975926
R13217 VDD.n845 VDD.n832 0.00975926
R13218 VDD.n850 VDD.n848 0.00975926
R13219 VDD.n709 VDD.n707 0.00975926
R13220 VDD.n716 VDD.n703 0.00975926
R13221 VDD.n721 VDD.n719 0.00975926
R13222 VDD.n558 VDD.n556 0.00975926
R13223 VDD.n565 VDD.n552 0.00975926
R13224 VDD.n570 VDD.n568 0.00975926
R13225 VDD.n429 VDD.n427 0.00975926
R13226 VDD.n436 VDD.n423 0.00975926
R13227 VDD.n441 VDD.n439 0.00975926
R13228 VDD.n300 VDD.n298 0.00975926
R13229 VDD.n307 VDD.n294 0.00975926
R13230 VDD.n312 VDD.n310 0.00975926
R13231 VDD.n171 VDD.n169 0.00975926
R13232 VDD.n178 VDD.n165 0.00975926
R13233 VDD.n183 VDD.n181 0.00975926
R13234 VDD.n2876 VDD.n2874 0.00975926
R13235 VDD.n2883 VDD.n2870 0.00975926
R13236 VDD.n2888 VDD.n2886 0.00975926
R13237 VDD.n682 VDD.n681 0.00788636
R13238 VDD.n1944 VDD.n1943 0.00754225
R13239 VDD VDD.n2693 0.0065307
R13240 VDD VDD.n2416 0.0065307
R13241 VDD VDD.n1745 0.0065307
R13242 VDD VDD.n1716 0.0065307
R13243 VDD VDD.n1766 0.0065307
R13244 VDD.n1840 VDD 0.0065307
R13245 VDD VDD.n1820 0.0065307
R13246 VDD.n1701 VDD 0.0065307
R13247 VDD.n1424 VDD 0.0065307
R13248 VDD VDD.n1494 0.0065307
R13249 VDD VDD.n1518 0.0065307
R13250 VDD VDD.n1542 0.0065307
R13251 VDD VDD.n1468 0.0065307
R13252 VDD VDD.n1391 0.0065307
R13253 VDD VDD.n2620 0.0065307
R13254 VDD VDD.n2436 0.0065307
R13255 VDD VDD.n2556 0.0065307
R13256 VDD VDD.n2456 0.0065307
R13257 VDD VDD.n2464 0.0065307
R13258 VDD VDD.n2471 0.0065307
R13259 VDD.n2855 VDD.n140 0.00639406
R13260 VDD.n2412 VDD.n2411 0.00613549
R13261 VDD.n2266 VDD.n2265 0.00597853
R13262 VDD.n1918 VDD.n1917 0.00578169
R13263 VDD.n2276 VDD 0.00570876
R13264 VDD.n689 VDD.n688 0.00497619
R13265 VDD.n1937 VDD.n1936 0.00460798
R13266 VDD.n1931 VDD.n1928 0.00460798
R13267 VDD.n1133 VDD 0.00368878
R13268 VDD VDD.n2532 0.00343427
R13269 VDD VDD.n2688 0.00343427
R13270 VDD VDD.n2706 0.00343427
R13271 VDD VDD.n1947 0.00343427
R13272 VDD.n1944 VDD 0.00343427
R13273 VDD.n1937 VDD 0.00343427
R13274 VDD.n1928 VDD 0.00343427
R13275 VDD.n1925 VDD 0.00343427
R13276 VDD.n1918 VDD 0.00343427
R13277 VDD.n1910 VDD 0.00343427
R13278 VDD.n1913 VDD.n1910 0.00343427
R13279 VDD.n1898 VDD 0.00343427
R13280 VDD VDD.n1739 0.00343427
R13281 VDD VDD.n1399 0.00343427
R13282 VDD VDD.n1779 0.00343427
R13283 VDD.n1762 VDD 0.00343427
R13284 VDD.n1848 VDD 0.00343427
R13285 VDD VDD.n1826 0.00343427
R13286 VDD.n1683 VDD 0.00343427
R13287 VDD.n1697 VDD 0.00343427
R13288 VDD.n1490 VDD 0.00343427
R13289 VDD.n1514 VDD 0.00343427
R13290 VDD VDD.n1555 0.00343427
R13291 VDD.n1538 VDD 0.00343427
R13292 VDD.n2616 VDD 0.00343427
R13293 VDD VDD.n2630 0.00343427
R13294 VDD.n2552 VDD 0.00343427
R13295 VDD VDD.n2566 0.00343427
R13296 VDD VDD.n2479 0.00343427
R13297 VDD.n682 VDD 0.00334091
R13298 VDD.n2696 VDD 0.00324123
R13299 VDD.n2673 VDD 0.00324123
R13300 VDD.n1748 VDD 0.00324123
R13301 VDD.n1719 VDD 0.00324123
R13302 VDD.n1769 VDD 0.00324123
R13303 VDD VDD.n1839 0.00324123
R13304 VDD.n1823 VDD 0.00324123
R13305 VDD VDD.n1700 0.00324123
R13306 VDD VDD.n1423 0.00324123
R13307 VDD.n1497 VDD 0.00324123
R13308 VDD.n1521 VDD 0.00324123
R13309 VDD.n1545 VDD 0.00324123
R13310 VDD.n1473 VDD 0.00324123
R13311 VDD.n1396 VDD 0.00324123
R13312 VDD.n2623 VDD 0.00324123
R13313 VDD.n2609 VDD 0.00324123
R13314 VDD.n2559 VDD 0.00324123
R13315 VDD.n2545 VDD 0.00324123
R13316 VDD.n2529 VDD 0.00324123
R13317 VDD.n2476 VDD 0.00324123
R13318 VDD.n1898 VDD.n1890 0.00284742
R13319 VDD.n1061 VDD.n1059 0.00282098
R13320 VDD.n932 VDD.n930 0.00282098
R13321 VDD.n803 VDD.n801 0.00282098
R13322 VDD.n652 VDD.n650 0.00282098
R13323 VDD.n523 VDD.n521 0.00282098
R13324 VDD.n394 VDD.n392 0.00282098
R13325 VDD.n265 VDD.n263 0.00282098
R13326 VDD.n127 VDD.n125 0.00282098
R13327 VDD.n2911 VDD.n2909 0.00282098
R13328 VDD.n687 VDD 0.0027381
R13329 VDD.n2538 VDD 0.00269298
R13330 VDD.n2682 VDD 0.00269298
R13331 VDD.n2700 VDD 0.00269298
R13332 VDD.n1709 VDD 0.00269298
R13333 VDD.n1773 VDD 0.00269298
R13334 VDD.n1752 VDD 0.00269298
R13335 VDD.n1833 VDD 0.00269298
R13336 VDD.n1687 VDD 0.00269298
R13337 VDD.n1813 VDD 0.00269298
R13338 VDD.n1852 VDD 0.00269298
R13339 VDD.n1501 VDD 0.00269298
R13340 VDD.n1549 VDD 0.00269298
R13341 VDD.n1525 VDD 0.00269298
R13342 VDD.n1477 VDD 0.00269298
R13343 VDD.n1733 VDD 0.00269298
R13344 VDD.n2666 VDD 0.00269298
R13345 VDD.n2433 VDD 0.00269298
R13346 VDD.n2602 VDD 0.00269298
R13347 VDD.n2453 VDD 0.00269298
R13348 VDD.n2522 VDD 0.00269298
R13349 VDD VDD.n1072 0.00258877
R13350 VDD VDD.n943 0.00258877
R13351 VDD VDD.n814 0.00258877
R13352 VDD VDD.n663 0.00258877
R13353 VDD VDD.n534 0.00258877
R13354 VDD VDD.n405 0.00258877
R13355 VDD VDD.n276 0.00258877
R13356 VDD VDD.n138 0.00258877
R13357 VDD VDD.n2922 0.00258877
R13358 VDD.n2045 VDD 0.00258333
R13359 VDD VDD.n2115 0.00258333
R13360 VDD.n2046 VDD 0.00258333
R13361 VDD.n2053 VDD 0.00258333
R13362 VDD.n2054 VDD 0.00258333
R13363 VDD VDD.n2057 0.00258333
R13364 VDD.n2058 VDD 0.00258333
R13365 VDD VDD.n2061 0.00258333
R13366 VDD.n2062 VDD 0.00258333
R13367 VDD VDD.n2065 0.00258333
R13368 VDD.n2066 VDD 0.00258333
R13369 VDD VDD.n2069 0.00258333
R13370 VDD.n2070 VDD 0.00258333
R13371 VDD VDD.n2073 0.00258333
R13372 VDD.n2074 VDD 0.00258333
R13373 VDD VDD.n2077 0.00258333
R13374 VDD.n2392 VDD 0.00226056
R13375 VDD.n2403 VDD 0.00226056
R13376 VDD.n2410 VDD 0.00226056
R13377 VDD.n2374 VDD 0.00226056
R13378 VDD.n1925 VDD.n1924 0.00226056
R13379 VDD.n1305 VDD 0.00226056
R13380 VDD.n1317 VDD 0.00226056
R13381 VDD.n1281 VDD 0.00226056
R13382 VDD.n1293 VDD 0.00226056
R13383 VDD.n1257 VDD 0.00226056
R13384 VDD.n1269 VDD 0.00226056
R13385 VDD.n1233 VDD 0.00226056
R13386 VDD.n1245 VDD 0.00226056
R13387 VDD.n1209 VDD 0.00226056
R13388 VDD.n1221 VDD 0.00226056
R13389 VDD.n1196 VDD 0.00226056
R13390 VDD.n1192 VDD 0.00226056
R13391 VDD.n2347 VDD.n2346 0.00219369
R13392 VDD.n2395 VDD.n2392 0.00167371
R13393 VDD.n2403 VDD.n2402 0.00167371
R13394 VDD.n2410 VDD.n2409 0.00167371
R13395 VDD.n2377 VDD.n2374 0.00167371
R13396 VDD.n1948 VDD 0.00167371
R13397 VDD.n1308 VDD.n1305 0.00167371
R13398 VDD.n1320 VDD.n1317 0.00167371
R13399 VDD.n1284 VDD.n1281 0.00167371
R13400 VDD.n1296 VDD.n1293 0.00167371
R13401 VDD.n1260 VDD.n1257 0.00167371
R13402 VDD.n1272 VDD.n1269 0.00167371
R13403 VDD.n1236 VDD.n1233 0.00167371
R13404 VDD.n1248 VDD.n1245 0.00167371
R13405 VDD.n1212 VDD.n1209 0.00167371
R13406 VDD.n1224 VDD.n1221 0.00167371
R13407 VDD.n1199 VDD.n1196 0.00167371
R13408 VDD.n1192 VDD.n1191 0.00167371
R13409 VDD.n150 VDD.n149 0.00157759
R13410 VDD.n2124 VDD 0.00154167
R13411 VDD.n2193 VDD 0.00154167
R13412 VDD VDD.n2127 0.00154167
R13413 VDD.n2185 VDD 0.00154167
R13414 VDD VDD.n2130 0.00154167
R13415 VDD.n2180 VDD 0.00154167
R13416 VDD VDD.n2133 0.00154167
R13417 VDD.n2150 VDD 0.00154167
R13418 VDD VDD.n2136 0.00154167
R13419 VDD.n2149 VDD 0.00154167
R13420 VDD VDD.n2139 0.00154167
R13421 VDD.n2148 VDD 0.00154167
R13422 VDD VDD.n2142 0.00154167
R13423 VDD.n2147 VDD 0.00154167
R13424 VDD VDD.n2145 0.00154167
R13425 VDD.n2146 VDD 0.00154167
R13426 VDD.n1137 VDD 0.00154022
R13427 VDD.n667 VDD 0.00116138
R13428 VDD.n2541 VDD.n2538 0.00104825
R13429 VDD.n2685 VDD.n2682 0.00104825
R13430 VDD.n2703 VDD.n2700 0.00104825
R13431 VDD.n1712 VDD.n1709 0.00104825
R13432 VDD.n1776 VDD.n1773 0.00104825
R13433 VDD.n1752 VDD.n1751 0.00104825
R13434 VDD.n1836 VDD.n1833 0.00104825
R13435 VDD.n1690 VDD.n1687 0.00104825
R13436 VDD.n1816 VDD.n1813 0.00104825
R13437 VDD.n1852 VDD.n1851 0.00104825
R13438 VDD.n1504 VDD.n1501 0.00104825
R13439 VDD.n1552 VDD.n1549 0.00104825
R13440 VDD.n1528 VDD.n1525 0.00104825
R13441 VDD.n1480 VDD.n1477 0.00104825
R13442 VDD.n1736 VDD.n1733 0.00104825
R13443 VDD.n2669 VDD.n2666 0.00104825
R13444 VDD.n2627 VDD.n2433 0.00104825
R13445 VDD.n2605 VDD.n2602 0.00104825
R13446 VDD.n2563 VDD.n2453 0.00104825
R13447 VDD.n2525 VDD.n2522 0.00104825
R13448 VDD.n685 VDD 0.000820513
R13449 mux8_2.NAND4F_0.Y.n1 mux8_2.NAND4F_0.Y.t10 1388.16
R13450 mux8_2.NAND4F_0.Y.n1 mux8_2.NAND4F_0.Y.t9 350.839
R13451 mux8_2.NAND4F_0.Y.n2 mux8_2.NAND4F_0.Y.t11 308.481
R13452 mux8_2.NAND4F_0.Y.n0 mux8_2.NAND4F_0.Y.n3 187.373
R13453 mux8_2.NAND4F_0.Y.n0 mux8_2.NAND4F_0.Y.n4 187.192
R13454 mux8_2.NAND4F_0.Y.n0 mux8_2.NAND4F_0.Y.n5 187.192
R13455 mux8_2.NAND4F_0.Y mux8_2.NAND4F_0.Y.n6 187.192
R13456 mux8_2.NAND4F_0.Y mux8_2.NAND4F_0.Y.n2 161.492
R13457 mux8_2.NAND4F_0.Y.n2 mux8_2.NAND4F_0.Y.n1 27.752
R13458 mux8_2.NAND4F_0.Y mux8_2.NAND4F_0.Y.t2 23.5085
R13459 mux8_2.NAND4F_0.Y.n3 mux8_2.NAND4F_0.Y.t6 20.1899
R13460 mux8_2.NAND4F_0.Y.n3 mux8_2.NAND4F_0.Y.t5 20.1899
R13461 mux8_2.NAND4F_0.Y.n4 mux8_2.NAND4F_0.Y.t8 20.1899
R13462 mux8_2.NAND4F_0.Y.n4 mux8_2.NAND4F_0.Y.t7 20.1899
R13463 mux8_2.NAND4F_0.Y.n5 mux8_2.NAND4F_0.Y.t3 20.1899
R13464 mux8_2.NAND4F_0.Y.n5 mux8_2.NAND4F_0.Y.t4 20.1899
R13465 mux8_2.NAND4F_0.Y.n6 mux8_2.NAND4F_0.Y.t1 20.1899
R13466 mux8_2.NAND4F_0.Y.n6 mux8_2.NAND4F_0.Y.t0 20.1899
R13467 mux8_2.NAND4F_0.Y mux8_2.NAND4F_0.Y.n0 0.358709
R13468 a_n12446_n11709.n2 a_n12446_n11709.t3 541.395
R13469 a_n12446_n11709.n3 a_n12446_n11709.t7 527.402
R13470 a_n12446_n11709.n2 a_n12446_n11709.t6 491.64
R13471 a_n12446_n11709.n5 a_n12446_n11709.t0 281.906
R13472 a_n12446_n11709.t1 a_n12446_n11709.n5 204.359
R13473 a_n12446_n11709.n0 a_n12446_n11709.t2 180.73
R13474 a_n12446_n11709.n1 a_n12446_n11709.t4 179.45
R13475 a_n12446_n11709.n0 a_n12446_n11709.t5 139.78
R13476 a_n12446_n11709.n4 a_n12446_n11709.n1 105.635
R13477 a_n12446_n11709.n4 a_n12446_n11709.n3 76.0005
R13478 a_n12446_n11709.n5 a_n12446_n11709.n4 67.9685
R13479 a_n12446_n11709.n3 a_n12446_n11709.n2 13.994
R13480 a_n12446_n11709.n1 a_n12446_n11709.n0 1.28015
R13481 a_n12416_n11683.n2 a_n12416_n11683.n1 121.353
R13482 a_n12416_n11683.n3 a_n12416_n11683.n2 121.001
R13483 a_n12416_n11683.n2 a_n12416_n11683.n0 120.977
R13484 a_n12416_n11683.n1 a_n12416_n11683.t0 30.462
R13485 a_n12416_n11683.n1 a_n12416_n11683.t1 30.462
R13486 a_n12416_n11683.n0 a_n12416_n11683.t4 30.462
R13487 a_n12416_n11683.n0 a_n12416_n11683.t5 30.462
R13488 a_n12416_n11683.n3 a_n12416_n11683.t3 30.462
R13489 a_n12416_n11683.t2 a_n12416_n11683.n3 30.462
R13490 mux8_5.NAND4F_8.Y.n1 mux8_5.NAND4F_8.Y.t13 379.173
R13491 mux8_5.NAND4F_8.Y.n2 mux8_5.NAND4F_8.Y.t12 312.599
R13492 mux8_5.NAND4F_8.Y.n1 mux8_5.NAND4F_8.Y.t14 247.428
R13493 mux8_5.NAND4F_8.Y.n4 mux8_5.NAND4F_8.Y.t9 247.428
R13494 mux8_5.NAND4F_8.Y.n3 mux8_5.NAND4F_8.Y.t11 247.428
R13495 mux8_5.NAND4F_8.Y.n2 mux8_5.NAND4F_8.Y.t10 247.428
R13496 mux8_5.NAND4F_8.Y.n0 mux8_5.NAND4F_8.Y.n6 187.373
R13497 mux8_5.NAND4F_8.Y.n0 mux8_5.NAND4F_8.Y.n7 187.192
R13498 mux8_5.NAND4F_8.Y.n0 mux8_5.NAND4F_8.Y.n8 187.192
R13499 mux8_5.NAND4F_8.Y.n10 mux8_5.NAND4F_8.Y.n9 187.192
R13500 mux8_5.NAND4F_8.Y mux8_5.NAND4F_8.Y.n5 162.139
R13501 mux8_5.NAND4F_8.Y.n4 mux8_5.NAND4F_8.Y.n3 65.1723
R13502 mux8_5.NAND4F_8.Y.n3 mux8_5.NAND4F_8.Y.n2 65.1723
R13503 mux8_5.NAND4F_8.Y.n5 mux8_5.NAND4F_8.Y.n4 33.2653
R13504 mux8_5.NAND4F_8.Y.n5 mux8_5.NAND4F_8.Y.n1 31.9075
R13505 mux8_5.NAND4F_8.Y mux8_5.NAND4F_8.Y.t2 22.6141
R13506 mux8_5.NAND4F_8.Y.n6 mux8_5.NAND4F_8.Y.t6 20.1899
R13507 mux8_5.NAND4F_8.Y.n6 mux8_5.NAND4F_8.Y.t5 20.1899
R13508 mux8_5.NAND4F_8.Y.n7 mux8_5.NAND4F_8.Y.t7 20.1899
R13509 mux8_5.NAND4F_8.Y.n7 mux8_5.NAND4F_8.Y.t8 20.1899
R13510 mux8_5.NAND4F_8.Y.n8 mux8_5.NAND4F_8.Y.t3 20.1899
R13511 mux8_5.NAND4F_8.Y.n8 mux8_5.NAND4F_8.Y.t4 20.1899
R13512 mux8_5.NAND4F_8.Y.n9 mux8_5.NAND4F_8.Y.t0 20.1899
R13513 mux8_5.NAND4F_8.Y.n9 mux8_5.NAND4F_8.Y.t1 20.1899
R13514 mux8_5.NAND4F_8.Y mux8_5.NAND4F_8.Y.n10 0.452586
R13515 mux8_5.NAND4F_8.Y.n10 mux8_5.NAND4F_8.Y.n0 0.358709
R13516 a_11865_n20887.n0 a_11865_n20887.n2 231.24
R13517 a_11865_n20887.n6 a_11865_n20887.n1 231.24
R13518 a_11865_n20887.n1 a_11865_n20887.n5 231.03
R13519 a_11865_n20887.n1 a_11865_n20887.n4 231.03
R13520 a_11865_n20887.n0 a_11865_n20887.n3 231.03
R13521 a_11865_n20887.n5 a_11865_n20887.t9 25.395
R13522 a_11865_n20887.n5 a_11865_n20887.t7 25.395
R13523 a_11865_n20887.n4 a_11865_n20887.t3 25.395
R13524 a_11865_n20887.n4 a_11865_n20887.t5 25.395
R13525 a_11865_n20887.n3 a_11865_n20887.t1 25.395
R13526 a_11865_n20887.n3 a_11865_n20887.t2 25.395
R13527 a_11865_n20887.n2 a_11865_n20887.t4 25.395
R13528 a_11865_n20887.n2 a_11865_n20887.t0 25.395
R13529 a_11865_n20887.t8 a_11865_n20887.n6 25.395
R13530 a_11865_n20887.n6 a_11865_n20887.t6 25.395
R13531 a_11865_n20887.n1 a_11865_n20887.n0 0.421553
R13532 mux8_1.NAND4F_8.Y.n1 mux8_1.NAND4F_8.Y.t14 379.173
R13533 mux8_1.NAND4F_8.Y.n2 mux8_1.NAND4F_8.Y.t10 312.599
R13534 mux8_1.NAND4F_8.Y.n1 mux8_1.NAND4F_8.Y.t9 247.428
R13535 mux8_1.NAND4F_8.Y.n4 mux8_1.NAND4F_8.Y.t13 247.428
R13536 mux8_1.NAND4F_8.Y.n3 mux8_1.NAND4F_8.Y.t12 247.428
R13537 mux8_1.NAND4F_8.Y.n2 mux8_1.NAND4F_8.Y.t11 247.428
R13538 mux8_1.NAND4F_8.Y.n0 mux8_1.NAND4F_8.Y.n6 187.373
R13539 mux8_1.NAND4F_8.Y.n0 mux8_1.NAND4F_8.Y.n7 187.192
R13540 mux8_1.NAND4F_8.Y.n0 mux8_1.NAND4F_8.Y.n8 187.192
R13541 mux8_1.NAND4F_8.Y.n10 mux8_1.NAND4F_8.Y.n9 187.192
R13542 mux8_1.NAND4F_8.Y mux8_1.NAND4F_8.Y.n5 162.139
R13543 mux8_1.NAND4F_8.Y.n4 mux8_1.NAND4F_8.Y.n3 65.1723
R13544 mux8_1.NAND4F_8.Y.n3 mux8_1.NAND4F_8.Y.n2 65.1723
R13545 mux8_1.NAND4F_8.Y.n5 mux8_1.NAND4F_8.Y.n4 33.2653
R13546 mux8_1.NAND4F_8.Y.n5 mux8_1.NAND4F_8.Y.n1 31.9075
R13547 mux8_1.NAND4F_8.Y mux8_1.NAND4F_8.Y.t5 22.6141
R13548 mux8_1.NAND4F_8.Y.n6 mux8_1.NAND4F_8.Y.t6 20.1899
R13549 mux8_1.NAND4F_8.Y.n6 mux8_1.NAND4F_8.Y.t7 20.1899
R13550 mux8_1.NAND4F_8.Y.n7 mux8_1.NAND4F_8.Y.t4 20.1899
R13551 mux8_1.NAND4F_8.Y.n7 mux8_1.NAND4F_8.Y.t3 20.1899
R13552 mux8_1.NAND4F_8.Y.n8 mux8_1.NAND4F_8.Y.t8 20.1899
R13553 mux8_1.NAND4F_8.Y.n8 mux8_1.NAND4F_8.Y.t2 20.1899
R13554 mux8_1.NAND4F_8.Y.n9 mux8_1.NAND4F_8.Y.t1 20.1899
R13555 mux8_1.NAND4F_8.Y.n9 mux8_1.NAND4F_8.Y.t0 20.1899
R13556 mux8_1.NAND4F_8.Y mux8_1.NAND4F_8.Y.n10 0.452586
R13557 mux8_1.NAND4F_8.Y.n10 mux8_1.NAND4F_8.Y.n0 0.358709
R13558 a_11865_n2775.n0 a_11865_n2775.n2 231.24
R13559 a_11865_n2775.n6 a_11865_n2775.n1 231.24
R13560 a_11865_n2775.n1 a_11865_n2775.n5 231.03
R13561 a_11865_n2775.n1 a_11865_n2775.n4 231.03
R13562 a_11865_n2775.n0 a_11865_n2775.n3 231.03
R13563 a_11865_n2775.n5 a_11865_n2775.t5 25.395
R13564 a_11865_n2775.n5 a_11865_n2775.t6 25.395
R13565 a_11865_n2775.n4 a_11865_n2775.t0 25.395
R13566 a_11865_n2775.n4 a_11865_n2775.t9 25.395
R13567 a_11865_n2775.n3 a_11865_n2775.t2 25.395
R13568 a_11865_n2775.n3 a_11865_n2775.t1 25.395
R13569 a_11865_n2775.n2 a_11865_n2775.t4 25.395
R13570 a_11865_n2775.n2 a_11865_n2775.t3 25.395
R13571 a_11865_n2775.n6 a_11865_n2775.t7 25.395
R13572 a_11865_n2775.t8 a_11865_n2775.n6 25.395
R13573 a_11865_n2775.n1 a_11865_n2775.n0 0.421553
R13574 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t7 485.221
R13575 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t8 367.928
R13576 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n3 227.526
R13577 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n5 227.266
R13578 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n4 227.266
R13579 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t10 224.478
R13580 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t9 213.688
R13581 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n1 84.5046
R13582 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n0 72.3005
R13583 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n2 61.0566
R13584 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t1 43.3573
R13585 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t2 30.379
R13586 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t4 30.379
R13587 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t6 30.379
R13588 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t0 30.379
R13589 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t3 30.379
R13590 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A.t5 30.379
R13591 a_n18305_n6187.t0 a_n18305_n6187.t1 19.8005
R13592 a_n20839_3190.n2 a_n20839_3190.t6 541.395
R13593 a_n20839_3190.n3 a_n20839_3190.t3 527.402
R13594 a_n20839_3190.n2 a_n20839_3190.t5 491.64
R13595 a_n20839_3190.n5 a_n20839_3190.t0 281.906
R13596 a_n20839_3190.t1 a_n20839_3190.n5 204.359
R13597 a_n20839_3190.n0 a_n20839_3190.t7 180.73
R13598 a_n20839_3190.n1 a_n20839_3190.t4 179.45
R13599 a_n20839_3190.n0 a_n20839_3190.t2 139.78
R13600 a_n20839_3190.n4 a_n20839_3190.n1 105.635
R13601 a_n20839_3190.n4 a_n20839_3190.n3 76.0005
R13602 a_n20839_3190.n5 a_n20839_3190.n4 67.9685
R13603 a_n20839_3190.n3 a_n20839_3190.n2 13.994
R13604 a_n20839_3190.n1 a_n20839_3190.n0 1.28015
R13605 a_n20083_3190.n3 a_n20083_3190.n2 121.353
R13606 a_n20083_3190.n2 a_n20083_3190.n1 121.001
R13607 a_n20083_3190.n2 a_n20083_3190.n0 120.977
R13608 a_n20083_3190.n0 a_n20083_3190.t3 30.462
R13609 a_n20083_3190.n0 a_n20083_3190.t5 30.462
R13610 a_n20083_3190.n1 a_n20083_3190.t0 30.462
R13611 a_n20083_3190.n1 a_n20083_3190.t4 30.462
R13612 a_n20083_3190.n3 a_n20083_3190.t1 30.462
R13613 a_n20083_3190.t2 a_n20083_3190.n3 30.462
R13614 MULT_0.inv_13.A.n4 MULT_0.inv_13.A.t9 291.829
R13615 MULT_0.inv_13.A.n4 MULT_0.inv_13.A.t7 291.829
R13616 MULT_0.inv_13.A.n0 MULT_0.inv_13.A.n1 227.526
R13617 MULT_0.inv_13.A.n0 MULT_0.inv_13.A.n3 227.266
R13618 MULT_0.inv_13.A.n0 MULT_0.inv_13.A.n2 227.266
R13619 MULT_0.inv_13.A.n4 MULT_0.inv_13.A.t10 221.72
R13620 MULT_0.inv_13.A.t8 MULT_0.inv_13.A.n0 393.897
R13621 MULT_0.inv_13.A.n3 MULT_0.inv_13.A.t3 30.379
R13622 MULT_0.inv_13.A.n3 MULT_0.inv_13.A.t4 30.379
R13623 MULT_0.inv_13.A.n1 MULT_0.inv_13.A.t1 30.379
R13624 MULT_0.inv_13.A.n1 MULT_0.inv_13.A.t2 30.379
R13625 MULT_0.inv_13.A.n2 MULT_0.inv_13.A.t5 30.379
R13626 MULT_0.inv_13.A.n2 MULT_0.inv_13.A.t0 30.379
R13627 MULT_0.inv_13.A.n4 MULT_0.inv_13.A.n0 53.491
R13628 MULT_0.inv_13.A.n0 MULT_0.inv_13.A.t6 43.3529
R13629 MULT_0.4bit_ADDER_1.A3.n3 MULT_0.4bit_ADDER_1.A3.t6 540.38
R13630 MULT_0.4bit_ADDER_1.A3.n4 MULT_0.4bit_ADDER_1.A3.t12 491.64
R13631 MULT_0.4bit_ADDER_1.A3.n4 MULT_0.4bit_ADDER_1.A3.t7 491.64
R13632 MULT_0.4bit_ADDER_1.A3.n4 MULT_0.4bit_ADDER_1.A3.t5 491.64
R13633 MULT_0.4bit_ADDER_1.A3.n4 MULT_0.4bit_ADDER_1.A3.t9 491.64
R13634 MULT_0.4bit_ADDER_1.A3.n1 MULT_0.4bit_ADDER_1.A3.t4 367.928
R13635 MULT_0.inv_13.Y MULT_0.4bit_ADDER_1.A3.t3 256.514
R13636 MULT_0.4bit_ADDER_1.A3.n2 MULT_0.4bit_ADDER_1.A3.t14 227.356
R13637 MULT_0.inv_13.Y MULT_0.4bit_ADDER_1.A3.n7 226.248
R13638 MULT_0.4bit_ADDER_1.A3.n1 MULT_0.4bit_ADDER_1.A3.t10 213.688
R13639 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_0.B MULT_0.4bit_ADDER_1.A3.n6 162.867
R13640 MULT_0.4bit_ADDER_1.A3.n3 MULT_0.4bit_ADDER_1.A3.n2 160.439
R13641 MULT_0.4bit_ADDER_1.A3.n5 MULT_0.4bit_ADDER_1.A3.t11 139.78
R13642 MULT_0.4bit_ADDER_1.A3.n5 MULT_0.4bit_ADDER_1.A3.t15 139.78
R13643 MULT_0.4bit_ADDER_1.A3.n5 MULT_0.4bit_ADDER_1.A3.t8 139.78
R13644 MULT_0.4bit_ADDER_1.A3.n5 MULT_0.4bit_ADDER_1.A3.t13 139.78
R13645 MULT_0.4bit_ADDER_1.A3.n2 MULT_0.4bit_ADDER_1.A3.n1 94.4341
R13646 MULT_0.inv_13.Y MULT_0.4bit_ADDER_1.A3.t0 83.8155
R13647 MULT_0.4bit_ADDER_1.A3.n6 MULT_0.4bit_ADDER_1.A3.n5 38.6833
R13648 MULT_0.4bit_ADDER_1.A3.n7 MULT_0.4bit_ADDER_1.A3.t2 30.379
R13649 MULT_0.4bit_ADDER_1.A3.n7 MULT_0.4bit_ADDER_1.A3.t1 30.379
R13650 MULT_0.4bit_ADDER_1.A3.n6 MULT_0.4bit_ADDER_1.A3.n4 28.3986
R13651 MULT_0.4bit_ADDER_1.A3.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_0.B 9.00496
R13652 MULT_0.4bit_ADDER_1.A3.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_0.B 3.87912
R13653 MULT_0.inv_13.Y MULT_0.4bit_ADDER_1.A3.n0 3.07356
R13654 MULT_0.4bit_ADDER_1.A3.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.A 1.47848
R13655 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_0.B MULT_0.4bit_ADDER_1.A3.n3 0.89693
R13656 SEL1.n176 SEL1.t8 978.795
R13657 SEL1.n173 SEL1.t80 978.795
R13658 SEL1.n169 SEL1.t33 978.795
R13659 SEL1.n167 SEL1.t110 978.795
R13660 SEL1.n155 SEL1.t26 978.795
R13661 SEL1.n152 SEL1.t89 978.795
R13662 SEL1.n148 SEL1.t45 978.795
R13663 SEL1.n146 SEL1.t123 978.795
R13664 SEL1.n134 SEL1.t83 978.795
R13665 SEL1.n131 SEL1.t124 978.795
R13666 SEL1.n127 SEL1.t42 978.795
R13667 SEL1.n125 SEL1.t143 978.795
R13668 SEL1.n113 SEL1.t13 978.795
R13669 SEL1.n110 SEL1.t57 978.795
R13670 SEL1.n106 SEL1.t107 978.795
R13671 SEL1.n104 SEL1.t72 978.795
R13672 SEL1.n92 SEL1.t3 978.795
R13673 SEL1.n89 SEL1.t50 978.795
R13674 SEL1.n85 SEL1.t139 978.795
R13675 SEL1.n83 SEL1.t106 978.795
R13676 SEL1.n71 SEL1.t119 978.795
R13677 SEL1.n68 SEL1.t7 978.795
R13678 SEL1.n64 SEL1.t76 978.795
R13679 SEL1.n62 SEL1.t40 978.795
R13680 SEL1.n50 SEL1.t131 978.795
R13681 SEL1.n47 SEL1.t21 978.795
R13682 SEL1.n43 SEL1.t109 978.795
R13683 SEL1.n41 SEL1.t75 978.795
R13684 SEL1.n30 SEL1.t85 978.795
R13685 SEL1.n27 SEL1.t129 978.795
R13686 SEL1.n23 SEL1.t79 978.795
R13687 SEL1.n21 SEL1.t41 978.795
R13688 SEL1.n11 SEL1.t67 978.795
R13689 SEL1.n8 SEL1.t90 978.795
R13690 SEL1.n4 SEL1.t53 978.795
R13691 SEL1.n2 SEL1.t134 978.795
R13692 SEL1.n181 SEL1.t118 385.697
R13693 SEL1.n160 SEL1.t125 385.697
R13694 SEL1.n139 SEL1.t94 385.697
R13695 SEL1.n118 SEL1.t18 385.697
R13696 SEL1.n97 SEL1.t133 385.697
R13697 SEL1.n76 SEL1.t24 385.697
R13698 SEL1.n55 SEL1.t97 385.697
R13699 SEL1.n35 SEL1.t91 385.697
R13700 SEL1.n16 SEL1.t35 385.697
R13701 SEL1.n175 SEL1.t30 308.481
R13702 SEL1.n175 SEL1.t82 308.481
R13703 SEL1.n172 SEL1.t141 308.481
R13704 SEL1.n172 SEL1.t56 308.481
R13705 SEL1.n168 SEL1.t61 308.481
R13706 SEL1.n168 SEL1.t1 308.481
R13707 SEL1.n166 SEL1.t84 308.481
R13708 SEL1.n166 SEL1.t37 308.481
R13709 SEL1.n154 SEL1.t138 308.481
R13710 SEL1.n154 SEL1.t54 308.481
R13711 SEL1.n151 SEL1.t113 308.481
R13712 SEL1.n151 SEL1.t17 308.481
R13713 SEL1.n147 SEL1.t27 308.481
R13714 SEL1.n147 SEL1.t116 308.481
R13715 SEL1.n145 SEL1.t59 308.481
R13716 SEL1.n145 SEL1.t0 308.481
R13717 SEL1.n133 SEL1.t23 308.481
R13718 SEL1.n133 SEL1.t108 308.481
R13719 SEL1.n130 SEL1.t44 308.481
R13720 SEL1.n130 SEL1.t132 308.481
R13721 SEL1.n126 SEL1.t137 308.481
R13722 SEL1.n126 SEL1.t58 308.481
R13723 SEL1.n124 SEL1.t121 308.481
R13724 SEL1.n124 SEL1.t36 308.481
R13725 SEL1.n112 SEL1.t96 308.481
R13726 SEL1.n112 SEL1.t43 308.481
R13727 SEL1.n109 SEL1.t117 308.481
R13728 SEL1.n109 SEL1.t63 308.481
R13729 SEL1.n105 SEL1.t66 308.481
R13730 SEL1.n105 SEL1.t122 308.481
R13731 SEL1.n103 SEL1.t48 308.481
R13732 SEL1.n103 SEL1.t100 308.481
R13733 SEL1.n91 SEL1.t60 308.481
R13734 SEL1.n91 SEL1.t140 308.481
R13735 SEL1.n88 SEL1.t77 308.481
R13736 SEL1.n88 SEL1.t20 308.481
R13737 SEL1.n84 SEL1.t68 308.481
R13738 SEL1.n84 SEL1.t127 308.481
R13739 SEL1.n82 SEL1.t49 308.481
R13740 SEL1.n82 SEL1.t101 308.481
R13741 SEL1.n70 SEL1.t98 308.481
R13742 SEL1.n70 SEL1.t46 308.481
R13743 SEL1.n67 SEL1.t120 308.481
R13744 SEL1.n67 SEL1.t64 308.481
R13745 SEL1.n63 SEL1.t34 308.481
R13746 SEL1.n63 SEL1.t88 308.481
R13747 SEL1.n61 SEL1.t5 308.481
R13748 SEL1.n61 SEL1.t70 308.481
R13749 SEL1.n49 SEL1.t11 308.481
R13750 SEL1.n49 SEL1.t102 308.481
R13751 SEL1.n46 SEL1.t39 308.481
R13752 SEL1.n46 SEL1.t128 308.481
R13753 SEL1.n42 SEL1.t71 308.481
R13754 SEL1.n42 SEL1.t130 308.481
R13755 SEL1.n40 SEL1.t51 308.481
R13756 SEL1.n40 SEL1.t103 308.481
R13757 SEL1.n29 SEL1.t25 308.481
R13758 SEL1.n29 SEL1.t111 308.481
R13759 SEL1.n26 SEL1.t47 308.481
R13760 SEL1.n26 SEL1.t135 308.481
R13761 SEL1.n22 SEL1.t38 308.481
R13762 SEL1.n22 SEL1.t92 308.481
R13763 SEL1.n20 SEL1.t10 308.481
R13764 SEL1.n20 SEL1.t73 308.481
R13765 SEL1.n10 SEL1.t87 308.481
R13766 SEL1.n10 SEL1.t19 308.481
R13767 SEL1.n7 SEL1.t78 308.481
R13768 SEL1.n7 SEL1.t2 308.481
R13769 SEL1.n3 SEL1.t4 308.481
R13770 SEL1.n3 SEL1.t105 308.481
R13771 SEL1.n1 SEL1.t29 308.481
R13772 SEL1.n1 SEL1.t126 308.481
R13773 SEL1.n165 SEL1.t55 291.829
R13774 SEL1.n165 SEL1.t104 291.829
R13775 SEL1.n144 SEL1.t112 291.829
R13776 SEL1.n144 SEL1.t22 291.829
R13777 SEL1.n123 SEL1.t28 291.829
R13778 SEL1.n123 SEL1.t81 291.829
R13779 SEL1.n102 SEL1.t86 291.829
R13780 SEL1.n102 SEL1.t136 291.829
R13781 SEL1.n81 SEL1.t114 291.829
R13782 SEL1.n81 SEL1.t74 291.829
R13783 SEL1.n60 SEL1.t6 291.829
R13784 SEL1.n60 SEL1.t65 291.829
R13785 SEL1.n39 SEL1.t115 291.829
R13786 SEL1.n39 SEL1.t31 291.829
R13787 SEL1.n19 SEL1.t9 291.829
R13788 SEL1.n19 SEL1.t69 291.829
R13789 SEL1.n0 SEL1.t95 291.829
R13790 SEL1.n0 SEL1.t142 291.829
R13791 SEL1.n165 SEL1.t99 221.72
R13792 SEL1.n144 SEL1.t12 221.72
R13793 SEL1.n123 SEL1.t32 221.72
R13794 SEL1.n102 SEL1.t93 221.72
R13795 SEL1.n81 SEL1.t14 221.72
R13796 SEL1.n60 SEL1.t62 221.72
R13797 SEL1.n39 SEL1.t15 221.72
R13798 SEL1.n19 SEL1.t16 221.72
R13799 SEL1.n0 SEL1.t52 221.72
R13800 SEL1 SEL1.n167 161.911
R13801 SEL1 SEL1.n146 161.911
R13802 SEL1 SEL1.n125 161.911
R13803 SEL1 SEL1.n104 161.911
R13804 SEL1 SEL1.n83 161.911
R13805 SEL1 SEL1.n62 161.911
R13806 SEL1 SEL1.n41 161.911
R13807 SEL1 SEL1.n21 161.911
R13808 SEL1 SEL1.n2 161.911
R13809 SEL1.n174 SEL1.n173 161.869
R13810 SEL1.n153 SEL1.n152 161.869
R13811 SEL1.n132 SEL1.n131 161.869
R13812 SEL1.n111 SEL1.n110 161.869
R13813 SEL1.n90 SEL1.n89 161.869
R13814 SEL1.n69 SEL1.n68 161.869
R13815 SEL1.n48 SEL1.n47 161.869
R13816 SEL1.n28 SEL1.n27 161.869
R13817 SEL1.n9 SEL1.n8 161.869
R13818 SEL1.n177 SEL1.n176 161.862
R13819 SEL1.n156 SEL1.n155 161.862
R13820 SEL1.n135 SEL1.n134 161.862
R13821 SEL1.n114 SEL1.n113 161.862
R13822 SEL1.n93 SEL1.n92 161.862
R13823 SEL1.n72 SEL1.n71 161.862
R13824 SEL1.n51 SEL1.n50 161.862
R13825 SEL1.n31 SEL1.n30 161.862
R13826 SEL1.n12 SEL1.n11 161.862
R13827 SEL1.n170 SEL1.n169 161.827
R13828 SEL1.n149 SEL1.n148 161.827
R13829 SEL1.n128 SEL1.n127 161.827
R13830 SEL1.n107 SEL1.n106 161.827
R13831 SEL1.n86 SEL1.n85 161.827
R13832 SEL1.n65 SEL1.n64 161.827
R13833 SEL1.n44 SEL1.n43 161.827
R13834 SEL1.n24 SEL1.n23 161.827
R13835 SEL1.n5 SEL1.n4 161.827
R13836 SEL1.n182 SEL1.n181 89.6005
R13837 SEL1.n161 SEL1.n160 89.6005
R13838 SEL1.n140 SEL1.n139 89.6005
R13839 SEL1.n119 SEL1.n118 89.6005
R13840 SEL1.n98 SEL1.n97 89.6005
R13841 SEL1.n77 SEL1.n76 89.6005
R13842 SEL1.n56 SEL1.n55 89.6005
R13843 SEL1.n36 SEL1.n35 89.6005
R13844 SEL1.n17 SEL1.n16 89.6005
R13845 SEL1.n182 SEL1.n165 50.6672
R13846 SEL1.n161 SEL1.n144 50.6672
R13847 SEL1.n140 SEL1.n123 50.6672
R13848 SEL1.n119 SEL1.n102 50.6672
R13849 SEL1.n98 SEL1.n81 50.6672
R13850 SEL1.n77 SEL1.n60 50.6672
R13851 SEL1.n56 SEL1.n39 50.6672
R13852 SEL1.n36 SEL1.n19 50.6672
R13853 SEL1.n17 SEL1.n0 50.6672
R13854 SEL1.n171 SEL1.n170 21.7997
R13855 SEL1.n150 SEL1.n149 21.7997
R13856 SEL1.n129 SEL1.n128 21.7997
R13857 SEL1.n108 SEL1.n107 21.7997
R13858 SEL1.n87 SEL1.n86 21.7997
R13859 SEL1.n66 SEL1.n65 21.7997
R13860 SEL1.n45 SEL1.n44 21.7997
R13861 SEL1.n25 SEL1.n24 21.7997
R13862 SEL1.n6 SEL1.n5 21.7997
R13863 SEL1.n179 SEL1.n178 11.3222
R13864 SEL1.n158 SEL1.n157 11.3222
R13865 SEL1.n137 SEL1.n136 11.3222
R13866 SEL1.n116 SEL1.n115 11.3222
R13867 SEL1.n95 SEL1.n94 11.3222
R13868 SEL1.n74 SEL1.n73 11.3222
R13869 SEL1.n53 SEL1.n52 11.3222
R13870 SEL1.n33 SEL1.n32 11.3222
R13871 SEL1.n14 SEL1.n13 11.3222
R13872 SEL1.n176 SEL1.n175 11.0463
R13873 SEL1.n173 SEL1.n172 11.0463
R13874 SEL1.n169 SEL1.n168 11.0463
R13875 SEL1.n167 SEL1.n166 11.0463
R13876 SEL1.n155 SEL1.n154 11.0463
R13877 SEL1.n152 SEL1.n151 11.0463
R13878 SEL1.n148 SEL1.n147 11.0463
R13879 SEL1.n146 SEL1.n145 11.0463
R13880 SEL1.n134 SEL1.n133 11.0463
R13881 SEL1.n131 SEL1.n130 11.0463
R13882 SEL1.n127 SEL1.n126 11.0463
R13883 SEL1.n125 SEL1.n124 11.0463
R13884 SEL1.n113 SEL1.n112 11.0463
R13885 SEL1.n110 SEL1.n109 11.0463
R13886 SEL1.n106 SEL1.n105 11.0463
R13887 SEL1.n104 SEL1.n103 11.0463
R13888 SEL1.n92 SEL1.n91 11.0463
R13889 SEL1.n89 SEL1.n88 11.0463
R13890 SEL1.n85 SEL1.n84 11.0463
R13891 SEL1.n83 SEL1.n82 11.0463
R13892 SEL1.n71 SEL1.n70 11.0463
R13893 SEL1.n68 SEL1.n67 11.0463
R13894 SEL1.n64 SEL1.n63 11.0463
R13895 SEL1.n62 SEL1.n61 11.0463
R13896 SEL1.n50 SEL1.n49 11.0463
R13897 SEL1.n47 SEL1.n46 11.0463
R13898 SEL1.n43 SEL1.n42 11.0463
R13899 SEL1.n41 SEL1.n40 11.0463
R13900 SEL1.n30 SEL1.n29 11.0463
R13901 SEL1.n27 SEL1.n26 11.0463
R13902 SEL1.n23 SEL1.n22 11.0463
R13903 SEL1.n21 SEL1.n20 11.0463
R13904 SEL1.n11 SEL1.n10 11.0463
R13905 SEL1.n8 SEL1.n7 11.0463
R13906 SEL1.n4 SEL1.n3 11.0463
R13907 SEL1.n2 SEL1.n1 11.0463
R13908 SEL1.n178 SEL1.n174 11.0005
R13909 SEL1.n157 SEL1.n153 11.0005
R13910 SEL1.n136 SEL1.n132 11.0005
R13911 SEL1.n115 SEL1.n111 11.0005
R13912 SEL1.n94 SEL1.n90 11.0005
R13913 SEL1.n73 SEL1.n69 11.0005
R13914 SEL1.n52 SEL1.n48 11.0005
R13915 SEL1.n32 SEL1.n28 11.0005
R13916 SEL1.n13 SEL1.n9 11.0005
R13917 SEL1 SEL1.n183 9.57444
R13918 SEL1.n185 SEL1.n18 9.55995
R13919 SEL1.n121 SEL1.n120 9.53096
R13920 SEL1.n79 SEL1.n78 9.53096
R13921 SEL1.n163 SEL1.n162 9.52734
R13922 SEL1.n100 SEL1.n99 9.50922
R13923 SEL1.n58 SEL1.n57 9.50017
R13924 SEL1.n38 SEL1.n37 9.49835
R13925 SEL1.n142 SEL1.n141 9.49111
R13926 SEL1.n181 SEL1.n180 9.3005
R13927 SEL1.n160 SEL1.n159 9.3005
R13928 SEL1.n139 SEL1.n138 9.3005
R13929 SEL1.n118 SEL1.n117 9.3005
R13930 SEL1.n97 SEL1.n96 9.3005
R13931 SEL1.n76 SEL1.n75 9.3005
R13932 SEL1.n55 SEL1.n54 9.3005
R13933 SEL1.n35 SEL1.n34 9.3005
R13934 SEL1.n16 SEL1.n15 9.3005
R13935 SEL1.n178 SEL1.n177 9.0005
R13936 SEL1.n157 SEL1.n156 9.0005
R13937 SEL1.n136 SEL1.n135 9.0005
R13938 SEL1.n115 SEL1.n114 9.0005
R13939 SEL1.n94 SEL1.n93 9.0005
R13940 SEL1.n73 SEL1.n72 9.0005
R13941 SEL1.n52 SEL1.n51 9.0005
R13942 SEL1.n32 SEL1.n31 9.0005
R13943 SEL1.n13 SEL1.n12 9.0005
R13944 SEL1.n59 SEL1.n38 6.49547
R13945 SEL1.n185 SEL1.n184 6.48453
R13946 SEL1.n179 SEL1.n171 4.08298
R13947 SEL1.n158 SEL1.n150 4.08298
R13948 SEL1.n137 SEL1.n129 4.08298
R13949 SEL1.n116 SEL1.n108 4.08298
R13950 SEL1.n95 SEL1.n87 4.08298
R13951 SEL1.n74 SEL1.n66 4.08298
R13952 SEL1.n53 SEL1.n45 4.08298
R13953 SEL1.n33 SEL1.n25 4.08298
R13954 SEL1.n14 SEL1.n6 4.08298
R13955 SEL1.n184 SEL1 3.41412
R13956 SEL1.n59 SEL1.n58 3.4105
R13957 SEL1.n80 SEL1.n79 3.4105
R13958 SEL1.n101 SEL1.n100 3.4105
R13959 SEL1.n122 SEL1.n121 3.4105
R13960 SEL1.n143 SEL1.n142 3.4105
R13961 SEL1.n164 SEL1.n163 3.4105
R13962 SEL1.n164 SEL1.n143 3.16653
R13963 SEL1.n183 SEL1.n182 3.1005
R13964 SEL1.n162 SEL1.n161 3.1005
R13965 SEL1.n141 SEL1.n140 3.1005
R13966 SEL1.n120 SEL1.n119 3.1005
R13967 SEL1.n99 SEL1.n98 3.1005
R13968 SEL1.n78 SEL1.n77 3.1005
R13969 SEL1.n57 SEL1.n56 3.1005
R13970 SEL1.n37 SEL1.n36 3.1005
R13971 SEL1.n18 SEL1.n17 3.1005
R13972 SEL1.n80 SEL1.n59 3.09637
R13973 SEL1.n122 SEL1.n101 3.09296
R13974 SEL1.n101 SEL1.n80 3.07662
R13975 SEL1.n143 SEL1.n122 3.0698
R13976 SEL1.n184 SEL1.n164 3.03575
R13977 SEL1.n171 SEL1 1.92095
R13978 SEL1.n150 SEL1 1.92095
R13979 SEL1.n129 SEL1 1.92095
R13980 SEL1.n108 SEL1 1.92095
R13981 SEL1.n87 SEL1 1.92095
R13982 SEL1.n66 SEL1 1.92095
R13983 SEL1.n45 SEL1 1.92095
R13984 SEL1.n25 SEL1 1.92095
R13985 SEL1.n6 SEL1 1.92095
R13986 SEL1.n180 SEL1.n179 1.18515
R13987 SEL1.n159 SEL1.n158 1.18515
R13988 SEL1.n138 SEL1.n137 1.18515
R13989 SEL1.n117 SEL1.n116 1.18515
R13990 SEL1.n96 SEL1.n95 1.18515
R13991 SEL1.n75 SEL1.n74 1.18515
R13992 SEL1.n54 SEL1.n53 1.18515
R13993 SEL1.n34 SEL1.n33 1.18515
R13994 SEL1.n15 SEL1.n14 1.18515
R13995 SEL1.n180 SEL1 0.397239
R13996 SEL1.n159 SEL1 0.397239
R13997 SEL1.n138 SEL1 0.397239
R13998 SEL1.n117 SEL1 0.397239
R13999 SEL1.n96 SEL1 0.397239
R14000 SEL1.n75 SEL1 0.397239
R14001 SEL1.n54 SEL1 0.397239
R14002 SEL1.n34 SEL1 0.397239
R14003 SEL1.n15 SEL1 0.397239
R14004 SEL1.n183 SEL1 0.237819
R14005 SEL1.n162 SEL1 0.237819
R14006 SEL1.n141 SEL1 0.237819
R14007 SEL1.n120 SEL1 0.237819
R14008 SEL1.n99 SEL1 0.237819
R14009 SEL1.n78 SEL1 0.237819
R14010 SEL1.n57 SEL1 0.237819
R14011 SEL1.n37 SEL1 0.237819
R14012 SEL1.n18 SEL1 0.237819
R14013 SEL1.n170 SEL1 0.0838333
R14014 SEL1.n149 SEL1 0.0838333
R14015 SEL1.n128 SEL1 0.0838333
R14016 SEL1.n142 SEL1 0.0838333
R14017 SEL1.n107 SEL1 0.0838333
R14018 SEL1.n86 SEL1 0.0838333
R14019 SEL1.n65 SEL1 0.0838333
R14020 SEL1.n44 SEL1 0.0838333
R14021 SEL1.n24 SEL1 0.0838333
R14022 SEL1.n5 SEL1 0.0838333
R14023 SEL1.n38 SEL1 0.076587
R14024 SEL1.n58 SEL1 0.0747754
R14025 SEL1.n100 SEL1 0.0657174
R14026 SEL1.n177 SEL1 0.0497424
R14027 SEL1.n156 SEL1 0.0497424
R14028 SEL1.n135 SEL1 0.0497424
R14029 SEL1.n114 SEL1 0.0497424
R14030 SEL1.n93 SEL1 0.0497424
R14031 SEL1.n72 SEL1 0.0497424
R14032 SEL1.n51 SEL1 0.0497424
R14033 SEL1.n31 SEL1 0.0497424
R14034 SEL1.n12 SEL1 0.0497424
R14035 SEL1.n163 SEL1 0.0476014
R14036 SEL1.n121 SEL1 0.0439783
R14037 SEL1.n79 SEL1 0.0439783
R14038 SEL1.n174 SEL1 0.0421667
R14039 SEL1.n153 SEL1 0.0421667
R14040 SEL1.n132 SEL1 0.0421667
R14041 SEL1.n111 SEL1 0.0421667
R14042 SEL1.n90 SEL1 0.0421667
R14043 SEL1.n69 SEL1 0.0421667
R14044 SEL1.n48 SEL1 0.0421667
R14045 SEL1.n28 SEL1 0.0421667
R14046 SEL1.n9 SEL1 0.0421667
R14047 SEL1 SEL1.n185 0.0113696
R14048 mux8_2.NAND4F_5.Y.n1 mux8_2.NAND4F_5.Y.t11 1032.02
R14049 mux8_2.NAND4F_5.Y.n1 mux8_2.NAND4F_5.Y.t10 336.962
R14050 mux8_2.NAND4F_5.Y.n1 mux8_2.NAND4F_5.Y.t9 326.154
R14051 mux8_2.NAND4F_5.Y.n0 mux8_2.NAND4F_5.Y.n3 187.373
R14052 mux8_2.NAND4F_5.Y.n0 mux8_2.NAND4F_5.Y.n4 187.192
R14053 mux8_2.NAND4F_5.Y.n0 mux8_2.NAND4F_5.Y.n5 187.192
R14054 mux8_2.NAND4F_5.Y.n7 mux8_2.NAND4F_5.Y.n6 187.192
R14055 mux8_2.NAND4F_5.Y mux8_2.NAND4F_5.Y.n1 162.94
R14056 mux8_2.NAND4F_5.Y.n2 mux8_2.NAND4F_5.Y 24.4721
R14057 mux8_2.NAND4F_5.Y.n2 mux8_2.NAND4F_5.Y.t1 22.6141
R14058 mux8_2.NAND4F_5.Y.n3 mux8_2.NAND4F_5.Y.t8 20.1899
R14059 mux8_2.NAND4F_5.Y.n3 mux8_2.NAND4F_5.Y.t7 20.1899
R14060 mux8_2.NAND4F_5.Y.n4 mux8_2.NAND4F_5.Y.t3 20.1899
R14061 mux8_2.NAND4F_5.Y.n4 mux8_2.NAND4F_5.Y.t4 20.1899
R14062 mux8_2.NAND4F_5.Y.n5 mux8_2.NAND4F_5.Y.t6 20.1899
R14063 mux8_2.NAND4F_5.Y.n5 mux8_2.NAND4F_5.Y.t5 20.1899
R14064 mux8_2.NAND4F_5.Y.n6 mux8_2.NAND4F_5.Y.t0 20.1899
R14065 mux8_2.NAND4F_5.Y.n6 mux8_2.NAND4F_5.Y.t2 20.1899
R14066 mux8_2.NAND4F_5.Y mux8_2.NAND4F_5.Y.n2 0.950576
R14067 mux8_2.NAND4F_5.Y mux8_2.NAND4F_5.Y.n7 0.396904
R14068 mux8_2.NAND4F_5.Y.n7 mux8_2.NAND4F_5.Y.n0 0.358709
R14069 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n9 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t18 540.38
R14070 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t9 491.64
R14071 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t12 491.64
R14072 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t10 491.64
R14073 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t13 491.64
R14074 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t16 367.928
R14075 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n1 227.526
R14076 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n8 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t11 227.356
R14077 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n3 227.266
R14078 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n2 227.266
R14079 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t7 213.688
R14080 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n6 162.852
R14081 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n9 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n8 160.439
R14082 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t15 139.78
R14083 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t8 139.78
R14084 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t14 139.78
R14085 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t17 139.78
R14086 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n8 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n7 94.4341
R14087 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t6 42.7831
R14088 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n5 38.6833
R14089 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t3 30.379
R14090 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t4 30.379
R14091 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t0 30.379
R14092 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t1 30.379
R14093 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t5 30.379
R14094 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t2 30.379
R14095 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n4 28.3986
R14096 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n0 18.8832
R14097 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n10 11.2587
R14098 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n10 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT 5.09176
R14099 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n10 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT 4.19292
R14100 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n9 0.794268
R14101 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t7 485.221
R14102 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t8 367.928
R14103 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n4 227.526
R14104 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n5 227.266
R14105 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n6 227.266
R14106 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t10 224.478
R14107 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t9 213.688
R14108 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n2 84.5046
R14109 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n1 72.3005
R14110 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n3 61.0566
R14111 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t0 42.7747
R14112 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t5 30.379
R14113 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t6 30.379
R14114 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t2 30.379
R14115 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t4 30.379
R14116 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t1 30.379
R14117 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.t3 30.379
R14118 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A.n0 0.583137
R14119 mux8_7.NAND4F_2.Y.n6 mux8_7.NAND4F_2.Y.t10 933.563
R14120 mux8_7.NAND4F_2.Y.n6 mux8_7.NAND4F_2.Y.t11 367.635
R14121 mux8_7.NAND4F_2.Y.n7 mux8_7.NAND4F_2.Y.t9 308.481
R14122 mux8_7.NAND4F_2.Y.n0 mux8_7.NAND4F_2.Y.n1 187.373
R14123 mux8_7.NAND4F_2.Y.n0 mux8_7.NAND4F_2.Y.n2 187.192
R14124 mux8_7.NAND4F_2.Y.n0 mux8_7.NAND4F_2.Y.n3 187.192
R14125 mux8_7.NAND4F_2.Y.n5 mux8_7.NAND4F_2.Y.n4 187.192
R14126 mux8_7.NAND4F_2.Y mux8_7.NAND4F_2.Y.n7 162.102
R14127 mux8_7.NAND4F_2.Y.n8 mux8_7.NAND4F_2.Y.t1 22.7096
R14128 mux8_7.NAND4F_2.Y.n8 mux8_7.NAND4F_2.Y 22.4285
R14129 mux8_7.NAND4F_2.Y.n1 mux8_7.NAND4F_2.Y.t7 20.1899
R14130 mux8_7.NAND4F_2.Y.n1 mux8_7.NAND4F_2.Y.t8 20.1899
R14131 mux8_7.NAND4F_2.Y.n2 mux8_7.NAND4F_2.Y.t3 20.1899
R14132 mux8_7.NAND4F_2.Y.n2 mux8_7.NAND4F_2.Y.t2 20.1899
R14133 mux8_7.NAND4F_2.Y.n3 mux8_7.NAND4F_2.Y.t5 20.1899
R14134 mux8_7.NAND4F_2.Y.n3 mux8_7.NAND4F_2.Y.t6 20.1899
R14135 mux8_7.NAND4F_2.Y.n4 mux8_7.NAND4F_2.Y.t0 20.1899
R14136 mux8_7.NAND4F_2.Y.n4 mux8_7.NAND4F_2.Y.t4 20.1899
R14137 mux8_7.NAND4F_2.Y.n7 mux8_7.NAND4F_2.Y.n6 10.955
R14138 mux8_7.NAND4F_2.Y mux8_7.NAND4F_2.Y.n8 0.799394
R14139 mux8_7.NAND4F_2.Y mux8_7.NAND4F_2.Y.n5 0.452586
R14140 mux8_7.NAND4F_2.Y.n5 mux8_7.NAND4F_2.Y.n0 0.358709
R14141 mux8_7.NAND4F_8.Y.n1 mux8_7.NAND4F_8.Y.t10 379.173
R14142 mux8_7.NAND4F_8.Y.n2 mux8_7.NAND4F_8.Y.t14 312.599
R14143 mux8_7.NAND4F_8.Y.n1 mux8_7.NAND4F_8.Y.t9 247.428
R14144 mux8_7.NAND4F_8.Y.n4 mux8_7.NAND4F_8.Y.t11 247.428
R14145 mux8_7.NAND4F_8.Y.n3 mux8_7.NAND4F_8.Y.t13 247.428
R14146 mux8_7.NAND4F_8.Y.n2 mux8_7.NAND4F_8.Y.t12 247.428
R14147 mux8_7.NAND4F_8.Y.n0 mux8_7.NAND4F_8.Y.n6 187.373
R14148 mux8_7.NAND4F_8.Y.n0 mux8_7.NAND4F_8.Y.n7 187.192
R14149 mux8_7.NAND4F_8.Y.n0 mux8_7.NAND4F_8.Y.n8 187.192
R14150 mux8_7.NAND4F_8.Y.n10 mux8_7.NAND4F_8.Y.n9 187.192
R14151 mux8_7.NAND4F_8.Y mux8_7.NAND4F_8.Y.n5 162.139
R14152 mux8_7.NAND4F_8.Y.n4 mux8_7.NAND4F_8.Y.n3 65.1723
R14153 mux8_7.NAND4F_8.Y.n3 mux8_7.NAND4F_8.Y.n2 65.1723
R14154 mux8_7.NAND4F_8.Y.n5 mux8_7.NAND4F_8.Y.n4 33.2653
R14155 mux8_7.NAND4F_8.Y.n5 mux8_7.NAND4F_8.Y.n1 31.9075
R14156 mux8_7.NAND4F_8.Y mux8_7.NAND4F_8.Y.t2 22.6141
R14157 mux8_7.NAND4F_8.Y.n6 mux8_7.NAND4F_8.Y.t4 20.1899
R14158 mux8_7.NAND4F_8.Y.n6 mux8_7.NAND4F_8.Y.t3 20.1899
R14159 mux8_7.NAND4F_8.Y.n7 mux8_7.NAND4F_8.Y.t5 20.1899
R14160 mux8_7.NAND4F_8.Y.n7 mux8_7.NAND4F_8.Y.t6 20.1899
R14161 mux8_7.NAND4F_8.Y.n8 mux8_7.NAND4F_8.Y.t7 20.1899
R14162 mux8_7.NAND4F_8.Y.n8 mux8_7.NAND4F_8.Y.t8 20.1899
R14163 mux8_7.NAND4F_8.Y.n9 mux8_7.NAND4F_8.Y.t0 20.1899
R14164 mux8_7.NAND4F_8.Y.n9 mux8_7.NAND4F_8.Y.t1 20.1899
R14165 mux8_7.NAND4F_8.Y mux8_7.NAND4F_8.Y.n10 0.452586
R14166 mux8_7.NAND4F_8.Y.n10 mux8_7.NAND4F_8.Y.n0 0.358709
R14167 mux8_5.NAND4F_6.Y.n1 mux8_5.NAND4F_6.Y.t10 933.563
R14168 mux8_5.NAND4F_6.Y.n1 mux8_5.NAND4F_6.Y.t11 367.635
R14169 mux8_5.NAND4F_6.Y.n2 mux8_5.NAND4F_6.Y.t9 308.481
R14170 mux8_5.NAND4F_6.Y.n0 mux8_5.NAND4F_6.Y.n4 187.373
R14171 mux8_5.NAND4F_6.Y.n0 mux8_5.NAND4F_6.Y.n5 187.192
R14172 mux8_5.NAND4F_6.Y.n0 mux8_5.NAND4F_6.Y.n6 187.192
R14173 mux8_5.NAND4F_6.Y.n8 mux8_5.NAND4F_6.Y.n7 187.192
R14174 mux8_5.NAND4F_6.Y mux8_5.NAND4F_6.Y.n2 162.047
R14175 mux8_5.NAND4F_6.Y.n3 mux8_5.NAND4F_6.Y.t0 22.7831
R14176 mux8_5.NAND4F_6.Y.n3 mux8_5.NAND4F_6.Y 22.171
R14177 mux8_5.NAND4F_6.Y.n4 mux8_5.NAND4F_6.Y.t7 20.1899
R14178 mux8_5.NAND4F_6.Y.n4 mux8_5.NAND4F_6.Y.t8 20.1899
R14179 mux8_5.NAND4F_6.Y.n5 mux8_5.NAND4F_6.Y.t4 20.1899
R14180 mux8_5.NAND4F_6.Y.n5 mux8_5.NAND4F_6.Y.t3 20.1899
R14181 mux8_5.NAND4F_6.Y.n6 mux8_5.NAND4F_6.Y.t6 20.1899
R14182 mux8_5.NAND4F_6.Y.n6 mux8_5.NAND4F_6.Y.t5 20.1899
R14183 mux8_5.NAND4F_6.Y.n7 mux8_5.NAND4F_6.Y.t1 20.1899
R14184 mux8_5.NAND4F_6.Y.n7 mux8_5.NAND4F_6.Y.t2 20.1899
R14185 mux8_5.NAND4F_6.Y.n2 mux8_5.NAND4F_6.Y.n1 10.955
R14186 mux8_5.NAND4F_6.Y mux8_5.NAND4F_6.Y.n3 0.781576
R14187 mux8_5.NAND4F_6.Y mux8_5.NAND4F_6.Y.n8 0.396904
R14188 mux8_5.NAND4F_6.Y.n8 mux8_5.NAND4F_6.Y.n0 0.358709
R14189 a_n4385_3190.n2 a_n4385_3190.t7 541.395
R14190 a_n4385_3190.n3 a_n4385_3190.t3 527.402
R14191 a_n4385_3190.n2 a_n4385_3190.t6 491.64
R14192 a_n4385_3190.n5 a_n4385_3190.t1 281.906
R14193 a_n4385_3190.t0 a_n4385_3190.n5 204.359
R14194 a_n4385_3190.n0 a_n4385_3190.t2 180.73
R14195 a_n4385_3190.n1 a_n4385_3190.t5 179.45
R14196 a_n4385_3190.n0 a_n4385_3190.t4 139.78
R14197 a_n4385_3190.n4 a_n4385_3190.n1 105.635
R14198 a_n4385_3190.n4 a_n4385_3190.n3 76.0005
R14199 a_n4385_3190.n5 a_n4385_3190.n4 67.9685
R14200 a_n4385_3190.n3 a_n4385_3190.n2 13.994
R14201 a_n4385_3190.n1 a_n4385_3190.n0 1.28015
R14202 a_n3629_3190.n2 a_n3629_3190.n0 121.353
R14203 a_n3629_3190.n3 a_n3629_3190.n2 121.001
R14204 a_n3629_3190.n2 a_n3629_3190.n1 120.977
R14205 a_n3629_3190.n1 a_n3629_3190.t3 30.462
R14206 a_n3629_3190.n1 a_n3629_3190.t5 30.462
R14207 a_n3629_3190.n0 a_n3629_3190.t0 30.462
R14208 a_n3629_3190.n0 a_n3629_3190.t1 30.462
R14209 a_n3629_3190.t2 a_n3629_3190.n3 30.462
R14210 a_n3629_3190.n3 a_n3629_3190.t4 30.462
R14211 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n9 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t8 540.38
R14212 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t7 491.64
R14213 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t13 491.64
R14214 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t17 491.64
R14215 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t15 491.64
R14216 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n7 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t10 367.928
R14217 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n1 227.526
R14218 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n8 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t11 227.356
R14219 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n3 227.266
R14220 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n2 227.266
R14221 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n7 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t12 213.688
R14222 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n6 162.852
R14223 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n9 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n8 160.439
R14224 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t14 139.78
R14225 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t9 139.78
R14226 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t16 139.78
R14227 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t18 139.78
R14228 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n8 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n7 94.4341
R14229 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t4 42.7831
R14230 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n6 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n5 38.6833
R14231 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n3 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t6 30.379
R14232 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n3 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t5 30.379
R14233 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n1 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t0 30.379
R14234 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n1 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t2 30.379
R14235 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n2 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t3 30.379
R14236 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n2 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t1 30.379
R14237 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n6 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n4 28.3986
R14238 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n0 18.8832
R14239 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n10 11.2587
R14240 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n10 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 5.09176
R14241 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n10 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 4.19292
R14242 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n9 0.794268
R14243 a_n13192_2026.n0 a_n13192_2026.n2 81.2978
R14244 a_n13192_2026.n0 a_n13192_2026.n3 81.1637
R14245 a_n13192_2026.n0 a_n13192_2026.n4 81.1637
R14246 a_n13192_2026.n1 a_n13192_2026.n5 81.1637
R14247 a_n13192_2026.n1 a_n13192_2026.n6 81.1637
R14248 a_n13192_2026.n7 a_n13192_2026.n1 80.9213
R14249 a_n13192_2026.n2 a_n13192_2026.t0 11.8205
R14250 a_n13192_2026.n2 a_n13192_2026.t2 11.8205
R14251 a_n13192_2026.n3 a_n13192_2026.t11 11.8205
R14252 a_n13192_2026.n3 a_n13192_2026.t1 11.8205
R14253 a_n13192_2026.n4 a_n13192_2026.t6 11.8205
R14254 a_n13192_2026.n4 a_n13192_2026.t10 11.8205
R14255 a_n13192_2026.n5 a_n13192_2026.t5 11.8205
R14256 a_n13192_2026.n5 a_n13192_2026.t4 11.8205
R14257 a_n13192_2026.n6 a_n13192_2026.t8 11.8205
R14258 a_n13192_2026.n6 a_n13192_2026.t3 11.8205
R14259 a_n13192_2026.t9 a_n13192_2026.n7 11.8205
R14260 a_n13192_2026.n7 a_n13192_2026.t7 11.8205
R14261 a_n13192_2026.n1 a_n13192_2026.n0 0.402735
R14262 A1.n13 A1.t9 540.38
R14263 A1.n19 A1.t6 540.38
R14264 A1.n16 A1.t32 540.38
R14265 A1.n10 A1.t2 540.38
R14266 A1.n2 A1.t13 540.38
R14267 A1.n26 A1.t27 540.375
R14268 A1.n3 A1.t10 491.64
R14269 A1.n3 A1.t39 491.64
R14270 A1.n3 A1.t34 491.64
R14271 A1.n3 A1.t31 491.64
R14272 A1.n36 A1.t7 491.64
R14273 A1.n36 A1.t5 491.64
R14274 A1.n36 A1.t38 491.64
R14275 A1.n36 A1.t23 491.64
R14276 A1.n11 A1.t28 367.928
R14277 A1.n17 A1.t33 367.928
R14278 A1.n14 A1.t0 367.928
R14279 A1.n8 A1.t20 367.928
R14280 A1.n0 A1.t18 367.928
R14281 A1.n24 A1.t44 343.827
R14282 A1.n29 A1.t35 312.599
R14283 A1.n32 A1.t25 247.428
R14284 A1.n31 A1.t11 247.428
R14285 A1.n30 A1.t8 247.428
R14286 A1.n29 A1.t40 247.428
R14287 A1.n24 A1.t1 237.787
R14288 A1.n33 A1.t24 229.754
R14289 A1.n25 A1.t19 227.356
R14290 A1.n12 A1.t41 227.356
R14291 A1.n18 A1.t3 227.356
R14292 A1.n15 A1.t45 227.356
R14293 A1.n9 A1.t36 227.356
R14294 A1.n1 A1.t15 227.356
R14295 A1.n11 A1.t42 213.688
R14296 A1.n17 A1.t4 213.688
R14297 A1.n14 A1.t29 213.688
R14298 A1.n8 A1.t21 213.688
R14299 A1.n0 A1.t16 213.688
R14300 A1 A1.n37 163.036
R14301 A1.n6 A1.n5 162.867
R14302 A1 A1.n33 162.409
R14303 A1.n13 A1.n12 160.439
R14304 A1.n19 A1.n18 160.439
R14305 A1.n16 A1.n15 160.439
R14306 A1.n10 A1.n9 160.439
R14307 A1.n2 A1.n1 160.439
R14308 A1.n26 A1.n25 160.433
R14309 A1.n4 A1.t17 139.78
R14310 A1.n4 A1.t12 139.78
R14311 A1.n4 A1.t37 139.78
R14312 A1.n4 A1.t22 139.78
R14313 A1.n35 A1.t14 139.78
R14314 A1.n35 A1.t43 139.78
R14315 A1.n35 A1.t30 139.78
R14316 A1.n35 A1.t26 139.78
R14317 A1.n12 A1.n11 94.4341
R14318 A1.n18 A1.n17 94.4341
R14319 A1.n15 A1.n14 94.4341
R14320 A1.n9 A1.n8 94.4341
R14321 A1.n1 A1.n0 94.4341
R14322 A1.n33 A1.n32 91.5805
R14323 A1.n25 A1.n24 70.3341
R14324 A1.n30 A1.n29 65.1723
R14325 A1.n31 A1.n30 65.1723
R14326 A1.n32 A1.n31 65.1723
R14327 A1.n37 A1.n35 38.8368
R14328 A1.n5 A1.n4 38.6833
R14329 A1.n23 A1 30.3458
R14330 A1.n5 A1.n3 28.3986
R14331 A1.n37 A1.n36 28.2451
R14332 A1 A1.n7 18.1883
R14333 A1.n38 A1.n34 15.973
R14334 A1.n34 A1 12.5318
R14335 A1.n28 A1.n27 12.4105
R14336 A1.n7 A1.n6 9.00496
R14337 A1 A1.n23 5.72922
R14338 A1.n23 A1.n22 4.83222
R14339 A1.n7 A1 3.87912
R14340 A1.n34 A1.n28 3.66175
R14341 A1.n20 A1 3.24541
R14342 A1.n21 A1 2.59446
R14343 A1.n20 A1 2.44812
R14344 A1.n38 A1 1.92708
R14345 A1.n22 A1.n21 1.7055
R14346 A1.n27 A1 1.36134
R14347 A1 A1.n26 0.905186
R14348 A1 A1.n13 0.900886
R14349 A1 A1.n19 0.900886
R14350 A1 A1.n16 0.900886
R14351 A1 A1.n10 0.900886
R14352 A1 A1.n2 0.89693
R14353 A1.n21 A1.n20 0.651689
R14354 A1.n22 A1 0.374163
R14355 A1.n27 A1 0.0594888
R14356 A1.n6 A1 0.0590664
R14357 A1 A1.n38 0.0186554
R14358 A1.n28 A1 0.012118
R14359 MULT_0.NAND2_9.Y.n5 MULT_0.NAND2_9.Y.t8 291.829
R14360 MULT_0.NAND2_9.Y.n5 MULT_0.NAND2_9.Y.t10 291.829
R14361 MULT_0.NAND2_9.Y.n0 MULT_0.NAND2_9.Y.n2 227.526
R14362 MULT_0.NAND2_9.Y.n0 MULT_0.NAND2_9.Y.n3 227.266
R14363 MULT_0.NAND2_9.Y.n0 MULT_0.NAND2_9.Y.n4 227.266
R14364 MULT_0.NAND2_9.Y.n5 MULT_0.NAND2_9.Y.t9 221.72
R14365 MULT_0.NAND2_9.Y.t7 MULT_0.NAND2_9.Y.n1 393.897
R14366 MULT_0.NAND2_9.Y.n0 MULT_0.NAND2_9.Y.t0 42.7333
R14367 MULT_0.NAND2_9.Y.n2 MULT_0.NAND2_9.Y.t6 30.379
R14368 MULT_0.NAND2_9.Y.n2 MULT_0.NAND2_9.Y.t5 30.379
R14369 MULT_0.NAND2_9.Y.n3 MULT_0.NAND2_9.Y.t1 30.379
R14370 MULT_0.NAND2_9.Y.n3 MULT_0.NAND2_9.Y.t4 30.379
R14371 MULT_0.NAND2_9.Y.n4 MULT_0.NAND2_9.Y.t3 30.379
R14372 MULT_0.NAND2_9.Y.n4 MULT_0.NAND2_9.Y.t2 30.379
R14373 MULT_0.NAND2_9.Y.n5 MULT_0.NAND2_9.Y.n1 53.4911
R14374 MULT_0.NAND2_9.Y.n0 MULT_0.NAND2_9.Y.n1 0.620447
R14375 mux8_3.NAND4F_8.Y.n1 mux8_3.NAND4F_8.Y.t9 379.173
R14376 mux8_3.NAND4F_8.Y.n2 mux8_3.NAND4F_8.Y.t13 312.599
R14377 mux8_3.NAND4F_8.Y.n1 mux8_3.NAND4F_8.Y.t14 247.428
R14378 mux8_3.NAND4F_8.Y.n4 mux8_3.NAND4F_8.Y.t10 247.428
R14379 mux8_3.NAND4F_8.Y.n3 mux8_3.NAND4F_8.Y.t12 247.428
R14380 mux8_3.NAND4F_8.Y.n2 mux8_3.NAND4F_8.Y.t11 247.428
R14381 mux8_3.NAND4F_8.Y.n0 mux8_3.NAND4F_8.Y.n6 187.373
R14382 mux8_3.NAND4F_8.Y.n0 mux8_3.NAND4F_8.Y.n7 187.192
R14383 mux8_3.NAND4F_8.Y.n0 mux8_3.NAND4F_8.Y.n8 187.192
R14384 mux8_3.NAND4F_8.Y.n10 mux8_3.NAND4F_8.Y.n9 187.192
R14385 mux8_3.NAND4F_8.Y mux8_3.NAND4F_8.Y.n5 162.139
R14386 mux8_3.NAND4F_8.Y.n4 mux8_3.NAND4F_8.Y.n3 65.1723
R14387 mux8_3.NAND4F_8.Y.n3 mux8_3.NAND4F_8.Y.n2 65.1723
R14388 mux8_3.NAND4F_8.Y.n5 mux8_3.NAND4F_8.Y.n4 33.2653
R14389 mux8_3.NAND4F_8.Y.n5 mux8_3.NAND4F_8.Y.n1 31.9075
R14390 mux8_3.NAND4F_8.Y mux8_3.NAND4F_8.Y.t5 22.6141
R14391 mux8_3.NAND4F_8.Y.n6 mux8_3.NAND4F_8.Y.t3 20.1899
R14392 mux8_3.NAND4F_8.Y.n6 mux8_3.NAND4F_8.Y.t2 20.1899
R14393 mux8_3.NAND4F_8.Y.n7 mux8_3.NAND4F_8.Y.t0 20.1899
R14394 mux8_3.NAND4F_8.Y.n7 mux8_3.NAND4F_8.Y.t1 20.1899
R14395 mux8_3.NAND4F_8.Y.n8 mux8_3.NAND4F_8.Y.t7 20.1899
R14396 mux8_3.NAND4F_8.Y.n8 mux8_3.NAND4F_8.Y.t8 20.1899
R14397 mux8_3.NAND4F_8.Y.n9 mux8_3.NAND4F_8.Y.t6 20.1899
R14398 mux8_3.NAND4F_8.Y.n9 mux8_3.NAND4F_8.Y.t4 20.1899
R14399 mux8_3.NAND4F_8.Y mux8_3.NAND4F_8.Y.n10 0.452586
R14400 mux8_3.NAND4F_8.Y.n10 mux8_3.NAND4F_8.Y.n0 0.358709
R14401 mux8_3.inv_0.A.n1 mux8_3.inv_0.A.t7 291.829
R14402 mux8_3.inv_0.A.n1 mux8_3.inv_0.A.t9 291.829
R14403 mux8_3.inv_0.A.n0 mux8_3.inv_0.A.t1 256.425
R14404 mux8_3.inv_0.A.n0 mux8_3.inv_0.A.n2 231.24
R14405 mux8_3.inv_0.A.n0 mux8_3.inv_0.A.n3 231.03
R14406 mux8_3.inv_0.A.n1 mux8_3.inv_0.A.t8 221.72
R14407 mux8_3.inv_0.A.t10 mux8_3.inv_0.A.n0 393.959
R14408 mux8_3.inv_0.A.n4 mux8_3.inv_0.A.n0 66.6316
R14409 mux8_3.inv_0.A.n0 mux8_3.inv_0.A.n1 54.1444
R14410 mux8_3.inv_0.A.n2 mux8_3.inv_0.A.t4 25.395
R14411 mux8_3.inv_0.A.n2 mux8_3.inv_0.A.t5 25.395
R14412 mux8_3.inv_0.A.n3 mux8_3.inv_0.A.t2 25.395
R14413 mux8_3.inv_0.A.n3 mux8_3.inv_0.A.t3 25.395
R14414 mux8_3.inv_0.A.n4 mux8_3.inv_0.A.t6 19.8005
R14415 mux8_3.inv_0.A.n4 mux8_3.inv_0.A.t0 19.8005
R14416 a_n18222_1406.n0 a_n18222_1406.t6 539.788
R14417 a_n18222_1406.n1 a_n18222_1406.t2 531.496
R14418 a_n18222_1406.n0 a_n18222_1406.t3 490.034
R14419 a_n18222_1406.n5 a_n18222_1406.t0 283.788
R14420 a_n18222_1406.t1 a_n18222_1406.n5 205.489
R14421 a_n18222_1406.n2 a_n18222_1406.t4 182.625
R14422 a_n18222_1406.n3 a_n18222_1406.t5 179.054
R14423 a_n18222_1406.n2 a_n18222_1406.t7 139.78
R14424 a_n18222_1406.n4 a_n18222_1406.n3 101.368
R14425 a_n18222_1406.n5 a_n18222_1406.n4 77.9135
R14426 a_n18222_1406.n4 a_n18222_1406.n1 76.1557
R14427 a_n18222_1406.n1 a_n18222_1406.n0 8.29297
R14428 a_n18222_1406.n3 a_n18222_1406.n2 3.57087
R14429 a_n18042_2026.n6 a_n18042_2026.n0 81.3236
R14430 a_n18042_2026.n0 a_n18042_2026.n1 81.2978
R14431 a_n18042_2026.n0 a_n18042_2026.n2 81.1637
R14432 a_n18042_2026.n0 a_n18042_2026.n3 81.1637
R14433 a_n18042_2026.n0 a_n18042_2026.n4 81.1637
R14434 a_n18042_2026.n0 a_n18042_2026.n5 81.1637
R14435 a_n18042_2026.n1 a_n18042_2026.t9 11.8205
R14436 a_n18042_2026.n1 a_n18042_2026.t10 11.8205
R14437 a_n18042_2026.n2 a_n18042_2026.t5 11.8205
R14438 a_n18042_2026.n2 a_n18042_2026.t11 11.8205
R14439 a_n18042_2026.n3 a_n18042_2026.t3 11.8205
R14440 a_n18042_2026.n3 a_n18042_2026.t4 11.8205
R14441 a_n18042_2026.n4 a_n18042_2026.t6 11.8205
R14442 a_n18042_2026.n4 a_n18042_2026.t8 11.8205
R14443 a_n18042_2026.n5 a_n18042_2026.t2 11.8205
R14444 a_n18042_2026.n5 a_n18042_2026.t7 11.8205
R14445 a_n18042_2026.n6 a_n18042_2026.t1 11.8205
R14446 a_n18042_2026.t0 a_n18042_2026.n6 11.8205
R14447 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t17 491.64
R14448 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t14 491.64
R14449 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t23 491.64
R14450 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t15 491.64
R14451 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t19 485.221
R14452 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t20 367.928
R14453 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t13 255.588
R14454 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t21 224.478
R14455 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t22 213.688
R14456 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n0 209.19
R14457 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t16 139.78
R14458 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t18 139.78
R14459 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t12 139.78
R14460 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n10 120.999
R14461 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n9 120.999
R14462 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n22 104.489
R14463 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n12 92.5005
R14464 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n18 86.2638
R14465 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n17 85.8873
R14466 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n15 85.724
R14467 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n7 84.5046
R14468 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n23 83.8907
R14469 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n17 75.0672
R14470 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n20 75.0672
R14471 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n15 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n14 73.1255
R14472 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n17 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n16 73.1255
R14473 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n19 73.1255
R14474 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n6 72.3005
R14475 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n15 68.8946
R14476 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n8 60.9797
R14477 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n13 41.9827
R14478 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t9 30.462
R14479 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t1 30.462
R14480 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t5 30.462
R14481 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t0 30.462
R14482 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t11 30.462
R14483 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t10 30.462
R14484 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n11 28.124
R14485 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n5 19.963
R14486 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n1 17.8661
R14487 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n2 17.8661
R14488 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n3 17.1217
R14489 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t7 11.8205
R14490 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t6 11.8205
R14491 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t8 11.8205
R14492 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t2 11.8205
R14493 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t3 11.8205
R14494 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t4 11.8205
R14495 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n21 9.3005
R14496 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n4 1.8615
R14497 a_n24654_1380.n2 a_n24654_1380.t4 541.395
R14498 a_n24654_1380.n3 a_n24654_1380.t6 527.402
R14499 a_n24654_1380.n2 a_n24654_1380.t5 491.64
R14500 a_n24654_1380.n5 a_n24654_1380.t0 281.906
R14501 a_n24654_1380.t1 a_n24654_1380.n5 204.359
R14502 a_n24654_1380.n0 a_n24654_1380.t7 180.73
R14503 a_n24654_1380.n1 a_n24654_1380.t2 179.45
R14504 a_n24654_1380.n0 a_n24654_1380.t3 139.78
R14505 a_n24654_1380.n4 a_n24654_1380.n1 105.635
R14506 a_n24654_1380.n4 a_n24654_1380.n3 76.0005
R14507 a_n24654_1380.n5 a_n24654_1380.n4 67.9685
R14508 a_n24654_1380.n3 a_n24654_1380.n2 13.994
R14509 a_n24654_1380.n1 a_n24654_1380.n0 1.28015
R14510 a_n24624_1406.n3 a_n24624_1406.n2 121.353
R14511 a_n24624_1406.n2 a_n24624_1406.n1 121.001
R14512 a_n24624_1406.n2 a_n24624_1406.n0 120.977
R14513 a_n24624_1406.n1 a_n24624_1406.t5 30.462
R14514 a_n24624_1406.n1 a_n24624_1406.t1 30.462
R14515 a_n24624_1406.n0 a_n24624_1406.t4 30.462
R14516 a_n24624_1406.n0 a_n24624_1406.t0 30.462
R14517 a_n24624_1406.n3 a_n24624_1406.t2 30.462
R14518 a_n24624_1406.t3 a_n24624_1406.n3 30.462
R14519 a_n14155_n8419.n0 a_n14155_n8419.t6 539.788
R14520 a_n14155_n8419.n1 a_n14155_n8419.t3 531.496
R14521 a_n14155_n8419.n0 a_n14155_n8419.t2 490.034
R14522 a_n14155_n8419.n5 a_n14155_n8419.t0 283.788
R14523 a_n14155_n8419.t1 a_n14155_n8419.n5 205.489
R14524 a_n14155_n8419.n2 a_n14155_n8419.t4 182.625
R14525 a_n14155_n8419.n3 a_n14155_n8419.t7 179.054
R14526 a_n14155_n8419.n2 a_n14155_n8419.t5 139.78
R14527 a_n14155_n8419.n4 a_n14155_n8419.n3 101.368
R14528 a_n14155_n8419.n5 a_n14155_n8419.n4 77.9135
R14529 a_n14155_n8419.n4 a_n14155_n8419.n1 76.1557
R14530 a_n14155_n8419.n1 a_n14155_n8419.n0 8.29297
R14531 a_n14155_n8419.n3 a_n14155_n8419.n2 3.57087
R14532 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t21 491.64
R14533 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t12 491.64
R14534 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t13 491.64
R14535 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t22 491.64
R14536 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n8 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t15 485.221
R14537 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t18 367.928
R14538 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t16 255.588
R14539 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t23 224.478
R14540 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t19 213.688
R14541 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n0 209.19
R14542 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t17 139.78
R14543 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t14 139.78
R14544 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t20 139.78
R14545 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n11 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n10 120.999
R14546 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n11 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n9 120.999
R14547 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n23 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n22 104.489
R14548 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n13 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n12 92.5005
R14549 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n20 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n18 86.2638
R14550 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n18 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n17 85.8873
R14551 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n18 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n15 85.724
R14552 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n8 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n7 84.5046
R14553 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n23 83.8907
R14554 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n21 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n20 75.0672
R14555 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n21 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n17 75.0672
R14556 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n20 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n19 73.1255
R14557 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n17 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n16 73.1255
R14558 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n15 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n14 73.1255
R14559 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n6 72.3005
R14560 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n22 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n15 68.8946
R14561 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n8 60.9797
R14562 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n23 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n13 41.9827
R14563 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n12 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t6 30.462
R14564 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n12 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t0 30.462
R14565 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n10 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t1 30.462
R14566 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n10 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t2 30.462
R14567 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n9 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t7 30.462
R14568 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n9 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t8 30.462
R14569 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n13 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n11 28.124
R14570 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n5 19.963
R14571 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n1 17.8661
R14572 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n2 17.8661
R14573 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n3 17.1217
R14574 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n16 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t9 11.8205
R14575 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n16 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t10 11.8205
R14576 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n19 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t5 11.8205
R14577 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n19 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t4 11.8205
R14578 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n14 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t11 11.8205
R14579 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n14 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t3 11.8205
R14580 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n22 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n21 9.3005
R14581 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n4 1.8615
R14582 a_n13975_n7799.n1 a_n13975_n7799.n5 81.2978
R14583 a_n13975_n7799.n1 a_n13975_n7799.n6 81.1637
R14584 a_n13975_n7799.n0 a_n13975_n7799.n4 81.1637
R14585 a_n13975_n7799.n0 a_n13975_n7799.n3 81.1637
R14586 a_n13975_n7799.n7 a_n13975_n7799.n1 81.1637
R14587 a_n13975_n7799.n0 a_n13975_n7799.n2 80.9213
R14588 a_n13975_n7799.n5 a_n13975_n7799.t8 11.8205
R14589 a_n13975_n7799.n5 a_n13975_n7799.t7 11.8205
R14590 a_n13975_n7799.n6 a_n13975_n7799.t4 11.8205
R14591 a_n13975_n7799.n6 a_n13975_n7799.t6 11.8205
R14592 a_n13975_n7799.n4 a_n13975_n7799.t10 11.8205
R14593 a_n13975_n7799.n4 a_n13975_n7799.t11 11.8205
R14594 a_n13975_n7799.n3 a_n13975_n7799.t2 11.8205
R14595 a_n13975_n7799.n3 a_n13975_n7799.t9 11.8205
R14596 a_n13975_n7799.n2 a_n13975_n7799.t1 11.8205
R14597 a_n13975_n7799.n2 a_n13975_n7799.t0 11.8205
R14598 a_n13975_n7799.n7 a_n13975_n7799.t3 11.8205
R14599 a_n13975_n7799.t5 a_n13975_n7799.n7 11.8205
R14600 a_n13975_n7799.n1 a_n13975_n7799.n0 0.402735
R14601 a_n12347_n15041.n2 a_n12347_n15041.t3 539.788
R14602 a_n12347_n15041.n3 a_n12347_n15041.t7 531.496
R14603 a_n12347_n15041.n2 a_n12347_n15041.t5 490.034
R14604 a_n12347_n15041.n5 a_n12347_n15041.t1 283.788
R14605 a_n12347_n15041.t0 a_n12347_n15041.n5 205.489
R14606 a_n12347_n15041.n0 a_n12347_n15041.t6 182.625
R14607 a_n12347_n15041.n1 a_n12347_n15041.t4 179.054
R14608 a_n12347_n15041.n0 a_n12347_n15041.t2 139.78
R14609 a_n12347_n15041.n4 a_n12347_n15041.n1 101.368
R14610 a_n12347_n15041.n5 a_n12347_n15041.n4 77.9135
R14611 a_n12347_n15041.n4 a_n12347_n15041.n3 76.1557
R14612 a_n12347_n15041.n3 a_n12347_n15041.n2 8.29297
R14613 a_n12347_n15041.n1 a_n12347_n15041.n0 3.57087
R14614 XOR8_0.S0.n0 XOR8_0.S0.t14 1032.02
R14615 XOR8_0.S0.n0 XOR8_0.S0.t13 336.962
R14616 XOR8_0.S0.n0 XOR8_0.S0.t12 326.154
R14617 XOR8_0.S0 XOR8_0.S0.n0 162.946
R14618 XOR8_0.S0.n3 XOR8_0.S0.n1 120.999
R14619 XOR8_0.S0.n3 XOR8_0.S0.n2 120.999
R14620 XOR8_0.S0.n15 XOR8_0.S0.n14 104.865
R14621 XOR8_0.S0.n5 XOR8_0.S0.n4 92.5005
R14622 XOR8_0.S0.n12 XOR8_0.S0.n10 86.2638
R14623 XOR8_0.S0.n10 XOR8_0.S0.n9 85.8873
R14624 XOR8_0.S0.n10 XOR8_0.S0.n7 85.724
R14625 XOR8_0.S0 XOR8_0.S0.n15 83.8907
R14626 XOR8_0.S0.n13 XOR8_0.S0.n9 75.0672
R14627 XOR8_0.S0.n13 XOR8_0.S0.n12 75.0672
R14628 XOR8_0.S0.n9 XOR8_0.S0.n8 73.1255
R14629 XOR8_0.S0.n12 XOR8_0.S0.n11 73.1255
R14630 XOR8_0.S0.n7 XOR8_0.S0.n6 73.1255
R14631 XOR8_0.S0.n14 XOR8_0.S0.n7 68.5181
R14632 XOR8_0.S0.n15 XOR8_0.S0.n5 41.9827
R14633 XOR8_0.S0.n4 XOR8_0.S0.t2 30.462
R14634 XOR8_0.S0.n4 XOR8_0.S0.t10 30.462
R14635 XOR8_0.S0.n1 XOR8_0.S0.t0 30.462
R14636 XOR8_0.S0.n1 XOR8_0.S0.t1 30.462
R14637 XOR8_0.S0.n2 XOR8_0.S0.t11 30.462
R14638 XOR8_0.S0.n2 XOR8_0.S0.t9 30.462
R14639 XOR8_0.S0.n5 XOR8_0.S0.n3 28.124
R14640 XOR8_0.S0.n11 XOR8_0.S0.t7 11.8205
R14641 XOR8_0.S0.n11 XOR8_0.S0.t6 11.8205
R14642 XOR8_0.S0.n8 XOR8_0.S0.t4 11.8205
R14643 XOR8_0.S0.n8 XOR8_0.S0.t5 11.8205
R14644 XOR8_0.S0.n6 XOR8_0.S0.t3 11.8205
R14645 XOR8_0.S0.n6 XOR8_0.S0.t8 11.8205
R14646 XOR8_0.S0.n14 XOR8_0.S0.n13 9.3005
R14647 a_n11276_n15299.n2 a_n11276_n15299.n1 121.353
R14648 a_n11276_n15299.n3 a_n11276_n15299.n2 121.001
R14649 a_n11276_n15299.n2 a_n11276_n15299.n0 120.977
R14650 a_n11276_n15299.n0 a_n11276_n15299.t3 30.462
R14651 a_n11276_n15299.n0 a_n11276_n15299.t5 30.462
R14652 a_n11276_n15299.n1 a_n11276_n15299.t1 30.462
R14653 a_n11276_n15299.n1 a_n11276_n15299.t2 30.462
R14654 a_n11276_n15299.t4 a_n11276_n15299.n3 30.462
R14655 a_n11276_n15299.n3 a_n11276_n15299.t0 30.462
R14656 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t7 540.38
R14657 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t8 367.928
R14658 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n4 227.526
R14659 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t10 227.356
R14660 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n6 227.266
R14661 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n5 227.266
R14662 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t9 213.688
R14663 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n2 160.439
R14664 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n1 94.4341
R14665 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t3 42.7943
R14666 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t0 30.379
R14667 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t1 30.379
R14668 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t5 30.379
R14669 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t6 30.379
R14670 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t2 30.379
R14671 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.t4 30.379
R14672 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n0 13.4358
R14673 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B.n3 0.821842
R14674 a_n11723_n9452.t0 a_n11723_n9452.t1 19.8005
R14675 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n9 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t9 540.38
R14676 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t12 491.64
R14677 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t18 491.64
R14678 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t16 491.64
R14679 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t8 491.64
R14680 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t11 367.928
R14681 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n1 227.526
R14682 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n8 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t17 227.356
R14683 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n2 227.266
R14684 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n3 227.266
R14685 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n7 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t14 213.688
R14686 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n6 162.852
R14687 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n9 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n8 160.439
R14688 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t10 139.78
R14689 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t15 139.78
R14690 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t7 139.78
R14691 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t13 139.78
R14692 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n8 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n7 94.4341
R14693 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t0 42.7831
R14694 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n5 38.6833
R14695 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t5 30.379
R14696 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t4 30.379
R14697 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t1 30.379
R14698 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t6 30.379
R14699 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t3 30.379
R14700 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t2 30.379
R14701 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n4 28.3986
R14702 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n0 18.8832
R14703 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n10 10.7052
R14704 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n10 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT 5.09176
R14705 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n10 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT 4.19292
R14706 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n9 0.794268
R14707 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t14 491.64
R14708 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t12 491.64
R14709 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t13 491.64
R14710 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t20 491.64
R14711 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t16 485.221
R14712 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t19 367.928
R14713 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t17 255.588
R14714 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n7 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t15 224.478
R14715 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t18 213.688
R14716 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n0 209.19
R14717 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t22 139.78
R14718 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t23 139.78
R14719 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t21 139.78
R14720 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n11 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n10 120.999
R14721 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n11 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n9 120.999
R14722 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n23 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n22 104.489
R14723 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n13 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n12 92.5005
R14724 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n20 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n18 86.2638
R14725 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n18 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n17 85.8873
R14726 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n18 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n15 85.724
R14727 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n7 84.5046
R14728 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n23 83.8907
R14729 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n21 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n20 75.0672
R14730 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n21 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n17 75.0672
R14731 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n20 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n19 73.1255
R14732 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n17 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n16 73.1255
R14733 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n15 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n14 73.1255
R14734 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n7 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n6 72.3005
R14735 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n22 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n15 68.8946
R14736 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n8 60.9797
R14737 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n23 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n13 41.9827
R14738 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n12 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t9 30.462
R14739 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n12 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t8 30.462
R14740 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t7 30.462
R14741 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t5 30.462
R14742 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t11 30.462
R14743 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t10 30.462
R14744 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n13 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n11 28.124
R14745 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n5 19.963
R14746 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n1 17.8661
R14747 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n2 17.8661
R14748 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n3 17.1217
R14749 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n16 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t2 11.8205
R14750 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n16 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t1 11.8205
R14751 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n19 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t3 11.8205
R14752 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n19 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t6 11.8205
R14753 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n14 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t0 11.8205
R14754 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n14 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t4 11.8205
R14755 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n22 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n21 9.3005
R14756 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n4 1.8615
R14757 a_n18998_n11063.n7 a_n18998_n11063.n1 81.2978
R14758 a_n18998_n11063.n1 a_n18998_n11063.n6 81.1637
R14759 a_n18998_n11063.n1 a_n18998_n11063.n5 81.1637
R14760 a_n18998_n11063.n0 a_n18998_n11063.n4 81.1637
R14761 a_n18998_n11063.n0 a_n18998_n11063.n3 81.1637
R14762 a_n18998_n11063.n0 a_n18998_n11063.n2 80.9213
R14763 a_n18998_n11063.n6 a_n18998_n11063.t8 11.8205
R14764 a_n18998_n11063.n6 a_n18998_n11063.t5 11.8205
R14765 a_n18998_n11063.n5 a_n18998_n11063.t4 11.8205
R14766 a_n18998_n11063.n5 a_n18998_n11063.t3 11.8205
R14767 a_n18998_n11063.n4 a_n18998_n11063.t10 11.8205
R14768 a_n18998_n11063.n4 a_n18998_n11063.t9 11.8205
R14769 a_n18998_n11063.n3 a_n18998_n11063.t0 11.8205
R14770 a_n18998_n11063.n3 a_n18998_n11063.t11 11.8205
R14771 a_n18998_n11063.n2 a_n18998_n11063.t1 11.8205
R14772 a_n18998_n11063.n2 a_n18998_n11063.t2 11.8205
R14773 a_n18998_n11063.t7 a_n18998_n11063.n7 11.8205
R14774 a_n18998_n11063.n7 a_n18998_n11063.t6 11.8205
R14775 a_n18998_n11063.n1 a_n18998_n11063.n0 0.402735
R14776 a_n24130_3190.n2 a_n24130_3190.t2 541.395
R14777 a_n24130_3190.n3 a_n24130_3190.t6 527.402
R14778 a_n24130_3190.n2 a_n24130_3190.t7 491.64
R14779 a_n24130_3190.n5 a_n24130_3190.t0 281.906
R14780 a_n24130_3190.t1 a_n24130_3190.n5 204.359
R14781 a_n24130_3190.n0 a_n24130_3190.t3 180.73
R14782 a_n24130_3190.n1 a_n24130_3190.t5 179.45
R14783 a_n24130_3190.n0 a_n24130_3190.t4 139.78
R14784 a_n24130_3190.n4 a_n24130_3190.n1 105.635
R14785 a_n24130_3190.n4 a_n24130_3190.n3 76.0005
R14786 a_n24130_3190.n5 a_n24130_3190.n4 67.9685
R14787 a_n24130_3190.n3 a_n24130_3190.n2 13.994
R14788 a_n24130_3190.n1 a_n24130_3190.n0 1.28015
R14789 a_n23950_3810.n0 a_n23950_3810.n2 81.3236
R14790 a_n23950_3810.n0 a_n23950_3810.n1 81.2978
R14791 a_n23950_3810.n0 a_n23950_3810.n3 81.1637
R14792 a_n23950_3810.n0 a_n23950_3810.n4 81.1637
R14793 a_n23950_3810.n0 a_n23950_3810.n5 81.1637
R14794 a_n23950_3810.n6 a_n23950_3810.n0 81.1637
R14795 a_n23950_3810.n2 a_n23950_3810.t8 11.8205
R14796 a_n23950_3810.n2 a_n23950_3810.t7 11.8205
R14797 a_n23950_3810.n3 a_n23950_3810.t4 11.8205
R14798 a_n23950_3810.n3 a_n23950_3810.t6 11.8205
R14799 a_n23950_3810.n4 a_n23950_3810.t5 11.8205
R14800 a_n23950_3810.n4 a_n23950_3810.t3 11.8205
R14801 a_n23950_3810.n5 a_n23950_3810.t10 11.8205
R14802 a_n23950_3810.n5 a_n23950_3810.t9 11.8205
R14803 a_n23950_3810.n1 a_n23950_3810.t2 11.8205
R14804 a_n23950_3810.n1 a_n23950_3810.t1 11.8205
R14805 a_n23950_3810.t0 a_n23950_3810.n6 11.8205
R14806 a_n23950_3810.n6 a_n23950_3810.t11 11.8205
R14807 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t12 491.64
R14808 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t18 491.64
R14809 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t14 491.64
R14810 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t22 491.64
R14811 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t15 485.221
R14812 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t17 367.928
R14813 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t16 255.588
R14814 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t19 224.478
R14815 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t20 213.688
R14816 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n18 209.19
R14817 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t23 139.78
R14818 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t13 139.78
R14819 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t21 139.78
R14820 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n1 120.999
R14821 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n0 120.999
R14822 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n13 104.489
R14823 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y 103.258
R14824 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n3 92.5005
R14825 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n8 86.2638
R14826 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n9 85.8873
R14827 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n6 85.724
R14828 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n16 84.5046
R14829 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n14 84.0545
R14830 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n11 75.0672
R14831 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n8 75.0672
R14832 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n10 73.1255
R14833 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n8 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n7 73.1255
R14834 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n6 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n5 73.1255
R14835 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n15 72.3005
R14836 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n6 68.8946
R14837 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n17 60.9816
R14838 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n4 41.9827
R14839 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t0 30.462
R14840 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t1 30.462
R14841 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t3 30.462
R14842 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t2 30.462
R14843 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t10 30.462
R14844 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t8 30.462
R14845 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n2 28.124
R14846 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n19 17.8661
R14847 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n20 17.8661
R14848 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n21 17.1217
R14849 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n23 15.6329
R14850 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t11 11.8205
R14851 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t9 11.8205
R14852 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t4 11.8205
R14853 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t5 11.8205
R14854 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t7 11.8205
R14855 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t6 11.8205
R14856 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y 10.8165
R14857 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n12 9.3005
R14858 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n24 2.50602
R14859 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n22 1.8615
R14860 MULT_0.4bit_ADDER_1.B2.n4 MULT_0.4bit_ADDER_1.B2.t22 491.64
R14861 MULT_0.4bit_ADDER_1.B2.n5 MULT_0.4bit_ADDER_1.B2.t23 491.64
R14862 MULT_0.4bit_ADDER_1.B2.n6 MULT_0.4bit_ADDER_1.B2.t14 491.64
R14863 MULT_0.4bit_ADDER_1.B2.n7 MULT_0.4bit_ADDER_1.B2.t19 491.64
R14864 MULT_0.4bit_ADDER_1.B2.n2 MULT_0.4bit_ADDER_1.B2.t20 485.221
R14865 MULT_0.4bit_ADDER_1.B2.n0 MULT_0.4bit_ADDER_1.B2.t13 367.928
R14866 MULT_0.4bit_ADDER_1.B2.n8 MULT_0.4bit_ADDER_1.B2.t15 255.588
R14867 MULT_0.4bit_ADDER_1.B2.n1 MULT_0.4bit_ADDER_1.B2.t16 224.478
R14868 MULT_0.4bit_ADDER_1.B2.n0 MULT_0.4bit_ADDER_1.B2.t12 213.688
R14869 MULT_0.4bit_ADDER_1.B2.n4 MULT_0.4bit_ADDER_1.B2.n3 209.19
R14870 MULT_0.4bit_ADDER_1.B2.n3 MULT_0.4bit_ADDER_1.B2.t18 139.78
R14871 MULT_0.4bit_ADDER_1.B2.n3 MULT_0.4bit_ADDER_1.B2.t17 139.78
R14872 MULT_0.4bit_ADDER_1.B2.n3 MULT_0.4bit_ADDER_1.B2.t21 139.78
R14873 MULT_0.4bit_ADDER_1.B2.n12 MULT_0.4bit_ADDER_1.B2.n11 120.999
R14874 MULT_0.4bit_ADDER_1.B2.n12 MULT_0.4bit_ADDER_1.B2.n10 120.999
R14875 MULT_0.4bit_ADDER_1.B2.n24 MULT_0.4bit_ADDER_1.B2.n23 104.489
R14876 MULT_0.4bit_ADDER_1.B2.n9 MULT_0.4bit_ADDER_1.B2 103.258
R14877 MULT_0.4bit_ADDER_1.B2.n14 MULT_0.4bit_ADDER_1.B2.n13 92.5005
R14878 MULT_0.4bit_ADDER_1.B2.n21 MULT_0.4bit_ADDER_1.B2.n19 86.2638
R14879 MULT_0.4bit_ADDER_1.B2.n19 MULT_0.4bit_ADDER_1.B2.n18 85.8873
R14880 MULT_0.4bit_ADDER_1.B2.n19 MULT_0.4bit_ADDER_1.B2.n16 85.724
R14881 MULT_0.4bit_ADDER_1.B2.n2 MULT_0.4bit_ADDER_1.B2.n1 84.5046
R14882 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_1.B2.n24 83.8907
R14883 MULT_0.4bit_ADDER_1.B2.n22 MULT_0.4bit_ADDER_1.B2.n21 75.0672
R14884 MULT_0.4bit_ADDER_1.B2.n22 MULT_0.4bit_ADDER_1.B2.n18 75.0672
R14885 MULT_0.4bit_ADDER_1.B2.n21 MULT_0.4bit_ADDER_1.B2.n20 73.1255
R14886 MULT_0.4bit_ADDER_1.B2.n18 MULT_0.4bit_ADDER_1.B2.n17 73.1255
R14887 MULT_0.4bit_ADDER_1.B2.n16 MULT_0.4bit_ADDER_1.B2.n15 73.1255
R14888 MULT_0.4bit_ADDER_1.B2.n1 MULT_0.4bit_ADDER_1.B2.n0 72.3005
R14889 MULT_0.4bit_ADDER_1.B2.n23 MULT_0.4bit_ADDER_1.B2.n16 68.8946
R14890 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_1.B2.n2 60.9816
R14891 MULT_0.4bit_ADDER_1.B2.n24 MULT_0.4bit_ADDER_1.B2.n14 41.9827
R14892 MULT_0.4bit_ADDER_1.B2.n13 MULT_0.4bit_ADDER_1.B2.t1 30.462
R14893 MULT_0.4bit_ADDER_1.B2.n13 MULT_0.4bit_ADDER_1.B2.t2 30.462
R14894 MULT_0.4bit_ADDER_1.B2.n11 MULT_0.4bit_ADDER_1.B2.t3 30.462
R14895 MULT_0.4bit_ADDER_1.B2.n11 MULT_0.4bit_ADDER_1.B2.t6 30.462
R14896 MULT_0.4bit_ADDER_1.B2.n10 MULT_0.4bit_ADDER_1.B2.t8 30.462
R14897 MULT_0.4bit_ADDER_1.B2.n10 MULT_0.4bit_ADDER_1.B2.t0 30.462
R14898 MULT_0.4bit_ADDER_1.B2.n14 MULT_0.4bit_ADDER_1.B2.n12 28.124
R14899 MULT_0.4bit_ADDER_1.B2.n5 MULT_0.4bit_ADDER_1.B2.n4 17.8661
R14900 MULT_0.4bit_ADDER_1.B2.n6 MULT_0.4bit_ADDER_1.B2.n5 17.8661
R14901 MULT_0.4bit_ADDER_1.B2.n7 MULT_0.4bit_ADDER_1.B2.n6 17.1217
R14902 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_1.B2.n8 15.6329
R14903 MULT_0.4bit_ADDER_1.B2.n17 MULT_0.4bit_ADDER_1.B2.t9 11.8205
R14904 MULT_0.4bit_ADDER_1.B2.n17 MULT_0.4bit_ADDER_1.B2.t10 11.8205
R14905 MULT_0.4bit_ADDER_1.B2.n20 MULT_0.4bit_ADDER_1.B2.t5 11.8205
R14906 MULT_0.4bit_ADDER_1.B2.n20 MULT_0.4bit_ADDER_1.B2.t7 11.8205
R14907 MULT_0.4bit_ADDER_1.B2.n15 MULT_0.4bit_ADDER_1.B2.t11 11.8205
R14908 MULT_0.4bit_ADDER_1.B2.n15 MULT_0.4bit_ADDER_1.B2.t4 11.8205
R14909 MULT_0.4bit_ADDER_1.B2.n9 MULT_0.4bit_ADDER_1.B2 10.8165
R14910 MULT_0.4bit_ADDER_1.B2.n23 MULT_0.4bit_ADDER_1.B2.n22 9.3005
R14911 MULT_0.4bit_ADDER_1.B2.n8 MULT_0.4bit_ADDER_1.B2.n7 1.8615
R14912 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_1.B2.n9 0.840348
R14913 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t8 540.38
R14914 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t9 367.928
R14915 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n5 227.526
R14916 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t7 227.356
R14917 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n6 227.266
R14918 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n4 227.266
R14919 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t10 213.688
R14920 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n2 160.439
R14921 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n1 94.4341
R14922 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t0 42.7944
R14923 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t3 30.379
R14924 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t5 30.379
R14925 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t1 30.379
R14926 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t2 30.379
R14927 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t6 30.379
R14928 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.t4 30.379
R14929 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n0 13.4358
R14930 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B.n3 0.821842
R14931 SEL2.n147 SEL2.t41 1388.16
R14932 SEL2.n149 SEL2.t73 1388.16
R14933 SEL2.n156 SEL2.t115 1388.16
R14934 SEL2.n152 SEL2.t94 1388.16
R14935 SEL2.n126 SEL2.t47 1388.16
R14936 SEL2.n128 SEL2.t89 1388.16
R14937 SEL2.n135 SEL2.t134 1388.16
R14938 SEL2.n131 SEL2.t109 1388.16
R14939 SEL2.n105 SEL2.t40 1388.16
R14940 SEL2.n107 SEL2.t29 1388.16
R14941 SEL2.n114 SEL2.t78 1388.16
R14942 SEL2.n110 SEL2.t2 1388.16
R14943 SEL2.n84 SEL2.t117 1388.16
R14944 SEL2.n86 SEL2.t93 1388.16
R14945 SEL2.n93 SEL2.t14 1388.16
R14946 SEL2.n89 SEL2.t52 1388.16
R14947 SEL2.n63 SEL2.t10 1388.16
R14948 SEL2.n65 SEL2.t140 1388.16
R14949 SEL2.n72 SEL2.t38 1388.16
R14950 SEL2.n68 SEL2.t98 1388.16
R14951 SEL2.n42 SEL2.t74 1388.16
R14952 SEL2.n44 SEL2.t55 1388.16
R14953 SEL2.n51 SEL2.t126 1388.16
R14954 SEL2.n47 SEL2.t31 1388.16
R14955 SEL2.n21 SEL2.t123 1388.16
R14956 SEL2.n23 SEL2.t99 1388.16
R14957 SEL2.n30 SEL2.t17 1388.16
R14958 SEL2.n26 SEL2.t60 1388.16
R14959 SEL2.n1 SEL2.t77 1388.16
R14960 SEL2.n3 SEL2.t58 1388.16
R14961 SEL2.n10 SEL2.t130 1388.16
R14962 SEL2.n6 SEL2.t33 1388.16
R14963 SEL2.n169 SEL2.t118 1388.16
R14964 SEL2.n171 SEL2.t86 1388.16
R14965 SEL2.n178 SEL2.t34 1388.16
R14966 SEL2.n174 SEL2.t133 1388.16
R14967 SEL2.n162 SEL2.t28 385.697
R14968 SEL2.n141 SEL2.t32 385.697
R14969 SEL2.n120 SEL2.t84 385.697
R14970 SEL2.n99 SEL2.t19 385.697
R14971 SEL2.n78 SEL2.t132 385.697
R14972 SEL2.n57 SEL2.t21 385.697
R14973 SEL2.n36 SEL2.t85 385.697
R14974 SEL2.n16 SEL2.t75 385.697
R14975 SEL2.n185 SEL2.t4 385.697
R14976 SEL2.n147 SEL2.t13 350.839
R14977 SEL2.n149 SEL2.t44 350.839
R14978 SEL2.n156 SEL2.t131 350.839
R14979 SEL2.n152 SEL2.t23 350.839
R14980 SEL2.n126 SEL2.t127 350.839
R14981 SEL2.n128 SEL2.t25 350.839
R14982 SEL2.n135 SEL2.t87 350.839
R14983 SEL2.n131 SEL2.t142 350.839
R14984 SEL2.n105 SEL2.t30 350.839
R14985 SEL2.n107 SEL2.t5 350.839
R14986 SEL2.n114 SEL2.t42 350.839
R14987 SEL2.n110 SEL2.t27 350.839
R14988 SEL2.n84 SEL2.t95 350.839
R14989 SEL2.n86 SEL2.t112 350.839
R14990 SEL2.n93 SEL2.t119 350.839
R14991 SEL2.n89 SEL2.t90 350.839
R14992 SEL2.n63 SEL2.t97 350.839
R14993 SEL2.n65 SEL2.t114 350.839
R14994 SEL2.n72 SEL2.t124 350.839
R14995 SEL2.n68 SEL2.t92 350.839
R14996 SEL2.n42 SEL2.t56 350.839
R14997 SEL2.n44 SEL2.t70 350.839
R14998 SEL2.n51 SEL2.t80 350.839
R14999 SEL2.n47 SEL2.t51 350.839
R15000 SEL2.n21 SEL2.t101 350.839
R15001 SEL2.n23 SEL2.t116 350.839
R15002 SEL2.n30 SEL2.t128 350.839
R15003 SEL2.n26 SEL2.t96 350.839
R15004 SEL2.n1 SEL2.t59 350.839
R15005 SEL2.n3 SEL2.t36 350.839
R15006 SEL2.n10 SEL2.t83 350.839
R15007 SEL2.n6 SEL2.t53 350.839
R15008 SEL2.n169 SEL2.t138 350.839
R15009 SEL2.n171 SEL2.t49 350.839
R15010 SEL2.n178 SEL2.t113 350.839
R15011 SEL2.n174 SEL2.t76 350.839
R15012 SEL2.n148 SEL2.t8 308.481
R15013 SEL2.n150 SEL2.t37 308.481
R15014 SEL2.n157 SEL2.t108 308.481
R15015 SEL2.n153 SEL2.t7 308.481
R15016 SEL2.n127 SEL2.t122 308.481
R15017 SEL2.n129 SEL2.t12 308.481
R15018 SEL2.n136 SEL2.t68 308.481
R15019 SEL2.n132 SEL2.t121 308.481
R15020 SEL2.n106 SEL2.t63 308.481
R15021 SEL2.n108 SEL2.t11 308.481
R15022 SEL2.n115 SEL2.t45 308.481
R15023 SEL2.n111 SEL2.t35 308.481
R15024 SEL2.n85 SEL2.t0 308.481
R15025 SEL2.n87 SEL2.t120 308.481
R15026 SEL2.n94 SEL2.t135 308.481
R15027 SEL2.n90 SEL2.t102 308.481
R15028 SEL2.n64 SEL2.t1 308.481
R15029 SEL2.n66 SEL2.t125 308.481
R15030 SEL2.n73 SEL2.t136 308.481
R15031 SEL2.n69 SEL2.t103 308.481
R15032 SEL2.n43 SEL2.t104 308.481
R15033 SEL2.n45 SEL2.t82 308.481
R15034 SEL2.n52 SEL2.t88 308.481
R15035 SEL2.n48 SEL2.t61 308.481
R15036 SEL2.n22 SEL2.t3 308.481
R15037 SEL2.n24 SEL2.t129 308.481
R15038 SEL2.n31 SEL2.t139 308.481
R15039 SEL2.n27 SEL2.t105 308.481
R15040 SEL2.n2 SEL2.t107 308.481
R15041 SEL2.n4 SEL2.t39 308.481
R15042 SEL2.n11 SEL2.t91 308.481
R15043 SEL2.n7 SEL2.t65 308.481
R15044 SEL2.n170 SEL2.t66 308.481
R15045 SEL2.n172 SEL2.t69 308.481
R15046 SEL2.n179 SEL2.t137 308.481
R15047 SEL2.n175 SEL2.t100 308.481
R15048 SEL2.n146 SEL2.t22 291.829
R15049 SEL2.n146 SEL2.t62 291.829
R15050 SEL2.n125 SEL2.t24 291.829
R15051 SEL2.n125 SEL2.t67 291.829
R15052 SEL2.n104 SEL2.t71 291.829
R15053 SEL2.n104 SEL2.t143 291.829
R15054 SEL2.n83 SEL2.t72 291.829
R15055 SEL2.n83 SEL2.t141 291.829
R15056 SEL2.n62 SEL2.t106 291.829
R15057 SEL2.n62 SEL2.t57 291.829
R15058 SEL2.n41 SEL2.t6 291.829
R15059 SEL2.n41 SEL2.t46 291.829
R15060 SEL2.n20 SEL2.t110 291.829
R15061 SEL2.n20 SEL2.t26 291.829
R15062 SEL2.n0 SEL2.t9 291.829
R15063 SEL2.n0 SEL2.t48 291.829
R15064 SEL2.n183 SEL2.t50 291.829
R15065 SEL2.n183 SEL2.t111 291.829
R15066 SEL2.n146 SEL2.t54 221.72
R15067 SEL2.n125 SEL2.t64 221.72
R15068 SEL2.n104 SEL2.t79 221.72
R15069 SEL2.n83 SEL2.t81 221.72
R15070 SEL2.n62 SEL2.t15 221.72
R15071 SEL2.n41 SEL2.t43 221.72
R15072 SEL2.n20 SEL2.t16 221.72
R15073 SEL2.n0 SEL2.t18 221.72
R15074 SEL2.n183 SEL2.t20 221.72
R15075 SEL2 SEL2.n148 161.492
R15076 SEL2 SEL2.n127 161.492
R15077 SEL2 SEL2.n106 161.492
R15078 SEL2 SEL2.n85 161.492
R15079 SEL2 SEL2.n64 161.492
R15080 SEL2 SEL2.n43 161.492
R15081 SEL2 SEL2.n22 161.492
R15082 SEL2 SEL2.n2 161.492
R15083 SEL2 SEL2.n170 161.492
R15084 SEL2.n154 SEL2.n153 161.442
R15085 SEL2.n133 SEL2.n132 161.442
R15086 SEL2.n112 SEL2.n111 161.442
R15087 SEL2.n91 SEL2.n90 161.442
R15088 SEL2.n70 SEL2.n69 161.442
R15089 SEL2.n49 SEL2.n48 161.442
R15090 SEL2.n28 SEL2.n27 161.442
R15091 SEL2.n8 SEL2.n7 161.442
R15092 SEL2.n176 SEL2.n175 161.442
R15093 SEL2.n158 SEL2.n157 161.429
R15094 SEL2.n137 SEL2.n136 161.429
R15095 SEL2.n116 SEL2.n115 161.429
R15096 SEL2.n95 SEL2.n94 161.429
R15097 SEL2.n74 SEL2.n73 161.429
R15098 SEL2.n53 SEL2.n52 161.429
R15099 SEL2.n32 SEL2.n31 161.429
R15100 SEL2.n12 SEL2.n11 161.429
R15101 SEL2.n180 SEL2.n179 161.429
R15102 SEL2.n151 SEL2.n150 161.389
R15103 SEL2.n130 SEL2.n129 161.389
R15104 SEL2.n109 SEL2.n108 161.389
R15105 SEL2.n88 SEL2.n87 161.389
R15106 SEL2.n67 SEL2.n66 161.389
R15107 SEL2.n46 SEL2.n45 161.389
R15108 SEL2.n25 SEL2.n24 161.389
R15109 SEL2.n5 SEL2.n4 161.389
R15110 SEL2.n173 SEL2.n172 161.389
R15111 SEL2.n163 SEL2.n162 89.6005
R15112 SEL2.n142 SEL2.n141 89.6005
R15113 SEL2.n121 SEL2.n120 89.6005
R15114 SEL2.n100 SEL2.n99 89.6005
R15115 SEL2.n79 SEL2.n78 89.6005
R15116 SEL2.n58 SEL2.n57 89.6005
R15117 SEL2.n37 SEL2.n36 89.6005
R15118 SEL2.n17 SEL2.n16 89.6005
R15119 SEL2.n185 SEL2.n184 89.6005
R15120 SEL2.n163 SEL2.n146 50.6672
R15121 SEL2.n142 SEL2.n125 50.6672
R15122 SEL2.n121 SEL2.n104 50.6672
R15123 SEL2.n100 SEL2.n83 50.6672
R15124 SEL2.n79 SEL2.n62 50.6672
R15125 SEL2.n58 SEL2.n41 50.6672
R15126 SEL2.n37 SEL2.n20 50.6672
R15127 SEL2.n17 SEL2.n0 50.6672
R15128 SEL2.n184 SEL2.n183 50.6672
R15129 SEL2.n148 SEL2.n147 27.752
R15130 SEL2.n150 SEL2.n149 27.752
R15131 SEL2.n157 SEL2.n156 27.752
R15132 SEL2.n153 SEL2.n152 27.752
R15133 SEL2.n127 SEL2.n126 27.752
R15134 SEL2.n129 SEL2.n128 27.752
R15135 SEL2.n136 SEL2.n135 27.752
R15136 SEL2.n132 SEL2.n131 27.752
R15137 SEL2.n106 SEL2.n105 27.752
R15138 SEL2.n108 SEL2.n107 27.752
R15139 SEL2.n115 SEL2.n114 27.752
R15140 SEL2.n111 SEL2.n110 27.752
R15141 SEL2.n85 SEL2.n84 27.752
R15142 SEL2.n87 SEL2.n86 27.752
R15143 SEL2.n94 SEL2.n93 27.752
R15144 SEL2.n90 SEL2.n89 27.752
R15145 SEL2.n64 SEL2.n63 27.752
R15146 SEL2.n66 SEL2.n65 27.752
R15147 SEL2.n73 SEL2.n72 27.752
R15148 SEL2.n69 SEL2.n68 27.752
R15149 SEL2.n43 SEL2.n42 27.752
R15150 SEL2.n45 SEL2.n44 27.752
R15151 SEL2.n52 SEL2.n51 27.752
R15152 SEL2.n48 SEL2.n47 27.752
R15153 SEL2.n22 SEL2.n21 27.752
R15154 SEL2.n24 SEL2.n23 27.752
R15155 SEL2.n31 SEL2.n30 27.752
R15156 SEL2.n27 SEL2.n26 27.752
R15157 SEL2.n2 SEL2.n1 27.752
R15158 SEL2.n4 SEL2.n3 27.752
R15159 SEL2.n11 SEL2.n10 27.752
R15160 SEL2.n7 SEL2.n6 27.752
R15161 SEL2.n170 SEL2.n169 27.752
R15162 SEL2.n172 SEL2.n171 27.752
R15163 SEL2.n179 SEL2.n178 27.752
R15164 SEL2.n175 SEL2.n174 27.752
R15165 SEL2.n160 SEL2.n159 11.1236
R15166 SEL2.n139 SEL2.n138 11.1236
R15167 SEL2.n118 SEL2.n117 11.1236
R15168 SEL2.n97 SEL2.n96 11.1236
R15169 SEL2.n76 SEL2.n75 11.1236
R15170 SEL2.n55 SEL2.n54 11.1236
R15171 SEL2.n34 SEL2.n33 11.1236
R15172 SEL2.n14 SEL2.n13 11.1236
R15173 SEL2.n182 SEL2.n181 11.1236
R15174 SEL2.n155 SEL2.n151 10.8168
R15175 SEL2.n134 SEL2.n130 10.8168
R15176 SEL2.n113 SEL2.n109 10.8168
R15177 SEL2.n92 SEL2.n88 10.8168
R15178 SEL2.n71 SEL2.n67 10.8168
R15179 SEL2.n50 SEL2.n46 10.8168
R15180 SEL2.n29 SEL2.n25 10.8168
R15181 SEL2.n9 SEL2.n5 10.8168
R15182 SEL2.n177 SEL2.n173 10.8168
R15183 SEL2.n144 SEL2.n143 9.56357
R15184 SEL2.n168 SEL2.n167 9.55995
R15185 SEL2.n81 SEL2.n80 9.54183
R15186 SEL2.n165 SEL2.n164 9.53096
R15187 SEL2.n19 SEL2.n18 9.52553
R15188 SEL2.n60 SEL2.n59 9.51285
R15189 SEL2.n102 SEL2.n101 9.50198
R15190 SEL2.n123 SEL2.n122 9.50017
R15191 SEL2.n39 SEL2.n38 9.49111
R15192 SEL2.n162 SEL2.n161 9.3005
R15193 SEL2.n141 SEL2.n140 9.3005
R15194 SEL2.n120 SEL2.n119 9.3005
R15195 SEL2.n99 SEL2.n98 9.3005
R15196 SEL2.n78 SEL2.n77 9.3005
R15197 SEL2.n57 SEL2.n56 9.3005
R15198 SEL2.n36 SEL2.n35 9.3005
R15199 SEL2.n16 SEL2.n15 9.3005
R15200 SEL2.n186 SEL2.n185 9.3005
R15201 SEL2.n155 SEL2.n154 9.0005
R15202 SEL2.n159 SEL2.n158 9.0005
R15203 SEL2.n134 SEL2.n133 9.0005
R15204 SEL2.n138 SEL2.n137 9.0005
R15205 SEL2.n113 SEL2.n112 9.0005
R15206 SEL2.n117 SEL2.n116 9.0005
R15207 SEL2.n92 SEL2.n91 9.0005
R15208 SEL2.n96 SEL2.n95 9.0005
R15209 SEL2.n71 SEL2.n70 9.0005
R15210 SEL2.n75 SEL2.n74 9.0005
R15211 SEL2.n50 SEL2.n49 9.0005
R15212 SEL2.n54 SEL2.n53 9.0005
R15213 SEL2.n29 SEL2.n28 9.0005
R15214 SEL2.n33 SEL2.n32 9.0005
R15215 SEL2.n9 SEL2.n8 9.0005
R15216 SEL2.n13 SEL2.n12 9.0005
R15217 SEL2.n177 SEL2.n176 9.0005
R15218 SEL2.n181 SEL2.n180 9.0005
R15219 SEL2.n161 SEL2.n160 7.80174
R15220 SEL2.n140 SEL2.n139 7.80174
R15221 SEL2.n119 SEL2.n118 7.80174
R15222 SEL2.n98 SEL2.n97 7.80174
R15223 SEL2.n77 SEL2.n76 7.80174
R15224 SEL2.n56 SEL2.n55 7.80174
R15225 SEL2.n35 SEL2.n34 7.80174
R15226 SEL2.n15 SEL2.n14 7.80174
R15227 SEL2.n186 SEL2.n182 7.80174
R15228 SEL2.n167 SEL2.n166 6.50224
R15229 SEL2.n40 SEL2.n19 6.48185
R15230 SEL2.n40 SEL2.n39 3.4105
R15231 SEL2.n61 SEL2.n60 3.4105
R15232 SEL2.n82 SEL2.n81 3.4105
R15233 SEL2.n103 SEL2.n102 3.4105
R15234 SEL2.n124 SEL2.n123 3.4105
R15235 SEL2.n145 SEL2.n144 3.4105
R15236 SEL2.n166 SEL2.n165 3.4105
R15237 SEL2.n145 SEL2.n124 3.17675
R15238 SEL2.n164 SEL2.n163 3.1005
R15239 SEL2.n143 SEL2.n142 3.1005
R15240 SEL2.n122 SEL2.n121 3.1005
R15241 SEL2.n101 SEL2.n100 3.1005
R15242 SEL2.n80 SEL2.n79 3.1005
R15243 SEL2.n59 SEL2.n58 3.1005
R15244 SEL2.n38 SEL2.n37 3.1005
R15245 SEL2.n18 SEL2.n17 3.1005
R15246 SEL2.n184 SEL2.n168 3.1005
R15247 SEL2.n82 SEL2.n61 3.09569
R15248 SEL2.n61 SEL2.n40 3.09296
R15249 SEL2.n124 SEL2.n103 3.08411
R15250 SEL2.n103 SEL2.n82 3.0698
R15251 SEL2.n166 SEL2.n145 3.00441
R15252 SEL2.n159 SEL2.n155 1.75997
R15253 SEL2.n138 SEL2.n134 1.75997
R15254 SEL2.n117 SEL2.n113 1.75997
R15255 SEL2.n96 SEL2.n92 1.75997
R15256 SEL2.n75 SEL2.n71 1.75997
R15257 SEL2.n54 SEL2.n50 1.75997
R15258 SEL2.n33 SEL2.n29 1.75997
R15259 SEL2.n13 SEL2.n9 1.75997
R15260 SEL2.n181 SEL2.n177 1.75997
R15261 SEL2.n161 SEL2 0.393745
R15262 SEL2.n140 SEL2 0.393745
R15263 SEL2.n119 SEL2 0.393745
R15264 SEL2.n98 SEL2 0.393745
R15265 SEL2.n77 SEL2 0.393745
R15266 SEL2.n56 SEL2 0.393745
R15267 SEL2.n35 SEL2 0.393745
R15268 SEL2.n15 SEL2 0.393745
R15269 SEL2 SEL2.n186 0.393745
R15270 SEL2.n160 SEL2 0.265652
R15271 SEL2.n139 SEL2 0.265652
R15272 SEL2.n118 SEL2 0.265652
R15273 SEL2.n97 SEL2 0.265652
R15274 SEL2.n76 SEL2 0.265652
R15275 SEL2.n55 SEL2 0.265652
R15276 SEL2.n34 SEL2 0.265652
R15277 SEL2.n14 SEL2 0.265652
R15278 SEL2.n182 SEL2 0.265652
R15279 SEL2.n164 SEL2 0.237819
R15280 SEL2.n143 SEL2 0.237819
R15281 SEL2.n122 SEL2 0.237819
R15282 SEL2.n101 SEL2 0.237819
R15283 SEL2.n80 SEL2 0.237819
R15284 SEL2.n59 SEL2 0.237819
R15285 SEL2.n38 SEL2 0.237819
R15286 SEL2.n18 SEL2 0.237819
R15287 SEL2 SEL2.n168 0.237819
R15288 SEL2.n151 SEL2 0.102773
R15289 SEL2.n130 SEL2 0.102773
R15290 SEL2.n109 SEL2 0.102773
R15291 SEL2.n88 SEL2 0.102773
R15292 SEL2.n67 SEL2 0.102773
R15293 SEL2.n46 SEL2 0.102773
R15294 SEL2.n25 SEL2 0.102773
R15295 SEL2.n5 SEL2 0.102773
R15296 SEL2.n173 SEL2 0.102773
R15297 SEL2.n39 SEL2 0.0838333
R15298 SEL2.n123 SEL2 0.0747754
R15299 SEL2.n102 SEL2 0.0729638
R15300 SEL2.n158 SEL2 0.063
R15301 SEL2.n137 SEL2 0.063
R15302 SEL2.n116 SEL2 0.063
R15303 SEL2.n95 SEL2 0.063
R15304 SEL2.n74 SEL2 0.063
R15305 SEL2.n53 SEL2 0.063
R15306 SEL2.n32 SEL2 0.063
R15307 SEL2.n12 SEL2 0.063
R15308 SEL2.n180 SEL2 0.063
R15309 SEL2.n60 SEL2 0.0620942
R15310 SEL2.n154 SEL2 0.0497424
R15311 SEL2.n133 SEL2 0.0497424
R15312 SEL2.n112 SEL2 0.0497424
R15313 SEL2.n91 SEL2 0.0497424
R15314 SEL2.n70 SEL2 0.0497424
R15315 SEL2.n49 SEL2 0.0497424
R15316 SEL2.n28 SEL2 0.0497424
R15317 SEL2.n8 SEL2 0.0497424
R15318 SEL2.n176 SEL2 0.0497424
R15319 SEL2.n19 SEL2 0.049413
R15320 SEL2.n165 SEL2 0.0439783
R15321 SEL2.n81 SEL2 0.0331087
R15322 SEL2.n167 SEL2 0.0149928
R15323 SEL2.n144 SEL2 0.0113696
R15324 mux8_4.NAND4F_5.Y.n1 mux8_4.NAND4F_5.Y.t9 1032.02
R15325 mux8_4.NAND4F_5.Y.n1 mux8_4.NAND4F_5.Y.t10 336.962
R15326 mux8_4.NAND4F_5.Y.n1 mux8_4.NAND4F_5.Y.t11 326.154
R15327 mux8_4.NAND4F_5.Y.n0 mux8_4.NAND4F_5.Y.n3 187.373
R15328 mux8_4.NAND4F_5.Y.n0 mux8_4.NAND4F_5.Y.n4 187.192
R15329 mux8_4.NAND4F_5.Y.n0 mux8_4.NAND4F_5.Y.n5 187.192
R15330 mux8_4.NAND4F_5.Y.n7 mux8_4.NAND4F_5.Y.n6 187.192
R15331 mux8_4.NAND4F_5.Y mux8_4.NAND4F_5.Y.n1 162.94
R15332 mux8_4.NAND4F_5.Y.n2 mux8_4.NAND4F_5.Y 24.4721
R15333 mux8_4.NAND4F_5.Y.n2 mux8_4.NAND4F_5.Y.t2 22.6141
R15334 mux8_4.NAND4F_5.Y.n3 mux8_4.NAND4F_5.Y.t0 20.1899
R15335 mux8_4.NAND4F_5.Y.n3 mux8_4.NAND4F_5.Y.t1 20.1899
R15336 mux8_4.NAND4F_5.Y.n4 mux8_4.NAND4F_5.Y.t6 20.1899
R15337 mux8_4.NAND4F_5.Y.n4 mux8_4.NAND4F_5.Y.t5 20.1899
R15338 mux8_4.NAND4F_5.Y.n5 mux8_4.NAND4F_5.Y.t7 20.1899
R15339 mux8_4.NAND4F_5.Y.n5 mux8_4.NAND4F_5.Y.t8 20.1899
R15340 mux8_4.NAND4F_5.Y.n6 mux8_4.NAND4F_5.Y.t3 20.1899
R15341 mux8_4.NAND4F_5.Y.n6 mux8_4.NAND4F_5.Y.t4 20.1899
R15342 mux8_4.NAND4F_5.Y mux8_4.NAND4F_5.Y.n2 0.950576
R15343 mux8_4.NAND4F_5.Y mux8_4.NAND4F_5.Y.n7 0.396904
R15344 mux8_4.NAND4F_5.Y.n7 mux8_4.NAND4F_5.Y.n0 0.358709
R15345 MULT_0.inv_9.Y.n2 MULT_0.inv_9.Y.t5 540.38
R15346 MULT_0.inv_9.Y.n3 MULT_0.inv_9.Y.t15 491.64
R15347 MULT_0.inv_9.Y.n3 MULT_0.inv_9.Y.t10 491.64
R15348 MULT_0.inv_9.Y.n3 MULT_0.inv_9.Y.t11 491.64
R15349 MULT_0.inv_9.Y.n3 MULT_0.inv_9.Y.t12 491.64
R15350 MULT_0.inv_9.Y.n0 MULT_0.inv_9.Y.t7 367.928
R15351 MULT_0.inv_9.Y MULT_0.inv_9.Y.t1 256.514
R15352 MULT_0.inv_9.Y.n1 MULT_0.inv_9.Y.t14 227.356
R15353 MULT_0.inv_9.Y MULT_0.inv_9.Y.n7 226.136
R15354 MULT_0.inv_9.Y.n0 MULT_0.inv_9.Y.t4 213.688
R15355 MULT_0.inv_9.Y MULT_0.inv_9.Y.n5 162.867
R15356 MULT_0.inv_9.Y.n2 MULT_0.inv_9.Y.n1 160.439
R15357 MULT_0.inv_9.Y.n4 MULT_0.inv_9.Y.t8 139.78
R15358 MULT_0.inv_9.Y.n4 MULT_0.inv_9.Y.t9 139.78
R15359 MULT_0.inv_9.Y.n4 MULT_0.inv_9.Y.t13 139.78
R15360 MULT_0.inv_9.Y.n4 MULT_0.inv_9.Y.t6 139.78
R15361 MULT_0.inv_9.Y.n1 MULT_0.inv_9.Y.n0 94.4341
R15362 MULT_0.inv_9.Y MULT_0.inv_9.Y.t0 83.8039
R15363 MULT_0.inv_9.Y.n5 MULT_0.inv_9.Y.n4 38.6833
R15364 MULT_0.inv_9.Y.n7 MULT_0.inv_9.Y.t3 30.379
R15365 MULT_0.inv_9.Y.n7 MULT_0.inv_9.Y.t2 30.379
R15366 MULT_0.inv_9.Y.n5 MULT_0.inv_9.Y.n3 28.3986
R15367 MULT_0.inv_9.Y MULT_0.inv_9.Y.n6 16.8032
R15368 MULT_0.inv_9.Y.n6 MULT_0.inv_9.Y 9.00496
R15369 MULT_0.inv_9.Y.n6 MULT_0.inv_9.Y 3.87912
R15370 MULT_0.inv_9.Y MULT_0.inv_9.Y.n2 0.89693
R15371 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t9 540.38
R15372 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t10 367.928
R15373 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n4 227.526
R15374 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t7 227.356
R15375 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n5 227.266
R15376 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n6 227.266
R15377 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t8 213.688
R15378 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n2 160.439
R15379 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n1 94.4341
R15380 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t0 42.7944
R15381 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t5 30.379
R15382 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t4 30.379
R15383 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t1 30.379
R15384 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t6 30.379
R15385 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t2 30.379
R15386 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.t3 30.379
R15387 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n0 13.4358
R15388 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B.n3 0.821842
R15389 a_n13381_373.t0 a_n13381_373.t1 19.8005
R15390 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t7 485.221
R15391 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t10 367.928
R15392 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n4 227.526
R15393 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n5 227.266
R15394 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n6 227.266
R15395 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t8 224.478
R15396 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t9 213.688
R15397 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n2 84.5046
R15398 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n1 72.3005
R15399 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n3 61.0566
R15400 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t3 42.7747
R15401 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t2 30.379
R15402 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t1 30.379
R15403 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t5 30.379
R15404 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t0 30.379
R15405 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t6 30.379
R15406 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.t4 30.379
R15407 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A.n0 0.583137
R15408 a_n14005_n8445.n2 a_n14005_n8445.t7 541.395
R15409 a_n14005_n8445.n3 a_n14005_n8445.t3 527.402
R15410 a_n14005_n8445.n2 a_n14005_n8445.t6 491.64
R15411 a_n14005_n8445.n5 a_n14005_n8445.t1 281.906
R15412 a_n14005_n8445.t0 a_n14005_n8445.n5 204.359
R15413 a_n14005_n8445.n0 a_n14005_n8445.t2 180.73
R15414 a_n14005_n8445.n1 a_n14005_n8445.t4 179.45
R15415 a_n14005_n8445.n0 a_n14005_n8445.t5 139.78
R15416 a_n14005_n8445.n4 a_n14005_n8445.n1 105.635
R15417 a_n14005_n8445.n4 a_n14005_n8445.n3 76.0005
R15418 a_n14005_n8445.n5 a_n14005_n8445.n4 67.9685
R15419 a_n14005_n8445.n3 a_n14005_n8445.n2 13.994
R15420 a_n14005_n8445.n1 a_n14005_n8445.n0 1.28015
R15421 a_n13975_n8419.n2 a_n13975_n8419.n0 121.353
R15422 a_n13975_n8419.n2 a_n13975_n8419.n1 121.001
R15423 a_n13975_n8419.n3 a_n13975_n8419.n2 120.977
R15424 a_n13975_n8419.n0 a_n13975_n8419.t3 30.462
R15425 a_n13975_n8419.n0 a_n13975_n8419.t4 30.462
R15426 a_n13975_n8419.n1 a_n13975_n8419.t0 30.462
R15427 a_n13975_n8419.n1 a_n13975_n8419.t5 30.462
R15428 a_n13975_n8419.t2 a_n13975_n8419.n3 30.462
R15429 a_n13975_n8419.n3 a_n13975_n8419.t1 30.462
R15430 mux8_5.NAND4F_0.C.n6 mux8_5.NAND4F_0.C.t5 978.795
R15431 mux8_5.NAND4F_0.C.n4 mux8_5.NAND4F_0.C.t12 978.795
R15432 mux8_5.NAND4F_0.C.n11 mux8_5.NAND4F_0.C.t13 978.795
R15433 mux8_5.NAND4F_0.C.n2 mux8_5.NAND4F_0.C.t14 978.795
R15434 mux8_5.NAND4F_0.C.n5 mux8_5.NAND4F_0.C.t4 308.481
R15435 mux8_5.NAND4F_0.C.n5 mux8_5.NAND4F_0.C.t15 308.481
R15436 mux8_5.NAND4F_0.C.n3 mux8_5.NAND4F_0.C.t11 308.481
R15437 mux8_5.NAND4F_0.C.n3 mux8_5.NAND4F_0.C.t9 308.481
R15438 mux8_5.NAND4F_0.C.n10 mux8_5.NAND4F_0.C.t6 308.481
R15439 mux8_5.NAND4F_0.C.n10 mux8_5.NAND4F_0.C.t7 308.481
R15440 mux8_5.NAND4F_0.C.n1 mux8_5.NAND4F_0.C.t8 308.481
R15441 mux8_5.NAND4F_0.C.n1 mux8_5.NAND4F_0.C.t10 308.481
R15442 mux8_5.NAND4F_0.C.n0 mux8_5.NAND4F_0.C.t2 256.514
R15443 mux8_5.NAND4F_0.C.n0 mux8_5.NAND4F_0.C.n8 226.258
R15444 mux8_5.NAND4F_0.C mux8_5.NAND4F_0.C.n6 161.856
R15445 mux8_5.NAND4F_0.C mux8_5.NAND4F_0.C.n4 161.847
R15446 mux8_5.NAND4F_0.C mux8_5.NAND4F_0.C.n11 161.84
R15447 mux8_5.NAND4F_0.C mux8_5.NAND4F_0.C.n2 161.831
R15448 mux8_5.NAND4F_0.C.n0 mux8_5.NAND4F_0.C.t0 83.7172
R15449 mux8_5.NAND4F_0.C.n8 mux8_5.NAND4F_0.C.t1 30.379
R15450 mux8_5.NAND4F_0.C.n8 mux8_5.NAND4F_0.C.t3 30.379
R15451 mux8_5.NAND4F_0.C.n9 mux8_5.NAND4F_0.C.n0 13.5186
R15452 mux8_5.NAND4F_0.C mux8_5.NAND4F_0.C.n12 13.0862
R15453 mux8_5.NAND4F_0.C.n7 mux8_5.NAND4F_0.C 13.0435
R15454 mux8_5.NAND4F_0.C.n12 mux8_5.NAND4F_0.C 12.4135
R15455 mux8_5.NAND4F_0.C.n7 mux8_5.NAND4F_0.C 12.4105
R15456 mux8_5.NAND4F_0.C.n6 mux8_5.NAND4F_0.C.n5 11.0463
R15457 mux8_5.NAND4F_0.C.n4 mux8_5.NAND4F_0.C.n3 11.0463
R15458 mux8_5.NAND4F_0.C.n11 mux8_5.NAND4F_0.C.n10 11.0463
R15459 mux8_5.NAND4F_0.C.n2 mux8_5.NAND4F_0.C.n1 11.0463
R15460 mux8_5.NAND4F_0.C.n12 mux8_5.NAND4F_0.C.n9 3.46056
R15461 mux8_5.NAND4F_0.C.n9 mux8_5.NAND4F_0.C.n7 1.8134
R15462 mux8_5.NAND4F_3.Y.n7 mux8_5.NAND4F_3.Y.t11 978.795
R15463 mux8_5.NAND4F_3.Y.n6 mux8_5.NAND4F_3.Y.t10 308.481
R15464 mux8_5.NAND4F_3.Y.n6 mux8_5.NAND4F_3.Y.t9 308.481
R15465 mux8_5.NAND4F_3.Y.n0 mux8_5.NAND4F_3.Y.n1 187.373
R15466 mux8_5.NAND4F_3.Y.n0 mux8_5.NAND4F_3.Y.n2 187.192
R15467 mux8_5.NAND4F_3.Y.n0 mux8_5.NAND4F_3.Y.n3 187.192
R15468 mux8_5.NAND4F_3.Y.n5 mux8_5.NAND4F_3.Y.n4 187.192
R15469 mux8_5.NAND4F_3.Y mux8_5.NAND4F_3.Y.n7 161.839
R15470 mux8_5.NAND4F_3.Y mux8_5.NAND4F_3.Y.t8 23.4426
R15471 mux8_5.NAND4F_3.Y.n1 mux8_5.NAND4F_3.Y.t2 20.1899
R15472 mux8_5.NAND4F_3.Y.n1 mux8_5.NAND4F_3.Y.t3 20.1899
R15473 mux8_5.NAND4F_3.Y.n2 mux8_5.NAND4F_3.Y.t0 20.1899
R15474 mux8_5.NAND4F_3.Y.n2 mux8_5.NAND4F_3.Y.t1 20.1899
R15475 mux8_5.NAND4F_3.Y.n3 mux8_5.NAND4F_3.Y.t4 20.1899
R15476 mux8_5.NAND4F_3.Y.n3 mux8_5.NAND4F_3.Y.t5 20.1899
R15477 mux8_5.NAND4F_3.Y.n4 mux8_5.NAND4F_3.Y.t6 20.1899
R15478 mux8_5.NAND4F_3.Y.n4 mux8_5.NAND4F_3.Y.t7 20.1899
R15479 mux8_5.NAND4F_3.Y.n7 mux8_5.NAND4F_3.Y.n6 11.0463
R15480 mux8_5.NAND4F_3.Y mux8_5.NAND4F_3.Y.n5 0.518495
R15481 mux8_5.NAND4F_3.Y.n5 mux8_5.NAND4F_3.Y.n0 0.358709
R15482 NOT8_0.S3.n1 NOT8_0.S3.t5 1032.02
R15483 NOT8_0.S3.n1 NOT8_0.S3.t6 336.962
R15484 NOT8_0.S3.n1 NOT8_0.S3.t4 326.154
R15485 NOT8_0.S3.n0 NOT8_0.S3.t1 256.514
R15486 NOT8_0.S3.n0 NOT8_0.S3.n2 226.258
R15487 NOT8_0.S3 NOT8_0.S3.n1 162.952
R15488 NOT8_0.S3.n0 NOT8_0.S3.t3 83.7172
R15489 NOT8_0.S3.n2 NOT8_0.S3.t2 30.379
R15490 NOT8_0.S3.n2 NOT8_0.S3.t0 30.379
R15491 NOT8_0.S3 NOT8_0.S3.n0 1.9182
R15492 mux8_4.NAND4F_7.Y.n2 mux8_4.NAND4F_7.Y.t11 1388.16
R15493 mux8_4.NAND4F_7.Y.n2 mux8_4.NAND4F_7.Y.t10 350.839
R15494 mux8_4.NAND4F_7.Y.n3 mux8_4.NAND4F_7.Y.t9 308.481
R15495 mux8_4.NAND4F_7.Y.n1 mux8_4.NAND4F_7.Y.n4 187.373
R15496 mux8_4.NAND4F_7.Y.n1 mux8_4.NAND4F_7.Y.n5 187.192
R15497 mux8_4.NAND4F_7.Y.n1 mux8_4.NAND4F_7.Y.n6 187.192
R15498 mux8_4.NAND4F_7.Y.n0 mux8_4.NAND4F_7.Y.n7 187.192
R15499 mux8_4.NAND4F_7.Y mux8_4.NAND4F_7.Y.n3 161.492
R15500 mux8_4.NAND4F_7.Y.n3 mux8_4.NAND4F_7.Y.n2 27.752
R15501 mux8_4.NAND4F_7.Y mux8_4.NAND4F_7.Y.t2 23.5642
R15502 mux8_4.NAND4F_7.Y.n4 mux8_4.NAND4F_7.Y.t1 20.1899
R15503 mux8_4.NAND4F_7.Y.n4 mux8_4.NAND4F_7.Y.t0 20.1899
R15504 mux8_4.NAND4F_7.Y.n5 mux8_4.NAND4F_7.Y.t7 20.1899
R15505 mux8_4.NAND4F_7.Y.n5 mux8_4.NAND4F_7.Y.t8 20.1899
R15506 mux8_4.NAND4F_7.Y.n6 mux8_4.NAND4F_7.Y.t6 20.1899
R15507 mux8_4.NAND4F_7.Y.n6 mux8_4.NAND4F_7.Y.t5 20.1899
R15508 mux8_4.NAND4F_7.Y.n7 mux8_4.NAND4F_7.Y.t3 20.1899
R15509 mux8_4.NAND4F_7.Y.n7 mux8_4.NAND4F_7.Y.t4 20.1899
R15510 mux8_4.NAND4F_7.Y mux8_4.NAND4F_7.Y.n0 0.472662
R15511 mux8_4.NAND4F_7.Y.n0 mux8_4.NAND4F_7.Y.n1 0.358709
R15512 B4.n28 B4.t18 491.64
R15513 B4.n27 B4.t22 491.64
R15514 B4.n26 B4.t3 491.64
R15515 B4.n25 B4.t34 491.64
R15516 B4.n15 B4.t0 491.64
R15517 B4.n14 B4.t4 491.64
R15518 B4.n13 B4.t37 491.64
R15519 B4.n12 B4.t26 491.64
R15520 B4.n32 B4.t14 485.443
R15521 B4.n8 B4.t23 394.37
R15522 B4.n4 B4.t12 394.37
R15523 B4.n1 B4.t30 394.37
R15524 B4.n18 B4.t25 379.173
R15525 B4.n30 B4.t20 343.827
R15526 B4.n19 B4.t19 312.599
R15527 B4.n7 B4.t31 291.829
R15528 B4.n7 B4.t29 291.829
R15529 B4.n3 B4.t32 291.829
R15530 B4.n3 B4.t13 291.829
R15531 B4.n0 B4.t7 291.829
R15532 B4.n0 B4.t6 291.829
R15533 B4.n29 B4.t15 255.588
R15534 B4.n16 B4.t21 255.588
R15535 B4.n19 B4.t8 247.428
R15536 B4.n20 B4.t5 247.428
R15537 B4.n21 B4.t28 247.428
R15538 B4.n18 B4.t27 247.428
R15539 B4.n30 B4.t33 237.787
R15540 B4.n31 B4.t9 224.478
R15541 B4.n7 B4.t11 221.72
R15542 B4.n3 B4.t35 221.72
R15543 B4.n0 B4.t2 221.72
R15544 B4.n12 B4.n11 209.407
R15545 B4.n25 B4.n24 209.19
R15546 B4 B4.n22 162.139
R15547 B4.n24 B4.t10 139.78
R15548 B4.n24 B4.t16 139.78
R15549 B4.n24 B4.t24 139.78
R15550 B4.n11 B4.t1 139.78
R15551 B4.n11 B4.t17 139.78
R15552 B4.n11 B4.t36 139.78
R15553 B4.n32 B4.n31 83.8438
R15554 B4.n21 B4.n20 65.1723
R15555 B4.n20 B4.n19 65.1723
R15556 B4 B4.n32 61.0461
R15557 B4.n8 B4.n7 53.374
R15558 B4.n4 B4.n3 53.374
R15559 B4.n1 B4.n0 53.374
R15560 B4.n31 B4.n30 48.2005
R15561 B4.n34 B4 41.9747
R15562 B4.n22 B4.n21 33.2653
R15563 B4.n22 B4.n18 31.9075
R15564 B4 B4.n16 27.4136
R15565 B4.n27 B4.n26 17.8661
R15566 B4.n26 B4.n25 17.8661
R15567 B4.n13 B4.n12 17.8661
R15568 B4.n14 B4.n13 17.8661
R15569 B4.n28 B4.n27 17.1217
R15570 B4.n15 B4.n14 17.1217
R15571 B4.n6 B4.n2 14.4947
R15572 B4.n17 B4 12.626
R15573 B4.n10 B4.n9 12.4648
R15574 B4.n23 B4 12.4399
R15575 B4.n34 B4.n33 12.4105
R15576 B4.n6 B4.n5 12.4105
R15577 B4 B4.n29 11.1665
R15578 B4.n17 B4.n10 10.2068
R15579 B4.n23 B4.n17 8.35141
R15580 B4.n35 B4.n23 5.12664
R15581 B4.n10 B4.n6 2.82311
R15582 B4.n29 B4.n28 1.8615
R15583 B4.n16 B4.n15 1.8615
R15584 B4.n33 B4 1.27044
R15585 B4.n9 B4.n8 1.23221
R15586 B4.n2 B4.n1 0.748199
R15587 B4.n5 B4.n4 0.743681
R15588 B4.n5 B4 0.0750482
R15589 B4.n2 B4 0.0705301
R15590 B4.n9 B4 0.049413
R15591 B4.n33 B4 0.0393514
R15592 B4 B4.n35 0.0187778
R15593 B4.n35 B4 0.0165488
R15594 B4 B4.n34 0.00795122
R15595 a_n12345_n26161.n2 a_n12345_n26161.t7 539.788
R15596 a_n12345_n26161.n3 a_n12345_n26161.t5 531.496
R15597 a_n12345_n26161.n2 a_n12345_n26161.t3 490.034
R15598 a_n12345_n26161.n5 a_n12345_n26161.t0 283.788
R15599 a_n12345_n26161.t1 a_n12345_n26161.n5 205.489
R15600 a_n12345_n26161.n0 a_n12345_n26161.t4 182.625
R15601 a_n12345_n26161.n1 a_n12345_n26161.t2 179.054
R15602 a_n12345_n26161.n0 a_n12345_n26161.t6 139.78
R15603 a_n12345_n26161.n4 a_n12345_n26161.n1 101.368
R15604 a_n12345_n26161.n5 a_n12345_n26161.n4 77.9135
R15605 a_n12345_n26161.n4 a_n12345_n26161.n3 76.1557
R15606 a_n12345_n26161.n3 a_n12345_n26161.n2 8.29297
R15607 a_n12345_n26161.n1 a_n12345_n26161.n0 3.57087
R15608 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_0.B MULT_0.inv_8.Y.t12 540.38
R15609 MULT_0.inv_8.Y.n3 MULT_0.inv_8.Y.t5 491.64
R15610 MULT_0.inv_8.Y.n3 MULT_0.inv_8.Y.t11 491.64
R15611 MULT_0.inv_8.Y.n3 MULT_0.inv_8.Y.t4 491.64
R15612 MULT_0.inv_8.Y.n3 MULT_0.inv_8.Y.t9 491.64
R15613 MULT_0.inv_8.Y.n1 MULT_0.inv_8.Y.t13 367.928
R15614 MULT_0.inv_8.Y.n0 MULT_0.inv_8.Y.t3 256.514
R15615 MULT_0.inv_8.Y.n2 MULT_0.inv_8.Y.t7 227.356
R15616 MULT_0.inv_8.Y.n0 MULT_0.inv_8.Y.n7 226.136
R15617 MULT_0.inv_8.Y.n1 MULT_0.inv_8.Y.t10 213.688
R15618 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_0.B MULT_0.inv_8.Y.n5 162.867
R15619 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_0.B MULT_0.inv_8.Y.n2 160.439
R15620 MULT_0.inv_8.Y.n4 MULT_0.inv_8.Y.t14 139.78
R15621 MULT_0.inv_8.Y.n4 MULT_0.inv_8.Y.t6 139.78
R15622 MULT_0.inv_8.Y.n4 MULT_0.inv_8.Y.t15 139.78
R15623 MULT_0.inv_8.Y.n4 MULT_0.inv_8.Y.t8 139.78
R15624 MULT_0.inv_8.Y.n2 MULT_0.inv_8.Y.n1 94.4341
R15625 MULT_0.inv_8.Y.n0 MULT_0.inv_8.Y.t1 83.833
R15626 MULT_0.inv_8.Y.n5 MULT_0.inv_8.Y.n4 38.6833
R15627 MULT_0.inv_8.Y.n7 MULT_0.inv_8.Y.t0 30.379
R15628 MULT_0.inv_8.Y.n7 MULT_0.inv_8.Y.t2 30.379
R15629 MULT_0.inv_8.Y.n5 MULT_0.inv_8.Y.n3 28.3986
R15630 MULT_0.inv_8.Y.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.A 24.204
R15631 MULT_0.4bit_ADDER_2.FULL_ADDER_3.A MULT_0.inv_8.Y.n6 16.8273
R15632 MULT_0.inv_8.Y.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_0.B 9.00496
R15633 MULT_0.inv_8.Y.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_0.B 4.77555
R15634 a_n10684_n11063.n0 a_n10684_n11063.n2 81.2978
R15635 a_n10684_n11063.n0 a_n10684_n11063.n3 81.1637
R15636 a_n10684_n11063.n0 a_n10684_n11063.n4 81.1637
R15637 a_n10684_n11063.n1 a_n10684_n11063.n5 81.1637
R15638 a_n10684_n11063.n1 a_n10684_n11063.n6 81.1637
R15639 a_n10684_n11063.n7 a_n10684_n11063.n1 80.9213
R15640 a_n10684_n11063.n2 a_n10684_n11063.t8 11.8205
R15641 a_n10684_n11063.n2 a_n10684_n11063.t7 11.8205
R15642 a_n10684_n11063.n3 a_n10684_n11063.t2 11.8205
R15643 a_n10684_n11063.n3 a_n10684_n11063.t0 11.8205
R15644 a_n10684_n11063.n4 a_n10684_n11063.t1 11.8205
R15645 a_n10684_n11063.n4 a_n10684_n11063.t3 11.8205
R15646 a_n10684_n11063.n5 a_n10684_n11063.t10 11.8205
R15647 a_n10684_n11063.n5 a_n10684_n11063.t9 11.8205
R15648 a_n10684_n11063.n6 a_n10684_n11063.t4 11.8205
R15649 a_n10684_n11063.n6 a_n10684_n11063.t11 11.8205
R15650 a_n10684_n11063.n7 a_n10684_n11063.t5 11.8205
R15651 a_n10684_n11063.t6 a_n10684_n11063.n7 11.8205
R15652 a_n10684_n11063.n1 a_n10684_n11063.n0 0.402735
R15653 B6.n6 B6.t4 491.64
R15654 B6.n5 B6.t24 491.64
R15655 B6.n4 B6.t7 491.64
R15656 B6.n3 B6.t32 491.64
R15657 B6.n23 B6.t13 491.64
R15658 B6.n22 B6.t21 491.64
R15659 B6.n21 B6.t12 491.64
R15660 B6.n20 B6.t31 491.64
R15661 B6.n10 B6.t0 485.443
R15662 B6.n27 B6.t8 394.37
R15663 B6.n31 B6.t19 394.37
R15664 B6.n1 B6.t30 394.37
R15665 B6.n13 B6.t9 379.173
R15666 B6.n8 B6.t15 343.827
R15667 B6.n14 B6.t33 312.599
R15668 B6.n26 B6.t16 291.829
R15669 B6.n26 B6.t27 291.829
R15670 B6.n30 B6.t37 291.829
R15671 B6.n30 B6.t20 291.829
R15672 B6.n0 B6.t6 291.829
R15673 B6.n0 B6.t5 291.829
R15674 B6.n7 B6.t36 255.588
R15675 B6.n24 B6.t28 255.588
R15676 B6.n14 B6.t23 247.428
R15677 B6.n15 B6.t22 247.428
R15678 B6.n16 B6.t14 247.428
R15679 B6.n13 B6.t11 247.428
R15680 B6.n8 B6.t25 237.787
R15681 B6.n9 B6.t34 224.478
R15682 B6.n26 B6.t29 221.72
R15683 B6.n30 B6.t3 221.72
R15684 B6.n0 B6.t2 221.72
R15685 B6.n20 B6.n19 209.407
R15686 B6.n3 B6.n2 209.19
R15687 B6 B6.n17 162.139
R15688 B6.n2 B6.t18 139.78
R15689 B6.n2 B6.t26 139.78
R15690 B6.n2 B6.t10 139.78
R15691 B6.n19 B6.t1 139.78
R15692 B6.n19 B6.t17 139.78
R15693 B6.n19 B6.t35 139.78
R15694 B6.n10 B6.n9 83.8438
R15695 B6.n16 B6.n15 65.1723
R15696 B6.n15 B6.n14 65.1723
R15697 B6 B6.n10 61.0461
R15698 B6.n27 B6.n26 53.374
R15699 B6.n31 B6.n30 53.374
R15700 B6.n1 B6.n0 53.374
R15701 B6.n9 B6.n8 48.2005
R15702 B6.n17 B6.n16 33.2653
R15703 B6.n17 B6.n13 31.9075
R15704 B6 B6.n24 27.4136
R15705 B6.n5 B6.n4 17.8661
R15706 B6.n4 B6.n3 17.8661
R15707 B6.n21 B6.n20 17.8661
R15708 B6.n22 B6.n21 17.8661
R15709 B6.n6 B6.n5 17.1217
R15710 B6.n23 B6.n22 17.1217
R15711 B6.n34 B6.n33 14.1821
R15712 B6.n25 B6 12.5928
R15713 B6.n29 B6.n28 12.5228
R15714 B6.n18 B6 12.4904
R15715 B6.n12 B6.n11 12.4105
R15716 B6.n33 B6.n32 12.4105
R15717 B6.n29 B6.n25 11.4059
R15718 B6 B6.n7 11.1665
R15719 B6.n25 B6.n18 8.56599
R15720 B6.n18 B6.n12 5.19596
R15721 B6.n33 B6.n29 2.82994
R15722 B6.n7 B6.n6 1.8615
R15723 B6.n24 B6.n23 1.8615
R15724 B6.n11 B6 1.249
R15725 B6.n28 B6.n27 1.20685
R15726 B6.n34 B6.n1 0.767025
R15727 B6.n32 B6.n31 0.765519
R15728 B6.n11 B6 0.116819
R15729 B6.n32 B6 0.0532108
R15730 B6.n28 B6 0.0530362
R15731 B6 B6.n34 0.0517048
R15732 B6.n12 B6 0.0148293
R15733 a_n23960_n22530.t0 a_n23960_n22530.t1 19.8005
R15734 a_n14155_n5154.n0 a_n14155_n5154.t6 539.788
R15735 a_n14155_n5154.n1 a_n14155_n5154.t3 531.496
R15736 a_n14155_n5154.n0 a_n14155_n5154.t7 490.034
R15737 a_n14155_n5154.n5 a_n14155_n5154.t0 283.788
R15738 a_n14155_n5154.t1 a_n14155_n5154.n5 205.489
R15739 a_n14155_n5154.n2 a_n14155_n5154.t4 182.625
R15740 a_n14155_n5154.n3 a_n14155_n5154.t2 179.054
R15741 a_n14155_n5154.n2 a_n14155_n5154.t5 139.78
R15742 a_n14155_n5154.n4 a_n14155_n5154.n3 101.368
R15743 a_n14155_n5154.n5 a_n14155_n5154.n4 77.9135
R15744 a_n14155_n5154.n4 a_n14155_n5154.n1 76.1557
R15745 a_n14155_n5154.n1 a_n14155_n5154.n0 8.29297
R15746 a_n14155_n5154.n3 a_n14155_n5154.n2 3.57087
R15747 a_n13975_n5154.n2 a_n13975_n5154.n1 121.353
R15748 a_n13975_n5154.n3 a_n13975_n5154.n2 121.001
R15749 a_n13975_n5154.n2 a_n13975_n5154.n0 120.977
R15750 a_n13975_n5154.n1 a_n13975_n5154.t2 30.462
R15751 a_n13975_n5154.n1 a_n13975_n5154.t1 30.462
R15752 a_n13975_n5154.n0 a_n13975_n5154.t4 30.462
R15753 a_n13975_n5154.n0 a_n13975_n5154.t3 30.462
R15754 a_n13975_n5154.n3 a_n13975_n5154.t5 30.462
R15755 a_n13975_n5154.t0 a_n13975_n5154.n3 30.462
R15756 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t18 491.64
R15757 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t23 491.64
R15758 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t12 491.64
R15759 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t19 491.64
R15760 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n8 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t22 485.221
R15761 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t13 367.928
R15762 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t16 255.588
R15763 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t20 224.478
R15764 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t14 213.688
R15765 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n0 209.19
R15766 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t17 139.78
R15767 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t15 139.78
R15768 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t21 139.78
R15769 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n11 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n10 120.999
R15770 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n11 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n9 120.999
R15771 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n23 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n22 104.489
R15772 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n13 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n12 92.5005
R15773 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n20 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n18 86.2638
R15774 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n18 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n17 85.8873
R15775 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n18 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n15 85.724
R15776 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n8 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n7 84.5046
R15777 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n23 83.8907
R15778 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n21 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n20 75.0672
R15779 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n21 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n17 75.0672
R15780 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n20 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n19 73.1255
R15781 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n15 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n14 73.1255
R15782 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n17 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n16 73.1255
R15783 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n6 72.3005
R15784 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n22 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n15 68.8946
R15785 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n8 60.9797
R15786 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n23 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n13 41.9827
R15787 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n12 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t2 30.462
R15788 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n12 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t10 30.462
R15789 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n10 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t9 30.462
R15790 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n10 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t11 30.462
R15791 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n9 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t0 30.462
R15792 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n9 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t1 30.462
R15793 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n13 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n11 28.124
R15794 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n5 19.963
R15795 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n1 17.8661
R15796 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n2 17.8661
R15797 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n3 17.1217
R15798 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n14 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t5 11.8205
R15799 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n14 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t7 11.8205
R15800 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n19 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t6 11.8205
R15801 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n19 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t8 11.8205
R15802 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n16 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t3 11.8205
R15803 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n16 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t4 11.8205
R15804 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n22 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n21 9.3005
R15805 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n4 1.8615
R15806 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n9 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t16 540.38
R15807 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t9 491.64
R15808 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t14 491.64
R15809 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t13 491.64
R15810 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t17 491.64
R15811 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t8 367.928
R15812 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n2 227.526
R15813 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n8 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t10 227.356
R15814 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n1 227.266
R15815 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n3 227.266
R15816 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t11 213.688
R15817 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n6 162.852
R15818 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n9 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n8 160.439
R15819 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t18 139.78
R15820 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t12 139.78
R15821 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t15 139.78
R15822 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t7 139.78
R15823 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n8 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n7 94.4341
R15824 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t0 42.7831
R15825 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n5 38.6833
R15826 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t5 30.379
R15827 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t6 30.379
R15828 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t2 30.379
R15829 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t1 30.379
R15830 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t3 30.379
R15831 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t4 30.379
R15832 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n4 28.3986
R15833 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n0 18.8832
R15834 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n10 10.7052
R15835 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n10 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT 5.09176
R15836 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n10 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT 4.19292
R15837 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n9 0.794268
R15838 a_n4205_3810.n0 a_n4205_3810.n4 81.3236
R15839 a_n4205_3810.n0 a_n4205_3810.n1 81.2978
R15840 a_n4205_3810.n0 a_n4205_3810.n5 81.1637
R15841 a_n4205_3810.n0 a_n4205_3810.n3 81.1637
R15842 a_n4205_3810.n0 a_n4205_3810.n2 81.1637
R15843 a_n4205_3810.n6 a_n4205_3810.n0 81.1637
R15844 a_n4205_3810.n4 a_n4205_3810.t8 11.8205
R15845 a_n4205_3810.n4 a_n4205_3810.t7 11.8205
R15846 a_n4205_3810.n5 a_n4205_3810.t2 11.8205
R15847 a_n4205_3810.n5 a_n4205_3810.t6 11.8205
R15848 a_n4205_3810.n3 a_n4205_3810.t3 11.8205
R15849 a_n4205_3810.n3 a_n4205_3810.t5 11.8205
R15850 a_n4205_3810.n2 a_n4205_3810.t9 11.8205
R15851 a_n4205_3810.n2 a_n4205_3810.t4 11.8205
R15852 a_n4205_3810.n1 a_n4205_3810.t11 11.8205
R15853 a_n4205_3810.n1 a_n4205_3810.t10 11.8205
R15854 a_n4205_3810.t0 a_n4205_3810.n6 11.8205
R15855 a_n4205_3810.n6 a_n4205_3810.t1 11.8205
R15856 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t18 491.64
R15857 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t17 491.64
R15858 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t22 491.64
R15859 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t23 491.64
R15860 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t16 485.221
R15861 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t13 367.928
R15862 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t20 255.588
R15863 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t14 224.478
R15864 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t12 213.688
R15865 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n18 209.19
R15866 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t21 139.78
R15867 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t15 139.78
R15868 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t19 139.78
R15869 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n1 120.999
R15870 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n0 120.999
R15871 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n13 104.489
R15872 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 103.258
R15873 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n3 92.5005
R15874 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n8 86.2638
R15875 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n9 85.8873
R15876 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n6 85.724
R15877 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n16 84.5046
R15878 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n14 84.0545
R15879 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n8 75.0672
R15880 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n11 75.0672
R15881 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n6 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n5 73.1255
R15882 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n8 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n7 73.1255
R15883 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n10 73.1255
R15884 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n15 72.3005
R15885 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n6 68.8946
R15886 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n17 60.9816
R15887 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n4 41.9827
R15888 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t7 30.462
R15889 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t10 30.462
R15890 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t9 30.462
R15891 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t11 30.462
R15892 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t5 30.462
R15893 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t3 30.462
R15894 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n2 28.124
R15895 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n19 17.8661
R15896 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n20 17.8661
R15897 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n21 17.1217
R15898 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n23 15.6329
R15899 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t6 11.8205
R15900 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t4 11.8205
R15901 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t8 11.8205
R15902 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t0 11.8205
R15903 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t1 11.8205
R15904 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t2 11.8205
R15905 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 10.8165
R15906 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n12 9.3005
R15907 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n24 2.50602
R15908 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n22 1.8615
R15909 a_n11274_n25843.n2 a_n11274_n25843.n0 121.353
R15910 a_n11274_n25843.n2 a_n11274_n25843.n1 121.353
R15911 a_n11274_n25843.n3 a_n11274_n25843.n2 121.001
R15912 a_n11274_n25843.n0 a_n11274_n25843.t3 30.462
R15913 a_n11274_n25843.n0 a_n11274_n25843.t4 30.462
R15914 a_n11274_n25843.n1 a_n11274_n25843.t2 30.462
R15915 a_n11274_n25843.n1 a_n11274_n25843.t1 30.462
R15916 a_n11274_n25843.n3 a_n11274_n25843.t5 30.462
R15917 a_n11274_n25843.t0 a_n11274_n25843.n3 30.462
R15918 XOR8_0.S4.n0 XOR8_0.S4.t12 1032.02
R15919 XOR8_0.S4.n0 XOR8_0.S4.t13 336.962
R15920 XOR8_0.S4.n0 XOR8_0.S4.t14 326.154
R15921 XOR8_0.S4 XOR8_0.S4.n0 162.946
R15922 XOR8_0.S4.n3 XOR8_0.S4.n1 120.999
R15923 XOR8_0.S4.n3 XOR8_0.S4.n2 120.999
R15924 XOR8_0.S4.n15 XOR8_0.S4.n14 104.865
R15925 XOR8_0.S4.n5 XOR8_0.S4.n4 92.5005
R15926 XOR8_0.S4.n12 XOR8_0.S4.n10 86.2638
R15927 XOR8_0.S4.n10 XOR8_0.S4.n9 85.8873
R15928 XOR8_0.S4.n10 XOR8_0.S4.n7 85.724
R15929 XOR8_0.S4 XOR8_0.S4.n15 83.8907
R15930 XOR8_0.S4.n13 XOR8_0.S4.n12 75.0672
R15931 XOR8_0.S4.n13 XOR8_0.S4.n9 75.0672
R15932 XOR8_0.S4.n7 XOR8_0.S4.n6 73.1255
R15933 XOR8_0.S4.n12 XOR8_0.S4.n11 73.1255
R15934 XOR8_0.S4.n9 XOR8_0.S4.n8 73.1255
R15935 XOR8_0.S4.n14 XOR8_0.S4.n7 68.5181
R15936 XOR8_0.S4.n15 XOR8_0.S4.n5 41.9827
R15937 XOR8_0.S4.n4 XOR8_0.S4.t4 30.462
R15938 XOR8_0.S4.n4 XOR8_0.S4.t10 30.462
R15939 XOR8_0.S4.n1 XOR8_0.S4.t3 30.462
R15940 XOR8_0.S4.n1 XOR8_0.S4.t5 30.462
R15941 XOR8_0.S4.n2 XOR8_0.S4.t9 30.462
R15942 XOR8_0.S4.n2 XOR8_0.S4.t11 30.462
R15943 XOR8_0.S4.n5 XOR8_0.S4.n3 28.124
R15944 XOR8_0.S4.n11 XOR8_0.S4.t8 11.8205
R15945 XOR8_0.S4.n11 XOR8_0.S4.t7 11.8205
R15946 XOR8_0.S4.n6 XOR8_0.S4.t2 11.8205
R15947 XOR8_0.S4.n6 XOR8_0.S4.t6 11.8205
R15948 XOR8_0.S4.n8 XOR8_0.S4.t0 11.8205
R15949 XOR8_0.S4.n8 XOR8_0.S4.t1 11.8205
R15950 XOR8_0.S4.n14 XOR8_0.S4.n13 9.3005
R15951 a_5167_4886.n2 a_5167_4886.t2 541.395
R15952 a_5167_4886.n3 a_5167_4886.t4 527.402
R15953 a_5167_4886.n2 a_5167_4886.t6 491.64
R15954 a_5167_4886.n5 a_5167_4886.t1 281.906
R15955 a_5167_4886.t0 a_5167_4886.n5 204.359
R15956 a_5167_4886.n0 a_5167_4886.t7 180.73
R15957 a_5167_4886.n1 a_5167_4886.t5 179.45
R15958 a_5167_4886.n0 a_5167_4886.t3 139.78
R15959 a_5167_4886.n4 a_5167_4886.n1 105.635
R15960 a_5167_4886.n4 a_5167_4886.n3 76.0005
R15961 a_5167_4886.n5 a_5167_4886.n4 67.9685
R15962 a_5167_4886.n3 a_5167_4886.n2 13.994
R15963 a_5167_4886.n1 a_5167_4886.n0 1.28015
R15964 V_FLAG_0.XOR2_0.Y.n2 V_FLAG_0.XOR2_0.Y.t13 485.221
R15965 V_FLAG_0.XOR2_0.Y.n0 V_FLAG_0.XOR2_0.Y.t14 367.928
R15966 V_FLAG_0.XOR2_0.Y.n1 V_FLAG_0.XOR2_0.Y.t12 224.478
R15967 V_FLAG_0.XOR2_0.Y.n0 V_FLAG_0.XOR2_0.Y.t15 213.688
R15968 V_FLAG_0.XOR2_0.Y.n5 V_FLAG_0.XOR2_0.Y.n4 120.999
R15969 V_FLAG_0.XOR2_0.Y.n5 V_FLAG_0.XOR2_0.Y.n3 120.999
R15970 V_FLAG_0.XOR2_0.Y.n17 V_FLAG_0.XOR2_0.Y.n16 104.489
R15971 V_FLAG_0.XOR2_0.Y.n7 V_FLAG_0.XOR2_0.Y.n6 92.5005
R15972 V_FLAG_0.XOR2_0.Y.n14 V_FLAG_0.XOR2_0.Y.n12 86.2638
R15973 V_FLAG_0.XOR2_0.Y.n12 V_FLAG_0.XOR2_0.Y.n11 85.8873
R15974 V_FLAG_0.XOR2_0.Y.n12 V_FLAG_0.XOR2_0.Y.n9 85.724
R15975 V_FLAG_0.XOR2_0.Y.n2 V_FLAG_0.XOR2_0.Y.n1 84.5046
R15976 V_FLAG_0.XOR2_0.Y V_FLAG_0.XOR2_0.Y.n17 83.8907
R15977 V_FLAG_0.XOR2_0.Y.n15 V_FLAG_0.XOR2_0.Y.n11 75.0672
R15978 V_FLAG_0.XOR2_0.Y.n15 V_FLAG_0.XOR2_0.Y.n14 75.0672
R15979 V_FLAG_0.XOR2_0.Y.n9 V_FLAG_0.XOR2_0.Y.n8 73.1255
R15980 V_FLAG_0.XOR2_0.Y.n11 V_FLAG_0.XOR2_0.Y.n10 73.1255
R15981 V_FLAG_0.XOR2_0.Y.n14 V_FLAG_0.XOR2_0.Y.n13 73.1255
R15982 V_FLAG_0.XOR2_0.Y.n1 V_FLAG_0.XOR2_0.Y.n0 72.3005
R15983 V_FLAG_0.XOR2_0.Y.n16 V_FLAG_0.XOR2_0.Y.n9 68.8946
R15984 V_FLAG_0.XOR2_0.Y V_FLAG_0.XOR2_0.Y.n2 61.5676
R15985 V_FLAG_0.XOR2_0.Y.n17 V_FLAG_0.XOR2_0.Y.n7 41.9827
R15986 V_FLAG_0.XOR2_0.Y.n6 V_FLAG_0.XOR2_0.Y.t10 30.462
R15987 V_FLAG_0.XOR2_0.Y.n6 V_FLAG_0.XOR2_0.Y.t2 30.462
R15988 V_FLAG_0.XOR2_0.Y.n4 V_FLAG_0.XOR2_0.Y.t5 30.462
R15989 V_FLAG_0.XOR2_0.Y.n4 V_FLAG_0.XOR2_0.Y.t0 30.462
R15990 V_FLAG_0.XOR2_0.Y.n3 V_FLAG_0.XOR2_0.Y.t11 30.462
R15991 V_FLAG_0.XOR2_0.Y.n3 V_FLAG_0.XOR2_0.Y.t6 30.462
R15992 V_FLAG_0.XOR2_0.Y.n7 V_FLAG_0.XOR2_0.Y.n5 28.124
R15993 V_FLAG_0.XOR2_0.Y.n10 V_FLAG_0.XOR2_0.Y.t8 11.8205
R15994 V_FLAG_0.XOR2_0.Y.n10 V_FLAG_0.XOR2_0.Y.t7 11.8205
R15995 V_FLAG_0.XOR2_0.Y.n8 V_FLAG_0.XOR2_0.Y.t9 11.8205
R15996 V_FLAG_0.XOR2_0.Y.n8 V_FLAG_0.XOR2_0.Y.t4 11.8205
R15997 V_FLAG_0.XOR2_0.Y.n13 V_FLAG_0.XOR2_0.Y.t1 11.8205
R15998 V_FLAG_0.XOR2_0.Y.n13 V_FLAG_0.XOR2_0.Y.t3 11.8205
R15999 V_FLAG_0.XOR2_0.Y.n16 V_FLAG_0.XOR2_0.Y.n15 9.3005
R16000 a_5197_5532.n0 a_5197_5532.n4 81.2978
R16001 a_5197_5532.n0 a_5197_5532.n5 81.1637
R16002 a_5197_5532.n0 a_5197_5532.n6 81.1637
R16003 a_5197_5532.n1 a_5197_5532.n3 81.1637
R16004 a_5197_5532.n7 a_5197_5532.n1 81.1637
R16005 a_5197_5532.n1 a_5197_5532.n2 80.9213
R16006 a_5197_5532.n4 a_5197_5532.t10 11.8205
R16007 a_5197_5532.n4 a_5197_5532.t11 11.8205
R16008 a_5197_5532.n5 a_5197_5532.t1 11.8205
R16009 a_5197_5532.n5 a_5197_5532.t3 11.8205
R16010 a_5197_5532.n6 a_5197_5532.t2 11.8205
R16011 a_5197_5532.n6 a_5197_5532.t0 11.8205
R16012 a_5197_5532.n3 a_5197_5532.t7 11.8205
R16013 a_5197_5532.n3 a_5197_5532.t5 11.8205
R16014 a_5197_5532.n2 a_5197_5532.t8 11.8205
R16015 a_5197_5532.n2 a_5197_5532.t9 11.8205
R16016 a_5197_5532.n7 a_5197_5532.t4 11.8205
R16017 a_5197_5532.t6 a_5197_5532.n7 11.8205
R16018 a_5197_5532.n1 a_5197_5532.n0 0.402735
R16019 NOT8_0.S5.n1 NOT8_0.S5.t4 1032.02
R16020 NOT8_0.S5.n1 NOT8_0.S5.t5 336.962
R16021 NOT8_0.S5.n1 NOT8_0.S5.t6 326.154
R16022 NOT8_0.S5.n0 NOT8_0.S5.t3 256.514
R16023 NOT8_0.S5.n0 NOT8_0.S5.n2 226.258
R16024 NOT8_0.S5 NOT8_0.S5.n1 162.952
R16025 NOT8_0.S5.n0 NOT8_0.S5.t1 83.7172
R16026 NOT8_0.S5.n2 NOT8_0.S5.t0 30.379
R16027 NOT8_0.S5.n2 NOT8_0.S5.t2 30.379
R16028 NOT8_0.S5 NOT8_0.S5.n0 1.9182
R16029 a_10459_n26405.t0 a_10459_n26405.t1 9.9005
R16030 mux8_7.NAND4F_7.Y.n2 mux8_7.NAND4F_7.Y.t11 1388.16
R16031 mux8_7.NAND4F_7.Y.n2 mux8_7.NAND4F_7.Y.t10 350.839
R16032 mux8_7.NAND4F_7.Y.n3 mux8_7.NAND4F_7.Y.t9 308.481
R16033 mux8_7.NAND4F_7.Y.n1 mux8_7.NAND4F_7.Y.n4 187.373
R16034 mux8_7.NAND4F_7.Y.n1 mux8_7.NAND4F_7.Y.n5 187.192
R16035 mux8_7.NAND4F_7.Y.n1 mux8_7.NAND4F_7.Y.n6 187.192
R16036 mux8_7.NAND4F_7.Y.n0 mux8_7.NAND4F_7.Y.n7 187.192
R16037 mux8_7.NAND4F_7.Y mux8_7.NAND4F_7.Y.n3 161.492
R16038 mux8_7.NAND4F_7.Y.n3 mux8_7.NAND4F_7.Y.n2 27.752
R16039 mux8_7.NAND4F_7.Y mux8_7.NAND4F_7.Y.t4 23.5642
R16040 mux8_7.NAND4F_7.Y.n4 mux8_7.NAND4F_7.Y.t1 20.1899
R16041 mux8_7.NAND4F_7.Y.n4 mux8_7.NAND4F_7.Y.t0 20.1899
R16042 mux8_7.NAND4F_7.Y.n5 mux8_7.NAND4F_7.Y.t2 20.1899
R16043 mux8_7.NAND4F_7.Y.n5 mux8_7.NAND4F_7.Y.t3 20.1899
R16044 mux8_7.NAND4F_7.Y.n6 mux8_7.NAND4F_7.Y.t8 20.1899
R16045 mux8_7.NAND4F_7.Y.n6 mux8_7.NAND4F_7.Y.t7 20.1899
R16046 mux8_7.NAND4F_7.Y.n7 mux8_7.NAND4F_7.Y.t6 20.1899
R16047 mux8_7.NAND4F_7.Y.n7 mux8_7.NAND4F_7.Y.t5 20.1899
R16048 mux8_7.NAND4F_7.Y mux8_7.NAND4F_7.Y.n0 0.472662
R16049 mux8_7.NAND4F_7.Y.n0 mux8_7.NAND4F_7.Y.n1 0.358709
R16050 a_n12345_n23393.n2 a_n12345_n23393.t3 539.788
R16051 a_n12345_n23393.n3 a_n12345_n23393.t7 531.496
R16052 a_n12345_n23393.n2 a_n12345_n23393.t5 490.034
R16053 a_n12345_n23393.n5 a_n12345_n23393.t0 283.788
R16054 a_n12345_n23393.t1 a_n12345_n23393.n5 205.489
R16055 a_n12345_n23393.n0 a_n12345_n23393.t6 182.625
R16056 a_n12345_n23393.n1 a_n12345_n23393.t4 179.054
R16057 a_n12345_n23393.n0 a_n12345_n23393.t2 139.78
R16058 a_n12345_n23393.n4 a_n12345_n23393.n1 101.368
R16059 a_n12345_n23393.n5 a_n12345_n23393.n4 77.9135
R16060 a_n12345_n23393.n4 a_n12345_n23393.n3 76.1557
R16061 a_n12345_n23393.n3 a_n12345_n23393.n2 8.29297
R16062 a_n12345_n23393.n1 a_n12345_n23393.n0 3.57087
R16063 XOR8_0.S3.n0 XOR8_0.S3.t12 1032.02
R16064 XOR8_0.S3.n0 XOR8_0.S3.t13 336.962
R16065 XOR8_0.S3.n0 XOR8_0.S3.t14 326.154
R16066 XOR8_0.S3 XOR8_0.S3.n0 162.946
R16067 XOR8_0.S3.n3 XOR8_0.S3.n1 120.999
R16068 XOR8_0.S3.n3 XOR8_0.S3.n2 120.999
R16069 XOR8_0.S3.n15 XOR8_0.S3.n14 104.865
R16070 XOR8_0.S3.n5 XOR8_0.S3.n4 92.5005
R16071 XOR8_0.S3.n12 XOR8_0.S3.n10 86.2638
R16072 XOR8_0.S3.n10 XOR8_0.S3.n9 85.8873
R16073 XOR8_0.S3.n10 XOR8_0.S3.n7 85.724
R16074 XOR8_0.S3 XOR8_0.S3.n15 83.8907
R16075 XOR8_0.S3.n13 XOR8_0.S3.n9 75.0672
R16076 XOR8_0.S3.n13 XOR8_0.S3.n12 75.0672
R16077 XOR8_0.S3.n9 XOR8_0.S3.n8 73.1255
R16078 XOR8_0.S3.n7 XOR8_0.S3.n6 73.1255
R16079 XOR8_0.S3.n12 XOR8_0.S3.n11 73.1255
R16080 XOR8_0.S3.n14 XOR8_0.S3.n7 68.5181
R16081 XOR8_0.S3.n15 XOR8_0.S3.n5 41.9827
R16082 XOR8_0.S3.n4 XOR8_0.S3.t8 30.462
R16083 XOR8_0.S3.n4 XOR8_0.S3.t0 30.462
R16084 XOR8_0.S3.n1 XOR8_0.S3.t6 30.462
R16085 XOR8_0.S3.n1 XOR8_0.S3.t7 30.462
R16086 XOR8_0.S3.n2 XOR8_0.S3.t4 30.462
R16087 XOR8_0.S3.n2 XOR8_0.S3.t5 30.462
R16088 XOR8_0.S3.n5 XOR8_0.S3.n3 28.124
R16089 XOR8_0.S3.n6 XOR8_0.S3.t9 11.8205
R16090 XOR8_0.S3.n6 XOR8_0.S3.t3 11.8205
R16091 XOR8_0.S3.n8 XOR8_0.S3.t10 11.8205
R16092 XOR8_0.S3.n8 XOR8_0.S3.t11 11.8205
R16093 XOR8_0.S3.n11 XOR8_0.S3.t2 11.8205
R16094 XOR8_0.S3.n11 XOR8_0.S3.t1 11.8205
R16095 XOR8_0.S3.n14 XOR8_0.S3.n13 9.3005
R16096 a_n11274_n23651.n2 a_n11274_n23651.n0 121.353
R16097 a_n11274_n23651.n2 a_n11274_n23651.n1 121.001
R16098 a_n11274_n23651.n3 a_n11274_n23651.n2 120.977
R16099 a_n11274_n23651.n1 a_n11274_n23651.t1 30.462
R16100 a_n11274_n23651.n1 a_n11274_n23651.t4 30.462
R16101 a_n11274_n23651.n0 a_n11274_n23651.t5 30.462
R16102 a_n11274_n23651.n0 a_n11274_n23651.t3 30.462
R16103 a_n11274_n23651.n3 a_n11274_n23651.t0 30.462
R16104 a_n11274_n23651.t2 a_n11274_n23651.n3 30.462
R16105 mux8_2.NAND4F_8.Y.n1 mux8_2.NAND4F_8.Y.t14 379.173
R16106 mux8_2.NAND4F_8.Y.n2 mux8_2.NAND4F_8.Y.t9 312.599
R16107 mux8_2.NAND4F_8.Y.n1 mux8_2.NAND4F_8.Y.t13 247.428
R16108 mux8_2.NAND4F_8.Y.n4 mux8_2.NAND4F_8.Y.t12 247.428
R16109 mux8_2.NAND4F_8.Y.n3 mux8_2.NAND4F_8.Y.t11 247.428
R16110 mux8_2.NAND4F_8.Y.n2 mux8_2.NAND4F_8.Y.t10 247.428
R16111 mux8_2.NAND4F_8.Y.n0 mux8_2.NAND4F_8.Y.n6 187.373
R16112 mux8_2.NAND4F_8.Y.n0 mux8_2.NAND4F_8.Y.n7 187.192
R16113 mux8_2.NAND4F_8.Y.n0 mux8_2.NAND4F_8.Y.n8 187.192
R16114 mux8_2.NAND4F_8.Y.n10 mux8_2.NAND4F_8.Y.n9 187.192
R16115 mux8_2.NAND4F_8.Y mux8_2.NAND4F_8.Y.n5 162.139
R16116 mux8_2.NAND4F_8.Y.n4 mux8_2.NAND4F_8.Y.n3 65.1723
R16117 mux8_2.NAND4F_8.Y.n3 mux8_2.NAND4F_8.Y.n2 65.1723
R16118 mux8_2.NAND4F_8.Y.n5 mux8_2.NAND4F_8.Y.n4 33.2653
R16119 mux8_2.NAND4F_8.Y.n5 mux8_2.NAND4F_8.Y.n1 31.9075
R16120 mux8_2.NAND4F_8.Y mux8_2.NAND4F_8.Y.t3 22.6141
R16121 mux8_2.NAND4F_8.Y.n6 mux8_2.NAND4F_8.Y.t5 20.1899
R16122 mux8_2.NAND4F_8.Y.n6 mux8_2.NAND4F_8.Y.t4 20.1899
R16123 mux8_2.NAND4F_8.Y.n7 mux8_2.NAND4F_8.Y.t8 20.1899
R16124 mux8_2.NAND4F_8.Y.n7 mux8_2.NAND4F_8.Y.t0 20.1899
R16125 mux8_2.NAND4F_8.Y.n8 mux8_2.NAND4F_8.Y.t7 20.1899
R16126 mux8_2.NAND4F_8.Y.n8 mux8_2.NAND4F_8.Y.t6 20.1899
R16127 mux8_2.NAND4F_8.Y.n9 mux8_2.NAND4F_8.Y.t2 20.1899
R16128 mux8_2.NAND4F_8.Y.n9 mux8_2.NAND4F_8.Y.t1 20.1899
R16129 mux8_2.NAND4F_8.Y mux8_2.NAND4F_8.Y.n10 0.452586
R16130 mux8_2.NAND4F_8.Y.n10 mux8_2.NAND4F_8.Y.n0 0.358709
R16131 MULT_0.4bit_ADDER_1.A2 MULT_0.4bit_ADDER_1.A2.t8 540.38
R16132 MULT_0.4bit_ADDER_1.A2.n4 MULT_0.4bit_ADDER_1.A2.t7 491.64
R16133 MULT_0.4bit_ADDER_1.A2.n4 MULT_0.4bit_ADDER_1.A2.t12 491.64
R16134 MULT_0.4bit_ADDER_1.A2.n4 MULT_0.4bit_ADDER_1.A2.t10 491.64
R16135 MULT_0.4bit_ADDER_1.A2.n4 MULT_0.4bit_ADDER_1.A2.t13 491.64
R16136 MULT_0.4bit_ADDER_1.A2.n2 MULT_0.4bit_ADDER_1.A2.t9 367.928
R16137 MULT_0.4bit_ADDER_1.A2.n0 MULT_0.4bit_ADDER_1.A2.t3 256.529
R16138 MULT_0.4bit_ADDER_1.A2.n3 MULT_0.4bit_ADDER_1.A2.t15 227.356
R16139 MULT_0.4bit_ADDER_1.A2.n0 MULT_0.4bit_ADDER_1.A2.n1 226.292
R16140 MULT_0.4bit_ADDER_1.A2.n2 MULT_0.4bit_ADDER_1.A2.t11 213.688
R16141 MULT_0.4bit_ADDER_1.A2 MULT_0.4bit_ADDER_1.A2.n6 162.867
R16142 MULT_0.4bit_ADDER_1.A2 MULT_0.4bit_ADDER_1.A2.n3 160.439
R16143 MULT_0.4bit_ADDER_1.A2.n5 MULT_0.4bit_ADDER_1.A2.t4 139.78
R16144 MULT_0.4bit_ADDER_1.A2.n5 MULT_0.4bit_ADDER_1.A2.t6 139.78
R16145 MULT_0.4bit_ADDER_1.A2.n5 MULT_0.4bit_ADDER_1.A2.t14 139.78
R16146 MULT_0.4bit_ADDER_1.A2.n5 MULT_0.4bit_ADDER_1.A2.t5 139.78
R16147 MULT_0.4bit_ADDER_1.A2.n3 MULT_0.4bit_ADDER_1.A2.n2 94.4341
R16148 MULT_0.4bit_ADDER_1.A2.n0 MULT_0.4bit_ADDER_1.A2.t0 83.7616
R16149 MULT_0.4bit_ADDER_1.A2.n6 MULT_0.4bit_ADDER_1.A2.n5 38.6833
R16150 MULT_0.4bit_ADDER_1.A2.n1 MULT_0.4bit_ADDER_1.A2.t1 30.379
R16151 MULT_0.4bit_ADDER_1.A2.n1 MULT_0.4bit_ADDER_1.A2.t2 30.379
R16152 MULT_0.4bit_ADDER_1.A2.n6 MULT_0.4bit_ADDER_1.A2.n4 28.3986
R16153 MULT_0.4bit_ADDER_1.A2 MULT_0.4bit_ADDER_1.A2.n7 16.8169
R16154 MULT_0.4bit_ADDER_1.A2 MULT_0.4bit_ADDER_1.A2.n0 15.5384
R16155 MULT_0.4bit_ADDER_1.A2.n7 MULT_0.4bit_ADDER_1.A2 9.00496
R16156 MULT_0.4bit_ADDER_1.A2.n7 MULT_0.4bit_ADDER_1.A2 4.77555
R16157 a_n16690_n8419.n2 a_n16690_n8419.n1 121.353
R16158 a_n16690_n8419.n2 a_n16690_n8419.n0 121.353
R16159 a_n16690_n8419.n3 a_n16690_n8419.n2 121.001
R16160 a_n16690_n8419.n1 a_n16690_n8419.t1 30.462
R16161 a_n16690_n8419.n1 a_n16690_n8419.t0 30.462
R16162 a_n16690_n8419.n0 a_n16690_n8419.t3 30.462
R16163 a_n16690_n8419.n0 a_n16690_n8419.t5 30.462
R16164 a_n16690_n8419.t4 a_n16690_n8419.n3 30.462
R16165 a_n16690_n8419.n3 a_n16690_n8419.t2 30.462
R16166 MULT_0.4bit_ADDER_2.B3.n5 MULT_0.4bit_ADDER_2.B3.t18 491.64
R16167 MULT_0.4bit_ADDER_2.B3.n6 MULT_0.4bit_ADDER_2.B3.t17 491.64
R16168 MULT_0.4bit_ADDER_2.B3.n7 MULT_0.4bit_ADDER_2.B3.t12 491.64
R16169 MULT_0.4bit_ADDER_2.B3.n8 MULT_0.4bit_ADDER_2.B3.t7 491.64
R16170 MULT_0.4bit_ADDER_2.B3.n3 MULT_0.4bit_ADDER_2.B3.t9 485.221
R16171 MULT_0.4bit_ADDER_2.B3.n1 MULT_0.4bit_ADDER_2.B3.t15 367.928
R16172 MULT_0.4bit_ADDER_2.B3.n9 MULT_0.4bit_ADDER_2.B3.t16 255.588
R16173 MULT_0.4bit_ADDER_2.B3.n0 MULT_0.4bit_ADDER_2.B3.n11 227.526
R16174 MULT_0.4bit_ADDER_2.B3.n0 MULT_0.4bit_ADDER_2.B3.n13 227.266
R16175 MULT_0.4bit_ADDER_2.B3.n0 MULT_0.4bit_ADDER_2.B3.n12 227.266
R16176 MULT_0.4bit_ADDER_2.B3.n2 MULT_0.4bit_ADDER_2.B3.t8 224.478
R16177 MULT_0.4bit_ADDER_2.B3.n1 MULT_0.4bit_ADDER_2.B3.t13 213.688
R16178 MULT_0.4bit_ADDER_2.B3.n5 MULT_0.4bit_ADDER_2.B3.n4 209.19
R16179 MULT_0.4bit_ADDER_2.B3.n4 MULT_0.4bit_ADDER_2.B3.t11 139.78
R16180 MULT_0.4bit_ADDER_2.B3.n4 MULT_0.4bit_ADDER_2.B3.t14 139.78
R16181 MULT_0.4bit_ADDER_2.B3.n4 MULT_0.4bit_ADDER_2.B3.t10 139.78
R16182 MULT_0.4bit_ADDER_2.B3.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_0.A 103.258
R16183 MULT_0.4bit_ADDER_2.B3.n3 MULT_0.4bit_ADDER_2.B3.n2 84.5046
R16184 MULT_0.4bit_ADDER_2.B3.n2 MULT_0.4bit_ADDER_2.B3.n1 72.3005
R16185 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_0.A MULT_0.4bit_ADDER_2.B3.n3 60.9816
R16186 MULT_0.4bit_ADDER_2.B3.n0 MULT_0.4bit_ADDER_2.B3.t3 42.7831
R16187 MULT_0.4bit_ADDER_2.B3.n13 MULT_0.4bit_ADDER_2.B3.t5 30.379
R16188 MULT_0.4bit_ADDER_2.B3.n13 MULT_0.4bit_ADDER_2.B3.t4 30.379
R16189 MULT_0.4bit_ADDER_2.B3.n11 MULT_0.4bit_ADDER_2.B3.t2 30.379
R16190 MULT_0.4bit_ADDER_2.B3.n11 MULT_0.4bit_ADDER_2.B3.t0 30.379
R16191 MULT_0.4bit_ADDER_2.B3.n12 MULT_0.4bit_ADDER_2.B3.t6 30.379
R16192 MULT_0.4bit_ADDER_2.B3.n12 MULT_0.4bit_ADDER_2.B3.t1 30.379
R16193 MULT_0.4bit_ADDER_1.FULL_ADDER_0.COUT MULT_0.4bit_ADDER_2.B3.n0 18.8681
R16194 MULT_0.4bit_ADDER_2.B3.n6 MULT_0.4bit_ADDER_2.B3.n5 17.8661
R16195 MULT_0.4bit_ADDER_2.B3.n7 MULT_0.4bit_ADDER_2.B3.n6 17.8661
R16196 MULT_0.4bit_ADDER_2.B3.n8 MULT_0.4bit_ADDER_2.B3.n7 17.1217
R16197 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_0.A MULT_0.4bit_ADDER_2.B3.n9 15.6329
R16198 MULT_0.4bit_ADDER_2.B3.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_0.A 10.8165
R16199 MULT_0.4bit_ADDER_1.FULL_ADDER_0.COUT MULT_0.4bit_ADDER_1.Cout 5.31784
R16200 MULT_0.4bit_ADDER_2.B3.n9 MULT_0.4bit_ADDER_2.B3.n8 1.8615
R16201 MULT_0.4bit_ADDER_1.Cout MULT_0.4bit_ADDER_2.B3.n10 1.47503
R16202 a_n20737_n11683.n0 a_n20737_n11683.t3 539.788
R16203 a_n20737_n11683.n1 a_n20737_n11683.t5 531.496
R16204 a_n20737_n11683.n0 a_n20737_n11683.t2 490.034
R16205 a_n20737_n11683.n5 a_n20737_n11683.t0 283.788
R16206 a_n20737_n11683.t1 a_n20737_n11683.n5 205.489
R16207 a_n20737_n11683.n2 a_n20737_n11683.t7 182.625
R16208 a_n20737_n11683.n3 a_n20737_n11683.t4 179.054
R16209 a_n20737_n11683.n2 a_n20737_n11683.t6 139.78
R16210 a_n20737_n11683.n4 a_n20737_n11683.n3 101.368
R16211 a_n20737_n11683.n5 a_n20737_n11683.n4 77.9135
R16212 a_n20737_n11683.n4 a_n20737_n11683.n1 76.1557
R16213 a_n20737_n11683.n1 a_n20737_n11683.n0 8.29297
R16214 a_n20737_n11683.n3 a_n20737_n11683.n2 3.57087
R16215 a_n8549_n11683.n2 a_n8549_n11683.n1 121.353
R16216 a_n8549_n11683.n2 a_n8549_n11683.n0 121.353
R16217 a_n8549_n11683.n3 a_n8549_n11683.n2 121.001
R16218 a_n8549_n11683.n1 a_n8549_n11683.t4 30.462
R16219 a_n8549_n11683.n1 a_n8549_n11683.t3 30.462
R16220 a_n8549_n11683.n0 a_n8549_n11683.t0 30.462
R16221 a_n8549_n11683.n0 a_n8549_n11683.t1 30.462
R16222 a_n8549_n11683.t2 a_n8549_n11683.n3 30.462
R16223 a_n8549_n11683.n3 a_n8549_n11683.t5 30.462
R16224 a_n11274_n31085.n2 a_n11274_n31085.n0 121.353
R16225 a_n11274_n31085.n3 a_n11274_n31085.n2 121.353
R16226 a_n11274_n31085.n2 a_n11274_n31085.n1 121.001
R16227 a_n11274_n31085.n0 a_n11274_n31085.t3 30.462
R16228 a_n11274_n31085.n0 a_n11274_n31085.t4 30.462
R16229 a_n11274_n31085.n1 a_n11274_n31085.t5 30.462
R16230 a_n11274_n31085.n1 a_n11274_n31085.t2 30.462
R16231 a_n11274_n31085.t0 a_n11274_n31085.n3 30.462
R16232 a_n11274_n31085.n3 a_n11274_n31085.t1 30.462
R16233 XOR8_0.S6.n0 XOR8_0.S6.t12 1032.02
R16234 XOR8_0.S6.n0 XOR8_0.S6.t13 336.962
R16235 XOR8_0.S6.n0 XOR8_0.S6.t14 326.154
R16236 XOR8_0.S6 XOR8_0.S6.n0 162.946
R16237 XOR8_0.S6.n3 XOR8_0.S6.n1 120.999
R16238 XOR8_0.S6.n3 XOR8_0.S6.n2 120.999
R16239 XOR8_0.S6.n15 XOR8_0.S6.n14 104.865
R16240 XOR8_0.S6.n5 XOR8_0.S6.n4 92.5005
R16241 XOR8_0.S6.n12 XOR8_0.S6.n10 86.2638
R16242 XOR8_0.S6.n10 XOR8_0.S6.n9 85.8873
R16243 XOR8_0.S6.n10 XOR8_0.S6.n7 85.724
R16244 XOR8_0.S6 XOR8_0.S6.n15 83.8907
R16245 XOR8_0.S6.n13 XOR8_0.S6.n9 75.0672
R16246 XOR8_0.S6.n13 XOR8_0.S6.n12 75.0672
R16247 XOR8_0.S6.n9 XOR8_0.S6.n8 73.1255
R16248 XOR8_0.S6.n12 XOR8_0.S6.n11 73.1255
R16249 XOR8_0.S6.n7 XOR8_0.S6.n6 73.1255
R16250 XOR8_0.S6.n14 XOR8_0.S6.n7 68.5181
R16251 XOR8_0.S6.n15 XOR8_0.S6.n5 41.9827
R16252 XOR8_0.S6.n4 XOR8_0.S6.t1 30.462
R16253 XOR8_0.S6.n4 XOR8_0.S6.t7 30.462
R16254 XOR8_0.S6.n1 XOR8_0.S6.t0 30.462
R16255 XOR8_0.S6.n1 XOR8_0.S6.t2 30.462
R16256 XOR8_0.S6.n2 XOR8_0.S6.t8 30.462
R16257 XOR8_0.S6.n2 XOR8_0.S6.t3 30.462
R16258 XOR8_0.S6.n5 XOR8_0.S6.n3 28.124
R16259 XOR8_0.S6.n11 XOR8_0.S6.t5 11.8205
R16260 XOR8_0.S6.n11 XOR8_0.S6.t6 11.8205
R16261 XOR8_0.S6.n8 XOR8_0.S6.t9 11.8205
R16262 XOR8_0.S6.n8 XOR8_0.S6.t10 11.8205
R16263 XOR8_0.S6.n6 XOR8_0.S6.t11 11.8205
R16264 XOR8_0.S6.n6 XOR8_0.S6.t4 11.8205
R16265 XOR8_0.S6.n14 XOR8_0.S6.n13 9.3005
R16266 A7.n18 A7.t21 540.38
R16267 A7.n28 A7.t0 540.375
R16268 A7.n19 A7.t20 491.64
R16269 A7.n19 A7.t37 491.64
R16270 A7.n19 A7.t15 491.64
R16271 A7.n19 A7.t35 491.64
R16272 A7.n10 A7.t7 491.64
R16273 A7.n11 A7.t34 491.64
R16274 A7.n12 A7.t39 491.64
R16275 A7.n13 A7.t16 491.64
R16276 A7.n4 A7.t5 491.64
R16277 A7.n5 A7.t13 491.64
R16278 A7.n6 A7.t19 491.64
R16279 A7.n7 A7.t45 491.64
R16280 A7.n1 A7.t2 491.64
R16281 A7.n1 A7.t1 491.64
R16282 A7.n1 A7.t36 491.64
R16283 A7.n1 A7.t8 491.64
R16284 A7.n16 A7.t29 367.928
R16285 A7.n26 A7.t11 343.827
R16286 A7.n31 A7.t38 312.599
R16287 A7.n14 A7.t43 255.588
R16288 A7.n8 A7.t23 255.588
R16289 A7.n34 A7.t25 247.428
R16290 A7.n33 A7.t10 247.428
R16291 A7.n32 A7.t9 247.428
R16292 A7.n31 A7.t40 247.428
R16293 A7.n15 A7 245.512
R16294 A7.n26 A7.t14 237.787
R16295 A7.n35 A7.t22 229.754
R16296 A7.n27 A7.t30 227.356
R16297 A7.n17 A7.t31 227.356
R16298 A7.n16 A7.t27 213.688
R16299 A7.n10 A7.n9 209.19
R16300 A7.n4 A7.n3 209.19
R16301 A7.n15 A7 205.016
R16302 A7 A7.n2 163.036
R16303 A7.n22 A7.n21 162.867
R16304 A7 A7.n35 162.409
R16305 A7.n18 A7.n17 160.439
R16306 A7.n28 A7.n27 160.433
R16307 A7.n20 A7.t41 139.78
R16308 A7.n20 A7.t17 139.78
R16309 A7.n20 A7.t3 139.78
R16310 A7.n20 A7.t18 139.78
R16311 A7.n9 A7.t6 139.78
R16312 A7.n9 A7.t44 139.78
R16313 A7.n9 A7.t32 139.78
R16314 A7.n3 A7.t4 139.78
R16315 A7.n3 A7.t42 139.78
R16316 A7.n3 A7.t28 139.78
R16317 A7.n0 A7.t12 139.78
R16318 A7.n0 A7.t33 139.78
R16319 A7.n0 A7.t26 139.78
R16320 A7.n0 A7.t24 139.78
R16321 A7.n17 A7.n16 94.4341
R16322 A7.n35 A7.n34 91.5805
R16323 A7.n27 A7.n26 70.3341
R16324 A7.n32 A7.n31 65.1723
R16325 A7.n33 A7.n32 65.1723
R16326 A7.n34 A7.n33 65.1723
R16327 A7.n25 A7 44.763
R16328 A7.n2 A7.n0 38.8368
R16329 A7.n21 A7.n20 38.6833
R16330 A7 A7.n25 29.2084
R16331 A7.n21 A7.n19 28.3986
R16332 A7.n2 A7.n1 28.2451
R16333 A7 A7.n14 27.4136
R16334 A7 A7.n8 27.4136
R16335 A7 A7.n36 20.055
R16336 A7.n24 A7.n23 18.1644
R16337 A7.n11 A7.n10 17.8661
R16338 A7.n12 A7.n11 17.8661
R16339 A7.n5 A7.n4 17.8661
R16340 A7.n6 A7.n5 17.8661
R16341 A7.n13 A7.n12 17.1217
R16342 A7.n7 A7.n6 17.1217
R16343 A7.n36 A7 12.491
R16344 A7.n30 A7.n29 12.4105
R16345 A7 A7.n24 9.66053
R16346 A7.n23 A7.n22 9.00496
R16347 A7.n36 A7.n30 4.28731
R16348 A7.n23 A7 3.87912
R16349 A7.n25 A7 3.10438
R16350 A7.n14 A7.n13 1.8615
R16351 A7.n8 A7.n7 1.8615
R16352 A7.n29 A7 1.38462
R16353 A7 A7.n28 0.905186
R16354 A7 A7.n18 0.89693
R16355 A7 A7.n15 0.452335
R16356 A7.n29 A7 0.0664722
R16357 A7.n22 A7 0.0590664
R16358 A7.n24 A7 0.0268761
R16359 A7.n30 A7 0.0113796
R16360 AND8_0.NOT8_0.A7.n2 AND8_0.NOT8_0.A7.t8 394.37
R16361 AND8_0.NOT8_0.A7.n1 AND8_0.NOT8_0.A7.t10 291.829
R16362 AND8_0.NOT8_0.A7.n1 AND8_0.NOT8_0.A7.t7 291.829
R16363 AND8_0.NOT8_0.A7.n0 AND8_0.NOT8_0.A7.n3 227.526
R16364 AND8_0.NOT8_0.A7.n0 AND8_0.NOT8_0.A7.n4 227.266
R16365 AND8_0.NOT8_0.A7.n0 AND8_0.NOT8_0.A7.n5 227.266
R16366 AND8_0.NOT8_0.A7.n1 AND8_0.NOT8_0.A7.t9 221.72
R16367 AND8_0.NOT8_0.A7.n2 AND8_0.NOT8_0.A7.n1 53.374
R16368 AND8_0.NOT8_0.A7.n0 AND8_0.NOT8_0.A7.t3 42.7803
R16369 AND8_0.NOT8_0.A7.n4 AND8_0.NOT8_0.A7.t0 30.379
R16370 AND8_0.NOT8_0.A7.n4 AND8_0.NOT8_0.A7.t6 30.379
R16371 AND8_0.NOT8_0.A7.n3 AND8_0.NOT8_0.A7.t4 30.379
R16372 AND8_0.NOT8_0.A7.n3 AND8_0.NOT8_0.A7.t5 30.379
R16373 AND8_0.NOT8_0.A7.n5 AND8_0.NOT8_0.A7.t2 30.379
R16374 AND8_0.NOT8_0.A7.n5 AND8_0.NOT8_0.A7.t1 30.379
R16375 AND8_0.NOT8_0.A7 AND8_0.NOT8_0.A7.n0 2.04786
R16376 AND8_0.NOT8_0.A7 AND8_0.NOT8_0.A7.n2 1.26301
R16377 a_n23960_n23839.t0 a_n23960_n23839.t1 19.8005
R16378 mux8_1.NAND4F_6.Y.n1 mux8_1.NAND4F_6.Y.t9 933.563
R16379 mux8_1.NAND4F_6.Y.n1 mux8_1.NAND4F_6.Y.t11 367.635
R16380 mux8_1.NAND4F_6.Y.n2 mux8_1.NAND4F_6.Y.t10 308.481
R16381 mux8_1.NAND4F_6.Y.n0 mux8_1.NAND4F_6.Y.n4 187.373
R16382 mux8_1.NAND4F_6.Y.n0 mux8_1.NAND4F_6.Y.n5 187.192
R16383 mux8_1.NAND4F_6.Y.n0 mux8_1.NAND4F_6.Y.n6 187.192
R16384 mux8_1.NAND4F_6.Y.n8 mux8_1.NAND4F_6.Y.n7 187.192
R16385 mux8_1.NAND4F_6.Y mux8_1.NAND4F_6.Y.n2 162.047
R16386 mux8_1.NAND4F_6.Y.n3 mux8_1.NAND4F_6.Y.t3 22.7831
R16387 mux8_1.NAND4F_6.Y.n3 mux8_1.NAND4F_6.Y 22.171
R16388 mux8_1.NAND4F_6.Y.n4 mux8_1.NAND4F_6.Y.t0 20.1899
R16389 mux8_1.NAND4F_6.Y.n4 mux8_1.NAND4F_6.Y.t1 20.1899
R16390 mux8_1.NAND4F_6.Y.n5 mux8_1.NAND4F_6.Y.t5 20.1899
R16391 mux8_1.NAND4F_6.Y.n5 mux8_1.NAND4F_6.Y.t6 20.1899
R16392 mux8_1.NAND4F_6.Y.n6 mux8_1.NAND4F_6.Y.t7 20.1899
R16393 mux8_1.NAND4F_6.Y.n6 mux8_1.NAND4F_6.Y.t8 20.1899
R16394 mux8_1.NAND4F_6.Y.n7 mux8_1.NAND4F_6.Y.t2 20.1899
R16395 mux8_1.NAND4F_6.Y.n7 mux8_1.NAND4F_6.Y.t4 20.1899
R16396 mux8_1.NAND4F_6.Y.n2 mux8_1.NAND4F_6.Y.n1 10.955
R16397 mux8_1.NAND4F_6.Y mux8_1.NAND4F_6.Y.n3 0.781576
R16398 mux8_1.NAND4F_6.Y mux8_1.NAND4F_6.Y.n8 0.396904
R16399 mux8_1.NAND4F_6.Y.n8 mux8_1.NAND4F_6.Y.n0 0.358709
R16400 MULT_0.4bit_ADDER_0.A2 MULT_0.4bit_ADDER_0.A2.t9 540.38
R16401 MULT_0.4bit_ADDER_0.A2.n4 MULT_0.4bit_ADDER_0.A2.t8 491.64
R16402 MULT_0.4bit_ADDER_0.A2.n4 MULT_0.4bit_ADDER_0.A2.t12 491.64
R16403 MULT_0.4bit_ADDER_0.A2.n4 MULT_0.4bit_ADDER_0.A2.t11 491.64
R16404 MULT_0.4bit_ADDER_0.A2.n4 MULT_0.4bit_ADDER_0.A2.t15 491.64
R16405 MULT_0.4bit_ADDER_0.A2.n2 MULT_0.4bit_ADDER_0.A2.t6 367.928
R16406 MULT_0.4bit_ADDER_0.A2.n0 MULT_0.4bit_ADDER_0.A2.t3 256.529
R16407 MULT_0.4bit_ADDER_0.A2.n3 MULT_0.4bit_ADDER_0.A2.t14 227.356
R16408 MULT_0.4bit_ADDER_0.A2.n0 MULT_0.4bit_ADDER_0.A2.n1 226.292
R16409 MULT_0.4bit_ADDER_0.A2.n2 MULT_0.4bit_ADDER_0.A2.t10 213.688
R16410 MULT_0.4bit_ADDER_0.A2 MULT_0.4bit_ADDER_0.A2.n6 162.867
R16411 MULT_0.4bit_ADDER_0.A2 MULT_0.4bit_ADDER_0.A2.n3 160.439
R16412 MULT_0.4bit_ADDER_0.A2.n5 MULT_0.4bit_ADDER_0.A2.t5 139.78
R16413 MULT_0.4bit_ADDER_0.A2.n5 MULT_0.4bit_ADDER_0.A2.t13 139.78
R16414 MULT_0.4bit_ADDER_0.A2.n5 MULT_0.4bit_ADDER_0.A2.t4 139.78
R16415 MULT_0.4bit_ADDER_0.A2.n5 MULT_0.4bit_ADDER_0.A2.t7 139.78
R16416 MULT_0.4bit_ADDER_0.A2.n3 MULT_0.4bit_ADDER_0.A2.n2 94.4341
R16417 MULT_0.4bit_ADDER_0.A2.n0 MULT_0.4bit_ADDER_0.A2.t0 83.7616
R16418 MULT_0.4bit_ADDER_0.A2.n6 MULT_0.4bit_ADDER_0.A2.n5 38.6833
R16419 MULT_0.4bit_ADDER_0.A2.n1 MULT_0.4bit_ADDER_0.A2.t1 30.379
R16420 MULT_0.4bit_ADDER_0.A2.n1 MULT_0.4bit_ADDER_0.A2.t2 30.379
R16421 MULT_0.4bit_ADDER_0.A2.n6 MULT_0.4bit_ADDER_0.A2.n4 28.3986
R16422 MULT_0.4bit_ADDER_0.A2 MULT_0.4bit_ADDER_0.A2.n7 16.8169
R16423 MULT_0.4bit_ADDER_0.A2 MULT_0.4bit_ADDER_0.A2.n0 15.535
R16424 MULT_0.4bit_ADDER_0.A2.n7 MULT_0.4bit_ADDER_0.A2 9.00496
R16425 MULT_0.4bit_ADDER_0.A2.n7 MULT_0.4bit_ADDER_0.A2 4.77555
R16426 a_n16690_n5154.n2 a_n16690_n5154.n0 121.353
R16427 a_n16690_n5154.n3 a_n16690_n5154.n2 121.353
R16428 a_n16690_n5154.n2 a_n16690_n5154.n1 121.001
R16429 a_n16690_n5154.n0 a_n16690_n5154.t5 30.462
R16430 a_n16690_n5154.n0 a_n16690_n5154.t3 30.462
R16431 a_n16690_n5154.n1 a_n16690_n5154.t0 30.462
R16432 a_n16690_n5154.n1 a_n16690_n5154.t4 30.462
R16433 a_n16690_n5154.t2 a_n16690_n5154.n3 30.462
R16434 a_n16690_n5154.n3 a_n16690_n5154.t1 30.462
R16435 A2.n13 A2.t23 540.38
R16436 A2.n2 A2.t4 540.38
R16437 A2.n26 A2.t21 540.375
R16438 A2.n3 A2.t25 491.64
R16439 A2.n3 A2.t40 491.64
R16440 A2.n3 A2.t6 491.64
R16441 A2.n3 A2.t2 491.64
R16442 A2.n36 A2.t33 491.64
R16443 A2.n36 A2.t7 491.64
R16444 A2.n36 A2.t19 491.64
R16445 A2.n36 A2.t34 491.64
R16446 A2.n10 A2.t36 485.221
R16447 A2.n16 A2.t31 485.221
R16448 A2.n20 A2.t14 485.221
R16449 A2.n8 A2.t1 367.928
R16450 A2.n14 A2.t11 367.928
R16451 A2.n11 A2.t44 367.928
R16452 A2.n18 A2.t32 367.928
R16453 A2.n0 A2.t5 367.928
R16454 A2.n24 A2.t0 343.827
R16455 A2.n29 A2.t22 312.599
R16456 A2.n32 A2.t12 247.428
R16457 A2.n31 A2.t43 247.428
R16458 A2.n30 A2.t41 247.428
R16459 A2.n29 A2.t24 247.428
R16460 A2.n24 A2.t16 237.787
R16461 A2.n33 A2.t9 229.754
R16462 A2.n25 A2.t26 227.356
R16463 A2.n12 A2.t15 227.356
R16464 A2.n1 A2.t35 227.356
R16465 A2.n9 A2.t29 224.478
R16466 A2.n15 A2.t18 224.478
R16467 A2.n19 A2.t39 224.478
R16468 A2.n8 A2.t45 213.688
R16469 A2.n14 A2.t17 213.688
R16470 A2.n11 A2.t3 213.688
R16471 A2.n18 A2.t37 213.688
R16472 A2.n0 A2.t38 213.688
R16473 A2 A2.n37 163.036
R16474 A2.n6 A2.n5 162.867
R16475 A2 A2.n33 162.409
R16476 A2.n13 A2.n12 160.439
R16477 A2.n2 A2.n1 160.439
R16478 A2.n26 A2.n25 160.433
R16479 A2.n4 A2.t30 139.78
R16480 A2.n4 A2.t27 139.78
R16481 A2.n4 A2.t8 139.78
R16482 A2.n4 A2.t20 139.78
R16483 A2.n35 A2.t42 139.78
R16484 A2.n35 A2.t13 139.78
R16485 A2.n35 A2.t10 139.78
R16486 A2.n35 A2.t28 139.78
R16487 A2.n12 A2.n11 94.4341
R16488 A2.n1 A2.n0 94.4341
R16489 A2.n33 A2.n32 91.5805
R16490 A2.n10 A2.n9 84.5046
R16491 A2.n16 A2.n15 84.5046
R16492 A2.n20 A2.n19 84.5046
R16493 A2.n9 A2.n8 72.3005
R16494 A2.n15 A2.n14 72.3005
R16495 A2.n19 A2.n18 72.3005
R16496 A2.n25 A2.n24 70.3341
R16497 A2.n30 A2.n29 65.1723
R16498 A2.n31 A2.n30 65.1723
R16499 A2.n32 A2.n31 65.1723
R16500 A2 A2.n10 61.0566
R16501 A2 A2.n16 61.0566
R16502 A2 A2.n20 61.0566
R16503 A2.n37 A2.n35 38.8368
R16504 A2.n5 A2.n4 38.6833
R16505 A2.n23 A2 31.8838
R16506 A2.n5 A2.n3 28.3986
R16507 A2.n37 A2.n36 28.2451
R16508 A2 A2.n7 18.1883
R16509 A2.n38 A2.n34 16.7501
R16510 A2.n34 A2 12.5661
R16511 A2.n28 A2.n27 12.4105
R16512 A2.n7 A2.n6 9.00496
R16513 A2.n23 A2.n22 7.00398
R16514 A2.n17 A2 6.43387
R16515 A2.n21 A2 6.03372
R16516 A2 A2.n23 4.73128
R16517 A2.n17 A2 4.56448
R16518 A2 A2.n17 4.17188
R16519 A2.n7 A2 3.87912
R16520 A2.n34 A2.n28 3.70809
R16521 A2.n22 A2 3.39248
R16522 A2.n22 A2.n21 2.11645
R16523 A2.n38 A2 1.93857
R16524 A2.n27 A2 1.34697
R16525 A2 A2.n26 0.905186
R16526 A2 A2.n2 0.89693
R16527 A2 A2.n13 0.878165
R16528 A2.n21 A2 0.405967
R16529 A2.n27 A2 0.0679157
R16530 A2.n6 A2 0.0590664
R16531 A2 A2.n38 0.0171495
R16532 A2.n28 A2 0.0166414
R16533 AND8_0.NOT8_0.A2.n2 AND8_0.NOT8_0.A2.t10 394.37
R16534 AND8_0.NOT8_0.A2.n1 AND8_0.NOT8_0.A2.t9 291.829
R16535 AND8_0.NOT8_0.A2.n1 AND8_0.NOT8_0.A2.t7 291.829
R16536 AND8_0.NOT8_0.A2.n0 AND8_0.NOT8_0.A2.n3 227.526
R16537 AND8_0.NOT8_0.A2.n0 AND8_0.NOT8_0.A2.n4 227.266
R16538 AND8_0.NOT8_0.A2.n0 AND8_0.NOT8_0.A2.n5 227.266
R16539 AND8_0.NOT8_0.A2.n1 AND8_0.NOT8_0.A2.t8 221.72
R16540 AND8_0.NOT8_0.A2.n2 AND8_0.NOT8_0.A2.n1 53.374
R16541 AND8_0.NOT8_0.A2.n0 AND8_0.NOT8_0.A2.t2 42.7803
R16542 AND8_0.NOT8_0.A2.n4 AND8_0.NOT8_0.A2.t3 30.379
R16543 AND8_0.NOT8_0.A2.n4 AND8_0.NOT8_0.A2.t0 30.379
R16544 AND8_0.NOT8_0.A2.n3 AND8_0.NOT8_0.A2.t1 30.379
R16545 AND8_0.NOT8_0.A2.n3 AND8_0.NOT8_0.A2.t6 30.379
R16546 AND8_0.NOT8_0.A2.n5 AND8_0.NOT8_0.A2.t5 30.379
R16547 AND8_0.NOT8_0.A2.n5 AND8_0.NOT8_0.A2.t4 30.379
R16548 AND8_0.NOT8_0.A2 AND8_0.NOT8_0.A2.n0 2.08362
R16549 AND8_0.NOT8_0.A2 AND8_0.NOT8_0.A2.n2 1.28475
R16550 a_n24804_1406.n0 a_n24804_1406.t2 539.788
R16551 a_n24804_1406.n1 a_n24804_1406.t4 531.496
R16552 a_n24804_1406.n0 a_n24804_1406.t5 490.034
R16553 a_n24804_1406.n5 a_n24804_1406.t0 283.788
R16554 a_n24804_1406.t1 a_n24804_1406.n5 205.489
R16555 a_n24804_1406.n2 a_n24804_1406.t6 182.625
R16556 a_n24804_1406.n3 a_n24804_1406.t7 179.054
R16557 a_n24804_1406.n2 a_n24804_1406.t3 139.78
R16558 a_n24804_1406.n4 a_n24804_1406.n3 101.368
R16559 a_n24804_1406.n5 a_n24804_1406.n4 77.9135
R16560 a_n24804_1406.n4 a_n24804_1406.n1 76.1557
R16561 a_n24804_1406.n1 a_n24804_1406.n0 8.29297
R16562 a_n24804_1406.n3 a_n24804_1406.n2 3.57087
R16563 a_n24624_2026.n0 a_n24624_2026.n2 81.2978
R16564 a_n24624_2026.n0 a_n24624_2026.n3 81.1637
R16565 a_n24624_2026.n0 a_n24624_2026.n4 81.1637
R16566 a_n24624_2026.n1 a_n24624_2026.n5 81.1637
R16567 a_n24624_2026.n1 a_n24624_2026.n6 81.1637
R16568 a_n24624_2026.n7 a_n24624_2026.n1 80.9213
R16569 a_n24624_2026.n2 a_n24624_2026.t9 11.8205
R16570 a_n24624_2026.n2 a_n24624_2026.t10 11.8205
R16571 a_n24624_2026.n3 a_n24624_2026.t1 11.8205
R16572 a_n24624_2026.n3 a_n24624_2026.t11 11.8205
R16573 a_n24624_2026.n4 a_n24624_2026.t2 11.8205
R16574 a_n24624_2026.n4 a_n24624_2026.t0 11.8205
R16575 a_n24624_2026.n5 a_n24624_2026.t7 11.8205
R16576 a_n24624_2026.n5 a_n24624_2026.t8 11.8205
R16577 a_n24624_2026.n6 a_n24624_2026.t3 11.8205
R16578 a_n24624_2026.n6 a_n24624_2026.t6 11.8205
R16579 a_n24624_2026.n7 a_n24624_2026.t4 11.8205
R16580 a_n24624_2026.t5 a_n24624_2026.n7 11.8205
R16581 a_n24624_2026.n1 a_n24624_2026.n0 0.402735
R16582 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t20 491.64
R16583 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t15 491.64
R16584 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t17 491.64
R16585 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t12 491.64
R16586 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t16 485.221
R16587 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t18 367.928
R16588 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t22 255.588
R16589 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t19 224.478
R16590 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t21 213.688
R16591 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n0 209.19
R16592 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t23 139.78
R16593 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t13 139.78
R16594 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t14 139.78
R16595 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n10 120.999
R16596 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n9 120.999
R16597 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n22 104.489
R16598 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n12 92.5005
R16599 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n18 86.2638
R16600 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n17 85.8873
R16601 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n15 85.724
R16602 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n7 84.5046
R16603 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n23 83.8907
R16604 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n20 75.0672
R16605 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n17 75.0672
R16606 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n19 73.1255
R16607 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n17 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n16 73.1255
R16608 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n15 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n14 73.1255
R16609 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n6 72.3005
R16610 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n15 68.8946
R16611 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n8 60.9797
R16612 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n13 41.9827
R16613 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t10 30.462
R16614 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t4 30.462
R16615 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t5 30.462
R16616 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t3 30.462
R16617 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t11 30.462
R16618 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t9 30.462
R16619 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n11 28.124
R16620 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n5 19.963
R16621 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n1 17.8661
R16622 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n2 17.8661
R16623 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n3 17.1217
R16624 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t6 11.8205
R16625 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t7 11.8205
R16626 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t0 11.8205
R16627 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t1 11.8205
R16628 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t8 11.8205
R16629 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t2 11.8205
R16630 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n21 9.3005
R16631 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n4 1.8615
R16632 mux8_0.NAND4F_8.Y.n1 mux8_0.NAND4F_8.Y.t11 379.173
R16633 mux8_0.NAND4F_8.Y.n2 mux8_0.NAND4F_8.Y.t10 312.599
R16634 mux8_0.NAND4F_8.Y.n1 mux8_0.NAND4F_8.Y.t9 247.428
R16635 mux8_0.NAND4F_8.Y.n4 mux8_0.NAND4F_8.Y.t12 247.428
R16636 mux8_0.NAND4F_8.Y.n3 mux8_0.NAND4F_8.Y.t13 247.428
R16637 mux8_0.NAND4F_8.Y.n2 mux8_0.NAND4F_8.Y.t14 247.428
R16638 mux8_0.NAND4F_8.Y.n0 mux8_0.NAND4F_8.Y.n6 187.373
R16639 mux8_0.NAND4F_8.Y.n0 mux8_0.NAND4F_8.Y.n7 187.192
R16640 mux8_0.NAND4F_8.Y.n0 mux8_0.NAND4F_8.Y.n8 187.192
R16641 mux8_0.NAND4F_8.Y.n10 mux8_0.NAND4F_8.Y.n9 187.192
R16642 mux8_0.NAND4F_8.Y mux8_0.NAND4F_8.Y.n5 162.139
R16643 mux8_0.NAND4F_8.Y.n4 mux8_0.NAND4F_8.Y.n3 65.1723
R16644 mux8_0.NAND4F_8.Y.n3 mux8_0.NAND4F_8.Y.n2 65.1723
R16645 mux8_0.NAND4F_8.Y.n5 mux8_0.NAND4F_8.Y.n4 33.2653
R16646 mux8_0.NAND4F_8.Y.n5 mux8_0.NAND4F_8.Y.n1 31.9075
R16647 mux8_0.NAND4F_8.Y mux8_0.NAND4F_8.Y.t8 22.6141
R16648 mux8_0.NAND4F_8.Y.n6 mux8_0.NAND4F_8.Y.t2 20.1899
R16649 mux8_0.NAND4F_8.Y.n6 mux8_0.NAND4F_8.Y.t3 20.1899
R16650 mux8_0.NAND4F_8.Y.n7 mux8_0.NAND4F_8.Y.t0 20.1899
R16651 mux8_0.NAND4F_8.Y.n7 mux8_0.NAND4F_8.Y.t1 20.1899
R16652 mux8_0.NAND4F_8.Y.n8 mux8_0.NAND4F_8.Y.t5 20.1899
R16653 mux8_0.NAND4F_8.Y.n8 mux8_0.NAND4F_8.Y.t4 20.1899
R16654 mux8_0.NAND4F_8.Y.n9 mux8_0.NAND4F_8.Y.t6 20.1899
R16655 mux8_0.NAND4F_8.Y.n9 mux8_0.NAND4F_8.Y.t7 20.1899
R16656 mux8_0.NAND4F_8.Y mux8_0.NAND4F_8.Y.n10 0.452586
R16657 mux8_0.NAND4F_8.Y.n10 mux8_0.NAND4F_8.Y.n0 0.358709
R16658 a_11865_1753.n1 a_11865_1753.n4 231.24
R16659 a_11865_1753.n0 a_11865_1753.n2 231.24
R16660 a_11865_1753.n1 a_11865_1753.n5 231.03
R16661 a_11865_1753.n0 a_11865_1753.n3 231.03
R16662 a_11865_1753.n6 a_11865_1753.n1 231.03
R16663 a_11865_1753.n4 a_11865_1753.t0 25.395
R16664 a_11865_1753.n4 a_11865_1753.t3 25.395
R16665 a_11865_1753.n5 a_11865_1753.t2 25.395
R16666 a_11865_1753.n5 a_11865_1753.t1 25.395
R16667 a_11865_1753.n3 a_11865_1753.t5 25.395
R16668 a_11865_1753.n3 a_11865_1753.t6 25.395
R16669 a_11865_1753.n2 a_11865_1753.t7 25.395
R16670 a_11865_1753.n2 a_11865_1753.t9 25.395
R16671 a_11865_1753.n6 a_11865_1753.t8 25.395
R16672 a_11865_1753.t4 a_11865_1753.n6 25.395
R16673 a_11865_1753.n1 a_11865_1753.n0 0.421553
R16674 V_FLAG_0.NAND2_0.Y.n5 V_FLAG_0.NAND2_0.Y.t8 385.697
R16675 V_FLAG_0.NAND2_0.Y.n0 V_FLAG_0.NAND2_0.Y.t7 291.829
R16676 V_FLAG_0.NAND2_0.Y.n0 V_FLAG_0.NAND2_0.Y.t9 291.829
R16677 V_FLAG_0.inv_0.A V_FLAG_0.NAND2_0.Y.n2 227.526
R16678 V_FLAG_0.inv_0.A V_FLAG_0.NAND2_0.Y.n3 227.266
R16679 V_FLAG_0.inv_0.A V_FLAG_0.NAND2_0.Y.n1 227.266
R16680 V_FLAG_0.NAND2_0.Y.n0 V_FLAG_0.NAND2_0.Y.t10 221.72
R16681 V_FLAG_0.NAND2_0.Y.n5 V_FLAG_0.NAND2_0.Y.n4 89.6005
R16682 V_FLAG_0.NAND2_0.Y.n4 V_FLAG_0.NAND2_0.Y.n0 50.6672
R16683 V_FLAG_0.inv_0.A V_FLAG_0.NAND2_0.Y.t1 42.8112
R16684 V_FLAG_0.NAND2_0.Y.n3 V_FLAG_0.NAND2_0.Y.t2 30.379
R16685 V_FLAG_0.NAND2_0.Y.n3 V_FLAG_0.NAND2_0.Y.t5 30.379
R16686 V_FLAG_0.NAND2_0.Y.n1 V_FLAG_0.NAND2_0.Y.t3 30.379
R16687 V_FLAG_0.NAND2_0.Y.n1 V_FLAG_0.NAND2_0.Y.t0 30.379
R16688 V_FLAG_0.NAND2_0.Y.n2 V_FLAG_0.NAND2_0.Y.t4 30.379
R16689 V_FLAG_0.NAND2_0.Y.n2 V_FLAG_0.NAND2_0.Y.t6 30.379
R16690 V_FLAG_0.inv_0.A V_FLAG_0.NAND2_0.Y.n5 9.56753
R16691 V_FLAG_0.NAND2_0.Y.n4 V_FLAG_0.inv_0.A 3.47999
R16692 V.n1 V.t2 256.514
R16693 V.n1 V.n0 226.258
R16694 V V.t0 83.7284
R16695 V.n0 V.t3 30.379
R16696 V.n0 V.t1 30.379
R16697 V V.n1 0.0397628
R16698 a_n15737_n8445.n2 a_n15737_n8445.t6 541.395
R16699 a_n15737_n8445.n3 a_n15737_n8445.t4 527.402
R16700 a_n15737_n8445.n2 a_n15737_n8445.t3 491.64
R16701 a_n15737_n8445.n5 a_n15737_n8445.t0 281.906
R16702 a_n15737_n8445.t1 a_n15737_n8445.n5 204.359
R16703 a_n15737_n8445.n0 a_n15737_n8445.t7 180.73
R16704 a_n15737_n8445.n1 a_n15737_n8445.t5 179.45
R16705 a_n15737_n8445.n0 a_n15737_n8445.t2 139.78
R16706 a_n15737_n8445.n4 a_n15737_n8445.n1 105.635
R16707 a_n15737_n8445.n4 a_n15737_n8445.n3 76.0005
R16708 a_n15737_n8445.n5 a_n15737_n8445.n4 67.9685
R16709 a_n15737_n8445.n3 a_n15737_n8445.n2 13.994
R16710 a_n15737_n8445.n1 a_n15737_n8445.n0 1.28015
R16711 a_n15707_n8419.n3 a_n15707_n8419.n2 121.353
R16712 a_n15707_n8419.n2 a_n15707_n8419.n1 121.001
R16713 a_n15707_n8419.n2 a_n15707_n8419.n0 120.977
R16714 a_n15707_n8419.n1 a_n15707_n8419.t2 30.462
R16715 a_n15707_n8419.n1 a_n15707_n8419.t3 30.462
R16716 a_n15707_n8419.n0 a_n15707_n8419.t0 30.462
R16717 a_n15707_n8419.n0 a_n15707_n8419.t1 30.462
R16718 a_n15707_n8419.n3 a_n15707_n8419.t5 30.462
R16719 a_n15707_n8419.t4 a_n15707_n8419.n3 30.462
R16720 XOR8_0.S1.n0 XOR8_0.S1.t13 1032.02
R16721 XOR8_0.S1.n0 XOR8_0.S1.t14 336.962
R16722 XOR8_0.S1.n0 XOR8_0.S1.t12 326.154
R16723 XOR8_0.S1 XOR8_0.S1.n0 162.946
R16724 XOR8_0.S1.n3 XOR8_0.S1.n1 120.999
R16725 XOR8_0.S1.n3 XOR8_0.S1.n2 120.999
R16726 XOR8_0.S1.n15 XOR8_0.S1.n14 104.865
R16727 XOR8_0.S1.n5 XOR8_0.S1.n4 92.5005
R16728 XOR8_0.S1.n12 XOR8_0.S1.n10 86.2638
R16729 XOR8_0.S1.n10 XOR8_0.S1.n9 85.8873
R16730 XOR8_0.S1.n10 XOR8_0.S1.n7 85.724
R16731 XOR8_0.S1 XOR8_0.S1.n15 83.8907
R16732 XOR8_0.S1.n13 XOR8_0.S1.n12 75.0672
R16733 XOR8_0.S1.n13 XOR8_0.S1.n9 75.0672
R16734 XOR8_0.S1.n7 XOR8_0.S1.n6 73.1255
R16735 XOR8_0.S1.n12 XOR8_0.S1.n11 73.1255
R16736 XOR8_0.S1.n9 XOR8_0.S1.n8 73.1255
R16737 XOR8_0.S1.n14 XOR8_0.S1.n7 68.5181
R16738 XOR8_0.S1.n15 XOR8_0.S1.n5 41.9827
R16739 XOR8_0.S1.n4 XOR8_0.S1.t6 30.462
R16740 XOR8_0.S1.n4 XOR8_0.S1.t11 30.462
R16741 XOR8_0.S1.n1 XOR8_0.S1.t4 30.462
R16742 XOR8_0.S1.n1 XOR8_0.S1.t5 30.462
R16743 XOR8_0.S1.n2 XOR8_0.S1.t0 30.462
R16744 XOR8_0.S1.n2 XOR8_0.S1.t7 30.462
R16745 XOR8_0.S1.n5 XOR8_0.S1.n3 28.124
R16746 XOR8_0.S1.n11 XOR8_0.S1.t9 11.8205
R16747 XOR8_0.S1.n11 XOR8_0.S1.t10 11.8205
R16748 XOR8_0.S1.n6 XOR8_0.S1.t3 11.8205
R16749 XOR8_0.S1.n6 XOR8_0.S1.t8 11.8205
R16750 XOR8_0.S1.n8 XOR8_0.S1.t1 11.8205
R16751 XOR8_0.S1.n8 XOR8_0.S1.t2 11.8205
R16752 XOR8_0.S1.n14 XOR8_0.S1.n13 9.3005
R16753 mux8_2.NAND4F_1.Y.n2 mux8_2.NAND4F_1.Y.t11 978.795
R16754 mux8_2.NAND4F_1.Y.n1 mux8_2.NAND4F_1.Y.t10 308.481
R16755 mux8_2.NAND4F_1.Y.n1 mux8_2.NAND4F_1.Y.t9 308.481
R16756 mux8_2.NAND4F_1.Y.n0 mux8_2.NAND4F_1.Y.n3 187.373
R16757 mux8_2.NAND4F_1.Y.n0 mux8_2.NAND4F_1.Y.n4 187.192
R16758 mux8_2.NAND4F_1.Y.n0 mux8_2.NAND4F_1.Y.n5 187.192
R16759 mux8_2.NAND4F_1.Y.n7 mux8_2.NAND4F_1.Y.n6 187.192
R16760 mux8_2.NAND4F_1.Y mux8_2.NAND4F_1.Y.n2 161.84
R16761 mux8_2.NAND4F_1.Y mux8_2.NAND4F_1.Y.t4 23.4335
R16762 mux8_2.NAND4F_1.Y.n3 mux8_2.NAND4F_1.Y.t0 20.1899
R16763 mux8_2.NAND4F_1.Y.n3 mux8_2.NAND4F_1.Y.t1 20.1899
R16764 mux8_2.NAND4F_1.Y.n4 mux8_2.NAND4F_1.Y.t6 20.1899
R16765 mux8_2.NAND4F_1.Y.n4 mux8_2.NAND4F_1.Y.t5 20.1899
R16766 mux8_2.NAND4F_1.Y.n5 mux8_2.NAND4F_1.Y.t8 20.1899
R16767 mux8_2.NAND4F_1.Y.n5 mux8_2.NAND4F_1.Y.t7 20.1899
R16768 mux8_2.NAND4F_1.Y.n6 mux8_2.NAND4F_1.Y.t2 20.1899
R16769 mux8_2.NAND4F_1.Y.n6 mux8_2.NAND4F_1.Y.t3 20.1899
R16770 mux8_2.NAND4F_1.Y.n2 mux8_2.NAND4F_1.Y.n1 11.0463
R16771 mux8_2.NAND4F_1.Y mux8_2.NAND4F_1.Y.n7 0.527586
R16772 mux8_2.NAND4F_1.Y.n7 mux8_2.NAND4F_1.Y.n0 0.358709
R16773 mux8_0.NAND4F_0.C.n6 mux8_0.NAND4F_0.C.t7 978.795
R16774 mux8_0.NAND4F_0.C.n4 mux8_0.NAND4F_0.C.t5 978.795
R16775 mux8_0.NAND4F_0.C.n11 mux8_0.NAND4F_0.C.t14 978.795
R16776 mux8_0.NAND4F_0.C.n2 mux8_0.NAND4F_0.C.t9 978.795
R16777 mux8_0.NAND4F_0.C.n5 mux8_0.NAND4F_0.C.t6 308.481
R16778 mux8_0.NAND4F_0.C.n5 mux8_0.NAND4F_0.C.t4 308.481
R16779 mux8_0.NAND4F_0.C.n3 mux8_0.NAND4F_0.C.t11 308.481
R16780 mux8_0.NAND4F_0.C.n3 mux8_0.NAND4F_0.C.t8 308.481
R16781 mux8_0.NAND4F_0.C.n10 mux8_0.NAND4F_0.C.t13 308.481
R16782 mux8_0.NAND4F_0.C.n10 mux8_0.NAND4F_0.C.t15 308.481
R16783 mux8_0.NAND4F_0.C.n1 mux8_0.NAND4F_0.C.t10 308.481
R16784 mux8_0.NAND4F_0.C.n1 mux8_0.NAND4F_0.C.t12 308.481
R16785 mux8_0.NAND4F_0.C.n0 mux8_0.NAND4F_0.C.t1 256.514
R16786 mux8_0.NAND4F_0.C.n0 mux8_0.NAND4F_0.C.n8 226.258
R16787 mux8_0.NAND4F_0.C mux8_0.NAND4F_0.C.n6 161.856
R16788 mux8_0.NAND4F_0.C mux8_0.NAND4F_0.C.n4 161.847
R16789 mux8_0.NAND4F_0.C mux8_0.NAND4F_0.C.n11 161.84
R16790 mux8_0.NAND4F_0.C mux8_0.NAND4F_0.C.n2 161.831
R16791 mux8_0.NAND4F_0.C.n0 mux8_0.NAND4F_0.C.t0 83.7172
R16792 mux8_0.NAND4F_0.C.n8 mux8_0.NAND4F_0.C.t2 30.379
R16793 mux8_0.NAND4F_0.C.n8 mux8_0.NAND4F_0.C.t3 30.379
R16794 mux8_0.NAND4F_0.C.n9 mux8_0.NAND4F_0.C.n0 13.5186
R16795 mux8_0.NAND4F_0.C mux8_0.NAND4F_0.C.n12 13.0862
R16796 mux8_0.NAND4F_0.C.n7 mux8_0.NAND4F_0.C 13.0435
R16797 mux8_0.NAND4F_0.C.n12 mux8_0.NAND4F_0.C 12.4135
R16798 mux8_0.NAND4F_0.C.n7 mux8_0.NAND4F_0.C 12.4105
R16799 mux8_0.NAND4F_0.C.n6 mux8_0.NAND4F_0.C.n5 11.0463
R16800 mux8_0.NAND4F_0.C.n4 mux8_0.NAND4F_0.C.n3 11.0463
R16801 mux8_0.NAND4F_0.C.n11 mux8_0.NAND4F_0.C.n10 11.0463
R16802 mux8_0.NAND4F_0.C.n2 mux8_0.NAND4F_0.C.n1 11.0463
R16803 mux8_0.NAND4F_0.C.n12 mux8_0.NAND4F_0.C.n9 3.46056
R16804 mux8_0.NAND4F_0.C.n9 mux8_0.NAND4F_0.C.n7 1.8134
R16805 mux8_0.NAND4F_3.Y.n7 mux8_0.NAND4F_3.Y.t9 978.795
R16806 mux8_0.NAND4F_3.Y.n6 mux8_0.NAND4F_3.Y.t11 308.481
R16807 mux8_0.NAND4F_3.Y.n6 mux8_0.NAND4F_3.Y.t10 308.481
R16808 mux8_0.NAND4F_3.Y.n0 mux8_0.NAND4F_3.Y.n1 187.373
R16809 mux8_0.NAND4F_3.Y.n0 mux8_0.NAND4F_3.Y.n2 187.192
R16810 mux8_0.NAND4F_3.Y.n0 mux8_0.NAND4F_3.Y.n3 187.192
R16811 mux8_0.NAND4F_3.Y.n5 mux8_0.NAND4F_3.Y.n4 187.192
R16812 mux8_0.NAND4F_3.Y mux8_0.NAND4F_3.Y.n7 161.839
R16813 mux8_0.NAND4F_3.Y mux8_0.NAND4F_3.Y.t6 23.4426
R16814 mux8_0.NAND4F_3.Y.n1 mux8_0.NAND4F_3.Y.t7 20.1899
R16815 mux8_0.NAND4F_3.Y.n1 mux8_0.NAND4F_3.Y.t8 20.1899
R16816 mux8_0.NAND4F_3.Y.n2 mux8_0.NAND4F_3.Y.t3 20.1899
R16817 mux8_0.NAND4F_3.Y.n2 mux8_0.NAND4F_3.Y.t2 20.1899
R16818 mux8_0.NAND4F_3.Y.n3 mux8_0.NAND4F_3.Y.t0 20.1899
R16819 mux8_0.NAND4F_3.Y.n3 mux8_0.NAND4F_3.Y.t1 20.1899
R16820 mux8_0.NAND4F_3.Y.n4 mux8_0.NAND4F_3.Y.t5 20.1899
R16821 mux8_0.NAND4F_3.Y.n4 mux8_0.NAND4F_3.Y.t4 20.1899
R16822 mux8_0.NAND4F_3.Y.n7 mux8_0.NAND4F_3.Y.n6 11.0463
R16823 mux8_0.NAND4F_3.Y mux8_0.NAND4F_3.Y.n5 0.518495
R16824 mux8_0.NAND4F_3.Y.n5 mux8_0.NAND4F_3.Y.n0 0.358709
R16825 A5.n5 A5.t25 540.38
R16826 A5.n13 A5.t24 540.375
R16827 A5.n6 A5.t10 491.64
R16828 A5.n6 A5.t16 491.64
R16829 A5.n6 A5.t4 491.64
R16830 A5.n6 A5.t13 491.64
R16831 A5.n1 A5.t6 491.64
R16832 A5.n1 A5.t2 491.64
R16833 A5.n1 A5.t23 491.64
R16834 A5.n1 A5.t7 491.64
R16835 A5.n3 A5.t27 367.928
R16836 A5.n11 A5.t20 343.827
R16837 A5.n16 A5.t11 312.599
R16838 A5.n19 A5.t3 247.428
R16839 A5.n18 A5.t22 247.428
R16840 A5.n17 A5.t21 247.428
R16841 A5.n16 A5.t12 247.428
R16842 A5.n11 A5.t5 237.787
R16843 A5.n20 A5.t1 229.754
R16844 A5.n12 A5.t14 227.356
R16845 A5.n4 A5.t28 227.356
R16846 A5.n3 A5.t29 213.688
R16847 A5 A5.n2 163.036
R16848 A5.n9 A5.n8 162.867
R16849 A5 A5.n20 162.409
R16850 A5.n5 A5.n4 160.439
R16851 A5.n13 A5.n12 160.433
R16852 A5.n7 A5.t19 139.78
R16853 A5.n7 A5.t0 139.78
R16854 A5.n7 A5.t26 139.78
R16855 A5.n7 A5.t8 139.78
R16856 A5.n0 A5.t9 139.78
R16857 A5.n0 A5.t18 139.78
R16858 A5.n0 A5.t17 139.78
R16859 A5.n0 A5.t15 139.78
R16860 A5.n4 A5.n3 94.4341
R16861 A5.n20 A5.n19 91.5805
R16862 A5.n12 A5.n11 70.3341
R16863 A5.n17 A5.n16 65.1723
R16864 A5.n18 A5.n17 65.1723
R16865 A5.n19 A5.n18 65.1723
R16866 A5.n2 A5.n0 38.8368
R16867 A5.n8 A5.n7 38.6833
R16868 A5.n8 A5.n6 28.3986
R16869 A5.n2 A5.n1 28.2451
R16870 A5 A5.n21 18.8691
R16871 A5 A5.n10 18.1875
R16872 A5.n21 A5 12.5006
R16873 A5.n15 A5.n14 12.4105
R16874 A5.n10 A5.n9 9.00496
R16875 A5.n21 A5.n15 4.14228
R16876 A5.n10 A5 3.87912
R16877 A5.n14 A5 1.41844
R16878 A5 A5.n13 0.905186
R16879 A5 A5.n5 0.89693
R16880 A5.n14 A5 0.0749382
R16881 A5.n9 A5 0.0590664
R16882 A5.n15 A5 0.0166414
R16883 a_n18072_1380.n2 a_n18072_1380.t7 541.395
R16884 a_n18072_1380.n3 a_n18072_1380.t5 527.402
R16885 a_n18072_1380.n2 a_n18072_1380.t4 491.64
R16886 a_n18072_1380.n5 a_n18072_1380.t0 281.906
R16887 a_n18072_1380.t1 a_n18072_1380.n5 204.359
R16888 a_n18072_1380.n0 a_n18072_1380.t3 180.73
R16889 a_n18072_1380.n1 a_n18072_1380.t2 179.45
R16890 a_n18072_1380.n0 a_n18072_1380.t6 139.78
R16891 a_n18072_1380.n4 a_n18072_1380.n1 105.635
R16892 a_n18072_1380.n4 a_n18072_1380.n3 76.0005
R16893 a_n18072_1380.n5 a_n18072_1380.n4 67.9685
R16894 a_n18072_1380.n3 a_n18072_1380.n2 13.994
R16895 a_n18072_1380.n1 a_n18072_1380.n0 1.28015
R16896 mux8_7.NAND4F_4.B.n10 mux8_7.NAND4F_4.B.t14 933.563
R16897 mux8_7.NAND4F_4.B.n5 mux8_7.NAND4F_4.B.t8 933.563
R16898 mux8_7.NAND4F_4.B.n3 mux8_7.NAND4F_4.B.t11 933.563
R16899 mux8_7.NAND4F_4.B.n1 mux8_7.NAND4F_4.B.t6 933.563
R16900 mux8_7.NAND4F_4.B.n10 mux8_7.NAND4F_4.B.t9 367.635
R16901 mux8_7.NAND4F_4.B.n5 mux8_7.NAND4F_4.B.t12 367.635
R16902 mux8_7.NAND4F_4.B.n3 mux8_7.NAND4F_4.B.t5 367.635
R16903 mux8_7.NAND4F_4.B.n1 mux8_7.NAND4F_4.B.t15 367.635
R16904 mux8_7.NAND4F_4.B.n11 mux8_7.NAND4F_4.B.t10 308.481
R16905 mux8_7.NAND4F_4.B.n6 mux8_7.NAND4F_4.B.t13 308.481
R16906 mux8_7.NAND4F_4.B.n4 mux8_7.NAND4F_4.B.t7 308.481
R16907 mux8_7.NAND4F_4.B.n2 mux8_7.NAND4F_4.B.t4 308.481
R16908 mux8_7.NAND4F_4.B.n0 mux8_7.NAND4F_4.B.t1 256.514
R16909 mux8_7.NAND4F_4.B.n0 mux8_7.NAND4F_4.B.n8 226.258
R16910 mux8_7.NAND4F_4.B mux8_7.NAND4F_4.B.n2 162.173
R16911 mux8_7.NAND4F_4.B mux8_7.NAND4F_4.B.n6 162.137
R16912 mux8_7.NAND4F_4.B mux8_7.NAND4F_4.B.n11 162.117
R16913 mux8_7.NAND4F_4.B.n7 mux8_7.NAND4F_4.B.n4 161.703
R16914 mux8_7.NAND4F_4.B.n0 mux8_7.NAND4F_4.B.t0 83.7172
R16915 mux8_7.NAND4F_4.B.n8 mux8_7.NAND4F_4.B.t3 30.379
R16916 mux8_7.NAND4F_4.B.n8 mux8_7.NAND4F_4.B.t2 30.379
R16917 mux8_7.NAND4F_4.B.n12 mux8_7.NAND4F_4.B 24.8912
R16918 mux8_7.NAND4F_4.B.n7 mux8_7.NAND4F_4.B 21.6618
R16919 mux8_7.NAND4F_4.B.n11 mux8_7.NAND4F_4.B.n10 10.955
R16920 mux8_7.NAND4F_4.B.n6 mux8_7.NAND4F_4.B.n5 10.955
R16921 mux8_7.NAND4F_4.B.n4 mux8_7.NAND4F_4.B.n3 10.955
R16922 mux8_7.NAND4F_4.B.n2 mux8_7.NAND4F_4.B.n1 10.955
R16923 mux8_7.NAND4F_4.B.n12 mux8_7.NAND4F_4.B.n9 3.67985
R16924 mux8_7.NAND4F_4.B.n9 mux8_7.NAND4F_4.B.n0 1.46835
R16925 mux8_7.NAND4F_4.B mux8_7.NAND4F_4.B.n12 0.502677
R16926 mux8_7.NAND4F_4.B.n9 mux8_7.NAND4F_4.B 0.498606
R16927 mux8_7.NAND4F_4.B mux8_7.NAND4F_4.B.n7 0.470197
R16928 mux8_7.NAND4F_5.Y.n1 mux8_7.NAND4F_5.Y.t9 1032.02
R16929 mux8_7.NAND4F_5.Y.n1 mux8_7.NAND4F_5.Y.t10 336.962
R16930 mux8_7.NAND4F_5.Y.n1 mux8_7.NAND4F_5.Y.t11 326.154
R16931 mux8_7.NAND4F_5.Y.n0 mux8_7.NAND4F_5.Y.n3 187.373
R16932 mux8_7.NAND4F_5.Y.n0 mux8_7.NAND4F_5.Y.n4 187.192
R16933 mux8_7.NAND4F_5.Y.n0 mux8_7.NAND4F_5.Y.n5 187.192
R16934 mux8_7.NAND4F_5.Y.n7 mux8_7.NAND4F_5.Y.n6 187.192
R16935 mux8_7.NAND4F_5.Y mux8_7.NAND4F_5.Y.n1 162.94
R16936 mux8_7.NAND4F_5.Y.n2 mux8_7.NAND4F_5.Y 24.4721
R16937 mux8_7.NAND4F_5.Y.n2 mux8_7.NAND4F_5.Y.t2 22.6141
R16938 mux8_7.NAND4F_5.Y.n3 mux8_7.NAND4F_5.Y.t1 20.1899
R16939 mux8_7.NAND4F_5.Y.n3 mux8_7.NAND4F_5.Y.t0 20.1899
R16940 mux8_7.NAND4F_5.Y.n4 mux8_7.NAND4F_5.Y.t5 20.1899
R16941 mux8_7.NAND4F_5.Y.n4 mux8_7.NAND4F_5.Y.t4 20.1899
R16942 mux8_7.NAND4F_5.Y.n5 mux8_7.NAND4F_5.Y.t6 20.1899
R16943 mux8_7.NAND4F_5.Y.n5 mux8_7.NAND4F_5.Y.t7 20.1899
R16944 mux8_7.NAND4F_5.Y.n6 mux8_7.NAND4F_5.Y.t3 20.1899
R16945 mux8_7.NAND4F_5.Y.n6 mux8_7.NAND4F_5.Y.t8 20.1899
R16946 mux8_7.NAND4F_5.Y mux8_7.NAND4F_5.Y.n2 0.950576
R16947 mux8_7.NAND4F_5.Y mux8_7.NAND4F_5.Y.n7 0.396904
R16948 mux8_7.NAND4F_5.Y.n7 mux8_7.NAND4F_5.Y.n0 0.358709
R16949 AND8_0.NOT8_0.A1.n2 AND8_0.NOT8_0.A1.t7 394.37
R16950 AND8_0.NOT8_0.A1.n1 AND8_0.NOT8_0.A1.t10 291.829
R16951 AND8_0.NOT8_0.A1.n1 AND8_0.NOT8_0.A1.t8 291.829
R16952 AND8_0.NOT8_0.A1.n0 AND8_0.NOT8_0.A1.n3 227.526
R16953 AND8_0.NOT8_0.A1.n0 AND8_0.NOT8_0.A1.n4 227.266
R16954 AND8_0.NOT8_0.A1.n0 AND8_0.NOT8_0.A1.n5 227.266
R16955 AND8_0.NOT8_0.A1.n1 AND8_0.NOT8_0.A1.t9 221.72
R16956 AND8_0.NOT8_0.A1.n2 AND8_0.NOT8_0.A1.n1 53.374
R16957 AND8_0.NOT8_0.A1.n0 AND8_0.NOT8_0.A1.t0 42.7824
R16958 AND8_0.NOT8_0.A1.n4 AND8_0.NOT8_0.A1.t2 30.379
R16959 AND8_0.NOT8_0.A1.n4 AND8_0.NOT8_0.A1.t5 30.379
R16960 AND8_0.NOT8_0.A1.n3 AND8_0.NOT8_0.A1.t6 30.379
R16961 AND8_0.NOT8_0.A1.n3 AND8_0.NOT8_0.A1.t4 30.379
R16962 AND8_0.NOT8_0.A1.n5 AND8_0.NOT8_0.A1.t1 30.379
R16963 AND8_0.NOT8_0.A1.n5 AND8_0.NOT8_0.A1.t3 30.379
R16964 AND8_0.NOT8_0.A1 AND8_0.NOT8_0.A1.n0 2.08054
R16965 AND8_0.NOT8_0.A1 AND8_0.NOT8_0.A1.n2 1.28475
R16966 OR8_0.S0.n1 OR8_0.S0.t6 1032.02
R16967 OR8_0.S0.n1 OR8_0.S0.t4 336.962
R16968 OR8_0.S0.n1 OR8_0.S0.t5 326.154
R16969 OR8_0.S0.n0 OR8_0.S0.t3 256.514
R16970 OR8_0.S0.n0 OR8_0.S0.n2 226.258
R16971 mux8_1.NAND4F_2.A OR8_0.S0.n1 162.952
R16972 OR8_0.NOT8_0.S0 mux8_1.A3 102.569
R16973 OR8_0.S0.n0 OR8_0.S0.t0 83.7172
R16974 OR8_0.S0.n2 OR8_0.S0.t2 30.379
R16975 OR8_0.S0.n2 OR8_0.S0.t1 30.379
R16976 mux8_1.A3 mux8_1.NAND4F_2.A 14.0763
R16977 OR8_0.NOT8_0.S0 OR8_0.S0.n0 1.88695
R16978 mux8_1.NAND4F_2.Y.n6 mux8_1.NAND4F_2.Y.t11 933.563
R16979 mux8_1.NAND4F_2.Y.n6 mux8_1.NAND4F_2.Y.t10 367.635
R16980 mux8_1.NAND4F_2.Y.n7 mux8_1.NAND4F_2.Y.t9 308.481
R16981 mux8_1.NAND4F_2.Y.n0 mux8_1.NAND4F_2.Y.n1 187.373
R16982 mux8_1.NAND4F_2.Y.n0 mux8_1.NAND4F_2.Y.n2 187.192
R16983 mux8_1.NAND4F_2.Y.n0 mux8_1.NAND4F_2.Y.n3 187.192
R16984 mux8_1.NAND4F_2.Y.n5 mux8_1.NAND4F_2.Y.n4 187.192
R16985 mux8_1.NAND4F_2.Y mux8_1.NAND4F_2.Y.n7 162.102
R16986 mux8_1.NAND4F_2.Y.n8 mux8_1.NAND4F_2.Y.t0 22.7096
R16987 mux8_1.NAND4F_2.Y.n8 mux8_1.NAND4F_2.Y 22.4285
R16988 mux8_1.NAND4F_2.Y.n1 mux8_1.NAND4F_2.Y.t4 20.1899
R16989 mux8_1.NAND4F_2.Y.n1 mux8_1.NAND4F_2.Y.t3 20.1899
R16990 mux8_1.NAND4F_2.Y.n2 mux8_1.NAND4F_2.Y.t6 20.1899
R16991 mux8_1.NAND4F_2.Y.n2 mux8_1.NAND4F_2.Y.t5 20.1899
R16992 mux8_1.NAND4F_2.Y.n3 mux8_1.NAND4F_2.Y.t7 20.1899
R16993 mux8_1.NAND4F_2.Y.n3 mux8_1.NAND4F_2.Y.t8 20.1899
R16994 mux8_1.NAND4F_2.Y.n4 mux8_1.NAND4F_2.Y.t2 20.1899
R16995 mux8_1.NAND4F_2.Y.n4 mux8_1.NAND4F_2.Y.t1 20.1899
R16996 mux8_1.NAND4F_2.Y.n7 mux8_1.NAND4F_2.Y.n6 10.955
R16997 mux8_1.NAND4F_2.Y mux8_1.NAND4F_2.Y.n8 0.799394
R16998 mux8_1.NAND4F_2.Y mux8_1.NAND4F_2.Y.n5 0.452586
R16999 mux8_1.NAND4F_2.Y.n5 mux8_1.NAND4F_2.Y.n0 0.358709
R17000 a_n15737_n5180.n2 a_n15737_n5180.t6 541.395
R17001 a_n15737_n5180.n3 a_n15737_n5180.t5 527.402
R17002 a_n15737_n5180.n2 a_n15737_n5180.t4 491.64
R17003 a_n15737_n5180.n5 a_n15737_n5180.t0 281.906
R17004 a_n15737_n5180.t1 a_n15737_n5180.n5 204.359
R17005 a_n15737_n5180.n0 a_n15737_n5180.t2 180.73
R17006 a_n15737_n5180.n1 a_n15737_n5180.t7 179.45
R17007 a_n15737_n5180.n0 a_n15737_n5180.t3 139.78
R17008 a_n15737_n5180.n4 a_n15737_n5180.n1 105.635
R17009 a_n15737_n5180.n4 a_n15737_n5180.n3 76.0005
R17010 a_n15737_n5180.n5 a_n15737_n5180.n4 67.9685
R17011 a_n15737_n5180.n3 a_n15737_n5180.n2 13.994
R17012 a_n15737_n5180.n1 a_n15737_n5180.n0 1.28015
R17013 a_n15707_n5154.n3 a_n15707_n5154.n2 121.353
R17014 a_n15707_n5154.n2 a_n15707_n5154.n1 121.001
R17015 a_n15707_n5154.n2 a_n15707_n5154.n0 120.977
R17016 a_n15707_n5154.n1 a_n15707_n5154.t0 30.462
R17017 a_n15707_n5154.n1 a_n15707_n5154.t5 30.462
R17018 a_n15707_n5154.n0 a_n15707_n5154.t2 30.462
R17019 a_n15707_n5154.n0 a_n15707_n5154.t1 30.462
R17020 a_n15707_n5154.t4 a_n15707_n5154.n3 30.462
R17021 a_n15707_n5154.n3 a_n15707_n5154.t3 30.462
R17022 right_shifter_0.buffer_4.inv_1.A.n0 right_shifter_0.buffer_4.inv_1.A.t4 393.921
R17023 right_shifter_0.buffer_4.inv_1.A.n2 right_shifter_0.buffer_4.inv_1.A.t7 291.829
R17024 right_shifter_0.buffer_4.inv_1.A.n2 right_shifter_0.buffer_4.inv_1.A.t6 291.829
R17025 right_shifter_0.buffer_4.inv_1.A.n0 right_shifter_0.buffer_4.inv_1.A.t1 256.514
R17026 right_shifter_0.buffer_4.inv_1.A.n0 right_shifter_0.buffer_4.inv_1.A.n1 226.162
R17027 right_shifter_0.buffer_4.inv_1.A.n2 right_shifter_0.buffer_4.inv_1.A.t5 221.72
R17028 right_shifter_0.buffer_4.inv_1.A.n0 right_shifter_0.buffer_4.inv_1.A.t0 83.795
R17029 right_shifter_0.buffer_4.inv_1.A.n0 right_shifter_0.buffer_4.inv_1.A.n2 53.7938
R17030 right_shifter_0.buffer_4.inv_1.A.n1 right_shifter_0.buffer_4.inv_1.A.t3 30.379
R17031 right_shifter_0.buffer_4.inv_1.A.n1 right_shifter_0.buffer_4.inv_1.A.t2 30.379
R17032 A3.n22 A3.t38 540.38
R17033 A3.n14 A3.t36 540.38
R17034 A3.n17 A3.t40 540.38
R17035 A3.n28 A3.t42 540.38
R17036 A3.n5 A3.t15 540.38
R17037 A3.n38 A3.t25 540.375
R17038 A3.n6 A3.t43 491.64
R17039 A3.n6 A3.t10 491.64
R17040 A3.n6 A3.t22 491.64
R17041 A3.n6 A3.t21 491.64
R17042 A3.n1 A3.t7 491.64
R17043 A3.n1 A3.t5 491.64
R17044 A3.n1 A3.t41 491.64
R17045 A3.n1 A3.t13 491.64
R17046 A3.n20 A3.t1 367.928
R17047 A3.n12 A3.t9 367.928
R17048 A3.n15 A3.t12 367.928
R17049 A3.n26 A3.t29 367.928
R17050 A3.n3 A3.t26 367.928
R17051 A3.n36 A3.t35 343.827
R17052 A3.n41 A3.t18 312.599
R17053 A3.n44 A3.t4 247.428
R17054 A3.n43 A3.t37 247.428
R17055 A3.n42 A3.t34 247.428
R17056 A3.n41 A3.t20 247.428
R17057 A3.n36 A3.t0 237.787
R17058 A3.n45 A3.t2 229.754
R17059 A3.n37 A3.t3 227.356
R17060 A3.n21 A3.t24 227.356
R17061 A3.n13 A3.t32 227.356
R17062 A3.n16 A3.t14 227.356
R17063 A3.n27 A3.t8 227.356
R17064 A3.n4 A3.t19 227.356
R17065 A3.n20 A3.t6 213.688
R17066 A3.n12 A3.t16 213.688
R17067 A3.n15 A3.t11 213.688
R17068 A3.n26 A3.t27 213.688
R17069 A3.n3 A3.t28 213.688
R17070 A3 A3.n2 163.036
R17071 A3.n9 A3.n8 162.867
R17072 A3 A3.n45 162.409
R17073 A3.n22 A3.n21 160.439
R17074 A3.n14 A3.n13 160.439
R17075 A3.n17 A3.n16 160.439
R17076 A3.n28 A3.n27 160.439
R17077 A3.n5 A3.n4 160.439
R17078 A3.n38 A3.n37 160.433
R17079 A3.n7 A3.t45 139.78
R17080 A3.n7 A3.t44 139.78
R17081 A3.n7 A3.t23 139.78
R17082 A3.n7 A3.t39 139.78
R17083 A3.n0 A3.t17 139.78
R17084 A3.n0 A3.t33 139.78
R17085 A3.n0 A3.t31 139.78
R17086 A3.n0 A3.t30 139.78
R17087 A3.n21 A3.n20 94.4341
R17088 A3.n13 A3.n12 94.4341
R17089 A3.n16 A3.n15 94.4341
R17090 A3.n27 A3.n26 94.4341
R17091 A3.n4 A3.n3 94.4341
R17092 A3.n45 A3.n44 91.5805
R17093 A3.n37 A3.n36 70.3341
R17094 A3.n42 A3.n41 65.1723
R17095 A3.n43 A3.n42 65.1723
R17096 A3.n44 A3.n43 65.1723
R17097 A3.n2 A3.n0 38.8368
R17098 A3.n8 A3.n7 38.6833
R17099 A3.n35 A3 31.6924
R17100 A3.n8 A3.n6 28.3986
R17101 A3.n2 A3.n1 28.2451
R17102 A3 A3.n46 18.6471
R17103 A3 A3.n10 18.1908
R17104 A3.n19 A3.n18 13.8236
R17105 A3.n46 A3 12.4204
R17106 A3.n40 A3.n39 12.4202
R17107 A3.n10 A3.n9 9.00496
R17108 A3.n35 A3.n34 6.14825
R17109 A3.n30 A3.n29 4.5005
R17110 A3 A3.n35 4.01029
R17111 A3.n46 A3.n40 3.97367
R17112 A3.n23 A3 3.91039
R17113 A3.n10 A3 3.87912
R17114 A3.n24 A3 3.67165
R17115 A3.n31 A3.n25 3.4105
R17116 A3.n33 A3.n32 3.4105
R17117 A3.n31 A3.n30 1.91502
R17118 A3.n39 A3 1.33698
R17119 A3 A3.n38 0.905186
R17120 A3 A3.n22 0.900886
R17121 A3 A3.n14 0.900886
R17122 A3 A3.n5 0.89693
R17123 A3.n29 A3.n28 0.878827
R17124 A3.n23 A3.n19 0.864715
R17125 A3.n24 A3.n23 0.825043
R17126 A3.n18 A3.n17 0.819085
R17127 A3.n25 A3.n24 0.774933
R17128 A3.n34 A3.n33 0.606532
R17129 A3.n34 A3.n11 0.18168
R17130 A3.n19 A3 0.135745
R17131 A3.n39 A3 0.11286
R17132 A3.n9 A3 0.0590664
R17133 A3.n29 A3 0.0225588
R17134 A3.n18 A3 0.012442
R17135 A3.n32 A3.n31 0.00760227
R17136 A3.n30 A3.n11 0.00735976
R17137 A3.n40 A3 0.0057809
R17138 A3.n32 A3.n11 0.00334091
R17139 A3.n33 A3.n25 0.00304054
R17140 AND8_0.NOT8_0.A3.n2 AND8_0.NOT8_0.A3.t8 394.37
R17141 AND8_0.NOT8_0.A3.n1 AND8_0.NOT8_0.A3.t7 291.829
R17142 AND8_0.NOT8_0.A3.n1 AND8_0.NOT8_0.A3.t9 291.829
R17143 AND8_0.NOT8_0.A3.n0 AND8_0.NOT8_0.A3.n3 227.526
R17144 AND8_0.NOT8_0.A3.n0 AND8_0.NOT8_0.A3.n4 227.266
R17145 AND8_0.NOT8_0.A3.n0 AND8_0.NOT8_0.A3.n5 227.266
R17146 AND8_0.NOT8_0.A3.n1 AND8_0.NOT8_0.A3.t10 221.72
R17147 AND8_0.NOT8_0.A3.n2 AND8_0.NOT8_0.A3.n1 53.374
R17148 AND8_0.NOT8_0.A3.n0 AND8_0.NOT8_0.A3.t6 42.8021
R17149 AND8_0.NOT8_0.A3.n4 AND8_0.NOT8_0.A3.t4 30.379
R17150 AND8_0.NOT8_0.A3.n4 AND8_0.NOT8_0.A3.t1 30.379
R17151 AND8_0.NOT8_0.A3.n3 AND8_0.NOT8_0.A3.t2 30.379
R17152 AND8_0.NOT8_0.A3.n3 AND8_0.NOT8_0.A3.t0 30.379
R17153 AND8_0.NOT8_0.A3.n5 AND8_0.NOT8_0.A3.t3 30.379
R17154 AND8_0.NOT8_0.A3.n5 AND8_0.NOT8_0.A3.t5 30.379
R17155 AND8_0.NOT8_0.A3 AND8_0.NOT8_0.A3.n0 2.14065
R17156 AND8_0.NOT8_0.A3 AND8_0.NOT8_0.A3.n2 1.28294
R17157 left_shifter_0.S0.n1 left_shifter_0.S0.t6 1032.02
R17158 left_shifter_0.S0.n1 left_shifter_0.S0.t5 336.962
R17159 left_shifter_0.S0.n1 left_shifter_0.S0.t4 326.154
R17160 left_shifter_0.S0.n0 left_shifter_0.S0.t2 256.89
R17161 left_shifter_0.S0.n0 left_shifter_0.S0.n2 226.635
R17162 left_shifter_0.S0 left_shifter_0.S0.n1 162.952
R17163 left_shifter_0.S0.n0 left_shifter_0.S0.t0 83.7172
R17164 left_shifter_0.S0.n2 left_shifter_0.S0.t3 30.379
R17165 left_shifter_0.S0.n2 left_shifter_0.S0.t1 30.379
R17166 left_shifter_0.S0 left_shifter_0.S0.n0 0.812762
R17167 a_n5059_1406.n0 a_n5059_1406.t5 539.788
R17168 a_n5059_1406.n1 a_n5059_1406.t2 531.496
R17169 a_n5059_1406.n0 a_n5059_1406.t4 490.034
R17170 a_n5059_1406.n5 a_n5059_1406.t0 283.788
R17171 a_n5059_1406.t1 a_n5059_1406.n5 205.489
R17172 a_n5059_1406.n2 a_n5059_1406.t3 182.625
R17173 a_n5059_1406.n3 a_n5059_1406.t6 179.054
R17174 a_n5059_1406.n2 a_n5059_1406.t7 139.78
R17175 a_n5059_1406.n4 a_n5059_1406.n3 101.368
R17176 a_n5059_1406.n5 a_n5059_1406.n4 77.9135
R17177 a_n5059_1406.n4 a_n5059_1406.n1 76.1557
R17178 a_n5059_1406.n1 a_n5059_1406.n0 8.29297
R17179 a_n5059_1406.n3 a_n5059_1406.n2 3.57087
R17180 a_n4879_2026.n7 a_n4879_2026.n1 81.2978
R17181 a_n4879_2026.n1 a_n4879_2026.n6 81.1637
R17182 a_n4879_2026.n1 a_n4879_2026.n5 81.1637
R17183 a_n4879_2026.n0 a_n4879_2026.n4 81.1637
R17184 a_n4879_2026.n0 a_n4879_2026.n3 81.1637
R17185 a_n4879_2026.n0 a_n4879_2026.n2 80.9213
R17186 a_n4879_2026.n6 a_n4879_2026.t2 11.8205
R17187 a_n4879_2026.n6 a_n4879_2026.t6 11.8205
R17188 a_n4879_2026.n5 a_n4879_2026.t0 11.8205
R17189 a_n4879_2026.n5 a_n4879_2026.t1 11.8205
R17190 a_n4879_2026.n4 a_n4879_2026.t3 11.8205
R17191 a_n4879_2026.n4 a_n4879_2026.t11 11.8205
R17192 a_n4879_2026.n3 a_n4879_2026.t8 11.8205
R17193 a_n4879_2026.n3 a_n4879_2026.t4 11.8205
R17194 a_n4879_2026.n2 a_n4879_2026.t10 11.8205
R17195 a_n4879_2026.n2 a_n4879_2026.t9 11.8205
R17196 a_n4879_2026.t7 a_n4879_2026.n7 11.8205
R17197 a_n4879_2026.n7 a_n4879_2026.t5 11.8205
R17198 a_n4879_2026.n1 a_n4879_2026.n0 0.402735
R17199 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t20 491.64
R17200 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t18 491.64
R17201 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t22 491.64
R17202 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t21 491.64
R17203 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t15 485.221
R17204 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t14 367.928
R17205 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t17 255.588
R17206 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t12 224.478
R17207 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t13 213.688
R17208 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n0 209.19
R17209 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t19 139.78
R17210 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t23 139.78
R17211 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t16 139.78
R17212 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n10 120.999
R17213 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n9 120.999
R17214 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n22 104.489
R17215 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n12 92.5005
R17216 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n18 86.2638
R17217 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n17 85.8873
R17218 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n15 85.724
R17219 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n7 84.5046
R17220 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n23 83.8907
R17221 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n17 75.0672
R17222 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n20 75.0672
R17223 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n15 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n14 73.1255
R17224 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n17 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n16 73.1255
R17225 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n19 73.1255
R17226 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n6 72.3005
R17227 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n15 68.8946
R17228 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n8 60.9797
R17229 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n13 41.9827
R17230 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t9 30.462
R17231 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t0 30.462
R17232 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t4 30.462
R17233 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t5 30.462
R17234 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t10 30.462
R17235 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t8 30.462
R17236 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n11 28.124
R17237 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n5 19.963
R17238 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n1 17.8661
R17239 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n2 17.8661
R17240 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n3 17.1217
R17241 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t7 11.8205
R17242 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t6 11.8205
R17243 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t11 11.8205
R17244 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t1 11.8205
R17245 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t2 11.8205
R17246 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t3 11.8205
R17247 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n21 9.3005
R17248 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n4 1.8615
R17249 mux8_5.NAND4F_5.Y.n1 mux8_5.NAND4F_5.Y.t9 1032.02
R17250 mux8_5.NAND4F_5.Y.n1 mux8_5.NAND4F_5.Y.t10 336.962
R17251 mux8_5.NAND4F_5.Y.n1 mux8_5.NAND4F_5.Y.t11 326.154
R17252 mux8_5.NAND4F_5.Y.n0 mux8_5.NAND4F_5.Y.n3 187.373
R17253 mux8_5.NAND4F_5.Y.n0 mux8_5.NAND4F_5.Y.n4 187.192
R17254 mux8_5.NAND4F_5.Y.n0 mux8_5.NAND4F_5.Y.n5 187.192
R17255 mux8_5.NAND4F_5.Y.n7 mux8_5.NAND4F_5.Y.n6 187.192
R17256 mux8_5.NAND4F_5.Y mux8_5.NAND4F_5.Y.n1 162.94
R17257 mux8_5.NAND4F_5.Y.n2 mux8_5.NAND4F_5.Y 24.4721
R17258 mux8_5.NAND4F_5.Y.n2 mux8_5.NAND4F_5.Y.t2 22.6141
R17259 mux8_5.NAND4F_5.Y.n3 mux8_5.NAND4F_5.Y.t0 20.1899
R17260 mux8_5.NAND4F_5.Y.n3 mux8_5.NAND4F_5.Y.t1 20.1899
R17261 mux8_5.NAND4F_5.Y.n4 mux8_5.NAND4F_5.Y.t8 20.1899
R17262 mux8_5.NAND4F_5.Y.n4 mux8_5.NAND4F_5.Y.t7 20.1899
R17263 mux8_5.NAND4F_5.Y.n5 mux8_5.NAND4F_5.Y.t5 20.1899
R17264 mux8_5.NAND4F_5.Y.n5 mux8_5.NAND4F_5.Y.t6 20.1899
R17265 mux8_5.NAND4F_5.Y.n6 mux8_5.NAND4F_5.Y.t3 20.1899
R17266 mux8_5.NAND4F_5.Y.n6 mux8_5.NAND4F_5.Y.t4 20.1899
R17267 mux8_5.NAND4F_5.Y mux8_5.NAND4F_5.Y.n2 0.950576
R17268 mux8_5.NAND4F_5.Y mux8_5.NAND4F_5.Y.n7 0.396904
R17269 mux8_5.NAND4F_5.Y.n7 mux8_5.NAND4F_5.Y.n0 0.358709
R17270 SEL3.n6 SEL3.t19 540.38
R17271 SEL3.n39 SEL3.t49 491.64
R17272 SEL3.n39 SEL3.t76 491.64
R17273 SEL3.n39 SEL3.t26 491.64
R17274 SEL3.n39 SEL3.t3 491.64
R17275 SEL3.n21 SEL3.t65 491.64
R17276 SEL3.n21 SEL3.t12 491.64
R17277 SEL3.n21 SEL3.t28 491.64
R17278 SEL3.n21 SEL3.t4 491.64
R17279 SEL3.n24 SEL3.t71 491.64
R17280 SEL3.n24 SEL3.t46 491.64
R17281 SEL3.n24 SEL3.t33 491.64
R17282 SEL3.n24 SEL3.t8 491.64
R17283 SEL3.n18 SEL3.t55 491.64
R17284 SEL3.n18 SEL3.t78 491.64
R17285 SEL3.n18 SEL3.t35 491.64
R17286 SEL3.n18 SEL3.t70 491.64
R17287 SEL3.n15 SEL3.t52 491.64
R17288 SEL3.n15 SEL3.t74 491.64
R17289 SEL3.n15 SEL3.t9 491.64
R17290 SEL3.n15 SEL3.t43 491.64
R17291 SEL3.n30 SEL3.t79 491.64
R17292 SEL3.n30 SEL3.t21 491.64
R17293 SEL3.n30 SEL3.t60 491.64
R17294 SEL3.n30 SEL3.t39 491.64
R17295 SEL3.n9 SEL3.t56 491.64
R17296 SEL3.n9 SEL3.t80 491.64
R17297 SEL3.n9 SEL3.t37 491.64
R17298 SEL3.n9 SEL3.t10 491.64
R17299 SEL3.n12 SEL3.t58 491.64
R17300 SEL3.n12 SEL3.t0 491.64
R17301 SEL3.n12 SEL3.t42 491.64
R17302 SEL3.n12 SEL3.t13 491.64
R17303 SEL3.n0 SEL3.t11 491.64
R17304 SEL3.n0 SEL3.t50 491.64
R17305 SEL3.n0 SEL3.t29 491.64
R17306 SEL3.n0 SEL3.t57 491.64
R17307 SEL3.n45 SEL3.t22 491.64
R17308 SEL3.n46 SEL3.t45 491.64
R17309 SEL3.n47 SEL3.t83 491.64
R17310 SEL3.n48 SEL3.t41 491.64
R17311 SEL3.n4 SEL3.t36 367.928
R17312 SEL3.n49 SEL3.t6 255.588
R17313 SEL3.n5 SEL3.t23 227.356
R17314 SEL3.n4 SEL3.t31 213.688
R17315 SEL3.n45 SEL3.n44 209.19
R17316 SEL3.n50 SEL3 197.833
R17317 SEL3 SEL3.n41 163.024
R17318 SEL3 SEL3.n23 163.024
R17319 SEL3 SEL3.n26 163.024
R17320 SEL3 SEL3.n20 163.024
R17321 SEL3 SEL3.n17 163.024
R17322 SEL3 SEL3.n32 163.024
R17323 SEL3 SEL3.n11 163.024
R17324 SEL3 SEL3.n14 163.024
R17325 SEL3.n3 SEL3.n2 162.852
R17326 SEL3.n6 SEL3.n5 160.439
R17327 SEL3.n40 SEL3.t16 139.78
R17328 SEL3.n40 SEL3.t75 139.78
R17329 SEL3.n40 SEL3.t40 139.78
R17330 SEL3.n40 SEL3.t66 139.78
R17331 SEL3.n22 SEL3.t17 139.78
R17332 SEL3.n22 SEL3.t77 139.78
R17333 SEL3.n22 SEL3.t59 139.78
R17334 SEL3.n22 SEL3.t5 139.78
R17335 SEL3.n25 SEL3.t20 139.78
R17336 SEL3.n25 SEL3.t82 139.78
R17337 SEL3.n25 SEL3.t63 139.78
R17338 SEL3.n25 SEL3.t38 139.78
R17339 SEL3.n19 SEL3.t24 139.78
R17340 SEL3.n19 SEL3.t62 139.78
R17341 SEL3.n19 SEL3.t47 139.78
R17342 SEL3.n19 SEL3.t68 139.78
R17343 SEL3.n16 SEL3.t1 139.78
R17344 SEL3.n16 SEL3.t32 139.78
R17345 SEL3.n16 SEL3.t44 139.78
R17346 SEL3.n16 SEL3.t64 139.78
R17347 SEL3.n31 SEL3.t54 139.78
R17348 SEL3.n31 SEL3.t27 139.78
R17349 SEL3.n31 SEL3.t69 139.78
R17350 SEL3.n31 SEL3.t14 139.78
R17351 SEL3.n10 SEL3.t25 139.78
R17352 SEL3.n10 SEL3.t2 139.78
R17353 SEL3.n10 SEL3.t48 139.78
R17354 SEL3.n10 SEL3.t72 139.78
R17355 SEL3.n13 SEL3.t30 139.78
R17356 SEL3.n13 SEL3.t7 139.78
R17357 SEL3.n13 SEL3.t51 139.78
R17358 SEL3.n13 SEL3.t73 139.78
R17359 SEL3.n1 SEL3.t81 139.78
R17360 SEL3.n1 SEL3.t18 139.78
R17361 SEL3.n1 SEL3.t61 139.78
R17362 SEL3.n1 SEL3.t15 139.78
R17363 SEL3.n44 SEL3.t53 139.78
R17364 SEL3.n44 SEL3.t34 139.78
R17365 SEL3.n44 SEL3.t67 139.78
R17366 SEL3.n5 SEL3.n4 94.4341
R17367 SEL3.n41 SEL3.n40 38.6833
R17368 SEL3.n23 SEL3.n22 38.6833
R17369 SEL3.n26 SEL3.n25 38.6833
R17370 SEL3.n20 SEL3.n19 38.6833
R17371 SEL3.n17 SEL3.n16 38.6833
R17372 SEL3.n32 SEL3.n31 38.6833
R17373 SEL3.n11 SEL3.n10 38.6833
R17374 SEL3.n14 SEL3.n13 38.6833
R17375 SEL3.n2 SEL3.n1 38.6833
R17376 SEL3.n41 SEL3.n39 28.3986
R17377 SEL3.n23 SEL3.n21 28.3986
R17378 SEL3.n26 SEL3.n24 28.3986
R17379 SEL3.n20 SEL3.n18 28.3986
R17380 SEL3.n17 SEL3.n15 28.3986
R17381 SEL3.n32 SEL3.n30 28.3986
R17382 SEL3.n11 SEL3.n9 28.3986
R17383 SEL3.n14 SEL3.n12 28.3986
R17384 SEL3.n2 SEL3.n0 28.3986
R17385 SEL3 SEL3.n49 27.4136
R17386 SEL3.n50 SEL3 18.4979
R17387 SEL3.n46 SEL3.n45 17.8661
R17388 SEL3.n47 SEL3.n46 17.8661
R17389 SEL3.n48 SEL3.n47 17.1217
R17390 SEL3 SEL3.n43 12.7036
R17391 SEL3 SEL3.n8 10.7052
R17392 SEL3.n8 SEL3.n3 5.09176
R17393 SEL3.n8 SEL3.n7 4.19292
R17394 SEL3.n43 SEL3 3.5788
R17395 SEL3.n27 SEL3 3.37473
R17396 SEL3.n35 SEL3 2.46517
R17397 SEL3.n29 SEL3 2.45291
R17398 SEL3.n36 SEL3 2.44378
R17399 SEL3.n28 SEL3 2.43697
R17400 SEL3.n37 SEL3.n36 2.38603
R17401 SEL3.n34 SEL3.n33 2.3781
R17402 SEL3.n36 SEL3.n35 2.35407
R17403 SEL3.n29 SEL3.n28 2.29921
R17404 SEL3.n28 SEL3.n27 2.27959
R17405 SEL3.n35 SEL3.n34 2.27907
R17406 SEL3.n34 SEL3.n29 2.27729
R17407 SEL3.n38 SEL3.n37 2.2505
R17408 SEL3.n49 SEL3.n48 1.8615
R17409 SEL3.n27 SEL3 1.17427
R17410 SEL3 SEL3.n50 1.01205
R17411 SEL3.n33 SEL3 0.903207
R17412 SEL3.n7 SEL3.n6 0.794268
R17413 SEL3.n43 SEL3.n42 0.556214
R17414 SEL3.n42 SEL3.n38 0.43225
R17415 SEL3.n42 SEL3 0.319636
R17416 SEL3.n38 SEL3 0.200821
R17417 SEL3.n37 SEL3 0.107331
R17418 SEL3.n7 SEL3 0.107118
R17419 SEL3.n3 SEL3 0.0730524
R17420 SEL3.n33 SEL3 0.0633571
R17421 a_n7676_3190.n2 a_n7676_3190.t3 541.395
R17422 a_n7676_3190.n3 a_n7676_3190.t5 527.402
R17423 a_n7676_3190.n2 a_n7676_3190.t7 491.64
R17424 a_n7676_3190.n5 a_n7676_3190.t0 281.906
R17425 a_n7676_3190.t1 a_n7676_3190.n5 204.359
R17426 a_n7676_3190.n0 a_n7676_3190.t2 180.73
R17427 a_n7676_3190.n1 a_n7676_3190.t6 179.45
R17428 a_n7676_3190.n0 a_n7676_3190.t4 139.78
R17429 a_n7676_3190.n4 a_n7676_3190.n1 105.635
R17430 a_n7676_3190.n4 a_n7676_3190.n3 76.0005
R17431 a_n7676_3190.n5 a_n7676_3190.n4 67.9685
R17432 a_n7676_3190.n3 a_n7676_3190.n2 13.994
R17433 a_n7676_3190.n1 a_n7676_3190.n0 1.28015
R17434 a_n8549_n5154.n2 a_n8549_n5154.n1 121.353
R17435 a_n8549_n5154.n2 a_n8549_n5154.n0 121.353
R17436 a_n8549_n5154.n3 a_n8549_n5154.n2 121.001
R17437 a_n8549_n5154.n1 a_n8549_n5154.t4 30.462
R17438 a_n8549_n5154.n1 a_n8549_n5154.t5 30.462
R17439 a_n8549_n5154.n0 a_n8549_n5154.t1 30.462
R17440 a_n8549_n5154.n0 a_n8549_n5154.t0 30.462
R17441 a_n8549_n5154.t2 a_n8549_n5154.n3 30.462
R17442 a_n8549_n5154.n3 a_n8549_n5154.t3 30.462
R17443 a_8496_n25478.t0 a_8496_n25478.t1 9.9005
R17444 a_8592_n25478.t0 a_8592_n25478.t1 9.9005
R17445 NOT8_0.S4.n1 NOT8_0.S4.t5 1032.02
R17446 NOT8_0.S4.n1 NOT8_0.S4.t6 336.962
R17447 NOT8_0.S4.n1 NOT8_0.S4.t4 326.154
R17448 NOT8_0.S4.n0 NOT8_0.S4.t1 256.514
R17449 NOT8_0.S4.n0 NOT8_0.S4.n2 226.258
R17450 NOT8_0.S4 NOT8_0.S4.n1 162.952
R17451 NOT8_0.S4.n0 NOT8_0.S4.t0 83.7172
R17452 NOT8_0.S4.n2 NOT8_0.S4.t3 30.379
R17453 NOT8_0.S4.n2 NOT8_0.S4.t2 30.379
R17454 NOT8_0.S4 NOT8_0.S4.n0 1.9182
R17455 mux8_5.NAND4F_7.Y.n2 mux8_5.NAND4F_7.Y.t11 1388.16
R17456 mux8_5.NAND4F_7.Y.n2 mux8_5.NAND4F_7.Y.t10 350.839
R17457 mux8_5.NAND4F_7.Y.n3 mux8_5.NAND4F_7.Y.t9 308.481
R17458 mux8_5.NAND4F_7.Y.n1 mux8_5.NAND4F_7.Y.n4 187.373
R17459 mux8_5.NAND4F_7.Y.n1 mux8_5.NAND4F_7.Y.n5 187.192
R17460 mux8_5.NAND4F_7.Y.n1 mux8_5.NAND4F_7.Y.n6 187.192
R17461 mux8_5.NAND4F_7.Y.n0 mux8_5.NAND4F_7.Y.n7 187.192
R17462 mux8_5.NAND4F_7.Y mux8_5.NAND4F_7.Y.n3 161.492
R17463 mux8_5.NAND4F_7.Y.n3 mux8_5.NAND4F_7.Y.n2 27.752
R17464 mux8_5.NAND4F_7.Y mux8_5.NAND4F_7.Y.t4 23.5642
R17465 mux8_5.NAND4F_7.Y.n4 mux8_5.NAND4F_7.Y.t1 20.1899
R17466 mux8_5.NAND4F_7.Y.n4 mux8_5.NAND4F_7.Y.t0 20.1899
R17467 mux8_5.NAND4F_7.Y.n5 mux8_5.NAND4F_7.Y.t3 20.1899
R17468 mux8_5.NAND4F_7.Y.n5 mux8_5.NAND4F_7.Y.t2 20.1899
R17469 mux8_5.NAND4F_7.Y.n6 mux8_5.NAND4F_7.Y.t8 20.1899
R17470 mux8_5.NAND4F_7.Y.n6 mux8_5.NAND4F_7.Y.t7 20.1899
R17471 mux8_5.NAND4F_7.Y.n7 mux8_5.NAND4F_7.Y.t5 20.1899
R17472 mux8_5.NAND4F_7.Y.n7 mux8_5.NAND4F_7.Y.t6 20.1899
R17473 mux8_5.NAND4F_7.Y mux8_5.NAND4F_7.Y.n0 0.472662
R17474 mux8_5.NAND4F_7.Y.n0 mux8_5.NAND4F_7.Y.n1 0.358709
R17475 mux8_4.NAND4F_6.Y.n1 mux8_4.NAND4F_6.Y.t10 933.563
R17476 mux8_4.NAND4F_6.Y.n1 mux8_4.NAND4F_6.Y.t11 367.635
R17477 mux8_4.NAND4F_6.Y.n2 mux8_4.NAND4F_6.Y.t9 308.481
R17478 mux8_4.NAND4F_6.Y.n0 mux8_4.NAND4F_6.Y.n4 187.373
R17479 mux8_4.NAND4F_6.Y.n0 mux8_4.NAND4F_6.Y.n5 187.192
R17480 mux8_4.NAND4F_6.Y.n0 mux8_4.NAND4F_6.Y.n6 187.192
R17481 mux8_4.NAND4F_6.Y.n8 mux8_4.NAND4F_6.Y.n7 187.192
R17482 mux8_4.NAND4F_6.Y mux8_4.NAND4F_6.Y.n2 162.047
R17483 mux8_4.NAND4F_6.Y.n3 mux8_4.NAND4F_6.Y.t2 22.7831
R17484 mux8_4.NAND4F_6.Y.n3 mux8_4.NAND4F_6.Y 22.171
R17485 mux8_4.NAND4F_6.Y.n4 mux8_4.NAND4F_6.Y.t1 20.1899
R17486 mux8_4.NAND4F_6.Y.n4 mux8_4.NAND4F_6.Y.t0 20.1899
R17487 mux8_4.NAND4F_6.Y.n5 mux8_4.NAND4F_6.Y.t6 20.1899
R17488 mux8_4.NAND4F_6.Y.n5 mux8_4.NAND4F_6.Y.t5 20.1899
R17489 mux8_4.NAND4F_6.Y.n6 mux8_4.NAND4F_6.Y.t7 20.1899
R17490 mux8_4.NAND4F_6.Y.n6 mux8_4.NAND4F_6.Y.t8 20.1899
R17491 mux8_4.NAND4F_6.Y.n7 mux8_4.NAND4F_6.Y.t3 20.1899
R17492 mux8_4.NAND4F_6.Y.n7 mux8_4.NAND4F_6.Y.t4 20.1899
R17493 mux8_4.NAND4F_6.Y.n2 mux8_4.NAND4F_6.Y.n1 10.955
R17494 mux8_4.NAND4F_6.Y mux8_4.NAND4F_6.Y.n3 0.781576
R17495 mux8_4.NAND4F_6.Y mux8_4.NAND4F_6.Y.n8 0.396904
R17496 mux8_4.NAND4F_6.Y.n8 mux8_4.NAND4F_6.Y.n0 0.358709
R17497 mux8_4.NAND4F_9.Y.n1 mux8_4.NAND4F_9.Y.t11 312.599
R17498 mux8_4.NAND4F_9.Y.n4 mux8_4.NAND4F_9.Y.t10 247.428
R17499 mux8_4.NAND4F_9.Y.n1 mux8_4.NAND4F_9.Y.t13 247.428
R17500 mux8_4.NAND4F_9.Y.n2 mux8_4.NAND4F_9.Y.t14 247.428
R17501 mux8_4.NAND4F_9.Y.n3 mux8_4.NAND4F_9.Y.t9 247.428
R17502 mux8_4.NAND4F_9.Y.n5 mux8_4.NAND4F_9.Y.t12 229.754
R17503 mux8_4.NAND4F_9.Y.n0 mux8_4.NAND4F_9.Y.n6 187.373
R17504 mux8_4.NAND4F_9.Y.n0 mux8_4.NAND4F_9.Y.n7 187.192
R17505 mux8_4.NAND4F_9.Y.n0 mux8_4.NAND4F_9.Y.n8 187.192
R17506 mux8_4.NAND4F_9.Y.n10 mux8_4.NAND4F_9.Y.n9 187.192
R17507 mux8_4.NAND4F_9.Y mux8_4.NAND4F_9.Y.n5 162.275
R17508 mux8_4.NAND4F_9.Y.n5 mux8_4.NAND4F_9.Y.n4 91.5805
R17509 mux8_4.NAND4F_9.Y.n2 mux8_4.NAND4F_9.Y.n1 65.1723
R17510 mux8_4.NAND4F_9.Y.n3 mux8_4.NAND4F_9.Y.n2 65.1723
R17511 mux8_4.NAND4F_9.Y.n4 mux8_4.NAND4F_9.Y.n3 65.1723
R17512 mux8_4.NAND4F_9.Y mux8_4.NAND4F_9.Y.t0 22.6141
R17513 mux8_4.NAND4F_9.Y.n6 mux8_4.NAND4F_9.Y.t5 20.1899
R17514 mux8_4.NAND4F_9.Y.n6 mux8_4.NAND4F_9.Y.t6 20.1899
R17515 mux8_4.NAND4F_9.Y.n7 mux8_4.NAND4F_9.Y.t7 20.1899
R17516 mux8_4.NAND4F_9.Y.n7 mux8_4.NAND4F_9.Y.t8 20.1899
R17517 mux8_4.NAND4F_9.Y.n8 mux8_4.NAND4F_9.Y.t3 20.1899
R17518 mux8_4.NAND4F_9.Y.n8 mux8_4.NAND4F_9.Y.t4 20.1899
R17519 mux8_4.NAND4F_9.Y.n9 mux8_4.NAND4F_9.Y.t2 20.1899
R17520 mux8_4.NAND4F_9.Y.n9 mux8_4.NAND4F_9.Y.t1 20.1899
R17521 mux8_4.NAND4F_9.Y mux8_4.NAND4F_9.Y.n10 0.396904
R17522 mux8_4.NAND4F_9.Y.n10 mux8_4.NAND4F_9.Y.n0 0.358709
R17523 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t7 540.38
R17524 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t13 491.64
R17525 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t12 491.64
R17526 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t14 491.64
R17527 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t15 491.64
R17528 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t17 367.928
R17529 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n1 227.526
R17530 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t18 227.356
R17531 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n3 227.266
R17532 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n2 227.266
R17533 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t16 213.688
R17534 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n6 162.852
R17535 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n8 160.439
R17536 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t10 139.78
R17537 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t11 139.78
R17538 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t9 139.78
R17539 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t8 139.78
R17540 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n7 94.4341
R17541 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t5 42.7831
R17542 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n5 38.6833
R17543 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t4 30.379
R17544 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t3 30.379
R17545 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t2 30.379
R17546 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t0 30.379
R17547 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t6 30.379
R17548 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t1 30.379
R17549 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n4 28.3986
R17550 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n0 18.8832
R17551 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n10 11.2587
R17552 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT 5.09176
R17553 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT 4.19292
R17554 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n9 0.794268
R17555 a_n19187_n12716.t0 a_n19187_n12716.t1 19.8005
R17556 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t8 485.221
R17557 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t10 367.928
R17558 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n5 227.526
R17559 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n6 227.266
R17560 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n4 227.266
R17561 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t7 224.478
R17562 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t9 213.688
R17563 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n2 84.5046
R17564 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n1 72.3005
R17565 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n3 61.0566
R17566 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t3 42.7747
R17567 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t4 30.379
R17568 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t0 30.379
R17569 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t5 30.379
R17570 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t6 30.379
R17571 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t1 30.379
R17572 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.t2 30.379
R17573 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A.n0 0.583137
R17574 a_n18422_n8419.n2 a_n18422_n8419.n0 121.353
R17575 a_n18422_n8419.n3 a_n18422_n8419.n2 121.353
R17576 a_n18422_n8419.n2 a_n18422_n8419.n1 121.001
R17577 a_n18422_n8419.n0 a_n18422_n8419.t1 30.462
R17578 a_n18422_n8419.n0 a_n18422_n8419.t2 30.462
R17579 a_n18422_n8419.n1 a_n18422_n8419.t5 30.462
R17580 a_n18422_n8419.n1 a_n18422_n8419.t0 30.462
R17581 a_n18422_n8419.t4 a_n18422_n8419.n3 30.462
R17582 a_n18422_n8419.n3 a_n18422_n8419.t3 30.462
R17583 B1.n17 B1.t9 540.38
R17584 B1.n10 B1.t40 540.38
R17585 B1.n6 B1.t53 491.64
R17586 B1.n5 B1.t28 491.64
R17587 B1.n4 B1.t18 491.64
R17588 B1.n3 B1.t4 491.64
R17589 B1.n39 B1.t1 491.64
R17590 B1.n38 B1.t21 491.64
R17591 B1.n37 B1.t0 491.64
R17592 B1.n36 B1.t51 491.64
R17593 B1.n26 B1.t10 485.443
R17594 B1.n20 B1.t15 485.221
R17595 B1.n13 B1.t43 485.221
R17596 B1.n43 B1.t41 394.37
R17597 B1.n46 B1.t44 394.37
R17598 B1.n1 B1.t47 394.37
R17599 B1.n29 B1.t45 379.173
R17600 B1.n15 B1.t14 367.928
R17601 B1.n18 B1.t3 367.928
R17602 B1.n8 B1.t37 367.928
R17603 B1.n11 B1.t30 367.928
R17604 B1.n24 B1.t35 343.827
R17605 B1.n30 B1.t34 312.599
R17606 B1.n42 B1.t20 291.829
R17607 B1.n42 B1.t17 291.829
R17608 B1.n45 B1.t5 291.829
R17609 B1.n45 B1.t29 291.829
R17610 B1.n0 B1.t12 291.829
R17611 B1.n0 B1.t11 291.829
R17612 B1.n7 B1.t48 255.588
R17613 B1.n40 B1.t26 255.588
R17614 B1.n30 B1.t16 247.428
R17615 B1.n31 B1.t13 247.428
R17616 B1.n32 B1.t50 247.428
R17617 B1.n29 B1.t46 247.428
R17618 B1.n24 B1.t38 237.787
R17619 B1.n16 B1.t32 227.356
R17620 B1.n9 B1.t6 227.356
R17621 B1.n25 B1.t2 224.478
R17622 B1.n19 B1.t27 224.478
R17623 B1.n12 B1.t39 224.478
R17624 B1.n42 B1.t23 221.72
R17625 B1.n45 B1.t8 221.72
R17626 B1.n0 B1.t7 221.72
R17627 B1.n15 B1.t33 213.688
R17628 B1.n18 B1.t25 213.688
R17629 B1.n8 B1.t42 213.688
R17630 B1.n11 B1.t36 213.688
R17631 B1.n36 B1.n35 209.407
R17632 B1.n3 B1.n2 209.19
R17633 B1 B1.n33 162.139
R17634 B1.n17 B1.n16 160.439
R17635 B1.n10 B1.n9 160.439
R17636 B1.n2 B1.t24 139.78
R17637 B1.n2 B1.t31 139.78
R17638 B1.n2 B1.t49 139.78
R17639 B1.n35 B1.t19 139.78
R17640 B1.n35 B1.t22 139.78
R17641 B1.n35 B1.t52 139.78
R17642 B1.n16 B1.n15 94.4341
R17643 B1.n9 B1.n8 94.4341
R17644 B1.n20 B1.n19 84.5046
R17645 B1.n13 B1.n12 84.5046
R17646 B1.n26 B1.n25 83.8438
R17647 B1.n19 B1.n18 72.3005
R17648 B1.n12 B1.n11 72.3005
R17649 B1.n32 B1.n31 65.1723
R17650 B1.n31 B1.n30 65.1723
R17651 B1 B1.n13 61.056
R17652 B1 B1.n20 61.0525
R17653 B1 B1.n26 61.0461
R17654 B1.n43 B1.n42 53.374
R17655 B1.n46 B1.n45 53.374
R17656 B1.n1 B1.n0 53.374
R17657 B1.n25 B1.n24 48.2005
R17658 B1.n23 B1 34.7047
R17659 B1.n33 B1.n32 33.2653
R17660 B1.n33 B1.n29 31.9075
R17661 B1 B1.n40 27.4136
R17662 B1.n5 B1.n4 17.8661
R17663 B1.n4 B1.n3 17.8661
R17664 B1.n37 B1.n36 17.8661
R17665 B1.n38 B1.n37 17.8661
R17666 B1.n6 B1.n5 17.1217
R17667 B1.n39 B1.n38 17.1217
R17668 B1.n49 B1.n48 14.1743
R17669 B1.n34 B1 12.5765
R17670 B1.n44 B1 12.4656
R17671 B1.n41 B1 12.4272
R17672 B1.n28 B1.n27 12.4105
R17673 B1.n48 B1.n47 12.4105
R17674 B1 B1.n7 11.1665
R17675 B1 B1.n23 8.01419
R17676 B1.n34 B1.n28 4.54318
R17677 B1.n23 B1 4.53613
R17678 B1.n41 B1.n34 4.41328
R17679 B1.n44 B1.n41 4.10256
R17680 B1.n22 B1.n14 3.84894
R17681 B1.n48 B1.n44 2.84792
R17682 B1.n22 B1.n21 2.2505
R17683 B1.n7 B1.n6 1.8615
R17684 B1.n40 B1.n39 1.8615
R17685 B1.n27 B1 1.19089
R17686 B1 B1.n43 1.18065
R17687 B1 B1.n17 0.900886
R17688 B1 B1.n10 0.900886
R17689 B1.n49 B1.n1 0.739916
R17690 B1.n21 B1 0.736713
R17691 B1.n14 B1 0.734379
R17692 B1.n47 B1.n46 0.729374
R17693 B1.n21 B1 0.379176
R17694 B1.n14 B1 0.369489
R17695 B1.n47 B1 0.0893554
R17696 B1.n27 B1 0.0890417
R17697 B1 B1.n49 0.0788133
R17698 B1 B1.n22 0.0490197
R17699 B1.n28 B1 0.0159756
R17700 a_n12314_n18115.n7 a_n12314_n18115.n1 81.2978
R17701 a_n12314_n18115.n0 a_n12314_n18115.n3 81.1637
R17702 a_n12314_n18115.n0 a_n12314_n18115.n4 81.1637
R17703 a_n12314_n18115.n1 a_n12314_n18115.n5 81.1637
R17704 a_n12314_n18115.n1 a_n12314_n18115.n6 81.1637
R17705 a_n12314_n18115.n0 a_n12314_n18115.n2 80.9213
R17706 a_n12314_n18115.n2 a_n12314_n18115.t6 11.8205
R17707 a_n12314_n18115.n2 a_n12314_n18115.t8 11.8205
R17708 a_n12314_n18115.n3 a_n12314_n18115.t7 11.8205
R17709 a_n12314_n18115.n3 a_n12314_n18115.t3 11.8205
R17710 a_n12314_n18115.n4 a_n12314_n18115.t4 11.8205
R17711 a_n12314_n18115.n4 a_n12314_n18115.t5 11.8205
R17712 a_n12314_n18115.n5 a_n12314_n18115.t9 11.8205
R17713 a_n12314_n18115.n5 a_n12314_n18115.t10 11.8205
R17714 a_n12314_n18115.n6 a_n12314_n18115.t11 11.8205
R17715 a_n12314_n18115.n6 a_n12314_n18115.t0 11.8205
R17716 a_n12314_n18115.t2 a_n12314_n18115.n7 11.8205
R17717 a_n12314_n18115.n7 a_n12314_n18115.t1 11.8205
R17718 a_n12314_n18115.n1 a_n12314_n18115.n0 0.402735
R17719 mux8_1.NAND4F_4.B.n10 mux8_1.NAND4F_4.B.t13 933.563
R17720 mux8_1.NAND4F_4.B.n5 mux8_1.NAND4F_4.B.t7 933.563
R17721 mux8_1.NAND4F_4.B.n3 mux8_1.NAND4F_4.B.t8 933.563
R17722 mux8_1.NAND4F_4.B.n1 mux8_1.NAND4F_4.B.t14 933.563
R17723 mux8_1.NAND4F_4.B.n10 mux8_1.NAND4F_4.B.t6 367.635
R17724 mux8_1.NAND4F_4.B.n5 mux8_1.NAND4F_4.B.t5 367.635
R17725 mux8_1.NAND4F_4.B.n3 mux8_1.NAND4F_4.B.t11 367.635
R17726 mux8_1.NAND4F_4.B.n1 mux8_1.NAND4F_4.B.t12 367.635
R17727 mux8_1.NAND4F_4.B.n11 mux8_1.NAND4F_4.B.t4 308.481
R17728 mux8_1.NAND4F_4.B.n6 mux8_1.NAND4F_4.B.t15 308.481
R17729 mux8_1.NAND4F_4.B.n4 mux8_1.NAND4F_4.B.t9 308.481
R17730 mux8_1.NAND4F_4.B.n2 mux8_1.NAND4F_4.B.t10 308.481
R17731 mux8_1.NAND4F_4.B.n0 mux8_1.NAND4F_4.B.t2 256.514
R17732 mux8_1.NAND4F_4.B.n0 mux8_1.NAND4F_4.B.n8 226.258
R17733 mux8_1.NAND4F_4.B mux8_1.NAND4F_4.B.n2 162.173
R17734 mux8_1.NAND4F_4.B mux8_1.NAND4F_4.B.n6 162.137
R17735 mux8_1.NAND4F_4.B mux8_1.NAND4F_4.B.n11 162.117
R17736 mux8_1.NAND4F_4.B.n7 mux8_1.NAND4F_4.B.n4 161.703
R17737 mux8_1.NAND4F_4.B.n0 mux8_1.NAND4F_4.B.t0 83.7172
R17738 mux8_1.NAND4F_4.B.n8 mux8_1.NAND4F_4.B.t1 30.379
R17739 mux8_1.NAND4F_4.B.n8 mux8_1.NAND4F_4.B.t3 30.379
R17740 mux8_1.NAND4F_4.B.n12 mux8_1.NAND4F_4.B 24.8912
R17741 mux8_1.NAND4F_4.B.n7 mux8_1.NAND4F_4.B 21.6618
R17742 mux8_1.NAND4F_4.B.n11 mux8_1.NAND4F_4.B.n10 10.955
R17743 mux8_1.NAND4F_4.B.n6 mux8_1.NAND4F_4.B.n5 10.955
R17744 mux8_1.NAND4F_4.B.n4 mux8_1.NAND4F_4.B.n3 10.955
R17745 mux8_1.NAND4F_4.B.n2 mux8_1.NAND4F_4.B.n1 10.955
R17746 mux8_1.NAND4F_4.B.n12 mux8_1.NAND4F_4.B.n9 3.67985
R17747 mux8_1.NAND4F_4.B.n9 mux8_1.NAND4F_4.B.n0 1.46835
R17748 mux8_1.NAND4F_4.B mux8_1.NAND4F_4.B.n12 0.502677
R17749 mux8_1.NAND4F_4.B.n9 mux8_1.NAND4F_4.B 0.498606
R17750 mux8_1.NAND4F_4.B mux8_1.NAND4F_4.B.n7 0.470197
R17751 mux8_1.NAND4F_1.Y.n2 mux8_1.NAND4F_1.Y.t9 978.795
R17752 mux8_1.NAND4F_1.Y.n1 mux8_1.NAND4F_1.Y.t11 308.481
R17753 mux8_1.NAND4F_1.Y.n1 mux8_1.NAND4F_1.Y.t10 308.481
R17754 mux8_1.NAND4F_1.Y.n0 mux8_1.NAND4F_1.Y.n3 187.373
R17755 mux8_1.NAND4F_1.Y.n0 mux8_1.NAND4F_1.Y.n4 187.192
R17756 mux8_1.NAND4F_1.Y.n0 mux8_1.NAND4F_1.Y.n5 187.192
R17757 mux8_1.NAND4F_1.Y.n7 mux8_1.NAND4F_1.Y.n6 187.192
R17758 mux8_1.NAND4F_1.Y mux8_1.NAND4F_1.Y.n2 161.84
R17759 mux8_1.NAND4F_1.Y mux8_1.NAND4F_1.Y.t4 23.4335
R17760 mux8_1.NAND4F_1.Y.n3 mux8_1.NAND4F_1.Y.t0 20.1899
R17761 mux8_1.NAND4F_1.Y.n3 mux8_1.NAND4F_1.Y.t1 20.1899
R17762 mux8_1.NAND4F_1.Y.n4 mux8_1.NAND4F_1.Y.t3 20.1899
R17763 mux8_1.NAND4F_1.Y.n4 mux8_1.NAND4F_1.Y.t2 20.1899
R17764 mux8_1.NAND4F_1.Y.n5 mux8_1.NAND4F_1.Y.t7 20.1899
R17765 mux8_1.NAND4F_1.Y.n5 mux8_1.NAND4F_1.Y.t8 20.1899
R17766 mux8_1.NAND4F_1.Y.n6 mux8_1.NAND4F_1.Y.t5 20.1899
R17767 mux8_1.NAND4F_1.Y.n6 mux8_1.NAND4F_1.Y.t6 20.1899
R17768 mux8_1.NAND4F_1.Y.n2 mux8_1.NAND4F_1.Y.n1 11.0463
R17769 mux8_1.NAND4F_1.Y mux8_1.NAND4F_1.Y.n7 0.527586
R17770 mux8_1.NAND4F_1.Y.n7 mux8_1.NAND4F_1.Y.n0 0.358709
R17771 mux8_1.NAND4F_7.Y.n2 mux8_1.NAND4F_7.Y.t10 1388.16
R17772 mux8_1.NAND4F_7.Y.n2 mux8_1.NAND4F_7.Y.t11 350.839
R17773 mux8_1.NAND4F_7.Y.n3 mux8_1.NAND4F_7.Y.t9 308.481
R17774 mux8_1.NAND4F_7.Y.n1 mux8_1.NAND4F_7.Y.n4 187.373
R17775 mux8_1.NAND4F_7.Y.n1 mux8_1.NAND4F_7.Y.n5 187.192
R17776 mux8_1.NAND4F_7.Y.n1 mux8_1.NAND4F_7.Y.n6 187.192
R17777 mux8_1.NAND4F_7.Y.n0 mux8_1.NAND4F_7.Y.n7 187.192
R17778 mux8_1.NAND4F_7.Y mux8_1.NAND4F_7.Y.n3 161.492
R17779 mux8_1.NAND4F_7.Y.n3 mux8_1.NAND4F_7.Y.n2 27.752
R17780 mux8_1.NAND4F_7.Y mux8_1.NAND4F_7.Y.t5 23.5642
R17781 mux8_1.NAND4F_7.Y.n4 mux8_1.NAND4F_7.Y.t0 20.1899
R17782 mux8_1.NAND4F_7.Y.n4 mux8_1.NAND4F_7.Y.t1 20.1899
R17783 mux8_1.NAND4F_7.Y.n5 mux8_1.NAND4F_7.Y.t3 20.1899
R17784 mux8_1.NAND4F_7.Y.n5 mux8_1.NAND4F_7.Y.t2 20.1899
R17785 mux8_1.NAND4F_7.Y.n6 mux8_1.NAND4F_7.Y.t8 20.1899
R17786 mux8_1.NAND4F_7.Y.n6 mux8_1.NAND4F_7.Y.t7 20.1899
R17787 mux8_1.NAND4F_7.Y.n7 mux8_1.NAND4F_7.Y.t6 20.1899
R17788 mux8_1.NAND4F_7.Y.n7 mux8_1.NAND4F_7.Y.t4 20.1899
R17789 mux8_1.NAND4F_7.Y mux8_1.NAND4F_7.Y.n0 0.472662
R17790 mux8_1.NAND4F_7.Y.n0 mux8_1.NAND4F_7.Y.n1 0.358709
R17791 mux8_1.NAND4F_9.Y.n1 mux8_1.NAND4F_9.Y.t13 312.599
R17792 mux8_1.NAND4F_9.Y.n4 mux8_1.NAND4F_9.Y.t9 247.428
R17793 mux8_1.NAND4F_9.Y.n1 mux8_1.NAND4F_9.Y.t12 247.428
R17794 mux8_1.NAND4F_9.Y.n2 mux8_1.NAND4F_9.Y.t11 247.428
R17795 mux8_1.NAND4F_9.Y.n3 mux8_1.NAND4F_9.Y.t10 247.428
R17796 mux8_1.NAND4F_9.Y.n5 mux8_1.NAND4F_9.Y.t14 229.754
R17797 mux8_1.NAND4F_9.Y.n0 mux8_1.NAND4F_9.Y.n6 187.373
R17798 mux8_1.NAND4F_9.Y.n0 mux8_1.NAND4F_9.Y.n7 187.192
R17799 mux8_1.NAND4F_9.Y.n0 mux8_1.NAND4F_9.Y.n8 187.192
R17800 mux8_1.NAND4F_9.Y.n10 mux8_1.NAND4F_9.Y.n9 187.192
R17801 mux8_1.NAND4F_9.Y mux8_1.NAND4F_9.Y.n5 162.275
R17802 mux8_1.NAND4F_9.Y.n5 mux8_1.NAND4F_9.Y.n4 91.5805
R17803 mux8_1.NAND4F_9.Y.n2 mux8_1.NAND4F_9.Y.n1 65.1723
R17804 mux8_1.NAND4F_9.Y.n3 mux8_1.NAND4F_9.Y.n2 65.1723
R17805 mux8_1.NAND4F_9.Y.n4 mux8_1.NAND4F_9.Y.n3 65.1723
R17806 mux8_1.NAND4F_9.Y mux8_1.NAND4F_9.Y.t4 22.6141
R17807 mux8_1.NAND4F_9.Y.n6 mux8_1.NAND4F_9.Y.t7 20.1899
R17808 mux8_1.NAND4F_9.Y.n6 mux8_1.NAND4F_9.Y.t8 20.1899
R17809 mux8_1.NAND4F_9.Y.n7 mux8_1.NAND4F_9.Y.t5 20.1899
R17810 mux8_1.NAND4F_9.Y.n7 mux8_1.NAND4F_9.Y.t6 20.1899
R17811 mux8_1.NAND4F_9.Y.n8 mux8_1.NAND4F_9.Y.t0 20.1899
R17812 mux8_1.NAND4F_9.Y.n8 mux8_1.NAND4F_9.Y.t1 20.1899
R17813 mux8_1.NAND4F_9.Y.n9 mux8_1.NAND4F_9.Y.t3 20.1899
R17814 mux8_1.NAND4F_9.Y.n9 mux8_1.NAND4F_9.Y.t2 20.1899
R17815 mux8_1.NAND4F_9.Y mux8_1.NAND4F_9.Y.n10 0.396904
R17816 mux8_1.NAND4F_9.Y.n10 mux8_1.NAND4F_9.Y.n0 0.358709
R17817 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n9 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t12 540.38
R17818 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t18 491.64
R17819 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t10 491.64
R17820 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t9 491.64
R17821 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t13 491.64
R17822 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t15 367.928
R17823 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n1 227.526
R17824 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n8 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t16 227.356
R17825 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n3 227.266
R17826 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n2 227.266
R17827 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t17 213.688
R17828 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n6 162.852
R17829 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n9 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n8 160.439
R17830 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t7 139.78
R17831 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t11 139.78
R17832 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t14 139.78
R17833 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t8 139.78
R17834 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n8 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n7 94.4341
R17835 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t0 42.7831
R17836 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n5 38.6833
R17837 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t1 30.379
R17838 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t5 30.379
R17839 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t2 30.379
R17840 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t3 30.379
R17841 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t6 30.379
R17842 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t4 30.379
R17843 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n4 28.3986
R17844 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n0 18.8832
R17845 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n10 11.2587
R17846 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n10 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT 5.09176
R17847 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n10 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT 4.19292
R17848 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n9 0.794268
R17849 a_n18422_n5154.n2 a_n18422_n5154.n0 121.353
R17850 a_n18422_n5154.n3 a_n18422_n5154.n2 121.353
R17851 a_n18422_n5154.n2 a_n18422_n5154.n1 121.001
R17852 a_n18422_n5154.n0 a_n18422_n5154.t0 30.462
R17853 a_n18422_n5154.n0 a_n18422_n5154.t1 30.462
R17854 a_n18422_n5154.n1 a_n18422_n5154.t3 30.462
R17855 a_n18422_n5154.n1 a_n18422_n5154.t5 30.462
R17856 a_n18422_n5154.n3 a_n18422_n5154.t2 30.462
R17857 a_n18422_n5154.t4 a_n18422_n5154.n3 30.462
R17858 mux8_8.NAND4F_6.Y.n1 mux8_8.NAND4F_6.Y.t10 933.563
R17859 mux8_8.NAND4F_6.Y.n1 mux8_8.NAND4F_6.Y.t11 367.635
R17860 mux8_8.NAND4F_6.Y.n2 mux8_8.NAND4F_6.Y.t9 308.481
R17861 mux8_8.NAND4F_6.Y.n0 mux8_8.NAND4F_6.Y.n4 187.373
R17862 mux8_8.NAND4F_6.Y.n0 mux8_8.NAND4F_6.Y.n5 187.192
R17863 mux8_8.NAND4F_6.Y.n0 mux8_8.NAND4F_6.Y.n6 187.192
R17864 mux8_8.NAND4F_6.Y.n8 mux8_8.NAND4F_6.Y.n7 187.192
R17865 mux8_8.NAND4F_6.Y mux8_8.NAND4F_6.Y.n2 162.047
R17866 mux8_8.NAND4F_6.Y.n3 mux8_8.NAND4F_6.Y.t2 22.7831
R17867 mux8_8.NAND4F_6.Y.n3 mux8_8.NAND4F_6.Y 22.171
R17868 mux8_8.NAND4F_6.Y.n4 mux8_8.NAND4F_6.Y.t1 20.1899
R17869 mux8_8.NAND4F_6.Y.n4 mux8_8.NAND4F_6.Y.t0 20.1899
R17870 mux8_8.NAND4F_6.Y.n5 mux8_8.NAND4F_6.Y.t6 20.1899
R17871 mux8_8.NAND4F_6.Y.n5 mux8_8.NAND4F_6.Y.t5 20.1899
R17872 mux8_8.NAND4F_6.Y.n6 mux8_8.NAND4F_6.Y.t8 20.1899
R17873 mux8_8.NAND4F_6.Y.n6 mux8_8.NAND4F_6.Y.t7 20.1899
R17874 mux8_8.NAND4F_6.Y.n7 mux8_8.NAND4F_6.Y.t3 20.1899
R17875 mux8_8.NAND4F_6.Y.n7 mux8_8.NAND4F_6.Y.t4 20.1899
R17876 mux8_8.NAND4F_6.Y.n2 mux8_8.NAND4F_6.Y.n1 10.955
R17877 mux8_8.NAND4F_6.Y mux8_8.NAND4F_6.Y.n3 0.781576
R17878 mux8_8.NAND4F_6.Y mux8_8.NAND4F_6.Y.n8 0.396904
R17879 mux8_8.NAND4F_6.Y.n8 mux8_8.NAND4F_6.Y.n0 0.358709
R17880 a_n14931_1406.n0 a_n14931_1406.t4 539.788
R17881 a_n14931_1406.n1 a_n14931_1406.t7 531.496
R17882 a_n14931_1406.n0 a_n14931_1406.t3 490.034
R17883 a_n14931_1406.n5 a_n14931_1406.t0 283.788
R17884 a_n14931_1406.t1 a_n14931_1406.n5 205.489
R17885 a_n14931_1406.n2 a_n14931_1406.t2 182.625
R17886 a_n14931_1406.n3 a_n14931_1406.t5 179.054
R17887 a_n14931_1406.n2 a_n14931_1406.t6 139.78
R17888 a_n14931_1406.n4 a_n14931_1406.n3 101.368
R17889 a_n14931_1406.n5 a_n14931_1406.n4 77.9135
R17890 a_n14931_1406.n4 a_n14931_1406.n1 76.1557
R17891 a_n14931_1406.n1 a_n14931_1406.n0 8.29297
R17892 a_n14931_1406.n3 a_n14931_1406.n2 3.57087
R17893 a_n14751_1406.n2 a_n14751_1406.n1 121.353
R17894 a_n14751_1406.n3 a_n14751_1406.n2 121.001
R17895 a_n14751_1406.n2 a_n14751_1406.n0 120.977
R17896 a_n14751_1406.n1 a_n14751_1406.t2 30.462
R17897 a_n14751_1406.n1 a_n14751_1406.t1 30.462
R17898 a_n14751_1406.n0 a_n14751_1406.t5 30.462
R17899 a_n14751_1406.n0 a_n14751_1406.t3 30.462
R17900 a_n14751_1406.n3 a_n14751_1406.t4 30.462
R17901 a_n14751_1406.t0 a_n14751_1406.n3 30.462
R17902 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t18 491.64
R17903 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t16 491.64
R17904 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t21 491.64
R17905 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t19 491.64
R17906 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t22 485.221
R17907 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t13 367.928
R17908 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t12 255.588
R17909 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t14 224.478
R17910 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t15 213.688
R17911 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n0 209.19
R17912 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t17 139.78
R17913 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t20 139.78
R17914 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t23 139.78
R17915 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n10 120.999
R17916 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n9 120.999
R17917 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n22 104.489
R17918 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n12 92.5005
R17919 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n18 86.2638
R17920 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n17 85.8873
R17921 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n15 85.724
R17922 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n7 84.5046
R17923 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n23 83.8907
R17924 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n20 75.0672
R17925 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n17 75.0672
R17926 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n19 73.1255
R17927 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n15 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n14 73.1255
R17928 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n17 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n16 73.1255
R17929 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n6 72.3005
R17930 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n15 68.8946
R17931 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n8 60.9797
R17932 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n13 41.9827
R17933 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t11 30.462
R17934 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t5 30.462
R17935 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t3 30.462
R17936 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t4 30.462
R17937 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t9 30.462
R17938 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t10 30.462
R17939 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n11 28.124
R17940 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n5 19.963
R17941 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n1 17.8661
R17942 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n2 17.8661
R17943 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n3 17.1217
R17944 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t1 11.8205
R17945 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t7 11.8205
R17946 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t8 11.8205
R17947 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t6 11.8205
R17948 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t0 11.8205
R17949 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t2 11.8205
R17950 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n21 9.3005
R17951 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n4 1.8615
R17952 mux8_4.NAND4F_4.B.n10 mux8_4.NAND4F_4.B.t6 933.563
R17953 mux8_4.NAND4F_4.B.n5 mux8_4.NAND4F_4.B.t11 933.563
R17954 mux8_4.NAND4F_4.B.n3 mux8_4.NAND4F_4.B.t4 933.563
R17955 mux8_4.NAND4F_4.B.n1 mux8_4.NAND4F_4.B.t10 933.563
R17956 mux8_4.NAND4F_4.B.n10 mux8_4.NAND4F_4.B.t13 367.635
R17957 mux8_4.NAND4F_4.B.n5 mux8_4.NAND4F_4.B.t12 367.635
R17958 mux8_4.NAND4F_4.B.n3 mux8_4.NAND4F_4.B.t5 367.635
R17959 mux8_4.NAND4F_4.B.n1 mux8_4.NAND4F_4.B.t7 367.635
R17960 mux8_4.NAND4F_4.B.n11 mux8_4.NAND4F_4.B.t15 308.481
R17961 mux8_4.NAND4F_4.B.n6 mux8_4.NAND4F_4.B.t14 308.481
R17962 mux8_4.NAND4F_4.B.n4 mux8_4.NAND4F_4.B.t8 308.481
R17963 mux8_4.NAND4F_4.B.n2 mux8_4.NAND4F_4.B.t9 308.481
R17964 mux8_4.NAND4F_4.B.n0 mux8_4.NAND4F_4.B.t1 256.514
R17965 mux8_4.NAND4F_4.B.n0 mux8_4.NAND4F_4.B.n8 226.258
R17966 mux8_4.NAND4F_4.B mux8_4.NAND4F_4.B.n2 162.173
R17967 mux8_4.NAND4F_4.B mux8_4.NAND4F_4.B.n6 162.137
R17968 mux8_4.NAND4F_4.B mux8_4.NAND4F_4.B.n11 162.117
R17969 mux8_4.NAND4F_4.B.n7 mux8_4.NAND4F_4.B.n4 161.703
R17970 mux8_4.NAND4F_4.B.n0 mux8_4.NAND4F_4.B.t0 83.7172
R17971 mux8_4.NAND4F_4.B.n8 mux8_4.NAND4F_4.B.t3 30.379
R17972 mux8_4.NAND4F_4.B.n8 mux8_4.NAND4F_4.B.t2 30.379
R17973 mux8_4.NAND4F_4.B.n12 mux8_4.NAND4F_4.B 24.8912
R17974 mux8_4.NAND4F_4.B.n7 mux8_4.NAND4F_4.B 21.6618
R17975 mux8_4.NAND4F_4.B.n11 mux8_4.NAND4F_4.B.n10 10.955
R17976 mux8_4.NAND4F_4.B.n6 mux8_4.NAND4F_4.B.n5 10.955
R17977 mux8_4.NAND4F_4.B.n4 mux8_4.NAND4F_4.B.n3 10.955
R17978 mux8_4.NAND4F_4.B.n2 mux8_4.NAND4F_4.B.n1 10.955
R17979 mux8_4.NAND4F_4.B.n12 mux8_4.NAND4F_4.B.n9 3.67985
R17980 mux8_4.NAND4F_4.B.n9 mux8_4.NAND4F_4.B.n0 1.46835
R17981 mux8_4.NAND4F_4.B mux8_4.NAND4F_4.B.n12 0.502677
R17982 mux8_4.NAND4F_4.B.n9 mux8_4.NAND4F_4.B 0.498606
R17983 mux8_4.NAND4F_4.B mux8_4.NAND4F_4.B.n7 0.470197
R17984 a_n14077_3810.n0 a_n14077_3810.n2 81.2978
R17985 a_n14077_3810.n1 a_n14077_3810.n6 81.1637
R17986 a_n14077_3810.n1 a_n14077_3810.n5 81.1637
R17987 a_n14077_3810.n0 a_n14077_3810.n4 81.1637
R17988 a_n14077_3810.n0 a_n14077_3810.n3 81.1637
R17989 a_n14077_3810.n7 a_n14077_3810.n1 80.9213
R17990 a_n14077_3810.n6 a_n14077_3810.t8 11.8205
R17991 a_n14077_3810.n6 a_n14077_3810.t1 11.8205
R17992 a_n14077_3810.n5 a_n14077_3810.t7 11.8205
R17993 a_n14077_3810.n5 a_n14077_3810.t6 11.8205
R17994 a_n14077_3810.n4 a_n14077_3810.t11 11.8205
R17995 a_n14077_3810.n4 a_n14077_3810.t9 11.8205
R17996 a_n14077_3810.n3 a_n14077_3810.t3 11.8205
R17997 a_n14077_3810.n3 a_n14077_3810.t10 11.8205
R17998 a_n14077_3810.n2 a_n14077_3810.t4 11.8205
R17999 a_n14077_3810.n2 a_n14077_3810.t5 11.8205
R18000 a_n14077_3810.n7 a_n14077_3810.t0 11.8205
R18001 a_n14077_3810.t2 a_n14077_3810.n7 11.8205
R18002 a_n14077_3810.n1 a_n14077_3810.n0 0.402735
R18003 V_FLAG_0.XOR2_2.Y.n2 V_FLAG_0.XOR2_2.Y.t13 540.38
R18004 V_FLAG_0.XOR2_2.Y.n0 V_FLAG_0.XOR2_2.Y.t15 367.928
R18005 V_FLAG_0.XOR2_2.Y.n1 V_FLAG_0.XOR2_2.Y.t14 227.356
R18006 V_FLAG_0.XOR2_2.Y.n0 V_FLAG_0.XOR2_2.Y.t12 213.688
R18007 V_FLAG_0.XOR2_2.Y.n2 V_FLAG_0.XOR2_2.Y.n1 160.439
R18008 V_FLAG_0.XOR2_2.Y.n5 V_FLAG_0.XOR2_2.Y.n4 120.999
R18009 V_FLAG_0.XOR2_2.Y.n5 V_FLAG_0.XOR2_2.Y.n3 120.999
R18010 V_FLAG_0.XOR2_2.Y.n17 V_FLAG_0.XOR2_2.Y.n16 104.489
R18011 V_FLAG_0.XOR2_2.Y.n1 V_FLAG_0.XOR2_2.Y.n0 94.4341
R18012 V_FLAG_0.XOR2_2.Y.n7 V_FLAG_0.XOR2_2.Y.n6 92.5005
R18013 V_FLAG_0.XOR2_2.Y.n14 V_FLAG_0.XOR2_2.Y.n12 86.2638
R18014 V_FLAG_0.XOR2_2.Y.n12 V_FLAG_0.XOR2_2.Y.n11 85.8873
R18015 V_FLAG_0.XOR2_2.Y.n12 V_FLAG_0.XOR2_2.Y.n9 85.724
R18016 V_FLAG_0.XOR2_2.Y V_FLAG_0.XOR2_2.Y.n17 83.9389
R18017 V_FLAG_0.XOR2_2.Y.n15 V_FLAG_0.XOR2_2.Y.n14 75.0672
R18018 V_FLAG_0.XOR2_2.Y.n15 V_FLAG_0.XOR2_2.Y.n11 75.0672
R18019 V_FLAG_0.XOR2_2.Y.n14 V_FLAG_0.XOR2_2.Y.n13 73.1255
R18020 V_FLAG_0.XOR2_2.Y.n9 V_FLAG_0.XOR2_2.Y.n8 73.1255
R18021 V_FLAG_0.XOR2_2.Y.n11 V_FLAG_0.XOR2_2.Y.n10 73.1255
R18022 V_FLAG_0.XOR2_2.Y.n16 V_FLAG_0.XOR2_2.Y.n9 68.8946
R18023 V_FLAG_0.XOR2_2.Y.n17 V_FLAG_0.XOR2_2.Y.n7 41.9827
R18024 V_FLAG_0.XOR2_2.Y.n6 V_FLAG_0.XOR2_2.Y.t0 30.462
R18025 V_FLAG_0.XOR2_2.Y.n6 V_FLAG_0.XOR2_2.Y.t11 30.462
R18026 V_FLAG_0.XOR2_2.Y.n4 V_FLAG_0.XOR2_2.Y.t7 30.462
R18027 V_FLAG_0.XOR2_2.Y.n4 V_FLAG_0.XOR2_2.Y.t10 30.462
R18028 V_FLAG_0.XOR2_2.Y.n3 V_FLAG_0.XOR2_2.Y.t2 30.462
R18029 V_FLAG_0.XOR2_2.Y.n3 V_FLAG_0.XOR2_2.Y.t1 30.462
R18030 V_FLAG_0.XOR2_2.Y.n7 V_FLAG_0.XOR2_2.Y.n5 28.124
R18031 V_FLAG_0.XOR2_2.Y.n8 V_FLAG_0.XOR2_2.Y.t4 11.8205
R18032 V_FLAG_0.XOR2_2.Y.n8 V_FLAG_0.XOR2_2.Y.t8 11.8205
R18033 V_FLAG_0.XOR2_2.Y.n13 V_FLAG_0.XOR2_2.Y.t9 11.8205
R18034 V_FLAG_0.XOR2_2.Y.n13 V_FLAG_0.XOR2_2.Y.t6 11.8205
R18035 V_FLAG_0.XOR2_2.Y.n10 V_FLAG_0.XOR2_2.Y.t5 11.8205
R18036 V_FLAG_0.XOR2_2.Y.n10 V_FLAG_0.XOR2_2.Y.t3 11.8205
R18037 V_FLAG_0.XOR2_2.Y.n16 V_FLAG_0.XOR2_2.Y.n15 9.3005
R18038 V_FLAG_0.XOR2_2.Y V_FLAG_0.XOR2_2.Y.n2 0.838386
R18039 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t21 491.64
R18040 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t22 491.64
R18041 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t20 491.64
R18042 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t17 491.64
R18043 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t13 485.221
R18044 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t16 367.928
R18045 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t15 255.588
R18046 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t23 224.478
R18047 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t12 213.688
R18048 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n0 209.19
R18049 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t18 139.78
R18050 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t19 139.78
R18051 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t14 139.78
R18052 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n11 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n10 120.999
R18053 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n11 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n9 120.999
R18054 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n23 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n22 104.489
R18055 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n13 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n12 92.5005
R18056 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n20 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n18 86.2638
R18057 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n18 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n17 85.8873
R18058 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n18 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n15 85.724
R18059 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n7 84.5046
R18060 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n23 83.8907
R18061 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n21 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n20 75.0672
R18062 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n21 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n17 75.0672
R18063 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n20 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n19 73.1255
R18064 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n17 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n16 73.1255
R18065 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n15 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n14 73.1255
R18066 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n6 72.3005
R18067 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n22 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n15 68.8946
R18068 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n8 60.9797
R18069 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n23 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n13 41.9827
R18070 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n12 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t0 30.462
R18071 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n12 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t6 30.462
R18072 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t3 30.462
R18073 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t2 30.462
R18074 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t8 30.462
R18075 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t7 30.462
R18076 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n13 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n11 28.124
R18077 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n5 19.963
R18078 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n1 17.8661
R18079 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n2 17.8661
R18080 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n3 17.1217
R18081 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n16 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t11 11.8205
R18082 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n16 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t10 11.8205
R18083 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n19 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t5 11.8205
R18084 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n19 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t4 11.8205
R18085 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n14 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t9 11.8205
R18086 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n14 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t1 11.8205
R18087 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n22 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n21 9.3005
R18088 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n4 1.8615
R18089 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t7 485.221
R18090 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t8 367.928
R18091 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n5 227.526
R18092 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n6 227.266
R18093 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n4 227.266
R18094 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t9 224.478
R18095 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t10 213.688
R18096 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n2 84.5046
R18097 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n1 72.3005
R18098 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n3 61.0566
R18099 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t3 42.7747
R18100 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t6 30.379
R18101 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t1 30.379
R18102 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t4 30.379
R18103 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t5 30.379
R18104 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t2 30.379
R18105 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.t0 30.379
R18106 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A.n0 0.583137
R18107 a_n3350_1380.n2 a_n3350_1380.t6 541.395
R18108 a_n3350_1380.n3 a_n3350_1380.t4 527.402
R18109 a_n3350_1380.n2 a_n3350_1380.t7 491.64
R18110 a_n3350_1380.n5 a_n3350_1380.t0 281.906
R18111 a_n3350_1380.t1 a_n3350_1380.n5 204.359
R18112 a_n3350_1380.n0 a_n3350_1380.t3 180.73
R18113 a_n3350_1380.n1 a_n3350_1380.t5 179.45
R18114 a_n3350_1380.n0 a_n3350_1380.t2 139.78
R18115 a_n3350_1380.n4 a_n3350_1380.n1 105.635
R18116 a_n3350_1380.n4 a_n3350_1380.n3 76.0005
R18117 a_n3350_1380.n5 a_n3350_1380.n4 67.9685
R18118 a_n3350_1380.n3 a_n3350_1380.n2 13.994
R18119 a_n3350_1380.n1 a_n3350_1380.n0 1.28015
R18120 a_n3320_1406.n3 a_n3320_1406.n2 121.353
R18121 a_n3320_1406.n2 a_n3320_1406.n1 121.001
R18122 a_n3320_1406.n2 a_n3320_1406.n0 120.977
R18123 a_n3320_1406.n1 a_n3320_1406.t4 30.462
R18124 a_n3320_1406.n1 a_n3320_1406.t1 30.462
R18125 a_n3320_1406.n0 a_n3320_1406.t5 30.462
R18126 a_n3320_1406.n0 a_n3320_1406.t3 30.462
R18127 a_n3320_1406.t2 a_n3320_1406.n3 30.462
R18128 a_n3320_1406.n3 a_n3320_1406.t0 30.462
R18129 a_n1768_1406.n0 a_n1768_1406.t5 539.788
R18130 a_n1768_1406.n1 a_n1768_1406.t6 531.496
R18131 a_n1768_1406.n0 a_n1768_1406.t3 490.034
R18132 a_n1768_1406.n5 a_n1768_1406.t1 283.788
R18133 a_n1768_1406.t0 a_n1768_1406.n5 205.489
R18134 a_n1768_1406.n2 a_n1768_1406.t2 182.625
R18135 a_n1768_1406.n3 a_n1768_1406.t4 179.054
R18136 a_n1768_1406.n2 a_n1768_1406.t7 139.78
R18137 a_n1768_1406.n4 a_n1768_1406.n3 101.368
R18138 a_n1768_1406.n5 a_n1768_1406.n4 77.9135
R18139 a_n1768_1406.n4 a_n1768_1406.n1 76.1557
R18140 a_n1768_1406.n1 a_n1768_1406.n0 8.29297
R18141 a_n1768_1406.n3 a_n1768_1406.n2 3.57087
R18142 a_n1588_1406.n2 a_n1588_1406.n0 121.353
R18143 a_n1588_1406.n2 a_n1588_1406.n1 121.001
R18144 a_n1588_1406.n3 a_n1588_1406.n2 120.977
R18145 a_n1588_1406.n0 a_n1588_1406.t5 30.462
R18146 a_n1588_1406.n0 a_n1588_1406.t4 30.462
R18147 a_n1588_1406.n1 a_n1588_1406.t1 30.462
R18148 a_n1588_1406.n1 a_n1588_1406.t3 30.462
R18149 a_n1588_1406.n3 a_n1588_1406.t2 30.462
R18150 a_n1588_1406.t0 a_n1588_1406.n3 30.462
R18151 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t21 491.64
R18152 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t19 491.64
R18153 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t23 491.64
R18154 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t22 491.64
R18155 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t16 485.221
R18156 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t13 367.928
R18157 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t18 255.588
R18158 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t14 224.478
R18159 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t12 213.688
R18160 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n0 209.19
R18161 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t20 139.78
R18162 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t17 139.78
R18163 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t15 139.78
R18164 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n10 120.999
R18165 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n9 120.999
R18166 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n22 104.489
R18167 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n12 92.5005
R18168 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n18 86.2638
R18169 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n17 85.8873
R18170 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n15 85.724
R18171 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n7 84.5046
R18172 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n23 83.8907
R18173 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n17 75.0672
R18174 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n20 75.0672
R18175 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n15 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n14 73.1255
R18176 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n17 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n16 73.1255
R18177 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n19 73.1255
R18178 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n6 72.3005
R18179 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n15 68.8946
R18180 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n8 60.9797
R18181 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n13 41.9827
R18182 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t9 30.462
R18183 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t5 30.462
R18184 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t3 30.462
R18185 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t4 30.462
R18186 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t11 30.462
R18187 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t10 30.462
R18188 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n11 28.124
R18189 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n5 19.963
R18190 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n1 17.8661
R18191 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n2 17.8661
R18192 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n3 17.1217
R18193 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t7 11.8205
R18194 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t6 11.8205
R18195 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t8 11.8205
R18196 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t2 11.8205
R18197 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t0 11.8205
R18198 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t1 11.8205
R18199 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n21 9.3005
R18200 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n4 1.8615
R18201 OR8_0.NOT8_0.A5.n3 OR8_0.NOT8_0.A5.t10 394.37
R18202 OR8_0.NOT8_0.A5.n2 OR8_0.NOT8_0.A5.t9 291.829
R18203 OR8_0.NOT8_0.A5.n2 OR8_0.NOT8_0.A5.t7 291.829
R18204 OR8_0.NOT8_0.A5.n0 OR8_0.NOT8_0.A5.t4 256.425
R18205 OR8_0.NOT8_0.A5.n0 OR8_0.NOT8_0.A5.n4 231.24
R18206 OR8_0.NOT8_0.A5.n0 OR8_0.NOT8_0.A5.n5 231.03
R18207 OR8_0.NOT8_0.A5.n2 OR8_0.NOT8_0.A5.t8 221.72
R18208 OR8_0.NOT8_0.A5.n0 OR8_0.NOT8_0.A5.n1 66.4681
R18209 OR8_0.NOT8_0.A5.n3 OR8_0.NOT8_0.A5.n2 53.374
R18210 OR8_0.NOT8_0.A5.n0 OR8_0.NOT8_0.A5 26.86
R18211 OR8_0.NOT8_0.A5.n5 OR8_0.NOT8_0.A5.t3 25.395
R18212 OR8_0.NOT8_0.A5.n5 OR8_0.NOT8_0.A5.t2 25.395
R18213 OR8_0.NOT8_0.A5.n4 OR8_0.NOT8_0.A5.t1 25.395
R18214 OR8_0.NOT8_0.A5.n4 OR8_0.NOT8_0.A5.t5 25.395
R18215 OR8_0.NOT8_0.A5.n1 OR8_0.NOT8_0.A5.t6 19.8005
R18216 OR8_0.NOT8_0.A5.n1 OR8_0.NOT8_0.A5.t0 19.8005
R18217 OR8_0.NOT8_0.A5 OR8_0.NOT8_0.A5.n3 1.27207
R18218 OR8_0.S5.n1 OR8_0.S5.t4 1032.02
R18219 OR8_0.S5.n1 OR8_0.S5.t5 336.962
R18220 OR8_0.S5.n1 OR8_0.S5.t6 326.154
R18221 OR8_0.S5.n0 OR8_0.S5.t1 256.514
R18222 OR8_0.S5.n0 OR8_0.S5.n2 226.258
R18223 mux8_7.NAND4F_2.A OR8_0.S5.n1 162.952
R18224 OR8_0.S5.n0 OR8_0.S5.t0 83.7172
R18225 OR8_0.NOT8_0.S5 mux8_7.A3 74.6063
R18226 OR8_0.S5.n2 OR8_0.S5.t2 30.379
R18227 OR8_0.S5.n2 OR8_0.S5.t3 30.379
R18228 mux8_7.A3 mux8_7.NAND4F_2.A 14.0763
R18229 OR8_0.NOT8_0.S5 OR8_0.S5.n0 1.9182
R18230 B0.n13 B0.t1 491.64
R18231 B0.n12 B0.t25 491.64
R18232 B0.n11 B0.t18 491.64
R18233 B0.n10 B0.t47 491.64
R18234 B0.n47 B0.t11 491.64
R18235 B0.n46 B0.t13 491.64
R18236 B0.n45 B0.t9 491.64
R18237 B0.n44 B0.t50 491.64
R18238 B0.n33 B0.t53 485.443
R18239 B0.n28 B0.t2 485.221
R18240 B0.n17 B0.t41 485.221
R18241 B0.n20 B0.t19 485.221
R18242 B0.n24 B0.t46 485.221
R18243 B0.n6 B0.t7 394.37
R18244 B0.n3 B0.t28 394.37
R18245 B0.n1 B0.t14 394.37
R18246 B0.n36 B0.t3 379.173
R18247 B0.n26 B0.t10 367.928
R18248 B0.n15 B0.t17 367.928
R18249 B0.n18 B0.t48 367.928
R18250 B0.n22 B0.t20 367.928
R18251 B0.n31 B0.t21 343.827
R18252 B0.n37 B0.t45 312.599
R18253 B0.n5 B0.t23 291.829
R18254 B0.n5 B0.t49 291.829
R18255 B0.n2 B0.t44 291.829
R18256 B0.n2 B0.t43 291.829
R18257 B0.n0 B0.t31 291.829
R18258 B0.n0 B0.t30 291.829
R18259 B0.n14 B0.t52 255.588
R18260 B0.n48 B0.t35 255.588
R18261 B0.n37 B0.t29 247.428
R18262 B0.n38 B0.t26 247.428
R18263 B0.n39 B0.t6 247.428
R18264 B0.n36 B0.t5 247.428
R18265 B0.n31 B0.t36 237.787
R18266 B0.n32 B0.t40 224.478
R18267 B0.n27 B0.t34 224.478
R18268 B0.n16 B0.t37 224.478
R18269 B0.n19 B0.t16 224.478
R18270 B0.n23 B0.t42 224.478
R18271 B0.n5 B0.t27 221.72
R18272 B0.n2 B0.t39 221.72
R18273 B0.n0 B0.t51 221.72
R18274 B0.n26 B0.t33 213.688
R18275 B0.n15 B0.t22 213.688
R18276 B0.n18 B0.t0 213.688
R18277 B0.n22 B0.t24 213.688
R18278 B0.n44 B0.n43 209.407
R18279 B0.n10 B0.n9 209.19
R18280 B0 B0.n40 162.139
R18281 B0.n9 B0.t15 139.78
R18282 B0.n9 B0.t38 139.78
R18283 B0.n9 B0.t4 139.78
R18284 B0.n43 B0.t12 139.78
R18285 B0.n43 B0.t32 139.78
R18286 B0.n43 B0.t8 139.78
R18287 B0.n28 B0.n27 84.5046
R18288 B0.n17 B0.n16 84.5046
R18289 B0.n20 B0.n19 84.5046
R18290 B0.n24 B0.n23 84.5046
R18291 B0.n33 B0.n32 83.8438
R18292 B0.n27 B0.n26 72.3005
R18293 B0.n16 B0.n15 72.3005
R18294 B0.n19 B0.n18 72.3005
R18295 B0.n23 B0.n22 72.3005
R18296 B0.n39 B0.n38 65.1723
R18297 B0.n38 B0.n37 65.1723
R18298 B0 B0.n24 61.0561
R18299 B0 B0.n17 61.0552
R18300 B0 B0.n20 61.0542
R18301 B0 B0.n28 61.0523
R18302 B0 B0.n33 61.0461
R18303 B0.n6 B0.n5 53.374
R18304 B0.n3 B0.n2 53.374
R18305 B0.n1 B0.n0 53.374
R18306 B0.n32 B0.n31 48.2005
R18307 B0.n30 B0 34.2079
R18308 B0.n40 B0.n39 33.2653
R18309 B0.n40 B0.n36 31.9075
R18310 B0 B0.n48 27.4136
R18311 B0.n12 B0.n11 17.8661
R18312 B0.n11 B0.n10 17.8661
R18313 B0.n45 B0.n44 17.8661
R18314 B0.n46 B0.n45 17.8661
R18315 B0.n13 B0.n12 17.1217
R18316 B0.n47 B0.n46 17.1217
R18317 B0.n8 B0.n4 14.1861
R18318 B0 B0.n50 12.6959
R18319 B0.n49 B0 12.5435
R18320 B0.n35 B0.n34 12.4105
R18321 B0.n42 B0.n41 12.4105
R18322 B0.n8 B0.n7 12.4105
R18323 B0 B0.n14 11.1665
R18324 B0 B0.n30 8.80378
R18325 B0.n21 B0 6.65761
R18326 B0.n42 B0.n35 4.53404
R18327 B0.n30 B0.n29 4.38057
R18328 B0.n21 B0 3.67532
R18329 B0.n49 B0.n42 3.41551
R18330 B0.n50 B0.n8 3.08789
R18331 B0.n50 B0.n49 2.61846
R18332 B0.n25 B0 2.58066
R18333 B0.n29 B0 2.46116
R18334 B0.n14 B0.n13 1.8615
R18335 B0.n48 B0.n47 1.8615
R18336 B0 B0.n25 1.81292
R18337 B0.n25 B0.n21 1.54977
R18338 B0 B0.n1 1.27074
R18339 B0.n34 B0 1.20397
R18340 B0.n41 B0 1.14949
R18341 B0.n7 B0.n6 0.761001
R18342 B0.n4 B0.n3 0.757989
R18343 B0.n29 B0 0.188437
R18344 B0.n34 B0 0.0682083
R18345 B0.n4 B0 0.060741
R18346 B0.n7 B0 0.0577289
R18347 B0.n41 B0 0.0255
R18348 B0.n35 B0 0.0165488
R18349 MULT_0.NAND2_2.Y.n5 MULT_0.NAND2_2.Y.t8 291.829
R18350 MULT_0.NAND2_2.Y.n5 MULT_0.NAND2_2.Y.t10 291.829
R18351 MULT_0.NAND2_2.Y.n0 MULT_0.NAND2_2.Y.n3 227.526
R18352 MULT_0.NAND2_2.Y.n0 MULT_0.NAND2_2.Y.n4 227.266
R18353 MULT_0.NAND2_2.Y.n0 MULT_0.NAND2_2.Y.n2 227.266
R18354 MULT_0.NAND2_2.Y.n5 MULT_0.NAND2_2.Y.t9 221.72
R18355 MULT_0.NAND2_2.Y.t7 MULT_0.NAND2_2.Y.n1 393.897
R18356 MULT_0.NAND2_2.Y.n0 MULT_0.NAND2_2.Y.t3 42.7333
R18357 MULT_0.NAND2_2.Y.n4 MULT_0.NAND2_2.Y.t4 30.379
R18358 MULT_0.NAND2_2.Y.n4 MULT_0.NAND2_2.Y.t0 30.379
R18359 MULT_0.NAND2_2.Y.n2 MULT_0.NAND2_2.Y.t6 30.379
R18360 MULT_0.NAND2_2.Y.n2 MULT_0.NAND2_2.Y.t5 30.379
R18361 MULT_0.NAND2_2.Y.n3 MULT_0.NAND2_2.Y.t2 30.379
R18362 MULT_0.NAND2_2.Y.n3 MULT_0.NAND2_2.Y.t1 30.379
R18363 MULT_0.NAND2_2.Y.n5 MULT_0.NAND2_2.Y.n1 53.4911
R18364 MULT_0.NAND2_2.Y.n0 MULT_0.NAND2_2.Y.n1 0.620447
R18365 a_n12345_n28506.n2 a_n12345_n28506.t7 541.395
R18366 a_n12345_n28506.n3 a_n12345_n28506.t4 527.402
R18367 a_n12345_n28506.n2 a_n12345_n28506.t5 491.64
R18368 a_n12345_n28506.n5 a_n12345_n28506.t0 281.906
R18369 a_n12345_n28506.t1 a_n12345_n28506.n5 204.359
R18370 a_n12345_n28506.n0 a_n12345_n28506.t3 180.73
R18371 a_n12345_n28506.n1 a_n12345_n28506.t2 179.45
R18372 a_n12345_n28506.n0 a_n12345_n28506.t6 139.78
R18373 a_n12345_n28506.n4 a_n12345_n28506.n1 105.635
R18374 a_n12345_n28506.n4 a_n12345_n28506.n3 76.0005
R18375 a_n12345_n28506.n5 a_n12345_n28506.n4 67.9685
R18376 a_n12345_n28506.n3 a_n12345_n28506.n2 13.994
R18377 a_n12345_n28506.n1 a_n12345_n28506.n0 1.28015
R18378 a_n11274_n29052.n3 a_n11274_n29052.n2 121.353
R18379 a_n11274_n29052.n2 a_n11274_n29052.n1 121.001
R18380 a_n11274_n29052.n2 a_n11274_n29052.n0 120.977
R18381 a_n11274_n29052.n0 a_n11274_n29052.t5 30.462
R18382 a_n11274_n29052.n0 a_n11274_n29052.t0 30.462
R18383 a_n11274_n29052.n1 a_n11274_n29052.t1 30.462
R18384 a_n11274_n29052.n1 a_n11274_n29052.t3 30.462
R18385 a_n11274_n29052.n3 a_n11274_n29052.t2 30.462
R18386 a_n11274_n29052.t4 a_n11274_n29052.n3 30.462
R18387 a_9336_n20950.t0 a_9336_n20950.t1 9.9005
R18388 a_9432_n20950.t0 a_9432_n20950.t1 9.9005
R18389 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t23 491.64
R18390 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t14 491.64
R18391 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t15 491.64
R18392 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t22 491.64
R18393 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n8 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t13 485.221
R18394 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t19 367.928
R18395 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t17 255.588
R18396 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n7 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t12 224.478
R18397 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t21 213.688
R18398 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n0 209.19
R18399 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t18 139.78
R18400 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t16 139.78
R18401 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t20 139.78
R18402 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n11 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n10 120.999
R18403 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n11 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n9 120.999
R18404 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n23 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n22 104.489
R18405 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n13 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n12 92.5005
R18406 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n20 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n18 86.2638
R18407 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n18 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n17 85.8873
R18408 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n18 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n15 85.724
R18409 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n8 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n7 84.5046
R18410 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n23 83.8907
R18411 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n21 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n20 75.0672
R18412 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n21 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n17 75.0672
R18413 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n20 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n19 73.1255
R18414 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n17 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n16 73.1255
R18415 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n15 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n14 73.1255
R18416 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n7 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n6 72.3005
R18417 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n22 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n15 68.8946
R18418 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n8 60.9797
R18419 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n23 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n13 41.9827
R18420 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n12 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t2 30.462
R18421 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n12 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t8 30.462
R18422 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n10 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t3 30.462
R18423 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n10 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t4 30.462
R18424 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n9 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t0 30.462
R18425 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n9 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t1 30.462
R18426 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n13 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n11 28.124
R18427 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n5 19.963
R18428 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n1 17.8661
R18429 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n2 17.8661
R18430 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n3 17.1217
R18431 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n16 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t10 11.8205
R18432 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n16 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t11 11.8205
R18433 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n19 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t6 11.8205
R18434 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n19 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t7 11.8205
R18435 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n14 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t9 11.8205
R18436 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n14 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t5 11.8205
R18437 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n22 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n21 9.3005
R18438 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n4 1.8615
R18439 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t8 485.221
R18440 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t9 367.928
R18441 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n5 227.526
R18442 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n6 227.266
R18443 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n4 227.266
R18444 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t7 224.478
R18445 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t10 213.688
R18446 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n2 84.5046
R18447 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n1 72.3005
R18448 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n3 61.0566
R18449 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t6 42.7747
R18450 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t4 30.379
R18451 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t1 30.379
R18452 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t5 30.379
R18453 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t3 30.379
R18454 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t0 30.379
R18455 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.t2 30.379
R18456 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A.n0 0.583137
R18457 MULT_0.4bit_ADDER_2.B2.n4 MULT_0.4bit_ADDER_2.B2.t22 491.64
R18458 MULT_0.4bit_ADDER_2.B2.n5 MULT_0.4bit_ADDER_2.B2.t19 491.64
R18459 MULT_0.4bit_ADDER_2.B2.n6 MULT_0.4bit_ADDER_2.B2.t17 491.64
R18460 MULT_0.4bit_ADDER_2.B2.n7 MULT_0.4bit_ADDER_2.B2.t12 491.64
R18461 MULT_0.4bit_ADDER_2.B2.n2 MULT_0.4bit_ADDER_2.B2.t16 485.221
R18462 MULT_0.4bit_ADDER_2.B2.n0 MULT_0.4bit_ADDER_2.B2.t15 367.928
R18463 MULT_0.4bit_ADDER_2.B2.n8 MULT_0.4bit_ADDER_2.B2.t21 255.588
R18464 MULT_0.4bit_ADDER_2.B2.n1 MULT_0.4bit_ADDER_2.B2.t14 224.478
R18465 MULT_0.4bit_ADDER_2.B2.n0 MULT_0.4bit_ADDER_2.B2.t18 213.688
R18466 MULT_0.4bit_ADDER_2.B2.n4 MULT_0.4bit_ADDER_2.B2.n3 209.19
R18467 MULT_0.4bit_ADDER_2.B2.n3 MULT_0.4bit_ADDER_2.B2.t23 139.78
R18468 MULT_0.4bit_ADDER_2.B2.n3 MULT_0.4bit_ADDER_2.B2.t13 139.78
R18469 MULT_0.4bit_ADDER_2.B2.n3 MULT_0.4bit_ADDER_2.B2.t20 139.78
R18470 MULT_0.4bit_ADDER_2.B2.n12 MULT_0.4bit_ADDER_2.B2.n11 120.999
R18471 MULT_0.4bit_ADDER_2.B2.n12 MULT_0.4bit_ADDER_2.B2.n10 120.999
R18472 MULT_0.4bit_ADDER_2.B2.n24 MULT_0.4bit_ADDER_2.B2.n23 104.489
R18473 MULT_0.4bit_ADDER_2.B2.n9 MULT_0.4bit_ADDER_2.B2 103.258
R18474 MULT_0.4bit_ADDER_2.B2.n14 MULT_0.4bit_ADDER_2.B2.n13 92.5005
R18475 MULT_0.4bit_ADDER_2.B2.n21 MULT_0.4bit_ADDER_2.B2.n19 86.2638
R18476 MULT_0.4bit_ADDER_2.B2.n19 MULT_0.4bit_ADDER_2.B2.n18 85.8873
R18477 MULT_0.4bit_ADDER_2.B2.n19 MULT_0.4bit_ADDER_2.B2.n16 85.724
R18478 MULT_0.4bit_ADDER_2.B2.n2 MULT_0.4bit_ADDER_2.B2.n1 84.5046
R18479 MULT_0.4bit_ADDER_2.B2 MULT_0.4bit_ADDER_2.B2.n24 83.8907
R18480 MULT_0.4bit_ADDER_2.B2.n22 MULT_0.4bit_ADDER_2.B2.n21 75.0672
R18481 MULT_0.4bit_ADDER_2.B2.n22 MULT_0.4bit_ADDER_2.B2.n18 75.0672
R18482 MULT_0.4bit_ADDER_2.B2.n21 MULT_0.4bit_ADDER_2.B2.n20 73.1255
R18483 MULT_0.4bit_ADDER_2.B2.n18 MULT_0.4bit_ADDER_2.B2.n17 73.1255
R18484 MULT_0.4bit_ADDER_2.B2.n16 MULT_0.4bit_ADDER_2.B2.n15 73.1255
R18485 MULT_0.4bit_ADDER_2.B2.n1 MULT_0.4bit_ADDER_2.B2.n0 72.3005
R18486 MULT_0.4bit_ADDER_2.B2.n23 MULT_0.4bit_ADDER_2.B2.n16 68.8946
R18487 MULT_0.4bit_ADDER_2.B2 MULT_0.4bit_ADDER_2.B2.n2 60.9816
R18488 MULT_0.4bit_ADDER_2.B2.n24 MULT_0.4bit_ADDER_2.B2.n14 41.9827
R18489 MULT_0.4bit_ADDER_2.B2.n13 MULT_0.4bit_ADDER_2.B2.t6 30.462
R18490 MULT_0.4bit_ADDER_2.B2.n13 MULT_0.4bit_ADDER_2.B2.t5 30.462
R18491 MULT_0.4bit_ADDER_2.B2.n11 MULT_0.4bit_ADDER_2.B2.t0 30.462
R18492 MULT_0.4bit_ADDER_2.B2.n11 MULT_0.4bit_ADDER_2.B2.t2 30.462
R18493 MULT_0.4bit_ADDER_2.B2.n10 MULT_0.4bit_ADDER_2.B2.t8 30.462
R18494 MULT_0.4bit_ADDER_2.B2.n10 MULT_0.4bit_ADDER_2.B2.t7 30.462
R18495 MULT_0.4bit_ADDER_2.B2.n14 MULT_0.4bit_ADDER_2.B2.n12 28.124
R18496 MULT_0.4bit_ADDER_2.B2.n5 MULT_0.4bit_ADDER_2.B2.n4 17.8661
R18497 MULT_0.4bit_ADDER_2.B2.n6 MULT_0.4bit_ADDER_2.B2.n5 17.8661
R18498 MULT_0.4bit_ADDER_2.B2.n7 MULT_0.4bit_ADDER_2.B2.n6 17.1217
R18499 MULT_0.4bit_ADDER_2.B2 MULT_0.4bit_ADDER_2.B2.n8 15.6329
R18500 MULT_0.4bit_ADDER_2.B2.n17 MULT_0.4bit_ADDER_2.B2.t10 11.8205
R18501 MULT_0.4bit_ADDER_2.B2.n17 MULT_0.4bit_ADDER_2.B2.t11 11.8205
R18502 MULT_0.4bit_ADDER_2.B2.n20 MULT_0.4bit_ADDER_2.B2.t3 11.8205
R18503 MULT_0.4bit_ADDER_2.B2.n20 MULT_0.4bit_ADDER_2.B2.t4 11.8205
R18504 MULT_0.4bit_ADDER_2.B2.n15 MULT_0.4bit_ADDER_2.B2.t9 11.8205
R18505 MULT_0.4bit_ADDER_2.B2.n15 MULT_0.4bit_ADDER_2.B2.t1 11.8205
R18506 MULT_0.4bit_ADDER_2.B2.n9 MULT_0.4bit_ADDER_2.B2 10.8165
R18507 MULT_0.4bit_ADDER_2.B2.n23 MULT_0.4bit_ADDER_2.B2.n22 9.3005
R18508 MULT_0.4bit_ADDER_2.B2.n8 MULT_0.4bit_ADDER_2.B2.n7 1.8615
R18509 MULT_0.4bit_ADDER_2.B2 MULT_0.4bit_ADDER_2.B2.n9 0.836623
R18510 a_n17446_n11683.n0 a_n17446_n11683.t7 539.788
R18511 a_n17446_n11683.n1 a_n17446_n11683.t6 531.496
R18512 a_n17446_n11683.n0 a_n17446_n11683.t5 490.034
R18513 a_n17446_n11683.n5 a_n17446_n11683.t0 283.788
R18514 a_n17446_n11683.t1 a_n17446_n11683.n5 205.489
R18515 a_n17446_n11683.n2 a_n17446_n11683.t4 182.625
R18516 a_n17446_n11683.n3 a_n17446_n11683.t3 179.054
R18517 a_n17446_n11683.n2 a_n17446_n11683.t2 139.78
R18518 a_n17446_n11683.n4 a_n17446_n11683.n3 101.368
R18519 a_n17446_n11683.n5 a_n17446_n11683.n4 77.9135
R18520 a_n17446_n11683.n4 a_n17446_n11683.n1 76.1557
R18521 a_n17446_n11683.n1 a_n17446_n11683.n0 8.29297
R18522 a_n17446_n11683.n3 a_n17446_n11683.n2 3.57087
R18523 mux8_3.NAND4F_4.Y.n6 mux8_3.NAND4F_4.Y.t10 1032.02
R18524 mux8_3.NAND4F_4.Y.n6 mux8_3.NAND4F_4.Y.t11 336.962
R18525 mux8_3.NAND4F_4.Y.n6 mux8_3.NAND4F_4.Y.t9 326.154
R18526 mux8_3.NAND4F_4.Y.n0 mux8_3.NAND4F_4.Y.n1 187.373
R18527 mux8_3.NAND4F_4.Y.n0 mux8_3.NAND4F_4.Y.n2 187.192
R18528 mux8_3.NAND4F_4.Y.n0 mux8_3.NAND4F_4.Y.n3 187.192
R18529 mux8_3.NAND4F_4.Y.n5 mux8_3.NAND4F_4.Y.n4 187.192
R18530 mux8_3.NAND4F_4.Y mux8_3.NAND4F_4.Y.n6 162.942
R18531 mux8_3.NAND4F_4.Y.n7 mux8_3.NAND4F_4.Y 24.5377
R18532 mux8_3.NAND4F_4.Y.n7 mux8_3.NAND4F_4.Y.t2 22.6141
R18533 mux8_3.NAND4F_4.Y.n1 mux8_3.NAND4F_4.Y.t7 20.1899
R18534 mux8_3.NAND4F_4.Y.n1 mux8_3.NAND4F_4.Y.t8 20.1899
R18535 mux8_3.NAND4F_4.Y.n2 mux8_3.NAND4F_4.Y.t3 20.1899
R18536 mux8_3.NAND4F_4.Y.n2 mux8_3.NAND4F_4.Y.t4 20.1899
R18537 mux8_3.NAND4F_4.Y.n3 mux8_3.NAND4F_4.Y.t5 20.1899
R18538 mux8_3.NAND4F_4.Y.n3 mux8_3.NAND4F_4.Y.t6 20.1899
R18539 mux8_3.NAND4F_4.Y.n4 mux8_3.NAND4F_4.Y.t0 20.1899
R18540 mux8_3.NAND4F_4.Y.n4 mux8_3.NAND4F_4.Y.t1 20.1899
R18541 mux8_3.NAND4F_4.Y mux8_3.NAND4F_4.Y.n7 0.894894
R18542 mux8_3.NAND4F_4.Y mux8_3.NAND4F_4.Y.n5 0.452586
R18543 mux8_3.NAND4F_4.Y.n5 mux8_3.NAND4F_4.Y.n0 0.358709
R18544 left_shifter_0.buffer_2.inv_1.A.n0 left_shifter_0.buffer_2.inv_1.A.t4 393.921
R18545 left_shifter_0.buffer_2.inv_1.A.n2 left_shifter_0.buffer_2.inv_1.A.t5 291.829
R18546 left_shifter_0.buffer_2.inv_1.A.n2 left_shifter_0.buffer_2.inv_1.A.t7 291.829
R18547 left_shifter_0.buffer_2.inv_1.A.n0 left_shifter_0.buffer_2.inv_1.A.t2 256.89
R18548 left_shifter_0.buffer_2.inv_1.A.n0 left_shifter_0.buffer_2.inv_1.A.n1 226.538
R18549 left_shifter_0.buffer_2.inv_1.A.n2 left_shifter_0.buffer_2.inv_1.A.t6 221.72
R18550 left_shifter_0.buffer_2.inv_1.A.n0 left_shifter_0.buffer_2.inv_1.A.t0 83.795
R18551 left_shifter_0.buffer_2.inv_1.A.n0 left_shifter_0.buffer_2.inv_1.A.n2 53.7938
R18552 left_shifter_0.buffer_2.inv_1.A.n1 left_shifter_0.buffer_2.inv_1.A.t3 30.379
R18553 left_shifter_0.buffer_2.inv_1.A.n1 left_shifter_0.buffer_2.inv_1.A.t1 30.379
R18554 left_shifter_0.S7.n1 left_shifter_0.S7.t4 1032.02
R18555 left_shifter_0.S7.n1 left_shifter_0.S7.t5 336.962
R18556 left_shifter_0.S7.n1 left_shifter_0.S7.t6 326.154
R18557 left_shifter_0.S7.n0 left_shifter_0.S7.t1 256.89
R18558 left_shifter_0.S7.n0 left_shifter_0.S7.n2 226.635
R18559 left_shifter_0.S7 left_shifter_0.S7.n1 162.952
R18560 left_shifter_0.S7.n0 left_shifter_0.S7.t0 83.7172
R18561 left_shifter_0.S7.n2 left_shifter_0.S7.t2 30.379
R18562 left_shifter_0.S7.n2 left_shifter_0.S7.t3 30.379
R18563 left_shifter_0.S7 left_shifter_0.S7.n0 0.755834
R18564 a_11865_n7203.n0 a_11865_n7203.n2 231.24
R18565 a_11865_n7203.n6 a_11865_n7203.n1 231.24
R18566 a_11865_n7203.n1 a_11865_n7203.n5 231.03
R18567 a_11865_n7203.n1 a_11865_n7203.n4 231.03
R18568 a_11865_n7203.n0 a_11865_n7203.n3 231.03
R18569 a_11865_n7203.n5 a_11865_n7203.t1 25.395
R18570 a_11865_n7203.n5 a_11865_n7203.t2 25.395
R18571 a_11865_n7203.n4 a_11865_n7203.t9 25.395
R18572 a_11865_n7203.n4 a_11865_n7203.t0 25.395
R18573 a_11865_n7203.n3 a_11865_n7203.t6 25.395
R18574 a_11865_n7203.n3 a_11865_n7203.t5 25.395
R18575 a_11865_n7203.n2 a_11865_n7203.t8 25.395
R18576 a_11865_n7203.n2 a_11865_n7203.t7 25.395
R18577 a_11865_n7203.n6 a_11865_n7203.t3 25.395
R18578 a_11865_n7203.t4 a_11865_n7203.n6 25.395
R18579 a_11865_n7203.n1 a_11865_n7203.n0 0.421553
R18580 a_3463_4888.n2 a_3463_4888.t4 541.395
R18581 a_3463_4888.n3 a_3463_4888.t6 527.402
R18582 a_3463_4888.n2 a_3463_4888.t2 491.64
R18583 a_3463_4888.n5 a_3463_4888.t0 281.906
R18584 a_3463_4888.t1 a_3463_4888.n5 204.359
R18585 a_3463_4888.n0 a_3463_4888.t7 180.73
R18586 a_3463_4888.n1 a_3463_4888.t5 179.45
R18587 a_3463_4888.n0 a_3463_4888.t3 139.78
R18588 a_3463_4888.n4 a_3463_4888.n1 105.635
R18589 a_3463_4888.n4 a_3463_4888.n3 76.0005
R18590 a_3463_4888.n5 a_3463_4888.n4 67.9685
R18591 a_3463_4888.n3 a_3463_4888.n2 13.994
R18592 a_3463_4888.n1 a_3463_4888.n0 1.28015
R18593 a_3493_5534.n1 a_3493_5534.n6 81.2978
R18594 a_3493_5534.n1 a_3493_5534.n5 81.1637
R18595 a_3493_5534.n0 a_3493_5534.n4 81.1637
R18596 a_3493_5534.n0 a_3493_5534.n3 81.1637
R18597 a_3493_5534.n7 a_3493_5534.n1 81.1637
R18598 a_3493_5534.n0 a_3493_5534.n2 80.9213
R18599 a_3493_5534.n6 a_3493_5534.t1 11.8205
R18600 a_3493_5534.n6 a_3493_5534.t0 11.8205
R18601 a_3493_5534.n5 a_3493_5534.t7 11.8205
R18602 a_3493_5534.n5 a_3493_5534.t8 11.8205
R18603 a_3493_5534.n4 a_3493_5534.t11 11.8205
R18604 a_3493_5534.n4 a_3493_5534.t10 11.8205
R18605 a_3493_5534.n3 a_3493_5534.t4 11.8205
R18606 a_3493_5534.n3 a_3493_5534.t9 11.8205
R18607 a_3493_5534.n2 a_3493_5534.t5 11.8205
R18608 a_3493_5534.n2 a_3493_5534.t3 11.8205
R18609 a_3493_5534.n7 a_3493_5534.t6 11.8205
R18610 a_3493_5534.t2 a_3493_5534.n7 11.8205
R18611 a_3493_5534.n1 a_3493_5534.n0 0.402735
R18612 NOT8_0.S7.n1 NOT8_0.S7.t4 1032.02
R18613 NOT8_0.S7.n1 NOT8_0.S7.t5 336.962
R18614 NOT8_0.S7.n1 NOT8_0.S7.t6 326.154
R18615 NOT8_0.S7.n0 NOT8_0.S7.t1 256.514
R18616 NOT8_0.S7.n0 NOT8_0.S7.n2 226.258
R18617 NOT8_0.S7 NOT8_0.S7.n1 162.952
R18618 NOT8_0.S7.n0 NOT8_0.S7.t3 83.7172
R18619 NOT8_0.S7.n2 NOT8_0.S7.t2 30.379
R18620 NOT8_0.S7.n2 NOT8_0.S7.t0 30.379
R18621 NOT8_0.S7 NOT8_0.S7.n0 1.94684
R18622 a_10459_n35461.t0 a_10459_n35461.t1 9.9005
R18623 mux8_6.NAND4F_7.Y.n2 mux8_6.NAND4F_7.Y.t11 1388.16
R18624 mux8_6.NAND4F_7.Y.n2 mux8_6.NAND4F_7.Y.t10 350.839
R18625 mux8_6.NAND4F_7.Y.n3 mux8_6.NAND4F_7.Y.t9 308.481
R18626 mux8_6.NAND4F_7.Y.n1 mux8_6.NAND4F_7.Y.n4 187.373
R18627 mux8_6.NAND4F_7.Y.n1 mux8_6.NAND4F_7.Y.n5 187.192
R18628 mux8_6.NAND4F_7.Y.n1 mux8_6.NAND4F_7.Y.n6 187.192
R18629 mux8_6.NAND4F_7.Y.n0 mux8_6.NAND4F_7.Y.n7 187.192
R18630 mux8_6.NAND4F_7.Y mux8_6.NAND4F_7.Y.n3 161.492
R18631 mux8_6.NAND4F_7.Y.n3 mux8_6.NAND4F_7.Y.n2 27.752
R18632 mux8_6.NAND4F_7.Y mux8_6.NAND4F_7.Y.t4 23.5642
R18633 mux8_6.NAND4F_7.Y.n4 mux8_6.NAND4F_7.Y.t1 20.1899
R18634 mux8_6.NAND4F_7.Y.n4 mux8_6.NAND4F_7.Y.t0 20.1899
R18635 mux8_6.NAND4F_7.Y.n5 mux8_6.NAND4F_7.Y.t2 20.1899
R18636 mux8_6.NAND4F_7.Y.n5 mux8_6.NAND4F_7.Y.t3 20.1899
R18637 mux8_6.NAND4F_7.Y.n6 mux8_6.NAND4F_7.Y.t8 20.1899
R18638 mux8_6.NAND4F_7.Y.n6 mux8_6.NAND4F_7.Y.t7 20.1899
R18639 mux8_6.NAND4F_7.Y.n7 mux8_6.NAND4F_7.Y.t6 20.1899
R18640 mux8_6.NAND4F_7.Y.n7 mux8_6.NAND4F_7.Y.t5 20.1899
R18641 mux8_6.NAND4F_7.Y mux8_6.NAND4F_7.Y.n0 0.472662
R18642 mux8_6.NAND4F_7.Y.n0 mux8_6.NAND4F_7.Y.n1 0.358709
R18643 a_n9125_n4534.n0 a_n9125_n4534.n2 81.2978
R18644 a_n9125_n4534.n0 a_n9125_n4534.n3 81.1637
R18645 a_n9125_n4534.n0 a_n9125_n4534.n4 81.1637
R18646 a_n9125_n4534.n1 a_n9125_n4534.n5 81.1637
R18647 a_n9125_n4534.n1 a_n9125_n4534.n6 81.1637
R18648 a_n9125_n4534.n7 a_n9125_n4534.n1 80.9213
R18649 a_n9125_n4534.n2 a_n9125_n4534.t11 11.8205
R18650 a_n9125_n4534.n2 a_n9125_n4534.t6 11.8205
R18651 a_n9125_n4534.n3 a_n9125_n4534.t5 11.8205
R18652 a_n9125_n4534.n3 a_n9125_n4534.t10 11.8205
R18653 a_n9125_n4534.n4 a_n9125_n4534.t3 11.8205
R18654 a_n9125_n4534.n4 a_n9125_n4534.t4 11.8205
R18655 a_n9125_n4534.n5 a_n9125_n4534.t2 11.8205
R18656 a_n9125_n4534.n5 a_n9125_n4534.t0 11.8205
R18657 a_n9125_n4534.n6 a_n9125_n4534.t7 11.8205
R18658 a_n9125_n4534.n6 a_n9125_n4534.t1 11.8205
R18659 a_n9125_n4534.t9 a_n9125_n4534.n7 11.8205
R18660 a_n9125_n4534.n7 a_n9125_n4534.t8 11.8205
R18661 a_n9125_n4534.n1 a_n9125_n4534.n0 0.402735
R18662 mux8_5.NAND4F_9.Y.n1 mux8_5.NAND4F_9.Y.t14 312.599
R18663 mux8_5.NAND4F_9.Y.n4 mux8_5.NAND4F_9.Y.t13 247.428
R18664 mux8_5.NAND4F_9.Y.n1 mux8_5.NAND4F_9.Y.t9 247.428
R18665 mux8_5.NAND4F_9.Y.n2 mux8_5.NAND4F_9.Y.t10 247.428
R18666 mux8_5.NAND4F_9.Y.n3 mux8_5.NAND4F_9.Y.t12 247.428
R18667 mux8_5.NAND4F_9.Y.n5 mux8_5.NAND4F_9.Y.t11 229.754
R18668 mux8_5.NAND4F_9.Y.n0 mux8_5.NAND4F_9.Y.n6 187.373
R18669 mux8_5.NAND4F_9.Y.n0 mux8_5.NAND4F_9.Y.n7 187.192
R18670 mux8_5.NAND4F_9.Y.n0 mux8_5.NAND4F_9.Y.n8 187.192
R18671 mux8_5.NAND4F_9.Y.n10 mux8_5.NAND4F_9.Y.n9 187.192
R18672 mux8_5.NAND4F_9.Y mux8_5.NAND4F_9.Y.n5 162.275
R18673 mux8_5.NAND4F_9.Y.n5 mux8_5.NAND4F_9.Y.n4 91.5805
R18674 mux8_5.NAND4F_9.Y.n2 mux8_5.NAND4F_9.Y.n1 65.1723
R18675 mux8_5.NAND4F_9.Y.n3 mux8_5.NAND4F_9.Y.n2 65.1723
R18676 mux8_5.NAND4F_9.Y.n4 mux8_5.NAND4F_9.Y.n3 65.1723
R18677 mux8_5.NAND4F_9.Y mux8_5.NAND4F_9.Y.t0 22.6141
R18678 mux8_5.NAND4F_9.Y.n6 mux8_5.NAND4F_9.Y.t3 20.1899
R18679 mux8_5.NAND4F_9.Y.n6 mux8_5.NAND4F_9.Y.t4 20.1899
R18680 mux8_5.NAND4F_9.Y.n7 mux8_5.NAND4F_9.Y.t7 20.1899
R18681 mux8_5.NAND4F_9.Y.n7 mux8_5.NAND4F_9.Y.t8 20.1899
R18682 mux8_5.NAND4F_9.Y.n8 mux8_5.NAND4F_9.Y.t5 20.1899
R18683 mux8_5.NAND4F_9.Y.n8 mux8_5.NAND4F_9.Y.t6 20.1899
R18684 mux8_5.NAND4F_9.Y.n9 mux8_5.NAND4F_9.Y.t2 20.1899
R18685 mux8_5.NAND4F_9.Y.n9 mux8_5.NAND4F_9.Y.t1 20.1899
R18686 mux8_5.NAND4F_9.Y mux8_5.NAND4F_9.Y.n10 0.396904
R18687 mux8_5.NAND4F_9.Y.n10 mux8_5.NAND4F_9.Y.n0 0.358709
R18688 a_10363_n30006.t0 a_10363_n30006.t1 9.9005
R18689 a_10459_n30006.t0 a_10459_n30006.t1 9.9005
R18690 a_n14077_3190.n2 a_n14077_3190.n0 121.353
R18691 a_n14077_3190.n3 a_n14077_3190.n2 121.353
R18692 a_n14077_3190.n2 a_n14077_3190.n1 121.001
R18693 a_n14077_3190.n1 a_n14077_3190.t3 30.462
R18694 a_n14077_3190.n1 a_n14077_3190.t1 30.462
R18695 a_n14077_3190.n0 a_n14077_3190.t4 30.462
R18696 a_n14077_3190.n0 a_n14077_3190.t5 30.462
R18697 a_n14077_3190.n3 a_n14077_3190.t0 30.462
R18698 a_n14077_3190.t2 a_n14077_3190.n3 30.462
R18699 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t15 491.64
R18700 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t22 491.64
R18701 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t21 491.64
R18702 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t18 491.64
R18703 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t12 485.221
R18704 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t17 367.928
R18705 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t14 255.588
R18706 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t23 224.478
R18707 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t16 213.688
R18708 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n0 209.19
R18709 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t19 139.78
R18710 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t20 139.78
R18711 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t13 139.78
R18712 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n11 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n10 120.999
R18713 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n11 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n9 120.999
R18714 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n23 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n22 104.489
R18715 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n13 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n12 92.5005
R18716 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n20 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n18 86.2638
R18717 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n18 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n17 85.8873
R18718 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n18 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n15 85.724
R18719 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n7 84.5046
R18720 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n23 83.8907
R18721 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n21 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n20 75.0672
R18722 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n21 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n17 75.0672
R18723 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n20 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n19 73.1255
R18724 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n17 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n16 73.1255
R18725 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n15 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n14 73.1255
R18726 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n6 72.3005
R18727 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n22 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n15 68.8946
R18728 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n8 60.9797
R18729 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n23 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n13 41.9827
R18730 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n12 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t3 30.462
R18731 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n12 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t7 30.462
R18732 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t6 30.462
R18733 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t10 30.462
R18734 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t5 30.462
R18735 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t4 30.462
R18736 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n13 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n11 28.124
R18737 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n5 19.963
R18738 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n1 17.8661
R18739 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n2 17.8661
R18740 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n3 17.1217
R18741 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n16 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t2 11.8205
R18742 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n16 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t1 11.8205
R18743 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n19 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t8 11.8205
R18744 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n19 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t11 11.8205
R18745 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n14 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t0 11.8205
R18746 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n14 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t9 11.8205
R18747 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n22 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n21 9.3005
R18748 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n4 1.8615
R18749 a_n12605_n12716.t0 a_n12605_n12716.t1 19.8005
R18750 a_n13714_n12716.t0 a_n13714_n12716.t1 19.8005
R18751 mux8_0.inv_0.A.n1 mux8_0.inv_0.A.t10 291.829
R18752 mux8_0.inv_0.A.n1 mux8_0.inv_0.A.t8 291.829
R18753 mux8_0.inv_0.A.n0 mux8_0.inv_0.A.t4 256.425
R18754 mux8_0.inv_0.A.n0 mux8_0.inv_0.A.n2 231.24
R18755 mux8_0.inv_0.A.n0 mux8_0.inv_0.A.n3 231.03
R18756 mux8_0.inv_0.A.n1 mux8_0.inv_0.A.t9 221.72
R18757 mux8_0.inv_0.A.t7 mux8_0.inv_0.A.n0 393.959
R18758 mux8_0.inv_0.A.n4 mux8_0.inv_0.A.n0 66.6316
R18759 mux8_0.inv_0.A.n0 mux8_0.inv_0.A.n1 54.1444
R18760 mux8_0.inv_0.A.n2 mux8_0.inv_0.A.t3 25.395
R18761 mux8_0.inv_0.A.n2 mux8_0.inv_0.A.t5 25.395
R18762 mux8_0.inv_0.A.n3 mux8_0.inv_0.A.t6 25.395
R18763 mux8_0.inv_0.A.n3 mux8_0.inv_0.A.t1 25.395
R18764 mux8_0.inv_0.A.n4 mux8_0.inv_0.A.t2 19.8005
R18765 mux8_0.inv_0.A.n4 mux8_0.inv_0.A.t0 19.8005
R18766 C.n1 C.t3 256.514
R18767 C.n1 C.n0 226.258
R18768 C C.t0 83.7296
R18769 C.n0 C.t1 30.379
R18770 C.n0 C.t2 30.379
R18771 C C.n1 0.0481763
R18772 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t10 540.38
R18773 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t7 367.928
R18774 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n4 227.526
R18775 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t9 227.356
R18776 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n6 227.266
R18777 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n5 227.266
R18778 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t8 213.688
R18779 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n2 160.439
R18780 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n1 94.4341
R18781 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t3 42.7943
R18782 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t4 30.379
R18783 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t5 30.379
R18784 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t2 30.379
R18785 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t0 30.379
R18786 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t6 30.379
R18787 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.t1 30.379
R18788 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n0 13.4358
R18789 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B.n3 0.821842
R18790 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n9 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t17 540.38
R18791 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t8 491.64
R18792 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t11 491.64
R18793 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t10 491.64
R18794 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t13 491.64
R18795 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t14 367.928
R18796 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n1 227.526
R18797 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n8 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t9 227.356
R18798 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n2 227.266
R18799 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n3 227.266
R18800 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t15 213.688
R18801 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n6 162.852
R18802 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n9 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n8 160.439
R18803 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t18 139.78
R18804 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t12 139.78
R18805 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t16 139.78
R18806 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t7 139.78
R18807 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n8 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n7 94.4341
R18808 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t0 42.7831
R18809 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n5 38.6833
R18810 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t6 30.379
R18811 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t4 30.379
R18812 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t1 30.379
R18813 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t5 30.379
R18814 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t3 30.379
R18815 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t2 30.379
R18816 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n4 28.3986
R18817 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n0 18.8832
R18818 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n10 10.7052
R18819 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n10 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT 5.09176
R18820 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n10 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT 4.19292
R18821 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n9 0.794268
R18822 MULT_0.NAND2_14.Y.n5 MULT_0.NAND2_14.Y.t8 291.829
R18823 MULT_0.NAND2_14.Y.n5 MULT_0.NAND2_14.Y.t7 291.829
R18824 MULT_0.NAND2_14.Y.n0 MULT_0.NAND2_14.Y.n3 227.526
R18825 MULT_0.NAND2_14.Y.n0 MULT_0.NAND2_14.Y.n2 227.266
R18826 MULT_0.NAND2_14.Y.n0 MULT_0.NAND2_14.Y.n4 227.266
R18827 MULT_0.NAND2_14.Y.n5 MULT_0.NAND2_14.Y.t10 221.72
R18828 MULT_0.NAND2_14.Y.t9 MULT_0.NAND2_14.Y.n1 393.897
R18829 MULT_0.NAND2_14.Y.n0 MULT_0.NAND2_14.Y.t6 42.7333
R18830 MULT_0.NAND2_14.Y.n3 MULT_0.NAND2_14.Y.t0 30.379
R18831 MULT_0.NAND2_14.Y.n3 MULT_0.NAND2_14.Y.t1 30.379
R18832 MULT_0.NAND2_14.Y.n2 MULT_0.NAND2_14.Y.t5 30.379
R18833 MULT_0.NAND2_14.Y.n2 MULT_0.NAND2_14.Y.t4 30.379
R18834 MULT_0.NAND2_14.Y.n4 MULT_0.NAND2_14.Y.t3 30.379
R18835 MULT_0.NAND2_14.Y.n4 MULT_0.NAND2_14.Y.t2 30.379
R18836 MULT_0.NAND2_14.Y.n5 MULT_0.NAND2_14.Y.n1 53.4913
R18837 MULT_0.NAND2_14.Y.n0 MULT_0.NAND2_14.Y.n1 0.621694
R18838 a_n12345_n17857.n2 a_n12345_n17857.t4 539.788
R18839 a_n12345_n17857.n3 a_n12345_n17857.t6 531.496
R18840 a_n12345_n17857.n2 a_n12345_n17857.t5 490.034
R18841 a_n12345_n17857.n5 a_n12345_n17857.t0 283.788
R18842 a_n12345_n17857.t1 a_n12345_n17857.n5 205.489
R18843 a_n12345_n17857.n0 a_n12345_n17857.t7 182.625
R18844 a_n12345_n17857.n1 a_n12345_n17857.t3 179.054
R18845 a_n12345_n17857.n0 a_n12345_n17857.t2 139.78
R18846 a_n12345_n17857.n4 a_n12345_n17857.n1 101.368
R18847 a_n12345_n17857.n5 a_n12345_n17857.n4 77.9135
R18848 a_n12345_n17857.n4 a_n12345_n17857.n3 76.1557
R18849 a_n12345_n17857.n3 a_n12345_n17857.n2 8.29297
R18850 a_n12345_n17857.n1 a_n12345_n17857.n0 3.57087
R18851 a_n4205_3190.n2 a_n4205_3190.n1 121.353
R18852 a_n4205_3190.n2 a_n4205_3190.n0 121.353
R18853 a_n4205_3190.n3 a_n4205_3190.n2 121.001
R18854 a_n4205_3190.n1 a_n4205_3190.t0 30.462
R18855 a_n4205_3190.n1 a_n4205_3190.t1 30.462
R18856 a_n4205_3190.n0 a_n4205_3190.t4 30.462
R18857 a_n4205_3190.n0 a_n4205_3190.t5 30.462
R18858 a_n4205_3190.n3 a_n4205_3190.t3 30.462
R18859 a_n4205_3190.t2 a_n4205_3190.n3 30.462
R18860 MULT_0.4bit_ADDER_0.B0.n6 MULT_0.4bit_ADDER_0.B0.t11 491.64
R18861 MULT_0.4bit_ADDER_0.B0.n7 MULT_0.4bit_ADDER_0.B0.t6 491.64
R18862 MULT_0.4bit_ADDER_0.B0.n8 MULT_0.4bit_ADDER_0.B0.t7 491.64
R18863 MULT_0.4bit_ADDER_0.B0.n9 MULT_0.4bit_ADDER_0.B0.t12 491.64
R18864 MULT_0.4bit_ADDER_0.B0.n4 MULT_0.4bit_ADDER_0.B0.t8 485.221
R18865 MULT_0.4bit_ADDER_0.B0.n2 MULT_0.4bit_ADDER_0.B0.t14 367.928
R18866 MULT_0.4bit_ADDER_0.B0.n0 MULT_0.4bit_ADDER_0.B0.t1 256.514
R18867 MULT_0.4bit_ADDER_0.B0.n10 MULT_0.4bit_ADDER_0.B0.t10 255.588
R18868 MULT_0.4bit_ADDER_0.B0.n0 MULT_0.4bit_ADDER_0.B0.n1 226.251
R18869 MULT_0.4bit_ADDER_0.B0.n3 MULT_0.4bit_ADDER_0.B0.t4 224.478
R18870 MULT_0.4bit_ADDER_0.B0.n2 MULT_0.4bit_ADDER_0.B0.t15 213.688
R18871 MULT_0.4bit_ADDER_0.B0.n6 MULT_0.4bit_ADDER_0.B0.n5 209.19
R18872 MULT_0.4bit_ADDER_0.B0.n5 MULT_0.4bit_ADDER_0.B0.t9 139.78
R18873 MULT_0.4bit_ADDER_0.B0.n5 MULT_0.4bit_ADDER_0.B0.t5 139.78
R18874 MULT_0.4bit_ADDER_0.B0.n5 MULT_0.4bit_ADDER_0.B0.t13 139.78
R18875 MULT_0.4bit_ADDER_0.B0.n11 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_0.A 103.258
R18876 MULT_0.4bit_ADDER_0.B0.n4 MULT_0.4bit_ADDER_0.B0.n3 84.5046
R18877 MULT_0.4bit_ADDER_0.B0.n0 MULT_0.4bit_ADDER_0.B0.t0 83.7599
R18878 MULT_0.4bit_ADDER_0.B0.n3 MULT_0.4bit_ADDER_0.B0.n2 72.3005
R18879 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_0.A MULT_0.4bit_ADDER_0.B0.n4 60.9816
R18880 MULT_0.4bit_ADDER_0.B0.n1 MULT_0.4bit_ADDER_0.B0.t3 30.379
R18881 MULT_0.4bit_ADDER_0.B0.n1 MULT_0.4bit_ADDER_0.B0.t2 30.379
R18882 MULT_0.4bit_ADDER_0.FULL_ADDER_3.B MULT_0.4bit_ADDER_0.B0.n0 19.8902
R18883 MULT_0.4bit_ADDER_0.B0.n7 MULT_0.4bit_ADDER_0.B0.n6 17.8661
R18884 MULT_0.4bit_ADDER_0.B0.n8 MULT_0.4bit_ADDER_0.B0.n7 17.8661
R18885 MULT_0.4bit_ADDER_0.B0.n9 MULT_0.4bit_ADDER_0.B0.n8 17.1217
R18886 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_0.A MULT_0.4bit_ADDER_0.B0.n10 15.6329
R18887 MULT_0.4bit_ADDER_0.B0.n11 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_0.A 10.8165
R18888 MULT_0.4bit_ADDER_0.B0.n10 MULT_0.4bit_ADDER_0.B0.n9 1.8615
R18889 MULT_0.4bit_ADDER_0.FULL_ADDER_3.B MULT_0.4bit_ADDER_0.B0.n11 0.868831
R18890 mux8_6.NAND4F_4.B.n10 mux8_6.NAND4F_4.B.t14 933.563
R18891 mux8_6.NAND4F_4.B.n5 mux8_6.NAND4F_4.B.t6 933.563
R18892 mux8_6.NAND4F_4.B.n3 mux8_6.NAND4F_4.B.t9 933.563
R18893 mux8_6.NAND4F_4.B.n1 mux8_6.NAND4F_4.B.t5 933.563
R18894 mux8_6.NAND4F_4.B.n10 mux8_6.NAND4F_4.B.t10 367.635
R18895 mux8_6.NAND4F_4.B.n5 mux8_6.NAND4F_4.B.t7 367.635
R18896 mux8_6.NAND4F_4.B.n3 mux8_6.NAND4F_4.B.t11 367.635
R18897 mux8_6.NAND4F_4.B.n1 mux8_6.NAND4F_4.B.t15 367.635
R18898 mux8_6.NAND4F_4.B.n11 mux8_6.NAND4F_4.B.t12 308.481
R18899 mux8_6.NAND4F_4.B.n6 mux8_6.NAND4F_4.B.t8 308.481
R18900 mux8_6.NAND4F_4.B.n4 mux8_6.NAND4F_4.B.t13 308.481
R18901 mux8_6.NAND4F_4.B.n2 mux8_6.NAND4F_4.B.t4 308.481
R18902 mux8_6.NAND4F_4.B.n0 mux8_6.NAND4F_4.B.t1 256.514
R18903 mux8_6.NAND4F_4.B.n0 mux8_6.NAND4F_4.B.n8 226.258
R18904 mux8_6.NAND4F_4.B mux8_6.NAND4F_4.B.n2 162.173
R18905 mux8_6.NAND4F_4.B mux8_6.NAND4F_4.B.n6 162.137
R18906 mux8_6.NAND4F_4.B mux8_6.NAND4F_4.B.n11 162.117
R18907 mux8_6.NAND4F_4.B.n7 mux8_6.NAND4F_4.B.n4 161.703
R18908 mux8_6.NAND4F_4.B.n0 mux8_6.NAND4F_4.B.t0 83.7172
R18909 mux8_6.NAND4F_4.B.n8 mux8_6.NAND4F_4.B.t3 30.379
R18910 mux8_6.NAND4F_4.B.n8 mux8_6.NAND4F_4.B.t2 30.379
R18911 mux8_6.NAND4F_4.B.n12 mux8_6.NAND4F_4.B 24.8912
R18912 mux8_6.NAND4F_4.B.n7 mux8_6.NAND4F_4.B 21.6618
R18913 mux8_6.NAND4F_4.B.n11 mux8_6.NAND4F_4.B.n10 10.955
R18914 mux8_6.NAND4F_4.B.n6 mux8_6.NAND4F_4.B.n5 10.955
R18915 mux8_6.NAND4F_4.B.n4 mux8_6.NAND4F_4.B.n3 10.955
R18916 mux8_6.NAND4F_4.B.n2 mux8_6.NAND4F_4.B.n1 10.955
R18917 mux8_6.NAND4F_4.B.n12 mux8_6.NAND4F_4.B.n9 3.67985
R18918 mux8_6.NAND4F_4.B.n9 mux8_6.NAND4F_4.B.n0 1.46835
R18919 mux8_6.NAND4F_4.B mux8_6.NAND4F_4.B.n12 0.502677
R18920 mux8_6.NAND4F_4.B.n9 mux8_6.NAND4F_4.B 0.498606
R18921 mux8_6.NAND4F_4.B mux8_6.NAND4F_4.B.n7 0.470197
R18922 mux8_6.NAND4F_5.Y.n1 mux8_6.NAND4F_5.Y.t9 1032.02
R18923 mux8_6.NAND4F_5.Y.n1 mux8_6.NAND4F_5.Y.t10 336.962
R18924 mux8_6.NAND4F_5.Y.n1 mux8_6.NAND4F_5.Y.t11 326.154
R18925 mux8_6.NAND4F_5.Y.n0 mux8_6.NAND4F_5.Y.n3 187.373
R18926 mux8_6.NAND4F_5.Y.n0 mux8_6.NAND4F_5.Y.n4 187.192
R18927 mux8_6.NAND4F_5.Y.n0 mux8_6.NAND4F_5.Y.n5 187.192
R18928 mux8_6.NAND4F_5.Y.n7 mux8_6.NAND4F_5.Y.n6 187.192
R18929 mux8_6.NAND4F_5.Y mux8_6.NAND4F_5.Y.n1 162.94
R18930 mux8_6.NAND4F_5.Y.n2 mux8_6.NAND4F_5.Y 24.4721
R18931 mux8_6.NAND4F_5.Y.n2 mux8_6.NAND4F_5.Y.t2 22.6141
R18932 mux8_6.NAND4F_5.Y.n3 mux8_6.NAND4F_5.Y.t1 20.1899
R18933 mux8_6.NAND4F_5.Y.n3 mux8_6.NAND4F_5.Y.t0 20.1899
R18934 mux8_6.NAND4F_5.Y.n4 mux8_6.NAND4F_5.Y.t6 20.1899
R18935 mux8_6.NAND4F_5.Y.n4 mux8_6.NAND4F_5.Y.t5 20.1899
R18936 mux8_6.NAND4F_5.Y.n5 mux8_6.NAND4F_5.Y.t7 20.1899
R18937 mux8_6.NAND4F_5.Y.n5 mux8_6.NAND4F_5.Y.t8 20.1899
R18938 mux8_6.NAND4F_5.Y.n6 mux8_6.NAND4F_5.Y.t4 20.1899
R18939 mux8_6.NAND4F_5.Y.n6 mux8_6.NAND4F_5.Y.t3 20.1899
R18940 mux8_6.NAND4F_5.Y mux8_6.NAND4F_5.Y.n2 0.950576
R18941 mux8_6.NAND4F_5.Y mux8_6.NAND4F_5.Y.n7 0.396904
R18942 mux8_6.NAND4F_5.Y.n7 mux8_6.NAND4F_5.Y.n0 0.358709
R18943 a_n11274_n18115.n2 a_n11274_n18115.n1 121.353
R18944 a_n11274_n18115.n3 a_n11274_n18115.n2 121.001
R18945 a_n11274_n18115.n2 a_n11274_n18115.n0 120.977
R18946 a_n11274_n18115.n0 a_n11274_n18115.t3 30.462
R18947 a_n11274_n18115.n0 a_n11274_n18115.t5 30.462
R18948 a_n11274_n18115.n1 a_n11274_n18115.t1 30.462
R18949 a_n11274_n18115.n1 a_n11274_n18115.t2 30.462
R18950 a_n11274_n18115.t4 a_n11274_n18115.n3 30.462
R18951 a_n11274_n18115.n3 a_n11274_n18115.t0 30.462
R18952 a_9336_n12822.t0 a_9336_n12822.t1 9.9005
R18953 a_n914_3810.n0 a_n914_3810.n2 81.2978
R18954 a_n914_3810.n1 a_n914_3810.n5 81.1637
R18955 a_n914_3810.n0 a_n914_3810.n4 81.1637
R18956 a_n914_3810.n0 a_n914_3810.n3 81.1637
R18957 a_n914_3810.n7 a_n914_3810.n1 81.1637
R18958 a_n914_3810.n1 a_n914_3810.n6 80.9213
R18959 a_n914_3810.n6 a_n914_3810.t0 11.8205
R18960 a_n914_3810.n6 a_n914_3810.t1 11.8205
R18961 a_n914_3810.n5 a_n914_3810.t5 11.8205
R18962 a_n914_3810.n5 a_n914_3810.t4 11.8205
R18963 a_n914_3810.n4 a_n914_3810.t10 11.8205
R18964 a_n914_3810.n4 a_n914_3810.t9 11.8205
R18965 a_n914_3810.n3 a_n914_3810.t6 11.8205
R18966 a_n914_3810.n3 a_n914_3810.t11 11.8205
R18967 a_n914_3810.n2 a_n914_3810.t7 11.8205
R18968 a_n914_3810.n2 a_n914_3810.t8 11.8205
R18969 a_n914_3810.n7 a_n914_3810.t3 11.8205
R18970 a_n914_3810.t2 a_n914_3810.n7 11.8205
R18971 a_n914_3810.n1 a_n914_3810.n0 0.402735
R18972 a_n11840_n5154.n2 a_n11840_n5154.n1 121.353
R18973 a_n11840_n5154.n2 a_n11840_n5154.n0 121.353
R18974 a_n11840_n5154.n3 a_n11840_n5154.n2 121.001
R18975 a_n11840_n5154.n1 a_n11840_n5154.t4 30.462
R18976 a_n11840_n5154.n1 a_n11840_n5154.t3 30.462
R18977 a_n11840_n5154.n0 a_n11840_n5154.t1 30.462
R18978 a_n11840_n5154.n0 a_n11840_n5154.t0 30.462
R18979 a_n11840_n5154.t2 a_n11840_n5154.n3 30.462
R18980 a_n11840_n5154.n3 a_n11840_n5154.t5 30.462
R18981 MULT_0.NAND2_11.Y.n5 MULT_0.NAND2_11.Y.t9 291.829
R18982 MULT_0.NAND2_11.Y.n5 MULT_0.NAND2_11.Y.t7 291.829
R18983 MULT_0.NAND2_11.Y.n0 MULT_0.NAND2_11.Y.n3 227.526
R18984 MULT_0.NAND2_11.Y.n0 MULT_0.NAND2_11.Y.n2 227.266
R18985 MULT_0.NAND2_11.Y.n0 MULT_0.NAND2_11.Y.n4 227.266
R18986 MULT_0.NAND2_11.Y.n5 MULT_0.NAND2_11.Y.t10 221.72
R18987 MULT_0.NAND2_11.Y.t8 MULT_0.NAND2_11.Y.n1 393.897
R18988 MULT_0.NAND2_11.Y.n0 MULT_0.NAND2_11.Y.t3 42.7333
R18989 MULT_0.NAND2_11.Y.n3 MULT_0.NAND2_11.Y.t1 30.379
R18990 MULT_0.NAND2_11.Y.n3 MULT_0.NAND2_11.Y.t0 30.379
R18991 MULT_0.NAND2_11.Y.n2 MULT_0.NAND2_11.Y.t6 30.379
R18992 MULT_0.NAND2_11.Y.n2 MULT_0.NAND2_11.Y.t5 30.379
R18993 MULT_0.NAND2_11.Y.n4 MULT_0.NAND2_11.Y.t4 30.379
R18994 MULT_0.NAND2_11.Y.n4 MULT_0.NAND2_11.Y.t2 30.379
R18995 MULT_0.NAND2_11.Y.n5 MULT_0.NAND2_11.Y.n1 53.4914
R18996 MULT_0.NAND2_11.Y.n0 MULT_0.NAND2_11.Y.n1 0.622011
R18997 mux8_8.NAND4F_5.Y.n1 mux8_8.NAND4F_5.Y.t9 1032.02
R18998 mux8_8.NAND4F_5.Y.n1 mux8_8.NAND4F_5.Y.t10 336.962
R18999 mux8_8.NAND4F_5.Y.n1 mux8_8.NAND4F_5.Y.t11 326.154
R19000 mux8_8.NAND4F_5.Y.n0 mux8_8.NAND4F_5.Y.n3 187.373
R19001 mux8_8.NAND4F_5.Y.n0 mux8_8.NAND4F_5.Y.n4 187.192
R19002 mux8_8.NAND4F_5.Y.n0 mux8_8.NAND4F_5.Y.n5 187.192
R19003 mux8_8.NAND4F_5.Y.n7 mux8_8.NAND4F_5.Y.n6 187.192
R19004 mux8_8.NAND4F_5.Y mux8_8.NAND4F_5.Y.n1 162.94
R19005 mux8_8.NAND4F_5.Y.n2 mux8_8.NAND4F_5.Y 24.4721
R19006 mux8_8.NAND4F_5.Y.n2 mux8_8.NAND4F_5.Y.t2 22.6141
R19007 mux8_8.NAND4F_5.Y.n3 mux8_8.NAND4F_5.Y.t0 20.1899
R19008 mux8_8.NAND4F_5.Y.n3 mux8_8.NAND4F_5.Y.t1 20.1899
R19009 mux8_8.NAND4F_5.Y.n4 mux8_8.NAND4F_5.Y.t6 20.1899
R19010 mux8_8.NAND4F_5.Y.n4 mux8_8.NAND4F_5.Y.t5 20.1899
R19011 mux8_8.NAND4F_5.Y.n5 mux8_8.NAND4F_5.Y.t7 20.1899
R19012 mux8_8.NAND4F_5.Y.n5 mux8_8.NAND4F_5.Y.t8 20.1899
R19013 mux8_8.NAND4F_5.Y.n6 mux8_8.NAND4F_5.Y.t3 20.1899
R19014 mux8_8.NAND4F_5.Y.n6 mux8_8.NAND4F_5.Y.t4 20.1899
R19015 mux8_8.NAND4F_5.Y mux8_8.NAND4F_5.Y.n2 0.950576
R19016 mux8_8.NAND4F_5.Y mux8_8.NAND4F_5.Y.n7 0.396904
R19017 mux8_8.NAND4F_5.Y.n7 mux8_8.NAND4F_5.Y.n0 0.358709
R19018 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t16 491.64
R19019 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t18 491.64
R19020 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t19 491.64
R19021 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t17 491.64
R19022 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n8 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t14 485.221
R19023 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t20 367.928
R19024 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t12 255.588
R19025 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t15 224.478
R19026 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t21 213.688
R19027 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n0 209.19
R19028 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t22 139.78
R19029 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t23 139.78
R19030 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t13 139.78
R19031 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n11 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n10 120.999
R19032 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n11 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n9 120.999
R19033 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n23 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n22 104.489
R19034 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n13 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n12 92.5005
R19035 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n20 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n18 86.2638
R19036 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n18 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n17 85.8873
R19037 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n18 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n15 85.724
R19038 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n8 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n7 84.5046
R19039 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n23 83.8907
R19040 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n21 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n20 75.0672
R19041 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n21 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n17 75.0672
R19042 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n20 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n19 73.1255
R19043 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n17 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n16 73.1255
R19044 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n15 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n14 73.1255
R19045 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n6 72.3005
R19046 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n22 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n15 68.8946
R19047 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n8 60.9797
R19048 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n23 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n13 41.9827
R19049 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n12 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t9 30.462
R19050 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n12 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t3 30.462
R19051 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n10 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t4 30.462
R19052 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n10 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t7 30.462
R19053 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n9 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t10 30.462
R19054 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n9 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t11 30.462
R19055 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n13 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n11 28.124
R19056 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n5 19.963
R19057 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n1 17.8661
R19058 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n2 17.8661
R19059 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n3 17.1217
R19060 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n16 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t1 11.8205
R19061 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n16 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t2 11.8205
R19062 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n19 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t6 11.8205
R19063 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n19 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t8 11.8205
R19064 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n14 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t0 11.8205
R19065 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n14 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t5 11.8205
R19066 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n22 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n21 9.3005
R19067 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n4 1.8615
R19068 a_n15887_n5154.n0 a_n15887_n5154.t5 539.788
R19069 a_n15887_n5154.n1 a_n15887_n5154.t2 531.496
R19070 a_n15887_n5154.n0 a_n15887_n5154.t6 490.034
R19071 a_n15887_n5154.n5 a_n15887_n5154.t0 283.788
R19072 a_n15887_n5154.t1 a_n15887_n5154.n5 205.489
R19073 a_n15887_n5154.n2 a_n15887_n5154.t3 182.625
R19074 a_n15887_n5154.n3 a_n15887_n5154.t7 179.054
R19075 a_n15887_n5154.n2 a_n15887_n5154.t4 139.78
R19076 a_n15887_n5154.n4 a_n15887_n5154.n3 101.368
R19077 a_n15887_n5154.n5 a_n15887_n5154.n4 77.9135
R19078 a_n15887_n5154.n4 a_n15887_n5154.n1 76.1557
R19079 a_n15887_n5154.n1 a_n15887_n5154.n0 8.29297
R19080 a_n15887_n5154.n3 a_n15887_n5154.n2 3.57087
R19081 B2.n10 B2.t46 540.38
R19082 B2.n17 B2.t3 540.38
R19083 B2.n6 B2.t1 491.64
R19084 B2.n5 B2.t25 491.64
R19085 B2.n4 B2.t15 491.64
R19086 B2.n3 B2.t5 491.64
R19087 B2.n38 B2.t45 491.64
R19088 B2.n37 B2.t50 491.64
R19089 B2.n36 B2.t30 491.64
R19090 B2.n35 B2.t11 491.64
R19091 B2.n25 B2.t19 485.443
R19092 B2.n13 B2.t0 485.221
R19093 B2.n20 B2.t21 485.221
R19094 B2.n43 B2.t48 394.37
R19095 B2.n47 B2.t20 394.37
R19096 B2.n1 B2.t22 394.37
R19097 B2.n28 B2.t26 379.173
R19098 B2.n8 B2.t9 367.928
R19099 B2.n11 B2.t34 367.928
R19100 B2.n15 B2.t18 367.928
R19101 B2.n18 B2.t8 367.928
R19102 B2.n23 B2.t49 343.827
R19103 B2.n29 B2.t17 312.599
R19104 B2.n42 B2.t7 291.829
R19105 B2.n42 B2.t6 291.829
R19106 B2.n46 B2.t35 291.829
R19107 B2.n46 B2.t10 291.829
R19108 B2.n0 B2.t44 291.829
R19109 B2.n0 B2.t42 291.829
R19110 B2.n7 B2.t47 255.588
R19111 B2.n39 B2.t16 255.588
R19112 B2.n29 B2.t4 247.428
R19113 B2.n30 B2.t2 247.428
R19114 B2.n31 B2.t31 247.428
R19115 B2.n28 B2.t27 247.428
R19116 B2.n40 B2 237.934
R19117 B2.n23 B2.t52 237.787
R19118 B2.n9 B2.t32 227.356
R19119 B2.n16 B2.t39 227.356
R19120 B2.n24 B2.t14 224.478
R19121 B2.n12 B2.t43 224.478
R19122 B2.n19 B2.t29 224.478
R19123 B2.n42 B2.t23 221.72
R19124 B2.n46 B2.t38 221.72
R19125 B2.n0 B2.t37 221.72
R19126 B2.n8 B2.t13 213.688
R19127 B2.n11 B2.t41 213.688
R19128 B2.n15 B2.t40 213.688
R19129 B2.n18 B2.t24 213.688
R19130 B2.n35 B2.n34 209.407
R19131 B2.n3 B2.n2 209.19
R19132 B2 B2.n32 162.139
R19133 B2.n10 B2.n9 160.439
R19134 B2.n17 B2.n16 160.439
R19135 B2.n2 B2.t36 139.78
R19136 B2.n2 B2.t51 139.78
R19137 B2.n2 B2.t12 139.78
R19138 B2.n34 B2.t33 139.78
R19139 B2.n34 B2.t53 139.78
R19140 B2.n34 B2.t28 139.78
R19141 B2.n9 B2.n8 94.4341
R19142 B2.n16 B2.n15 94.4341
R19143 B2.n13 B2.n12 84.5046
R19144 B2.n20 B2.n19 84.5046
R19145 B2.n25 B2.n24 83.8438
R19146 B2.n12 B2.n11 72.3005
R19147 B2.n19 B2.n18 72.3005
R19148 B2.n31 B2.n30 65.1723
R19149 B2.n30 B2.n29 65.1723
R19150 B2 B2.n13 61.0566
R19151 B2 B2.n20 61.0566
R19152 B2 B2.n25 61.0461
R19153 B2.n43 B2.n42 53.374
R19154 B2.n47 B2.n46 53.374
R19155 B2.n1 B2.n0 53.374
R19156 B2.n24 B2.n23 48.2005
R19157 B2.n22 B2 36.6239
R19158 B2.n32 B2.n31 33.2653
R19159 B2.n32 B2.n28 31.9075
R19160 B2 B2.n39 27.4136
R19161 B2.n5 B2.n4 17.8661
R19162 B2.n4 B2.n3 17.8661
R19163 B2.n36 B2.n35 17.8661
R19164 B2.n37 B2.n36 17.8661
R19165 B2.n6 B2.n5 17.1217
R19166 B2.n38 B2.n37 17.1217
R19167 B2.n50 B2.n49 14.2301
R19168 B2.n45 B2.n44 12.5554
R19169 B2.n33 B2 12.443
R19170 B2.n27 B2.n26 12.4105
R19171 B2.n41 B2.n40 12.4105
R19172 B2.n49 B2.n48 12.4105
R19173 B2 B2.n7 11.1665
R19174 B2.n22 B2.n21 7.20514
R19175 B2 B2.n22 7.06326
R19176 B2.n45 B2.n41 5.81514
R19177 B2.n41 B2.n33 5.73181
R19178 B2.n21 B2 5.10536
R19179 B2.n33 B2.n27 4.8791
R19180 B2.n14 B2 3.60258
R19181 B2.n21 B2 3.33577
R19182 B2.n14 B2 3.32643
R19183 B2.n49 B2.n45 2.71605
R19184 B2.n7 B2.n6 1.8615
R19185 B2.n39 B2.n38 1.8615
R19186 B2 B2.n14 1.26161
R19187 B2.n26 B2 1.25791
R19188 B2.n44 B2.n43 1.22678
R19189 B2 B2.n17 0.900886
R19190 B2 B2.n10 0.898246
R19191 B2.n50 B2.n1 0.756483
R19192 B2.n48 B2.n47 0.751965
R19193 B2.n21 B2 0.17087
R19194 B2.n48 B2 0.0667651
R19195 B2.n26 B2 0.0665714
R19196 B2 B2.n50 0.062247
R19197 B2.n44 B2 0.058471
R19198 B2.n40 B2 0.0390638
R19199 B2.n27 B2 0.0146
R19200 a_n22426_n9284.t0 a_n22426_n9284.t1 19.8005
R19201 NOT8_0.S6.n1 NOT8_0.S6.t5 1032.02
R19202 NOT8_0.S6.n1 NOT8_0.S6.t6 336.962
R19203 NOT8_0.S6.n1 NOT8_0.S6.t4 326.154
R19204 NOT8_0.S6.n0 NOT8_0.S6.t3 256.514
R19205 NOT8_0.S6.n0 NOT8_0.S6.n2 226.258
R19206 NOT8_0.S6 NOT8_0.S6.n1 162.952
R19207 NOT8_0.S6.n0 NOT8_0.S6.t0 83.7172
R19208 NOT8_0.S6.n2 NOT8_0.S6.t1 30.379
R19209 NOT8_0.S6.n2 NOT8_0.S6.t2 30.379
R19210 NOT8_0.S6 NOT8_0.S6.n0 1.95466
R19211 mux8_8.NAND4F_7.Y.n2 mux8_8.NAND4F_7.Y.t11 1388.16
R19212 mux8_8.NAND4F_7.Y.n2 mux8_8.NAND4F_7.Y.t10 350.839
R19213 mux8_8.NAND4F_7.Y.n3 mux8_8.NAND4F_7.Y.t9 308.481
R19214 mux8_8.NAND4F_7.Y.n1 mux8_8.NAND4F_7.Y.n4 187.373
R19215 mux8_8.NAND4F_7.Y.n1 mux8_8.NAND4F_7.Y.n5 187.192
R19216 mux8_8.NAND4F_7.Y.n1 mux8_8.NAND4F_7.Y.n6 187.192
R19217 mux8_8.NAND4F_7.Y.n0 mux8_8.NAND4F_7.Y.n7 187.192
R19218 mux8_8.NAND4F_7.Y mux8_8.NAND4F_7.Y.n3 161.492
R19219 mux8_8.NAND4F_7.Y.n3 mux8_8.NAND4F_7.Y.n2 27.752
R19220 mux8_8.NAND4F_7.Y mux8_8.NAND4F_7.Y.t8 23.5642
R19221 mux8_8.NAND4F_7.Y.n4 mux8_8.NAND4F_7.Y.t1 20.1899
R19222 mux8_8.NAND4F_7.Y.n4 mux8_8.NAND4F_7.Y.t0 20.1899
R19223 mux8_8.NAND4F_7.Y.n5 mux8_8.NAND4F_7.Y.t2 20.1899
R19224 mux8_8.NAND4F_7.Y.n5 mux8_8.NAND4F_7.Y.t3 20.1899
R19225 mux8_8.NAND4F_7.Y.n6 mux8_8.NAND4F_7.Y.t5 20.1899
R19226 mux8_8.NAND4F_7.Y.n6 mux8_8.NAND4F_7.Y.t4 20.1899
R19227 mux8_8.NAND4F_7.Y.n7 mux8_8.NAND4F_7.Y.t6 20.1899
R19228 mux8_8.NAND4F_7.Y.n7 mux8_8.NAND4F_7.Y.t7 20.1899
R19229 mux8_8.NAND4F_7.Y mux8_8.NAND4F_7.Y.n0 0.472662
R19230 mux8_8.NAND4F_7.Y.n0 mux8_8.NAND4F_7.Y.n1 0.358709
R19231 right_shifter_0.buffer_2.inv_1.A.n0 right_shifter_0.buffer_2.inv_1.A.t4 393.921
R19232 right_shifter_0.buffer_2.inv_1.A.n2 right_shifter_0.buffer_2.inv_1.A.t7 291.829
R19233 right_shifter_0.buffer_2.inv_1.A.n2 right_shifter_0.buffer_2.inv_1.A.t6 291.829
R19234 right_shifter_0.buffer_2.inv_1.A.n0 right_shifter_0.buffer_2.inv_1.A.t1 256.514
R19235 right_shifter_0.buffer_2.inv_1.A.n0 right_shifter_0.buffer_2.inv_1.A.n1 226.162
R19236 right_shifter_0.buffer_2.inv_1.A.n2 right_shifter_0.buffer_2.inv_1.A.t5 221.72
R19237 right_shifter_0.buffer_2.inv_1.A.n0 right_shifter_0.buffer_2.inv_1.A.t0 83.795
R19238 right_shifter_0.buffer_2.inv_1.A.n0 right_shifter_0.buffer_2.inv_1.A.n2 53.7938
R19239 right_shifter_0.buffer_2.inv_1.A.n1 right_shifter_0.buffer_2.inv_1.A.t3 30.379
R19240 right_shifter_0.buffer_2.inv_1.A.n1 right_shifter_0.buffer_2.inv_1.A.t2 30.379
R19241 a_11386_n26406.t0 a_11386_n26406.t1 9.9005
R19242 mux8_7.NAND4F_9.Y.n1 mux8_7.NAND4F_9.Y.t12 312.599
R19243 mux8_7.NAND4F_9.Y.n4 mux8_7.NAND4F_9.Y.t10 247.428
R19244 mux8_7.NAND4F_9.Y.n1 mux8_7.NAND4F_9.Y.t13 247.428
R19245 mux8_7.NAND4F_9.Y.n2 mux8_7.NAND4F_9.Y.t14 247.428
R19246 mux8_7.NAND4F_9.Y.n3 mux8_7.NAND4F_9.Y.t9 247.428
R19247 mux8_7.NAND4F_9.Y.n5 mux8_7.NAND4F_9.Y.t11 229.754
R19248 mux8_7.NAND4F_9.Y.n0 mux8_7.NAND4F_9.Y.n6 187.373
R19249 mux8_7.NAND4F_9.Y.n0 mux8_7.NAND4F_9.Y.n7 187.192
R19250 mux8_7.NAND4F_9.Y.n0 mux8_7.NAND4F_9.Y.n8 187.192
R19251 mux8_7.NAND4F_9.Y.n10 mux8_7.NAND4F_9.Y.n9 187.192
R19252 mux8_7.NAND4F_9.Y mux8_7.NAND4F_9.Y.n5 162.275
R19253 mux8_7.NAND4F_9.Y.n5 mux8_7.NAND4F_9.Y.n4 91.5805
R19254 mux8_7.NAND4F_9.Y.n2 mux8_7.NAND4F_9.Y.n1 65.1723
R19255 mux8_7.NAND4F_9.Y.n3 mux8_7.NAND4F_9.Y.n2 65.1723
R19256 mux8_7.NAND4F_9.Y.n4 mux8_7.NAND4F_9.Y.n3 65.1723
R19257 mux8_7.NAND4F_9.Y mux8_7.NAND4F_9.Y.t4 22.6141
R19258 mux8_7.NAND4F_9.Y.n6 mux8_7.NAND4F_9.Y.t0 20.1899
R19259 mux8_7.NAND4F_9.Y.n6 mux8_7.NAND4F_9.Y.t1 20.1899
R19260 mux8_7.NAND4F_9.Y.n7 mux8_7.NAND4F_9.Y.t7 20.1899
R19261 mux8_7.NAND4F_9.Y.n7 mux8_7.NAND4F_9.Y.t8 20.1899
R19262 mux8_7.NAND4F_9.Y.n8 mux8_7.NAND4F_9.Y.t2 20.1899
R19263 mux8_7.NAND4F_9.Y.n8 mux8_7.NAND4F_9.Y.t3 20.1899
R19264 mux8_7.NAND4F_9.Y.n9 mux8_7.NAND4F_9.Y.t6 20.1899
R19265 mux8_7.NAND4F_9.Y.n9 mux8_7.NAND4F_9.Y.t5 20.1899
R19266 mux8_7.NAND4F_9.Y mux8_7.NAND4F_9.Y.n10 0.396904
R19267 mux8_7.NAND4F_9.Y.n10 mux8_7.NAND4F_9.Y.n0 0.358709
R19268 MULT_0.4bit_ADDER_1.B1.n4 MULT_0.4bit_ADDER_1.B1.t16 491.64
R19269 MULT_0.4bit_ADDER_1.B1.n5 MULT_0.4bit_ADDER_1.B1.t20 491.64
R19270 MULT_0.4bit_ADDER_1.B1.n6 MULT_0.4bit_ADDER_1.B1.t19 491.64
R19271 MULT_0.4bit_ADDER_1.B1.n7 MULT_0.4bit_ADDER_1.B1.t12 491.64
R19272 MULT_0.4bit_ADDER_1.B1.n2 MULT_0.4bit_ADDER_1.B1.t13 485.221
R19273 MULT_0.4bit_ADDER_1.B1.n0 MULT_0.4bit_ADDER_1.B1.t15 367.928
R19274 MULT_0.4bit_ADDER_1.B1.n8 MULT_0.4bit_ADDER_1.B1.t17 255.588
R19275 MULT_0.4bit_ADDER_1.B1.n1 MULT_0.4bit_ADDER_1.B1.t22 224.478
R19276 MULT_0.4bit_ADDER_1.B1.n0 MULT_0.4bit_ADDER_1.B1.t18 213.688
R19277 MULT_0.4bit_ADDER_1.B1.n4 MULT_0.4bit_ADDER_1.B1.n3 209.19
R19278 MULT_0.4bit_ADDER_1.B1.n3 MULT_0.4bit_ADDER_1.B1.t23 139.78
R19279 MULT_0.4bit_ADDER_1.B1.n3 MULT_0.4bit_ADDER_1.B1.t21 139.78
R19280 MULT_0.4bit_ADDER_1.B1.n3 MULT_0.4bit_ADDER_1.B1.t14 139.78
R19281 MULT_0.4bit_ADDER_1.B1.n12 MULT_0.4bit_ADDER_1.B1.n11 120.999
R19282 MULT_0.4bit_ADDER_1.B1.n12 MULT_0.4bit_ADDER_1.B1.n10 120.999
R19283 MULT_0.4bit_ADDER_1.B1.n24 MULT_0.4bit_ADDER_1.B1.n23 104.489
R19284 MULT_0.4bit_ADDER_1.B1.n9 MULT_0.4bit_ADDER_1.B1 103.258
R19285 MULT_0.4bit_ADDER_1.B1.n14 MULT_0.4bit_ADDER_1.B1.n13 92.5005
R19286 MULT_0.4bit_ADDER_1.B1.n21 MULT_0.4bit_ADDER_1.B1.n19 86.2638
R19287 MULT_0.4bit_ADDER_1.B1.n19 MULT_0.4bit_ADDER_1.B1.n18 85.8873
R19288 MULT_0.4bit_ADDER_1.B1.n19 MULT_0.4bit_ADDER_1.B1.n16 85.724
R19289 MULT_0.4bit_ADDER_1.B1.n2 MULT_0.4bit_ADDER_1.B1.n1 84.5046
R19290 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_1.B1.n24 83.8907
R19291 MULT_0.4bit_ADDER_1.B1.n22 MULT_0.4bit_ADDER_1.B1.n18 75.0672
R19292 MULT_0.4bit_ADDER_1.B1.n22 MULT_0.4bit_ADDER_1.B1.n21 75.0672
R19293 MULT_0.4bit_ADDER_1.B1.n16 MULT_0.4bit_ADDER_1.B1.n15 73.1255
R19294 MULT_0.4bit_ADDER_1.B1.n18 MULT_0.4bit_ADDER_1.B1.n17 73.1255
R19295 MULT_0.4bit_ADDER_1.B1.n21 MULT_0.4bit_ADDER_1.B1.n20 73.1255
R19296 MULT_0.4bit_ADDER_1.B1.n1 MULT_0.4bit_ADDER_1.B1.n0 72.3005
R19297 MULT_0.4bit_ADDER_1.B1.n23 MULT_0.4bit_ADDER_1.B1.n16 68.8946
R19298 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_1.B1.n2 60.9816
R19299 MULT_0.4bit_ADDER_1.B1.n24 MULT_0.4bit_ADDER_1.B1.n14 41.9827
R19300 MULT_0.4bit_ADDER_1.B1.n13 MULT_0.4bit_ADDER_1.B1.t2 30.462
R19301 MULT_0.4bit_ADDER_1.B1.n13 MULT_0.4bit_ADDER_1.B1.t8 30.462
R19302 MULT_0.4bit_ADDER_1.B1.n11 MULT_0.4bit_ADDER_1.B1.t7 30.462
R19303 MULT_0.4bit_ADDER_1.B1.n11 MULT_0.4bit_ADDER_1.B1.t6 30.462
R19304 MULT_0.4bit_ADDER_1.B1.n10 MULT_0.4bit_ADDER_1.B1.t0 30.462
R19305 MULT_0.4bit_ADDER_1.B1.n10 MULT_0.4bit_ADDER_1.B1.t1 30.462
R19306 MULT_0.4bit_ADDER_1.B1.n14 MULT_0.4bit_ADDER_1.B1.n12 28.124
R19307 MULT_0.4bit_ADDER_1.B1.n5 MULT_0.4bit_ADDER_1.B1.n4 17.8661
R19308 MULT_0.4bit_ADDER_1.B1.n6 MULT_0.4bit_ADDER_1.B1.n5 17.8661
R19309 MULT_0.4bit_ADDER_1.B1.n7 MULT_0.4bit_ADDER_1.B1.n6 17.1217
R19310 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_1.B1.n8 15.6329
R19311 MULT_0.4bit_ADDER_1.B1.n17 MULT_0.4bit_ADDER_1.B1.t10 11.8205
R19312 MULT_0.4bit_ADDER_1.B1.n17 MULT_0.4bit_ADDER_1.B1.t11 11.8205
R19313 MULT_0.4bit_ADDER_1.B1.n15 MULT_0.4bit_ADDER_1.B1.t9 11.8205
R19314 MULT_0.4bit_ADDER_1.B1.n15 MULT_0.4bit_ADDER_1.B1.t4 11.8205
R19315 MULT_0.4bit_ADDER_1.B1.n20 MULT_0.4bit_ADDER_1.B1.t3 11.8205
R19316 MULT_0.4bit_ADDER_1.B1.n20 MULT_0.4bit_ADDER_1.B1.t5 11.8205
R19317 MULT_0.4bit_ADDER_1.B1.n9 MULT_0.4bit_ADDER_1.B1 10.8165
R19318 MULT_0.4bit_ADDER_1.B1.n23 MULT_0.4bit_ADDER_1.B1.n22 9.3005
R19319 MULT_0.4bit_ADDER_1.B1.n8 MULT_0.4bit_ADDER_1.B1.n7 1.8615
R19320 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_1.B1.n9 0.838155
R19321 a_n12314_n26419.n7 a_n12314_n26419.n1 81.2978
R19322 a_n12314_n26419.n0 a_n12314_n26419.n3 81.1637
R19323 a_n12314_n26419.n0 a_n12314_n26419.n4 81.1637
R19324 a_n12314_n26419.n1 a_n12314_n26419.n5 81.1637
R19325 a_n12314_n26419.n1 a_n12314_n26419.n6 81.1637
R19326 a_n12314_n26419.n0 a_n12314_n26419.n2 80.9213
R19327 a_n12314_n26419.n2 a_n12314_n26419.t10 11.8205
R19328 a_n12314_n26419.n2 a_n12314_n26419.t11 11.8205
R19329 a_n12314_n26419.n3 a_n12314_n26419.t9 11.8205
R19330 a_n12314_n26419.n3 a_n12314_n26419.t0 11.8205
R19331 a_n12314_n26419.n4 a_n12314_n26419.t1 11.8205
R19332 a_n12314_n26419.n4 a_n12314_n26419.t2 11.8205
R19333 a_n12314_n26419.n5 a_n12314_n26419.t6 11.8205
R19334 a_n12314_n26419.n5 a_n12314_n26419.t8 11.8205
R19335 a_n12314_n26419.n6 a_n12314_n26419.t7 11.8205
R19336 a_n12314_n26419.n6 a_n12314_n26419.t4 11.8205
R19337 a_n12314_n26419.n7 a_n12314_n26419.t3 11.8205
R19338 a_n12314_n26419.t5 a_n12314_n26419.n7 11.8205
R19339 a_n12314_n26419.n1 a_n12314_n26419.n0 0.402735
R19340 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n9 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t11 540.38
R19341 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t13 491.64
R19342 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t16 491.64
R19343 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t17 491.64
R19344 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t15 491.64
R19345 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n7 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t12 367.928
R19346 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n1 227.526
R19347 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n8 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t7 227.356
R19348 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n3 227.266
R19349 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n2 227.266
R19350 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n7 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t8 213.688
R19351 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n6 162.852
R19352 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n9 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n8 160.439
R19353 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t14 139.78
R19354 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t9 139.78
R19355 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t18 139.78
R19356 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t10 139.78
R19357 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n8 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n7 94.4341
R19358 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t0 42.7831
R19359 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n6 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n5 38.6833
R19360 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n3 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t2 30.379
R19361 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n3 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t3 30.379
R19362 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n1 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t6 30.379
R19363 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n1 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t4 30.379
R19364 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n2 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t1 30.379
R19365 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n2 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t5 30.379
R19366 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n6 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n4 28.3986
R19367 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n0 18.8832
R19368 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n10 11.2587
R19369 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n10 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 5.09176
R19370 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n10 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 4.19292
R19371 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n9 0.794268
R19372 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t8 485.221
R19373 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t10 367.928
R19374 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n5 227.526
R19375 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n6 227.266
R19376 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n4 227.266
R19377 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t7 224.478
R19378 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t9 213.688
R19379 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n2 84.5046
R19380 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n1 72.3005
R19381 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n3 61.0566
R19382 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t3 42.7747
R19383 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t6 30.379
R19384 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t0 30.379
R19385 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t4 30.379
R19386 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t5 30.379
R19387 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t1 30.379
R19388 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.t2 30.379
R19389 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A.n0 0.583137
R19390 a_9528_n8194.t0 a_9528_n8194.t1 9.9005
R19391 AND8_0.NOT8_0.A0.n2 AND8_0.NOT8_0.A0.t8 394.37
R19392 AND8_0.NOT8_0.A0.n1 AND8_0.NOT8_0.A0.t7 291.829
R19393 AND8_0.NOT8_0.A0.n1 AND8_0.NOT8_0.A0.t9 291.829
R19394 AND8_0.NOT8_0.A0.n0 AND8_0.NOT8_0.A0.n4 227.526
R19395 AND8_0.NOT8_0.A0.n0 AND8_0.NOT8_0.A0.n3 227.266
R19396 AND8_0.NOT8_0.A0.n0 AND8_0.NOT8_0.A0.n5 227.266
R19397 AND8_0.NOT8_0.A0.n1 AND8_0.NOT8_0.A0.t10 221.72
R19398 AND8_0.NOT8_0.A0.n2 AND8_0.NOT8_0.A0.n1 53.374
R19399 AND8_0.NOT8_0.A0.n0 AND8_0.NOT8_0.A0.t4 42.7873
R19400 AND8_0.NOT8_0.A0.n4 AND8_0.NOT8_0.A0.t1 30.379
R19401 AND8_0.NOT8_0.A0.n4 AND8_0.NOT8_0.A0.t0 30.379
R19402 AND8_0.NOT8_0.A0.n3 AND8_0.NOT8_0.A0.t5 30.379
R19403 AND8_0.NOT8_0.A0.n3 AND8_0.NOT8_0.A0.t6 30.379
R19404 AND8_0.NOT8_0.A0.n5 AND8_0.NOT8_0.A0.t3 30.379
R19405 AND8_0.NOT8_0.A0.n5 AND8_0.NOT8_0.A0.t2 30.379
R19406 AND8_0.NOT8_0.A0 AND8_0.NOT8_0.A0.n0 2.10064
R19407 AND8_0.NOT8_0.A0 AND8_0.NOT8_0.A0.n2 1.27931
R19408 AND8_0.S0.n1 AND8_0.S0.t6 1032.02
R19409 AND8_0.S0.n1 AND8_0.S0.t5 336.962
R19410 AND8_0.S0.n1 AND8_0.S0.t4 326.154
R19411 AND8_0.S0.n0 AND8_0.S0.t3 256.514
R19412 AND8_0.S0.n0 AND8_0.S0.n2 226.258
R19413 AND8_0.S0 AND8_0.S0.n1 162.945
R19414 AND8_0.S0.n0 AND8_0.S0.t0 83.7172
R19415 AND8_0.S0.n2 AND8_0.S0.t1 30.379
R19416 AND8_0.S0.n2 AND8_0.S0.t2 30.379
R19417 AND8_0.S0 AND8_0.S0.n0 1.93382
R19418 a_n209_1406.n0 a_n209_1406.t7 539.788
R19419 a_n209_1406.n1 a_n209_1406.t4 531.496
R19420 a_n209_1406.n0 a_n209_1406.t3 490.034
R19421 a_n209_1406.n5 a_n209_1406.t0 283.788
R19422 a_n209_1406.t1 a_n209_1406.n5 205.489
R19423 a_n209_1406.n2 a_n209_1406.t5 182.625
R19424 a_n209_1406.n3 a_n209_1406.t2 179.054
R19425 a_n209_1406.n2 a_n209_1406.t6 139.78
R19426 a_n209_1406.n4 a_n209_1406.n3 101.368
R19427 a_n209_1406.n5 a_n209_1406.n4 77.9135
R19428 a_n209_1406.n4 a_n209_1406.n1 76.1557
R19429 a_n209_1406.n1 a_n209_1406.n0 8.29297
R19430 a_n209_1406.n3 a_n209_1406.n2 3.57087
R19431 a_n29_1406.n2 a_n29_1406.n0 121.353
R19432 a_n29_1406.n2 a_n29_1406.n1 121.001
R19433 a_n29_1406.n3 a_n29_1406.n2 120.977
R19434 a_n29_1406.n0 a_n29_1406.t5 30.462
R19435 a_n29_1406.n0 a_n29_1406.t4 30.462
R19436 a_n29_1406.n1 a_n29_1406.t2 30.462
R19437 a_n29_1406.n1 a_n29_1406.t3 30.462
R19438 a_n29_1406.n3 a_n29_1406.t1 30.462
R19439 a_n29_1406.t0 a_n29_1406.n3 30.462
R19440 8bit_ADDER_0.S0.n0 8bit_ADDER_0.S0.t13 1032.02
R19441 8bit_ADDER_0.S0.n0 8bit_ADDER_0.S0.t14 336.962
R19442 8bit_ADDER_0.S0.n0 8bit_ADDER_0.S0.t12 326.154
R19443 8bit_ADDER_0.S0 8bit_ADDER_0.S0.n0 162.952
R19444 8bit_ADDER_0.S0.n3 8bit_ADDER_0.S0.n2 120.999
R19445 8bit_ADDER_0.S0.n3 8bit_ADDER_0.S0.n1 120.999
R19446 8bit_ADDER_0.S0.n15 8bit_ADDER_0.S0.n14 104.489
R19447 8bit_ADDER_0.S0.n5 8bit_ADDER_0.S0.n4 92.5005
R19448 8bit_ADDER_0.S0.n12 8bit_ADDER_0.S0.n10 86.2638
R19449 8bit_ADDER_0.S0.n10 8bit_ADDER_0.S0.n9 85.8873
R19450 8bit_ADDER_0.S0.n10 8bit_ADDER_0.S0.n7 85.724
R19451 8bit_ADDER_0.S0 8bit_ADDER_0.S0.n15 83.8907
R19452 8bit_ADDER_0.S0.n13 8bit_ADDER_0.S0.n12 75.0672
R19453 8bit_ADDER_0.S0.n13 8bit_ADDER_0.S0.n9 75.0672
R19454 8bit_ADDER_0.S0.n12 8bit_ADDER_0.S0.n11 73.1255
R19455 8bit_ADDER_0.S0.n9 8bit_ADDER_0.S0.n8 73.1255
R19456 8bit_ADDER_0.S0.n7 8bit_ADDER_0.S0.n6 73.1255
R19457 8bit_ADDER_0.S0.n14 8bit_ADDER_0.S0.n7 68.8946
R19458 8bit_ADDER_0.S0.n15 8bit_ADDER_0.S0.n5 41.9827
R19459 8bit_ADDER_0.S0.n4 8bit_ADDER_0.S0.t10 30.462
R19460 8bit_ADDER_0.S0.n4 8bit_ADDER_0.S0.t1 30.462
R19461 8bit_ADDER_0.S0.n2 8bit_ADDER_0.S0.t0 30.462
R19462 8bit_ADDER_0.S0.n2 8bit_ADDER_0.S0.t2 30.462
R19463 8bit_ADDER_0.S0.n1 8bit_ADDER_0.S0.t9 30.462
R19464 8bit_ADDER_0.S0.n1 8bit_ADDER_0.S0.t8 30.462
R19465 8bit_ADDER_0.S0.n5 8bit_ADDER_0.S0.n3 28.124
R19466 8bit_ADDER_0.S0.n8 8bit_ADDER_0.S0.t7 11.8205
R19467 8bit_ADDER_0.S0.n8 8bit_ADDER_0.S0.t6 11.8205
R19468 8bit_ADDER_0.S0.n11 8bit_ADDER_0.S0.t5 11.8205
R19469 8bit_ADDER_0.S0.n11 8bit_ADDER_0.S0.t4 11.8205
R19470 8bit_ADDER_0.S0.n6 8bit_ADDER_0.S0.t11 11.8205
R19471 8bit_ADDER_0.S0.n6 8bit_ADDER_0.S0.t3 11.8205
R19472 8bit_ADDER_0.S0.n14 8bit_ADDER_0.S0.n13 9.3005
R19473 left_shifter_0.buffer_6.inv_1.A.n0 left_shifter_0.buffer_6.inv_1.A.t5 393.921
R19474 left_shifter_0.buffer_6.inv_1.A.n2 left_shifter_0.buffer_6.inv_1.A.t6 291.829
R19475 left_shifter_0.buffer_6.inv_1.A.n2 left_shifter_0.buffer_6.inv_1.A.t4 291.829
R19476 left_shifter_0.buffer_6.inv_1.A.n0 left_shifter_0.buffer_6.inv_1.A.t1 256.89
R19477 left_shifter_0.buffer_6.inv_1.A.n0 left_shifter_0.buffer_6.inv_1.A.n1 226.538
R19478 left_shifter_0.buffer_6.inv_1.A.n2 left_shifter_0.buffer_6.inv_1.A.t7 221.72
R19479 left_shifter_0.buffer_6.inv_1.A.n0 left_shifter_0.buffer_6.inv_1.A.t0 83.795
R19480 left_shifter_0.buffer_6.inv_1.A.n0 left_shifter_0.buffer_6.inv_1.A.n2 53.7938
R19481 left_shifter_0.buffer_6.inv_1.A.n1 left_shifter_0.buffer_6.inv_1.A.t2 30.379
R19482 left_shifter_0.buffer_6.inv_1.A.n1 left_shifter_0.buffer_6.inv_1.A.t3 30.379
R19483 left_shifter_0.S1.n1 left_shifter_0.S1.t5 1032.02
R19484 left_shifter_0.S1.n1 left_shifter_0.S1.t4 336.962
R19485 left_shifter_0.S1.n1 left_shifter_0.S1.t6 326.154
R19486 left_shifter_0.S1.n0 left_shifter_0.S1.t3 256.89
R19487 left_shifter_0.S1.n0 left_shifter_0.S1.n2 226.635
R19488 mux8_2.NAND4F_5.A left_shifter_0.S1.n1 162.952
R19489 left_shifter_0.S1.n0 left_shifter_0.S1.t0 83.7172
R19490 mux8_2.A6 left_shifter_0.S1.n0 51.9196
R19491 left_shifter_0.S1.n2 left_shifter_0.S1.t1 30.379
R19492 left_shifter_0.S1.n2 left_shifter_0.S1.t2 30.379
R19493 mux8_2.A6 mux8_2.NAND4F_5.A 11.8717
R19494 mux8_0.NAND4F_0.Y.n1 mux8_0.NAND4F_0.Y.t11 1388.16
R19495 mux8_0.NAND4F_0.Y.n1 mux8_0.NAND4F_0.Y.t9 350.839
R19496 mux8_0.NAND4F_0.Y.n2 mux8_0.NAND4F_0.Y.t10 308.481
R19497 mux8_0.NAND4F_0.Y.n0 mux8_0.NAND4F_0.Y.n3 187.373
R19498 mux8_0.NAND4F_0.Y.n0 mux8_0.NAND4F_0.Y.n4 187.192
R19499 mux8_0.NAND4F_0.Y.n0 mux8_0.NAND4F_0.Y.n5 187.192
R19500 mux8_0.NAND4F_0.Y mux8_0.NAND4F_0.Y.n6 187.192
R19501 mux8_0.NAND4F_0.Y mux8_0.NAND4F_0.Y.n2 161.492
R19502 mux8_0.NAND4F_0.Y.n2 mux8_0.NAND4F_0.Y.n1 27.752
R19503 mux8_0.NAND4F_0.Y mux8_0.NAND4F_0.Y.t2 23.5085
R19504 mux8_0.NAND4F_0.Y.n3 mux8_0.NAND4F_0.Y.t5 20.1899
R19505 mux8_0.NAND4F_0.Y.n3 mux8_0.NAND4F_0.Y.t6 20.1899
R19506 mux8_0.NAND4F_0.Y.n4 mux8_0.NAND4F_0.Y.t1 20.1899
R19507 mux8_0.NAND4F_0.Y.n4 mux8_0.NAND4F_0.Y.t0 20.1899
R19508 mux8_0.NAND4F_0.Y.n5 mux8_0.NAND4F_0.Y.t8 20.1899
R19509 mux8_0.NAND4F_0.Y.n5 mux8_0.NAND4F_0.Y.t7 20.1899
R19510 mux8_0.NAND4F_0.Y.n6 mux8_0.NAND4F_0.Y.t4 20.1899
R19511 mux8_0.NAND4F_0.Y.n6 mux8_0.NAND4F_0.Y.t3 20.1899
R19512 mux8_0.NAND4F_0.Y mux8_0.NAND4F_0.Y.n0 0.358709
R19513 MULT_0.NAND2_5.Y.n5 MULT_0.NAND2_5.Y.t10 291.829
R19514 MULT_0.NAND2_5.Y.n5 MULT_0.NAND2_5.Y.t8 291.829
R19515 MULT_0.NAND2_5.Y.n0 MULT_0.NAND2_5.Y.n3 227.526
R19516 MULT_0.NAND2_5.Y.n0 MULT_0.NAND2_5.Y.n2 227.266
R19517 MULT_0.NAND2_5.Y.n0 MULT_0.NAND2_5.Y.n4 227.266
R19518 MULT_0.NAND2_5.Y.n5 MULT_0.NAND2_5.Y.t7 221.72
R19519 MULT_0.NAND2_5.Y.t9 MULT_0.NAND2_5.Y.n1 393.897
R19520 MULT_0.NAND2_5.Y.n0 MULT_0.NAND2_5.Y.t3 42.7333
R19521 MULT_0.NAND2_5.Y.n3 MULT_0.NAND2_5.Y.t1 30.379
R19522 MULT_0.NAND2_5.Y.n3 MULT_0.NAND2_5.Y.t0 30.379
R19523 MULT_0.NAND2_5.Y.n2 MULT_0.NAND2_5.Y.t6 30.379
R19524 MULT_0.NAND2_5.Y.n2 MULT_0.NAND2_5.Y.t4 30.379
R19525 MULT_0.NAND2_5.Y.n4 MULT_0.NAND2_5.Y.t5 30.379
R19526 MULT_0.NAND2_5.Y.n4 MULT_0.NAND2_5.Y.t2 30.379
R19527 MULT_0.NAND2_5.Y.n5 MULT_0.NAND2_5.Y.n1 53.4912
R19528 MULT_0.NAND2_5.Y.n0 MULT_0.NAND2_5.Y.n1 0.621379
R19529 MULT_0.4bit_ADDER_0.A1.n3 MULT_0.4bit_ADDER_0.A1.t12 540.38
R19530 MULT_0.4bit_ADDER_0.A1.n4 MULT_0.4bit_ADDER_0.A1.t11 491.64
R19531 MULT_0.4bit_ADDER_0.A1.n4 MULT_0.4bit_ADDER_0.A1.t13 491.64
R19532 MULT_0.4bit_ADDER_0.A1.n4 MULT_0.4bit_ADDER_0.A1.t10 491.64
R19533 MULT_0.4bit_ADDER_0.A1.n4 MULT_0.4bit_ADDER_0.A1.t6 491.64
R19534 MULT_0.4bit_ADDER_0.A1.n1 MULT_0.4bit_ADDER_0.A1.t14 367.928
R19535 MULT_0.4bit_ADDER_0.A1.n0 MULT_0.4bit_ADDER_0.A1.t2 256.514
R19536 MULT_0.4bit_ADDER_0.A1.n2 MULT_0.4bit_ADDER_0.A1.t5 227.356
R19537 MULT_0.4bit_ADDER_0.A1.n0 MULT_0.4bit_ADDER_0.A1.n8 226.136
R19538 MULT_0.4bit_ADDER_0.A1.n1 MULT_0.4bit_ADDER_0.A1.t4 213.688
R19539 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_0.B MULT_0.4bit_ADDER_0.A1.n6 162.867
R19540 MULT_0.4bit_ADDER_0.A1.n3 MULT_0.4bit_ADDER_0.A1.n2 160.439
R19541 MULT_0.4bit_ADDER_0.A1.n5 MULT_0.4bit_ADDER_0.A1.t7 139.78
R19542 MULT_0.4bit_ADDER_0.A1.n5 MULT_0.4bit_ADDER_0.A1.t15 139.78
R19543 MULT_0.4bit_ADDER_0.A1.n5 MULT_0.4bit_ADDER_0.A1.t8 139.78
R19544 MULT_0.4bit_ADDER_0.A1.n5 MULT_0.4bit_ADDER_0.A1.t9 139.78
R19545 MULT_0.4bit_ADDER_0.A1.n2 MULT_0.4bit_ADDER_0.A1.n1 94.4341
R19546 MULT_0.4bit_ADDER_0.A1.n0 MULT_0.4bit_ADDER_0.A1.t0 83.8129
R19547 MULT_0.4bit_ADDER_0.A1.n6 MULT_0.4bit_ADDER_0.A1.n5 38.6833
R19548 MULT_0.4bit_ADDER_0.A1.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.A 34.387
R19549 MULT_0.4bit_ADDER_0.A1.n8 MULT_0.4bit_ADDER_0.A1.t1 30.379
R19550 MULT_0.4bit_ADDER_0.A1.n8 MULT_0.4bit_ADDER_0.A1.t3 30.379
R19551 MULT_0.4bit_ADDER_0.A1.n6 MULT_0.4bit_ADDER_0.A1.n4 28.3986
R19552 MULT_0.4bit_ADDER_0.FULL_ADDER_2.A MULT_0.4bit_ADDER_0.A1.n7 16.8032
R19553 MULT_0.4bit_ADDER_0.A1.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_0.B 9.00496
R19554 MULT_0.4bit_ADDER_0.A1.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_0.B 3.87912
R19555 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_0.B MULT_0.4bit_ADDER_0.A1.n3 0.89693
R19556 mux8_5.A1.n0 mux8_5.A1.t13 1032.02
R19557 mux8_5.A1.n0 mux8_5.A1.t14 336.962
R19558 mux8_5.A1.n0 mux8_5.A1.t12 326.154
R19559 mux8_5.A1 mux8_5.A1.n0 162.952
R19560 mux8_5.A1.n3 mux8_5.A1.n2 120.999
R19561 mux8_5.A1.n3 mux8_5.A1.n1 120.999
R19562 mux8_5.A1.n15 mux8_5.A1.n14 104.489
R19563 mux8_5.A1.n5 mux8_5.A1.n4 92.5005
R19564 mux8_5.A1.n12 mux8_5.A1.n10 86.2638
R19565 mux8_5.A1.n10 mux8_5.A1.n9 85.8873
R19566 mux8_5.A1.n10 mux8_5.A1.n7 85.724
R19567 mux8_5.A1 mux8_5.A1.n15 83.8907
R19568 mux8_5.A1.n13 mux8_5.A1.n12 75.0672
R19569 mux8_5.A1.n13 mux8_5.A1.n9 75.0672
R19570 mux8_5.A1.n12 mux8_5.A1.n11 73.1255
R19571 mux8_5.A1.n7 mux8_5.A1.n6 73.1255
R19572 mux8_5.A1.n9 mux8_5.A1.n8 73.1255
R19573 mux8_5.A1.n14 mux8_5.A1.n7 68.8946
R19574 mux8_5.A1.n15 mux8_5.A1.n5 41.9827
R19575 mux8_5.A1.n4 mux8_5.A1.t5 30.462
R19576 mux8_5.A1.n4 mux8_5.A1.t7 30.462
R19577 mux8_5.A1.n2 mux8_5.A1.t10 30.462
R19578 mux8_5.A1.n2 mux8_5.A1.t6 30.462
R19579 mux8_5.A1.n1 mux8_5.A1.t3 30.462
R19580 mux8_5.A1.n1 mux8_5.A1.t4 30.462
R19581 mux8_5.A1.n5 mux8_5.A1.n3 28.124
R19582 mux8_5.A1.n6 mux8_5.A1.t2 11.8205
R19583 mux8_5.A1.n6 mux8_5.A1.t9 11.8205
R19584 mux8_5.A1.n11 mux8_5.A1.t11 11.8205
R19585 mux8_5.A1.n11 mux8_5.A1.t8 11.8205
R19586 mux8_5.A1.n8 mux8_5.A1.t0 11.8205
R19587 mux8_5.A1.n8 mux8_5.A1.t1 11.8205
R19588 mux8_5.A1.n14 mux8_5.A1.n13 9.3005
R19589 mux8_5.NAND4F_0.Y.n1 mux8_5.NAND4F_0.Y.t11 1388.16
R19590 mux8_5.NAND4F_0.Y.n1 mux8_5.NAND4F_0.Y.t10 350.839
R19591 mux8_5.NAND4F_0.Y.n2 mux8_5.NAND4F_0.Y.t9 308.481
R19592 mux8_5.NAND4F_0.Y.n0 mux8_5.NAND4F_0.Y.n3 187.373
R19593 mux8_5.NAND4F_0.Y.n0 mux8_5.NAND4F_0.Y.n4 187.192
R19594 mux8_5.NAND4F_0.Y.n0 mux8_5.NAND4F_0.Y.n5 187.192
R19595 mux8_5.NAND4F_0.Y mux8_5.NAND4F_0.Y.n6 187.192
R19596 mux8_5.NAND4F_0.Y mux8_5.NAND4F_0.Y.n2 161.492
R19597 mux8_5.NAND4F_0.Y.n2 mux8_5.NAND4F_0.Y.n1 27.752
R19598 mux8_5.NAND4F_0.Y mux8_5.NAND4F_0.Y.t4 23.5085
R19599 mux8_5.NAND4F_0.Y.n3 mux8_5.NAND4F_0.Y.t5 20.1899
R19600 mux8_5.NAND4F_0.Y.n3 mux8_5.NAND4F_0.Y.t6 20.1899
R19601 mux8_5.NAND4F_0.Y.n4 mux8_5.NAND4F_0.Y.t1 20.1899
R19602 mux8_5.NAND4F_0.Y.n4 mux8_5.NAND4F_0.Y.t0 20.1899
R19603 mux8_5.NAND4F_0.Y.n5 mux8_5.NAND4F_0.Y.t8 20.1899
R19604 mux8_5.NAND4F_0.Y.n5 mux8_5.NAND4F_0.Y.t7 20.1899
R19605 mux8_5.NAND4F_0.Y.n6 mux8_5.NAND4F_0.Y.t2 20.1899
R19606 mux8_5.NAND4F_0.Y.n6 mux8_5.NAND4F_0.Y.t3 20.1899
R19607 mux8_5.NAND4F_0.Y mux8_5.NAND4F_0.Y.n0 0.358709
R19608 a_n14490_373.t0 a_n14490_373.t1 19.8005
R19609 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t8 485.221
R19610 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t9 367.928
R19611 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n5 227.526
R19612 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n6 227.266
R19613 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n4 227.266
R19614 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t10 224.478
R19615 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t7 213.688
R19616 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n2 84.5046
R19617 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n1 72.3005
R19618 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n3 61.0566
R19619 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t4 42.7747
R19620 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t3 30.379
R19621 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t1 30.379
R19622 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t6 30.379
R19623 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t5 30.379
R19624 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t2 30.379
R19625 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.t0 30.379
R19626 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A.n0 0.583137
R19627 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t10 540.38
R19628 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t7 491.64
R19629 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t14 491.64
R19630 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t15 491.64
R19631 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t8 491.64
R19632 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t11 367.928
R19633 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n2 227.526
R19634 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t17 227.356
R19635 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n1 227.266
R19636 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n3 227.266
R19637 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n7 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t9 213.688
R19638 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n6 162.852
R19639 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n8 160.439
R19640 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t13 139.78
R19641 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t18 139.78
R19642 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t16 139.78
R19643 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t12 139.78
R19644 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n7 94.4341
R19645 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t0 42.7831
R19646 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n5 38.6833
R19647 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t6 30.379
R19648 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t4 30.379
R19649 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t1 30.379
R19650 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t2 30.379
R19651 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t3 30.379
R19652 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t5 30.379
R19653 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n4 28.3986
R19654 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n0 18.8832
R19655 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n10 10.7052
R19656 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT 5.09176
R19657 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT 4.19292
R19658 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n9 0.794268
R19659 a_n18042_1406.n3 a_n18042_1406.n2 121.353
R19660 a_n18042_1406.n2 a_n18042_1406.n1 121.001
R19661 a_n18042_1406.n2 a_n18042_1406.n0 120.977
R19662 a_n18042_1406.n1 a_n18042_1406.t4 30.462
R19663 a_n18042_1406.n1 a_n18042_1406.t1 30.462
R19664 a_n18042_1406.n0 a_n18042_1406.t5 30.462
R19665 a_n18042_1406.n0 a_n18042_1406.t3 30.462
R19666 a_n18042_1406.n3 a_n18042_1406.t0 30.462
R19667 a_n18042_1406.t2 a_n18042_1406.n3 30.462
R19668 mux8_0.NAND4F_2.Y.n6 mux8_0.NAND4F_2.Y.t10 933.563
R19669 mux8_0.NAND4F_2.Y.n6 mux8_0.NAND4F_2.Y.t11 367.635
R19670 mux8_0.NAND4F_2.Y.n7 mux8_0.NAND4F_2.Y.t9 308.481
R19671 mux8_0.NAND4F_2.Y.n0 mux8_0.NAND4F_2.Y.n1 187.373
R19672 mux8_0.NAND4F_2.Y.n0 mux8_0.NAND4F_2.Y.n2 187.192
R19673 mux8_0.NAND4F_2.Y.n0 mux8_0.NAND4F_2.Y.n3 187.192
R19674 mux8_0.NAND4F_2.Y.n5 mux8_0.NAND4F_2.Y.n4 187.192
R19675 mux8_0.NAND4F_2.Y mux8_0.NAND4F_2.Y.n7 162.102
R19676 mux8_0.NAND4F_2.Y.n8 mux8_0.NAND4F_2.Y.t0 22.7096
R19677 mux8_0.NAND4F_2.Y.n8 mux8_0.NAND4F_2.Y 22.4285
R19678 mux8_0.NAND4F_2.Y.n1 mux8_0.NAND4F_2.Y.t5 20.1899
R19679 mux8_0.NAND4F_2.Y.n1 mux8_0.NAND4F_2.Y.t6 20.1899
R19680 mux8_0.NAND4F_2.Y.n2 mux8_0.NAND4F_2.Y.t4 20.1899
R19681 mux8_0.NAND4F_2.Y.n2 mux8_0.NAND4F_2.Y.t3 20.1899
R19682 mux8_0.NAND4F_2.Y.n3 mux8_0.NAND4F_2.Y.t8 20.1899
R19683 mux8_0.NAND4F_2.Y.n3 mux8_0.NAND4F_2.Y.t7 20.1899
R19684 mux8_0.NAND4F_2.Y.n4 mux8_0.NAND4F_2.Y.t1 20.1899
R19685 mux8_0.NAND4F_2.Y.n4 mux8_0.NAND4F_2.Y.t2 20.1899
R19686 mux8_0.NAND4F_2.Y.n7 mux8_0.NAND4F_2.Y.n6 10.955
R19687 mux8_0.NAND4F_2.Y mux8_0.NAND4F_2.Y.n8 0.799394
R19688 mux8_0.NAND4F_2.Y mux8_0.NAND4F_2.Y.n5 0.452586
R19689 mux8_0.NAND4F_2.Y.n5 mux8_0.NAND4F_2.Y.n0 0.358709
R19690 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n9 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t9 540.38
R19691 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t16 491.64
R19692 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t11 491.64
R19693 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t12 491.64
R19694 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t8 491.64
R19695 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n7 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t13 367.928
R19696 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n1 227.526
R19697 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n8 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t14 227.356
R19698 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n3 227.266
R19699 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n2 227.266
R19700 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n7 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t15 213.688
R19701 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n6 162.852
R19702 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n9 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n8 160.439
R19703 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t7 139.78
R19704 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t17 139.78
R19705 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t10 139.78
R19706 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t18 139.78
R19707 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n8 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n7 94.4341
R19708 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t0 42.7831
R19709 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n6 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n5 38.6833
R19710 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n3 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t3 30.379
R19711 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n3 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t2 30.379
R19712 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n1 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t5 30.379
R19713 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n1 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t4 30.379
R19714 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n2 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t1 30.379
R19715 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n2 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t6 30.379
R19716 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n6 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n4 28.3986
R19717 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n0 18.8832
R19718 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n10 11.2574
R19719 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n10 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 5.09176
R19720 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n10 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 4.19292
R19721 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n9 0.794268
R19722 a_n9325_1406.n2 a_n9325_1406.n0 121.353
R19723 a_n9325_1406.n3 a_n9325_1406.n2 121.353
R19724 a_n9325_1406.n2 a_n9325_1406.n1 121.001
R19725 a_n9325_1406.n0 a_n9325_1406.t5 30.462
R19726 a_n9325_1406.n0 a_n9325_1406.t3 30.462
R19727 a_n9325_1406.n1 a_n9325_1406.t0 30.462
R19728 a_n9325_1406.n1 a_n9325_1406.t4 30.462
R19729 a_n9325_1406.n3 a_n9325_1406.t1 30.462
R19730 a_n9325_1406.t2 a_n9325_1406.n3 30.462
R19731 Y1.n0 Y1.t4 883.668
R19732 Y1.n1 Y1.t6 740.381
R19733 Y1.n0 Y1.t5 729.428
R19734 Y1.n2 Y1.t7 700.508
R19735 Y1.n4 Y1.t0 256.514
R19736 Y1.n5 Y1.n3 226.251
R19737 Y1 Y1.n2 162.986
R19738 Y1.n4 Y1.t1 83.7599
R19739 Y1.n1 Y1.n0 72.3005
R19740 Y1.n3 Y1.t2 30.379
R19741 Y1.n3 Y1.t3 30.379
R19742 Y1.n2 Y1.n1 16.7975
R19743 Y1.n5 Y1 0.0415053
R19744 Y1.n5 Y1.n4 0.0323878
R19745 Y1 Y1.n5 0.0126173
R19746 a_16143_n18523.n2 a_16143_n18523.n1 140.65
R19747 a_16143_n18523.n2 a_16143_n18523.n0 140.65
R19748 a_16143_n18523.n3 a_16143_n18523.n2 140.587
R19749 a_16143_n18523.n1 a_16143_n18523.t4 7.59513
R19750 a_16143_n18523.n1 a_16143_n18523.t5 7.59513
R19751 a_16143_n18523.n0 a_16143_n18523.t2 7.59513
R19752 a_16143_n18523.n0 a_16143_n18523.t1 7.59513
R19753 a_16143_n18523.t0 a_16143_n18523.n3 7.59513
R19754 a_16143_n18523.n3 a_16143_n18523.t3 7.59513
R19755 a_16431_n18523.n2 a_16431_n18523.n0 140.274
R19756 a_16431_n18523.n3 a_16431_n18523.n2 140.274
R19757 a_16431_n18523.n2 a_16431_n18523.n1 140.21
R19758 a_16431_n18523.n1 a_16431_n18523.t2 7.59513
R19759 a_16431_n18523.n1 a_16431_n18523.t5 7.59513
R19760 a_16431_n18523.n0 a_16431_n18523.t0 7.59513
R19761 a_16431_n18523.n0 a_16431_n18523.t1 7.59513
R19762 a_16431_n18523.t4 a_16431_n18523.n3 7.59513
R19763 a_16431_n18523.n3 a_16431_n18523.t3 7.59513
R19764 mux8_8.NAND4F_9.Y.n1 mux8_8.NAND4F_9.Y.t9 312.599
R19765 mux8_8.NAND4F_9.Y.n4 mux8_8.NAND4F_9.Y.t14 247.428
R19766 mux8_8.NAND4F_9.Y.n1 mux8_8.NAND4F_9.Y.t10 247.428
R19767 mux8_8.NAND4F_9.Y.n2 mux8_8.NAND4F_9.Y.t11 247.428
R19768 mux8_8.NAND4F_9.Y.n3 mux8_8.NAND4F_9.Y.t13 247.428
R19769 mux8_8.NAND4F_9.Y.n5 mux8_8.NAND4F_9.Y.t12 229.754
R19770 mux8_8.NAND4F_9.Y.n0 mux8_8.NAND4F_9.Y.n6 187.373
R19771 mux8_8.NAND4F_9.Y.n0 mux8_8.NAND4F_9.Y.n7 187.192
R19772 mux8_8.NAND4F_9.Y.n0 mux8_8.NAND4F_9.Y.n8 187.192
R19773 mux8_8.NAND4F_9.Y.n10 mux8_8.NAND4F_9.Y.n9 187.192
R19774 mux8_8.NAND4F_9.Y mux8_8.NAND4F_9.Y.n5 162.275
R19775 mux8_8.NAND4F_9.Y.n5 mux8_8.NAND4F_9.Y.n4 91.5805
R19776 mux8_8.NAND4F_9.Y.n2 mux8_8.NAND4F_9.Y.n1 65.1723
R19777 mux8_8.NAND4F_9.Y.n3 mux8_8.NAND4F_9.Y.n2 65.1723
R19778 mux8_8.NAND4F_9.Y.n4 mux8_8.NAND4F_9.Y.n3 65.1723
R19779 mux8_8.NAND4F_9.Y mux8_8.NAND4F_9.Y.t0 22.6141
R19780 mux8_8.NAND4F_9.Y.n6 mux8_8.NAND4F_9.Y.t7 20.1899
R19781 mux8_8.NAND4F_9.Y.n6 mux8_8.NAND4F_9.Y.t8 20.1899
R19782 mux8_8.NAND4F_9.Y.n7 mux8_8.NAND4F_9.Y.t5 20.1899
R19783 mux8_8.NAND4F_9.Y.n7 mux8_8.NAND4F_9.Y.t6 20.1899
R19784 mux8_8.NAND4F_9.Y.n8 mux8_8.NAND4F_9.Y.t3 20.1899
R19785 mux8_8.NAND4F_9.Y.n8 mux8_8.NAND4F_9.Y.t4 20.1899
R19786 mux8_8.NAND4F_9.Y.n9 mux8_8.NAND4F_9.Y.t2 20.1899
R19787 mux8_8.NAND4F_9.Y.n9 mux8_8.NAND4F_9.Y.t1 20.1899
R19788 mux8_8.NAND4F_9.Y mux8_8.NAND4F_9.Y.n10 0.396904
R19789 mux8_8.NAND4F_9.Y.n10 mux8_8.NAND4F_9.Y.n0 0.358709
R19790 a_11865_n29943.n0 a_11865_n29943.n4 231.451
R19791 a_11865_n29943.n0 a_11865_n29943.n3 231.24
R19792 a_11865_n29943.n0 a_11865_n29943.n1 231.24
R19793 a_11865_n29943.n0 a_11865_n29943.n2 231.03
R19794 a_11865_n29943.n5 a_11865_n29943.n0 231.03
R19795 a_11865_n29943.n3 a_11865_n29943.t6 25.395
R19796 a_11865_n29943.n3 a_11865_n29943.t8 25.395
R19797 a_11865_n29943.n4 a_11865_n29943.t5 25.395
R19798 a_11865_n29943.n4 a_11865_n29943.t7 25.395
R19799 a_11865_n29943.n2 a_11865_n29943.t2 25.395
R19800 a_11865_n29943.n2 a_11865_n29943.t1 25.395
R19801 a_11865_n29943.n1 a_11865_n29943.t4 25.395
R19802 a_11865_n29943.n1 a_11865_n29943.t3 25.395
R19803 a_11865_n29943.t0 a_11865_n29943.n5 25.395
R19804 a_11865_n29943.n5 a_11865_n29943.t9 25.395
R19805 mux8_8.inv_0.A.n3 mux8_8.inv_0.A.t8 291.829
R19806 mux8_8.inv_0.A.n3 mux8_8.inv_0.A.t7 291.829
R19807 mux8_8.inv_0.A.n0 mux8_8.inv_0.A.t4 256.425
R19808 mux8_8.inv_0.A.n0 mux8_8.inv_0.A.n4 231.24
R19809 mux8_8.inv_0.A.n0 mux8_8.inv_0.A.n5 231.03
R19810 mux8_8.inv_0.A.n3 mux8_8.inv_0.A.t9 221.72
R19811 mux8_8.inv_0.A.t10 mux8_8.inv_0.A.n2 393.959
R19812 mux8_8.inv_0.A.n6 mux8_8.inv_0.A.n1 66.6316
R19813 mux8_8.inv_0.A.n2 mux8_8.inv_0.A.n3 53.4611
R19814 mux8_8.inv_0.A.n4 mux8_8.inv_0.A.t1 25.395
R19815 mux8_8.inv_0.A.n4 mux8_8.inv_0.A.t0 25.395
R19816 mux8_8.inv_0.A.n5 mux8_8.inv_0.A.t3 25.395
R19817 mux8_8.inv_0.A.n5 mux8_8.inv_0.A.t2 25.395
R19818 mux8_8.inv_0.A.n6 mux8_8.inv_0.A.t5 19.8005
R19819 mux8_8.inv_0.A.n6 mux8_8.inv_0.A.t6 19.8005
R19820 mux8_8.inv_0.A.n1 mux8_8.inv_0.A.n0 0.38953
R19821 mux8_8.inv_0.A.n1 mux8_8.inv_0.A.n2 0.294762
R19822 a_n17677_n21025.n0 a_n17677_n21025.n2 231.24
R19823 a_n17677_n21025.n1 a_n17677_n21025.n5 231.24
R19824 a_n17677_n21025.n0 a_n17677_n21025.n3 231.03
R19825 a_n17677_n21025.n1 a_n17677_n21025.n4 231.03
R19826 a_n17677_n21025.n6 a_n17677_n21025.n1 231.03
R19827 a_n17677_n21025.n2 a_n17677_n21025.t6 25.395
R19828 a_n17677_n21025.n2 a_n17677_n21025.t7 25.395
R19829 a_n17677_n21025.n3 a_n17677_n21025.t8 25.395
R19830 a_n17677_n21025.n3 a_n17677_n21025.t9 25.395
R19831 a_n17677_n21025.n4 a_n17677_n21025.t5 25.395
R19832 a_n17677_n21025.n4 a_n17677_n21025.t1 25.395
R19833 a_n17677_n21025.n5 a_n17677_n21025.t3 25.395
R19834 a_n17677_n21025.n5 a_n17677_n21025.t2 25.395
R19835 a_n17677_n21025.n6 a_n17677_n21025.t0 25.395
R19836 a_n17677_n21025.t4 a_n17677_n21025.n6 25.395
R19837 a_n17677_n21025.n1 a_n17677_n21025.n0 0.421553
R19838 a_n23245_1406.n0 a_n23245_1406.t5 539.788
R19839 a_n23245_1406.n1 a_n23245_1406.t6 531.496
R19840 a_n23245_1406.n0 a_n23245_1406.t3 490.034
R19841 a_n23245_1406.n5 a_n23245_1406.t0 283.788
R19842 a_n23245_1406.t1 a_n23245_1406.n5 205.489
R19843 a_n23245_1406.n2 a_n23245_1406.t2 182.625
R19844 a_n23245_1406.n3 a_n23245_1406.t4 179.054
R19845 a_n23245_1406.n2 a_n23245_1406.t7 139.78
R19846 a_n23245_1406.n4 a_n23245_1406.n3 101.368
R19847 a_n23245_1406.n5 a_n23245_1406.n4 77.9135
R19848 a_n23245_1406.n4 a_n23245_1406.n1 76.1557
R19849 a_n23245_1406.n1 a_n23245_1406.n0 8.29297
R19850 a_n23245_1406.n3 a_n23245_1406.n2 3.57087
R19851 a_7644_n8194.t0 a_7644_n8194.t1 9.9005
R19852 a_n19028_n11709.n2 a_n19028_n11709.t6 541.395
R19853 a_n19028_n11709.n3 a_n19028_n11709.t2 527.402
R19854 a_n19028_n11709.n2 a_n19028_n11709.t7 491.64
R19855 a_n19028_n11709.n5 a_n19028_n11709.t0 281.906
R19856 a_n19028_n11709.t1 a_n19028_n11709.n5 204.359
R19857 a_n19028_n11709.n0 a_n19028_n11709.t5 180.73
R19858 a_n19028_n11709.n1 a_n19028_n11709.t4 179.45
R19859 a_n19028_n11709.n0 a_n19028_n11709.t3 139.78
R19860 a_n19028_n11709.n4 a_n19028_n11709.n1 105.635
R19861 a_n19028_n11709.n4 a_n19028_n11709.n3 76.0005
R19862 a_n19028_n11709.n5 a_n19028_n11709.n4 67.9685
R19863 a_n19028_n11709.n3 a_n19028_n11709.n2 13.994
R19864 a_n19028_n11709.n1 a_n19028_n11709.n0 1.28015
R19865 mux8_8.A1.n0 mux8_8.A1.t14 1032.02
R19866 mux8_8.A1.n0 mux8_8.A1.t12 336.962
R19867 mux8_8.A1.n0 mux8_8.A1.t13 326.154
R19868 mux8_8.A1 mux8_8.A1.n0 162.952
R19869 mux8_8.A1.n3 mux8_8.A1.n2 120.999
R19870 mux8_8.A1.n3 mux8_8.A1.n1 120.999
R19871 mux8_8.A1.n15 mux8_8.A1.n14 104.489
R19872 mux8_8.A1.n5 mux8_8.A1.n4 92.5005
R19873 mux8_8.A1.n12 mux8_8.A1.n10 86.2638
R19874 mux8_8.A1.n10 mux8_8.A1.n9 85.8873
R19875 mux8_8.A1.n10 mux8_8.A1.n7 85.724
R19876 mux8_8.A1 mux8_8.A1.n15 83.8907
R19877 mux8_8.A1.n13 mux8_8.A1.n12 75.0672
R19878 mux8_8.A1.n13 mux8_8.A1.n9 75.0672
R19879 mux8_8.A1.n12 mux8_8.A1.n11 73.1255
R19880 mux8_8.A1.n7 mux8_8.A1.n6 73.1255
R19881 mux8_8.A1.n9 mux8_8.A1.n8 73.1255
R19882 mux8_8.A1.n14 mux8_8.A1.n7 68.8946
R19883 mux8_8.A1.n15 mux8_8.A1.n5 41.9827
R19884 mux8_8.A1.n4 mux8_8.A1.t4 30.462
R19885 mux8_8.A1.n4 mux8_8.A1.t0 30.462
R19886 mux8_8.A1.n2 mux8_8.A1.t11 30.462
R19887 mux8_8.A1.n2 mux8_8.A1.t3 30.462
R19888 mux8_8.A1.n1 mux8_8.A1.t5 30.462
R19889 mux8_8.A1.n1 mux8_8.A1.t6 30.462
R19890 mux8_8.A1.n5 mux8_8.A1.n3 28.124
R19891 mux8_8.A1.n6 mux8_8.A1.t8 11.8205
R19892 mux8_8.A1.n6 mux8_8.A1.t2 11.8205
R19893 mux8_8.A1.n11 mux8_8.A1.t1 11.8205
R19894 mux8_8.A1.n11 mux8_8.A1.t10 11.8205
R19895 mux8_8.A1.n8 mux8_8.A1.t9 11.8205
R19896 mux8_8.A1.n8 mux8_8.A1.t7 11.8205
R19897 mux8_8.A1.n14 mux8_8.A1.n13 9.3005
R19898 MULT_0.4bit_ADDER_1.B3.n5 MULT_0.4bit_ADDER_1.B3.t15 491.64
R19899 MULT_0.4bit_ADDER_1.B3.n6 MULT_0.4bit_ADDER_1.B3.t17 491.64
R19900 MULT_0.4bit_ADDER_1.B3.n7 MULT_0.4bit_ADDER_1.B3.t9 491.64
R19901 MULT_0.4bit_ADDER_1.B3.n8 MULT_0.4bit_ADDER_1.B3.t16 491.64
R19902 MULT_0.4bit_ADDER_1.B3.n3 MULT_0.4bit_ADDER_1.B3.t13 485.221
R19903 MULT_0.4bit_ADDER_1.B3.n1 MULT_0.4bit_ADDER_1.B3.t18 367.928
R19904 MULT_0.4bit_ADDER_1.B3.n9 MULT_0.4bit_ADDER_1.B3.t11 255.588
R19905 MULT_0.4bit_ADDER_1.B3.n0 MULT_0.4bit_ADDER_1.B3.n12 227.526
R19906 MULT_0.4bit_ADDER_1.B3.n0 MULT_0.4bit_ADDER_1.B3.n11 227.266
R19907 MULT_0.4bit_ADDER_1.B3.n0 MULT_0.4bit_ADDER_1.B3.n13 227.266
R19908 MULT_0.4bit_ADDER_1.B3.n2 MULT_0.4bit_ADDER_1.B3.t12 224.478
R19909 MULT_0.4bit_ADDER_1.B3.n1 MULT_0.4bit_ADDER_1.B3.t7 213.688
R19910 MULT_0.4bit_ADDER_1.B3.n5 MULT_0.4bit_ADDER_1.B3.n4 209.19
R19911 MULT_0.4bit_ADDER_1.B3.n4 MULT_0.4bit_ADDER_1.B3.t10 139.78
R19912 MULT_0.4bit_ADDER_1.B3.n4 MULT_0.4bit_ADDER_1.B3.t8 139.78
R19913 MULT_0.4bit_ADDER_1.B3.n4 MULT_0.4bit_ADDER_1.B3.t14 139.78
R19914 MULT_0.4bit_ADDER_1.B3.n10 MULT_0.4bit_ADDER_1.B3 103.258
R19915 MULT_0.4bit_ADDER_1.B3.n3 MULT_0.4bit_ADDER_1.B3.n2 84.5046
R19916 MULT_0.4bit_ADDER_1.B3.n2 MULT_0.4bit_ADDER_1.B3.n1 72.3005
R19917 MULT_0.4bit_ADDER_1.B3 MULT_0.4bit_ADDER_1.B3.n3 60.9816
R19918 MULT_0.4bit_ADDER_1.B3.n0 MULT_0.4bit_ADDER_1.B3.t3 42.7831
R19919 MULT_0.4bit_ADDER_1.B3.n12 MULT_0.4bit_ADDER_1.B3.t5 30.379
R19920 MULT_0.4bit_ADDER_1.B3.n12 MULT_0.4bit_ADDER_1.B3.t4 30.379
R19921 MULT_0.4bit_ADDER_1.B3.n11 MULT_0.4bit_ADDER_1.B3.t2 30.379
R19922 MULT_0.4bit_ADDER_1.B3.n11 MULT_0.4bit_ADDER_1.B3.t1 30.379
R19923 MULT_0.4bit_ADDER_1.B3.n13 MULT_0.4bit_ADDER_1.B3.t0 30.379
R19924 MULT_0.4bit_ADDER_1.B3.n13 MULT_0.4bit_ADDER_1.B3.t6 30.379
R19925 MULT_0.4bit_ADDER_1.B3 MULT_0.4bit_ADDER_1.B3.n0 18.8681
R19926 MULT_0.4bit_ADDER_1.B3.n6 MULT_0.4bit_ADDER_1.B3.n5 17.8661
R19927 MULT_0.4bit_ADDER_1.B3.n7 MULT_0.4bit_ADDER_1.B3.n6 17.8661
R19928 MULT_0.4bit_ADDER_1.B3.n8 MULT_0.4bit_ADDER_1.B3.n7 17.1217
R19929 MULT_0.4bit_ADDER_1.B3 MULT_0.4bit_ADDER_1.B3.n9 15.6329
R19930 MULT_0.4bit_ADDER_1.B3.n10 MULT_0.4bit_ADDER_1.B3 10.8165
R19931 MULT_0.4bit_ADDER_1.B3.n9 MULT_0.4bit_ADDER_1.B3.n8 1.8615
R19932 MULT_0.4bit_ADDER_1.B3 MULT_0.4bit_ADDER_1.B3.n10 0.862278
R19933 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t7 540.38
R19934 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t9 367.928
R19935 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n5 227.526
R19936 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t10 227.356
R19937 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n6 227.266
R19938 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n4 227.266
R19939 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t8 213.688
R19940 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n2 160.439
R19941 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n1 94.4341
R19942 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t3 42.7944
R19943 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t4 30.379
R19944 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t0 30.379
R19945 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t6 30.379
R19946 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t5 30.379
R19947 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t2 30.379
R19948 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.t1 30.379
R19949 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n0 13.4358
R19950 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B.n3 0.821842
R19951 mux8_7.inv_0.A.n1 mux8_7.inv_0.A.t8 291.829
R19952 mux8_7.inv_0.A.n1 mux8_7.inv_0.A.t10 291.829
R19953 mux8_7.inv_0.A.n0 mux8_7.inv_0.A.t3 256.425
R19954 mux8_7.inv_0.A.n0 mux8_7.inv_0.A.n2 231.24
R19955 mux8_7.inv_0.A.n0 mux8_7.inv_0.A.n3 231.03
R19956 mux8_7.inv_0.A.n1 mux8_7.inv_0.A.t9 221.72
R19957 mux8_7.inv_0.A.t7 mux8_7.inv_0.A.n0 393.959
R19958 mux8_7.inv_0.A.n4 mux8_7.inv_0.A.n0 66.6316
R19959 mux8_7.inv_0.A.n0 mux8_7.inv_0.A.n1 54.1444
R19960 mux8_7.inv_0.A.n2 mux8_7.inv_0.A.t5 25.395
R19961 mux8_7.inv_0.A.n2 mux8_7.inv_0.A.t4 25.395
R19962 mux8_7.inv_0.A.n3 mux8_7.inv_0.A.t2 25.395
R19963 mux8_7.inv_0.A.n3 mux8_7.inv_0.A.t1 25.395
R19964 mux8_7.inv_0.A.n4 mux8_7.inv_0.A.t0 19.8005
R19965 mux8_7.inv_0.A.n4 mux8_7.inv_0.A.t6 19.8005
R19966 a_11865_n25415.n0 a_11865_n25415.n2 231.24
R19967 a_11865_n25415.n5 a_11865_n25415.n1 231.24
R19968 a_11865_n25415.n0 a_11865_n25415.n3 231.03
R19969 a_11865_n25415.n0 a_11865_n25415.n4 231.03
R19970 a_11865_n25415.n6 a_11865_n25415.n5 231.03
R19971 a_11865_n25415.n2 a_11865_n25415.t7 25.395
R19972 a_11865_n25415.n2 a_11865_n25415.t5 25.395
R19973 a_11865_n25415.n3 a_11865_n25415.t8 25.395
R19974 a_11865_n25415.n3 a_11865_n25415.t6 25.395
R19975 a_11865_n25415.n4 a_11865_n25415.t3 25.395
R19976 a_11865_n25415.n4 a_11865_n25415.t9 25.395
R19977 a_11865_n25415.n1 a_11865_n25415.t2 25.395
R19978 a_11865_n25415.n1 a_11865_n25415.t1 25.395
R19979 a_11865_n25415.n6 a_11865_n25415.t0 25.395
R19980 a_11865_n25415.t4 a_11865_n25415.n6 25.395
R19981 a_11865_n25415.n5 a_11865_n25415.n0 0.421553
R19982 mux8_7.A0.n0 mux8_7.A0.t13 1032.02
R19983 mux8_7.A0.n0 mux8_7.A0.t12 336.962
R19984 mux8_7.A0.n0 mux8_7.A0.t14 326.154
R19985 mux8_7.A0 mux8_7.A0.n0 162.952
R19986 mux8_7.A0.n3 mux8_7.A0.n2 120.999
R19987 mux8_7.A0.n3 mux8_7.A0.n1 120.999
R19988 mux8_7.A0.n15 mux8_7.A0.n14 104.489
R19989 mux8_7.A0.n5 mux8_7.A0.n4 92.5005
R19990 mux8_7.A0.n12 mux8_7.A0.n10 86.2638
R19991 mux8_7.A0.n10 mux8_7.A0.n9 85.8873
R19992 mux8_7.A0.n10 mux8_7.A0.n7 85.724
R19993 mux8_7.A0 mux8_7.A0.n15 83.8907
R19994 mux8_7.A0.n13 mux8_7.A0.n9 75.0672
R19995 mux8_7.A0.n13 mux8_7.A0.n12 75.0672
R19996 mux8_7.A0.n7 mux8_7.A0.n6 73.1255
R19997 mux8_7.A0.n9 mux8_7.A0.n8 73.1255
R19998 mux8_7.A0.n12 mux8_7.A0.n11 73.1255
R19999 mux8_7.A0.n14 mux8_7.A0.n7 68.8946
R20000 mux8_7.A0.n15 mux8_7.A0.n5 41.9827
R20001 mux8_7.A0.n4 mux8_7.A0.t10 30.462
R20002 mux8_7.A0.n4 mux8_7.A0.t1 30.462
R20003 mux8_7.A0.n2 mux8_7.A0.t4 30.462
R20004 mux8_7.A0.n2 mux8_7.A0.t2 30.462
R20005 mux8_7.A0.n1 mux8_7.A0.t9 30.462
R20006 mux8_7.A0.n1 mux8_7.A0.t11 30.462
R20007 mux8_7.A0.n5 mux8_7.A0.n3 28.124
R20008 mux8_7.A0.n8 mux8_7.A0.t6 11.8205
R20009 mux8_7.A0.n8 mux8_7.A0.t8 11.8205
R20010 mux8_7.A0.n6 mux8_7.A0.t7 11.8205
R20011 mux8_7.A0.n6 mux8_7.A0.t3 11.8205
R20012 mux8_7.A0.n11 mux8_7.A0.t0 11.8205
R20013 mux8_7.A0.n11 mux8_7.A0.t5 11.8205
R20014 mux8_7.A0.n14 mux8_7.A0.n13 9.3005
R20015 a_n15907_1406.n2 a_n15907_1406.n0 121.353
R20016 a_n15907_1406.n3 a_n15907_1406.n2 121.353
R20017 a_n15907_1406.n2 a_n15907_1406.n1 121.001
R20018 a_n15907_1406.n1 a_n15907_1406.t5 30.462
R20019 a_n15907_1406.n1 a_n15907_1406.t0 30.462
R20020 a_n15907_1406.n0 a_n15907_1406.t4 30.462
R20021 a_n15907_1406.n0 a_n15907_1406.t3 30.462
R20022 a_n15907_1406.n3 a_n15907_1406.t1 30.462
R20023 a_n15907_1406.t2 a_n15907_1406.n3 30.462
R20024 mux8_7.NAND4F_3.Y.n7 mux8_7.NAND4F_3.Y.t9 978.795
R20025 mux8_7.NAND4F_3.Y.n6 mux8_7.NAND4F_3.Y.t11 308.481
R20026 mux8_7.NAND4F_3.Y.n6 mux8_7.NAND4F_3.Y.t10 308.481
R20027 mux8_7.NAND4F_3.Y.n0 mux8_7.NAND4F_3.Y.n1 187.373
R20028 mux8_7.NAND4F_3.Y.n0 mux8_7.NAND4F_3.Y.n2 187.192
R20029 mux8_7.NAND4F_3.Y.n0 mux8_7.NAND4F_3.Y.n3 187.192
R20030 mux8_7.NAND4F_3.Y.n5 mux8_7.NAND4F_3.Y.n4 187.192
R20031 mux8_7.NAND4F_3.Y mux8_7.NAND4F_3.Y.n7 161.839
R20032 mux8_7.NAND4F_3.Y mux8_7.NAND4F_3.Y.t2 23.4426
R20033 mux8_7.NAND4F_3.Y.n1 mux8_7.NAND4F_3.Y.t7 20.1899
R20034 mux8_7.NAND4F_3.Y.n1 mux8_7.NAND4F_3.Y.t8 20.1899
R20035 mux8_7.NAND4F_3.Y.n2 mux8_7.NAND4F_3.Y.t0 20.1899
R20036 mux8_7.NAND4F_3.Y.n2 mux8_7.NAND4F_3.Y.t1 20.1899
R20037 mux8_7.NAND4F_3.Y.n3 mux8_7.NAND4F_3.Y.t6 20.1899
R20038 mux8_7.NAND4F_3.Y.n3 mux8_7.NAND4F_3.Y.t5 20.1899
R20039 mux8_7.NAND4F_3.Y.n4 mux8_7.NAND4F_3.Y.t4 20.1899
R20040 mux8_7.NAND4F_3.Y.n4 mux8_7.NAND4F_3.Y.t3 20.1899
R20041 mux8_7.NAND4F_3.Y.n7 mux8_7.NAND4F_3.Y.n6 11.0463
R20042 mux8_7.NAND4F_3.Y mux8_7.NAND4F_3.Y.n5 0.518495
R20043 mux8_7.NAND4F_3.Y.n5 mux8_7.NAND4F_3.Y.n0 0.358709
R20044 a_11194_n25478.t0 a_11194_n25478.t1 9.9005
R20045 a_11290_n25478.t0 a_11290_n25478.t1 9.9005
R20046 a_n20113_3164.n0 a_n20113_3164.t3 539.788
R20047 a_n20113_3164.n1 a_n20113_3164.t7 531.496
R20048 a_n20113_3164.n0 a_n20113_3164.t5 490.034
R20049 a_n20113_3164.n5 a_n20113_3164.t0 283.788
R20050 a_n20113_3164.t1 a_n20113_3164.n5 205.489
R20051 a_n20113_3164.n2 a_n20113_3164.t2 182.625
R20052 a_n20113_3164.n3 a_n20113_3164.t6 179.054
R20053 a_n20113_3164.n2 a_n20113_3164.t4 139.78
R20054 a_n20113_3164.n4 a_n20113_3164.n3 101.368
R20055 a_n20113_3164.n5 a_n20113_3164.n4 77.9135
R20056 a_n20113_3164.n4 a_n20113_3164.n1 76.1557
R20057 a_n20113_3164.n1 a_n20113_3164.n0 8.29297
R20058 a_n20113_3164.n3 a_n20113_3164.n2 3.57087
R20059 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_0.B MULT_0.4bit_ADDER_1.A0.t5 540.38
R20060 MULT_0.4bit_ADDER_1.A0.n3 MULT_0.4bit_ADDER_1.A0.t13 491.64
R20061 MULT_0.4bit_ADDER_1.A0.n3 MULT_0.4bit_ADDER_1.A0.t7 491.64
R20062 MULT_0.4bit_ADDER_1.A0.n3 MULT_0.4bit_ADDER_1.A0.t15 491.64
R20063 MULT_0.4bit_ADDER_1.A0.n3 MULT_0.4bit_ADDER_1.A0.t6 491.64
R20064 MULT_0.4bit_ADDER_1.A0.n1 MULT_0.4bit_ADDER_1.A0.t10 367.928
R20065 MULT_0.4bit_ADDER_1.A0.n0 MULT_0.4bit_ADDER_1.A0.t3 256.514
R20066 MULT_0.4bit_ADDER_1.A0.n2 MULT_0.4bit_ADDER_1.A0.t4 227.356
R20067 MULT_0.4bit_ADDER_1.A0.n0 MULT_0.4bit_ADDER_1.A0.n7 226.136
R20068 MULT_0.4bit_ADDER_1.A0.n1 MULT_0.4bit_ADDER_1.A0.t11 213.688
R20069 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_0.B MULT_0.4bit_ADDER_1.A0.n5 162.867
R20070 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_0.B MULT_0.4bit_ADDER_1.A0.n2 160.439
R20071 MULT_0.4bit_ADDER_1.A0.n4 MULT_0.4bit_ADDER_1.A0.t9 139.78
R20072 MULT_0.4bit_ADDER_1.A0.n4 MULT_0.4bit_ADDER_1.A0.t12 139.78
R20073 MULT_0.4bit_ADDER_1.A0.n4 MULT_0.4bit_ADDER_1.A0.t8 139.78
R20074 MULT_0.4bit_ADDER_1.A0.n4 MULT_0.4bit_ADDER_1.A0.t14 139.78
R20075 MULT_0.4bit_ADDER_1.A0.n2 MULT_0.4bit_ADDER_1.A0.n1 94.4341
R20076 MULT_0.4bit_ADDER_1.A0.n0 MULT_0.4bit_ADDER_1.A0.t0 83.8326
R20077 MULT_0.4bit_ADDER_1.A0.n5 MULT_0.4bit_ADDER_1.A0.n4 38.6833
R20078 MULT_0.4bit_ADDER_1.A0.n7 MULT_0.4bit_ADDER_1.A0.t1 30.379
R20079 MULT_0.4bit_ADDER_1.A0.n7 MULT_0.4bit_ADDER_1.A0.t2 30.379
R20080 MULT_0.4bit_ADDER_1.A0.n5 MULT_0.4bit_ADDER_1.A0.n3 28.3986
R20081 MULT_0.4bit_ADDER_1.A0.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.A 24.1898
R20082 MULT_0.4bit_ADDER_1.FULL_ADDER_3.A MULT_0.4bit_ADDER_1.A0.n6 16.8273
R20083 MULT_0.4bit_ADDER_1.A0.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_0.B 9.00496
R20084 MULT_0.4bit_ADDER_1.A0.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_0.B 4.77555
R20085 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t10 540.38
R20086 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t7 367.928
R20087 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n5 227.526
R20088 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t9 227.356
R20089 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n4 227.266
R20090 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n6 227.266
R20091 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t8 213.688
R20092 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n2 160.439
R20093 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n1 94.4341
R20094 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t3 42.7944
R20095 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t1 30.379
R20096 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t2 30.379
R20097 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t5 30.379
R20098 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t4 30.379
R20099 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t6 30.379
R20100 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.t0 30.379
R20101 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n0 13.4358
R20102 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B.n3 0.821842
R20103 MULT_0.inv_14.Y.n4 MULT_0.inv_14.Y.t14 540.38
R20104 MULT_0.inv_14.Y.n5 MULT_0.inv_14.Y.t13 491.64
R20105 MULT_0.inv_14.Y.n5 MULT_0.inv_14.Y.t11 491.64
R20106 MULT_0.inv_14.Y.n5 MULT_0.inv_14.Y.t12 491.64
R20107 MULT_0.inv_14.Y.n5 MULT_0.inv_14.Y.t5 491.64
R20108 MULT_0.inv_14.Y.n2 MULT_0.inv_14.Y.t10 367.928
R20109 MULT_0.inv_14.Y.n0 MULT_0.inv_14.Y.t3 256.529
R20110 MULT_0.inv_14.Y.n3 MULT_0.inv_14.Y.t4 227.356
R20111 MULT_0.inv_14.Y.n0 MULT_0.inv_14.Y.n1 226.292
R20112 MULT_0.inv_14.Y.n2 MULT_0.inv_14.Y.t8 213.688
R20113 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_0.B MULT_0.inv_14.Y.n7 162.867
R20114 MULT_0.inv_14.Y.n4 MULT_0.inv_14.Y.n3 160.439
R20115 MULT_0.inv_14.Y.n6 MULT_0.inv_14.Y.t7 139.78
R20116 MULT_0.inv_14.Y.n6 MULT_0.inv_14.Y.t15 139.78
R20117 MULT_0.inv_14.Y.n6 MULT_0.inv_14.Y.t9 139.78
R20118 MULT_0.inv_14.Y.n6 MULT_0.inv_14.Y.t6 139.78
R20119 MULT_0.inv_14.Y.n3 MULT_0.inv_14.Y.n2 94.4341
R20120 MULT_0.inv_14.Y.n0 MULT_0.inv_14.Y.t0 83.7616
R20121 MULT_0.inv_14.Y.n7 MULT_0.inv_14.Y.n6 38.6833
R20122 MULT_0.inv_14.Y.n1 MULT_0.inv_14.Y.t2 30.379
R20123 MULT_0.inv_14.Y.n1 MULT_0.inv_14.Y.t1 30.379
R20124 MULT_0.inv_14.Y.n7 MULT_0.inv_14.Y.n5 28.3986
R20125 MULT_0.4bit_ADDER_2.A2 MULT_0.inv_14.Y.n8 16.8169
R20126 MULT_0.4bit_ADDER_2.A2 MULT_0.inv_14.Y.n0 15.5384
R20127 MULT_0.inv_14.Y.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_0.B 9.00496
R20128 MULT_0.inv_14.Y.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_0.B 3.87912
R20129 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_0.B MULT_0.inv_14.Y.n4 0.89693
R20130 a_n12416_n4534.n0 a_n12416_n4534.n2 81.2978
R20131 a_n12416_n4534.n0 a_n12416_n4534.n3 81.1637
R20132 a_n12416_n4534.n0 a_n12416_n4534.n4 81.1637
R20133 a_n12416_n4534.n1 a_n12416_n4534.n5 81.1637
R20134 a_n12416_n4534.n1 a_n12416_n4534.n6 81.1637
R20135 a_n12416_n4534.n7 a_n12416_n4534.n1 80.9213
R20136 a_n12416_n4534.n2 a_n12416_n4534.t6 11.8205
R20137 a_n12416_n4534.n2 a_n12416_n4534.t8 11.8205
R20138 a_n12416_n4534.n3 a_n12416_n4534.t0 11.8205
R20139 a_n12416_n4534.n3 a_n12416_n4534.t7 11.8205
R20140 a_n12416_n4534.n4 a_n12416_n4534.t5 11.8205
R20141 a_n12416_n4534.n4 a_n12416_n4534.t4 11.8205
R20142 a_n12416_n4534.n5 a_n12416_n4534.t10 11.8205
R20143 a_n12416_n4534.n5 a_n12416_n4534.t11 11.8205
R20144 a_n12416_n4534.n6 a_n12416_n4534.t1 11.8205
R20145 a_n12416_n4534.n6 a_n12416_n4534.t9 11.8205
R20146 a_n12416_n4534.t3 a_n12416_n4534.n7 11.8205
R20147 a_n12416_n4534.n7 a_n12416_n4534.t2 11.8205
R20148 a_n12416_n4534.n1 a_n12416_n4534.n0 0.402735
R20149 mux8_3.NAND4F_7.Y.n2 mux8_3.NAND4F_7.Y.t10 1388.16
R20150 mux8_3.NAND4F_7.Y.n2 mux8_3.NAND4F_7.Y.t9 350.839
R20151 mux8_3.NAND4F_7.Y.n3 mux8_3.NAND4F_7.Y.t11 308.481
R20152 mux8_3.NAND4F_7.Y.n1 mux8_3.NAND4F_7.Y.n4 187.373
R20153 mux8_3.NAND4F_7.Y.n1 mux8_3.NAND4F_7.Y.n5 187.192
R20154 mux8_3.NAND4F_7.Y.n1 mux8_3.NAND4F_7.Y.n6 187.192
R20155 mux8_3.NAND4F_7.Y.n0 mux8_3.NAND4F_7.Y.n7 187.192
R20156 mux8_3.NAND4F_7.Y mux8_3.NAND4F_7.Y.n3 161.492
R20157 mux8_3.NAND4F_7.Y.n3 mux8_3.NAND4F_7.Y.n2 27.752
R20158 mux8_3.NAND4F_7.Y mux8_3.NAND4F_7.Y.t3 23.5642
R20159 mux8_3.NAND4F_7.Y.n4 mux8_3.NAND4F_7.Y.t1 20.1899
R20160 mux8_3.NAND4F_7.Y.n4 mux8_3.NAND4F_7.Y.t0 20.1899
R20161 mux8_3.NAND4F_7.Y.n5 mux8_3.NAND4F_7.Y.t5 20.1899
R20162 mux8_3.NAND4F_7.Y.n5 mux8_3.NAND4F_7.Y.t6 20.1899
R20163 mux8_3.NAND4F_7.Y.n6 mux8_3.NAND4F_7.Y.t8 20.1899
R20164 mux8_3.NAND4F_7.Y.n6 mux8_3.NAND4F_7.Y.t7 20.1899
R20165 mux8_3.NAND4F_7.Y.n7 mux8_3.NAND4F_7.Y.t4 20.1899
R20166 mux8_3.NAND4F_7.Y.n7 mux8_3.NAND4F_7.Y.t2 20.1899
R20167 mux8_3.NAND4F_7.Y mux8_3.NAND4F_7.Y.n0 0.472662
R20168 mux8_3.NAND4F_7.Y.n0 mux8_3.NAND4F_7.Y.n1 0.358709
R20169 mux8_3.NAND4F_9.Y.n1 mux8_3.NAND4F_9.Y.t9 312.599
R20170 mux8_3.NAND4F_9.Y.n4 mux8_3.NAND4F_9.Y.t13 247.428
R20171 mux8_3.NAND4F_9.Y.n1 mux8_3.NAND4F_9.Y.t10 247.428
R20172 mux8_3.NAND4F_9.Y.n2 mux8_3.NAND4F_9.Y.t11 247.428
R20173 mux8_3.NAND4F_9.Y.n3 mux8_3.NAND4F_9.Y.t12 247.428
R20174 mux8_3.NAND4F_9.Y.n5 mux8_3.NAND4F_9.Y.t14 229.754
R20175 mux8_3.NAND4F_9.Y.n0 mux8_3.NAND4F_9.Y.n6 187.373
R20176 mux8_3.NAND4F_9.Y.n0 mux8_3.NAND4F_9.Y.n7 187.192
R20177 mux8_3.NAND4F_9.Y.n0 mux8_3.NAND4F_9.Y.n8 187.192
R20178 mux8_3.NAND4F_9.Y.n10 mux8_3.NAND4F_9.Y.n9 187.192
R20179 mux8_3.NAND4F_9.Y mux8_3.NAND4F_9.Y.n5 162.275
R20180 mux8_3.NAND4F_9.Y.n5 mux8_3.NAND4F_9.Y.n4 91.5805
R20181 mux8_3.NAND4F_9.Y.n2 mux8_3.NAND4F_9.Y.n1 65.1723
R20182 mux8_3.NAND4F_9.Y.n3 mux8_3.NAND4F_9.Y.n2 65.1723
R20183 mux8_3.NAND4F_9.Y.n4 mux8_3.NAND4F_9.Y.n3 65.1723
R20184 mux8_3.NAND4F_9.Y mux8_3.NAND4F_9.Y.t2 22.6141
R20185 mux8_3.NAND4F_9.Y.n6 mux8_3.NAND4F_9.Y.t6 20.1899
R20186 mux8_3.NAND4F_9.Y.n6 mux8_3.NAND4F_9.Y.t5 20.1899
R20187 mux8_3.NAND4F_9.Y.n7 mux8_3.NAND4F_9.Y.t7 20.1899
R20188 mux8_3.NAND4F_9.Y.n7 mux8_3.NAND4F_9.Y.t8 20.1899
R20189 mux8_3.NAND4F_9.Y.n8 mux8_3.NAND4F_9.Y.t3 20.1899
R20190 mux8_3.NAND4F_9.Y.n8 mux8_3.NAND4F_9.Y.t4 20.1899
R20191 mux8_3.NAND4F_9.Y.n9 mux8_3.NAND4F_9.Y.t0 20.1899
R20192 mux8_3.NAND4F_9.Y.n9 mux8_3.NAND4F_9.Y.t1 20.1899
R20193 mux8_3.NAND4F_9.Y mux8_3.NAND4F_9.Y.n10 0.396904
R20194 mux8_3.NAND4F_9.Y.n10 mux8_3.NAND4F_9.Y.n0 0.358709
R20195 mux8_6.A0.n0 mux8_6.A0.t13 1032.02
R20196 mux8_6.A0.n1 mux8_6.A0.t19 491.64
R20197 mux8_6.A0.n1 mux8_6.A0.t17 491.64
R20198 mux8_6.A0.n1 mux8_6.A0.t22 491.64
R20199 mux8_6.A0.n1 mux8_6.A0.t15 491.64
R20200 mux8_6.A0.n0 mux8_6.A0.t20 336.962
R20201 mux8_6.A0.n0 mux8_6.A0.t14 326.154
R20202 mux8_6.A0 mux8_6.A0.n0 162.952
R20203 mux8_6.A0 mux8_6.A0.n3 162.909
R20204 mux8_6.A0.n2 mux8_6.A0.t18 139.78
R20205 mux8_6.A0.n2 mux8_6.A0.t21 139.78
R20206 mux8_6.A0.n2 mux8_6.A0.t16 139.78
R20207 mux8_6.A0.n2 mux8_6.A0.t12 139.78
R20208 mux8_6.A0.n8 mux8_6.A0.n7 120.999
R20209 mux8_6.A0.n8 mux8_6.A0.n6 120.999
R20210 mux8_6.A0.n20 mux8_6.A0.n19 104.489
R20211 mux8_6.A0.n10 mux8_6.A0.n9 92.5005
R20212 mux8_6.A0.n17 mux8_6.A0.n15 86.2638
R20213 mux8_6.A0.n15 mux8_6.A0.n14 85.8873
R20214 mux8_6.A0.n15 mux8_6.A0.n12 85.724
R20215 mux8_6.A0 mux8_6.A0.n20 83.8907
R20216 mux8_6.A0.n5 mux8_6.A0 77.7751
R20217 mux8_6.A0.n18 mux8_6.A0.n17 75.0672
R20218 mux8_6.A0.n18 mux8_6.A0.n14 75.0672
R20219 mux8_6.A0.n17 mux8_6.A0.n16 73.1255
R20220 mux8_6.A0.n12 mux8_6.A0.n11 73.1255
R20221 mux8_6.A0.n14 mux8_6.A0.n13 73.1255
R20222 mux8_6.A0.n19 mux8_6.A0.n12 68.8946
R20223 mux8_6.A0 mux8_6.A0.n5 56.1975
R20224 mux8_6.A0.n5 mux8_6.A0.n4 45.3038
R20225 mux8_6.A0.n20 mux8_6.A0.n10 41.9827
R20226 mux8_6.A0.n3 mux8_6.A0.n2 38.6833
R20227 mux8_6.A0.n9 mux8_6.A0.t0 30.462
R20228 mux8_6.A0.n9 mux8_6.A0.t11 30.462
R20229 mux8_6.A0.n7 mux8_6.A0.t6 30.462
R20230 mux8_6.A0.n7 mux8_6.A0.t7 30.462
R20231 mux8_6.A0.n6 mux8_6.A0.t1 30.462
R20232 mux8_6.A0.n6 mux8_6.A0.t2 30.462
R20233 mux8_6.A0.n3 mux8_6.A0.n1 28.3986
R20234 mux8_6.A0.n10 mux8_6.A0.n8 28.124
R20235 mux8_6.A0.n11 mux8_6.A0.t5 11.8205
R20236 mux8_6.A0.n11 mux8_6.A0.t10 11.8205
R20237 mux8_6.A0.n16 mux8_6.A0.t8 11.8205
R20238 mux8_6.A0.n16 mux8_6.A0.t9 11.8205
R20239 mux8_6.A0.n13 mux8_6.A0.t4 11.8205
R20240 mux8_6.A0.n13 mux8_6.A0.t3 11.8205
R20241 mux8_6.A0.n4 mux8_6.A0 10.8551
R20242 mux8_6.A0.n19 mux8_6.A0.n18 9.3005
R20243 mux8_6.A0.n4 mux8_6.A0 4.5005
R20244 a_5773_4912.n2 a_5773_4912.n0 121.353
R20245 a_5773_4912.n3 a_5773_4912.n2 121.353
R20246 a_5773_4912.n2 a_5773_4912.n1 121.001
R20247 a_5773_4912.n1 a_5773_4912.t5 30.462
R20248 a_5773_4912.n1 a_5773_4912.t0 30.462
R20249 a_5773_4912.n0 a_5773_4912.t4 30.462
R20250 a_5773_4912.n0 a_5773_4912.t3 30.462
R20251 a_5773_4912.t2 a_5773_4912.n3 30.462
R20252 a_5773_4912.n3 a_5773_4912.t1 30.462
R20253 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t17 491.64
R20254 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t15 491.64
R20255 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t13 491.64
R20256 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t20 491.64
R20257 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t19 485.221
R20258 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t23 367.928
R20259 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t14 255.588
R20260 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t21 224.478
R20261 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t22 213.688
R20262 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n0 209.19
R20263 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t16 139.78
R20264 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t12 139.78
R20265 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t18 139.78
R20266 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n10 120.999
R20267 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n9 120.999
R20268 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n22 104.489
R20269 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n12 92.5005
R20270 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n18 86.2638
R20271 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n17 85.8873
R20272 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n15 85.724
R20273 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n7 84.5046
R20274 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n23 83.8907
R20275 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n17 75.0672
R20276 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n20 75.0672
R20277 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n15 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n14 73.1255
R20278 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n17 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n16 73.1255
R20279 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n19 73.1255
R20280 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n6 72.3005
R20281 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n15 68.8946
R20282 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n8 60.9797
R20283 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n13 41.9827
R20284 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t7 30.462
R20285 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t1 30.462
R20286 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t11 30.462
R20287 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t10 30.462
R20288 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t6 30.462
R20289 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t5 30.462
R20290 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n11 28.124
R20291 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n5 19.963
R20292 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n1 17.8661
R20293 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n2 17.8661
R20294 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n3 17.1217
R20295 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t3 11.8205
R20296 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t2 11.8205
R20297 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t4 11.8205
R20298 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t9 11.8205
R20299 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t8 11.8205
R20300 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t0 11.8205
R20301 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n21 9.3005
R20302 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n4 1.8615
R20303 8bit_ADDER_0.S2.n0 8bit_ADDER_0.S2.t12 1032.02
R20304 8bit_ADDER_0.S2.n0 8bit_ADDER_0.S2.t14 336.962
R20305 8bit_ADDER_0.S2.n0 8bit_ADDER_0.S2.t13 326.154
R20306 8bit_ADDER_0.S2 8bit_ADDER_0.S2.n0 162.952
R20307 8bit_ADDER_0.S2.n3 8bit_ADDER_0.S2.n2 120.999
R20308 8bit_ADDER_0.S2.n3 8bit_ADDER_0.S2.n1 120.999
R20309 8bit_ADDER_0.S2.n15 8bit_ADDER_0.S2.n14 104.489
R20310 8bit_ADDER_0.S2.n5 8bit_ADDER_0.S2.n4 92.5005
R20311 8bit_ADDER_0.S2.n12 8bit_ADDER_0.S2.n10 86.2638
R20312 8bit_ADDER_0.S2.n10 8bit_ADDER_0.S2.n9 85.8873
R20313 8bit_ADDER_0.S2.n10 8bit_ADDER_0.S2.n7 85.724
R20314 8bit_ADDER_0.S2 8bit_ADDER_0.S2.n15 83.8907
R20315 8bit_ADDER_0.S2.n13 8bit_ADDER_0.S2.n12 75.0672
R20316 8bit_ADDER_0.S2.n13 8bit_ADDER_0.S2.n9 75.0672
R20317 8bit_ADDER_0.S2.n12 8bit_ADDER_0.S2.n11 73.1255
R20318 8bit_ADDER_0.S2.n9 8bit_ADDER_0.S2.n8 73.1255
R20319 8bit_ADDER_0.S2.n7 8bit_ADDER_0.S2.n6 73.1255
R20320 8bit_ADDER_0.S2.n14 8bit_ADDER_0.S2.n7 68.8946
R20321 8bit_ADDER_0.S2.n15 8bit_ADDER_0.S2.n5 41.9827
R20322 8bit_ADDER_0.S2.n4 8bit_ADDER_0.S2.t4 30.462
R20323 8bit_ADDER_0.S2.n4 8bit_ADDER_0.S2.t11 30.462
R20324 8bit_ADDER_0.S2.n2 8bit_ADDER_0.S2.t0 30.462
R20325 8bit_ADDER_0.S2.n2 8bit_ADDER_0.S2.t9 30.462
R20326 8bit_ADDER_0.S2.n1 8bit_ADDER_0.S2.t6 30.462
R20327 8bit_ADDER_0.S2.n1 8bit_ADDER_0.S2.t5 30.462
R20328 8bit_ADDER_0.S2.n5 8bit_ADDER_0.S2.n3 28.124
R20329 8bit_ADDER_0.S2.n8 8bit_ADDER_0.S2.t2 11.8205
R20330 8bit_ADDER_0.S2.n8 8bit_ADDER_0.S2.t3 11.8205
R20331 8bit_ADDER_0.S2.n11 8bit_ADDER_0.S2.t10 11.8205
R20332 8bit_ADDER_0.S2.n11 8bit_ADDER_0.S2.t7 11.8205
R20333 8bit_ADDER_0.S2.n6 8bit_ADDER_0.S2.t1 11.8205
R20334 8bit_ADDER_0.S2.n6 8bit_ADDER_0.S2.t8 11.8205
R20335 8bit_ADDER_0.S2.n14 8bit_ADDER_0.S2.n13 9.3005
R20336 a_n6035_1406.n2 a_n6035_1406.n0 121.353
R20337 a_n6035_1406.n3 a_n6035_1406.n2 121.353
R20338 a_n6035_1406.n2 a_n6035_1406.n1 121.001
R20339 a_n6035_1406.n1 a_n6035_1406.t1 30.462
R20340 a_n6035_1406.n1 a_n6035_1406.t5 30.462
R20341 a_n6035_1406.n0 a_n6035_1406.t0 30.462
R20342 a_n6035_1406.n0 a_n6035_1406.t2 30.462
R20343 a_n6035_1406.t4 a_n6035_1406.n3 30.462
R20344 a_n6035_1406.n3 a_n6035_1406.t3 30.462
R20345 a_n17296_n8445.n2 a_n17296_n8445.t3 541.395
R20346 a_n17296_n8445.n3 a_n17296_n8445.t7 527.402
R20347 a_n17296_n8445.n2 a_n17296_n8445.t2 491.64
R20348 a_n17296_n8445.n5 a_n17296_n8445.t0 281.906
R20349 a_n17296_n8445.t1 a_n17296_n8445.n5 204.359
R20350 a_n17296_n8445.n0 a_n17296_n8445.t4 180.73
R20351 a_n17296_n8445.n1 a_n17296_n8445.t6 179.45
R20352 a_n17296_n8445.n0 a_n17296_n8445.t5 139.78
R20353 a_n17296_n8445.n4 a_n17296_n8445.n1 105.635
R20354 a_n17296_n8445.n4 a_n17296_n8445.n3 76.0005
R20355 a_n17296_n8445.n5 a_n17296_n8445.n4 67.9685
R20356 a_n17296_n8445.n3 a_n17296_n8445.n2 13.994
R20357 a_n17296_n8445.n1 a_n17296_n8445.n0 1.28015
R20358 a_n17266_n7799.n7 a_n17266_n7799.n1 81.2978
R20359 a_n17266_n7799.n1 a_n17266_n7799.n6 81.1637
R20360 a_n17266_n7799.n1 a_n17266_n7799.n5 81.1637
R20361 a_n17266_n7799.n0 a_n17266_n7799.n4 81.1637
R20362 a_n17266_n7799.n0 a_n17266_n7799.n3 81.1637
R20363 a_n17266_n7799.n0 a_n17266_n7799.n2 80.9213
R20364 a_n17266_n7799.n6 a_n17266_n7799.t8 11.8205
R20365 a_n17266_n7799.n6 a_n17266_n7799.t6 11.8205
R20366 a_n17266_n7799.n5 a_n17266_n7799.t3 11.8205
R20367 a_n17266_n7799.n5 a_n17266_n7799.t4 11.8205
R20368 a_n17266_n7799.n4 a_n17266_n7799.t2 11.8205
R20369 a_n17266_n7799.n4 a_n17266_n7799.t1 11.8205
R20370 a_n17266_n7799.n3 a_n17266_n7799.t9 11.8205
R20371 a_n17266_n7799.n3 a_n17266_n7799.t0 11.8205
R20372 a_n17266_n7799.n2 a_n17266_n7799.t11 11.8205
R20373 a_n17266_n7799.n2 a_n17266_n7799.t10 11.8205
R20374 a_n17266_n7799.n7 a_n17266_n7799.t5 11.8205
R20375 a_n17266_n7799.t7 a_n17266_n7799.n7 11.8205
R20376 a_n17266_n7799.n1 a_n17266_n7799.n0 0.402735
R20377 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t14 491.64
R20378 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t17 491.64
R20379 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t19 491.64
R20380 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t15 491.64
R20381 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n8 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t18 485.221
R20382 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t12 367.928
R20383 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t22 255.588
R20384 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t16 224.478
R20385 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t13 213.688
R20386 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n0 209.19
R20387 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t20 139.78
R20388 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t21 139.78
R20389 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t23 139.78
R20390 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n11 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n10 120.999
R20391 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n11 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n9 120.999
R20392 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n23 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n22 104.489
R20393 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n13 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n12 92.5005
R20394 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n20 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n18 86.2638
R20395 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n18 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n17 85.8873
R20396 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n18 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n15 85.724
R20397 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n8 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n7 84.5046
R20398 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n23 83.8907
R20399 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n21 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n20 75.0672
R20400 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n21 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n17 75.0672
R20401 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n20 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n19 73.1255
R20402 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n15 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n14 73.1255
R20403 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n17 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n16 73.1255
R20404 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n7 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n6 72.3005
R20405 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n22 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n15 68.8946
R20406 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n8 60.9797
R20407 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n23 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n13 41.9827
R20408 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n12 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t8 30.462
R20409 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n12 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t3 30.462
R20410 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n10 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t4 30.462
R20411 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n10 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t5 30.462
R20412 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n9 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t10 30.462
R20413 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n9 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t9 30.462
R20414 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n13 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n11 28.124
R20415 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n5 19.963
R20416 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n1 17.8661
R20417 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n2 17.8661
R20418 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n3 17.1217
R20419 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n14 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t1 11.8205
R20420 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n14 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t6 11.8205
R20421 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n19 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t7 11.8205
R20422 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n19 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t11 11.8205
R20423 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n16 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t0 11.8205
R20424 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n16 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t2 11.8205
R20425 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n22 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n21 9.3005
R20426 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n4 1.8615
R20427 a_n6950_3164.n0 a_n6950_3164.t7 539.788
R20428 a_n6950_3164.n1 a_n6950_3164.t5 531.496
R20429 a_n6950_3164.n0 a_n6950_3164.t3 490.034
R20430 a_n6950_3164.n5 a_n6950_3164.t0 283.788
R20431 a_n6950_3164.t1 a_n6950_3164.n5 205.489
R20432 a_n6950_3164.n2 a_n6950_3164.t6 182.625
R20433 a_n6950_3164.n3 a_n6950_3164.t4 179.054
R20434 a_n6950_3164.n2 a_n6950_3164.t2 139.78
R20435 a_n6950_3164.n4 a_n6950_3164.n3 101.368
R20436 a_n6950_3164.n5 a_n6950_3164.n4 77.9135
R20437 a_n6950_3164.n4 a_n6950_3164.n1 76.1557
R20438 a_n6950_3164.n1 a_n6950_3164.n0 8.29297
R20439 a_n6950_3164.n3 a_n6950_3164.n2 3.57087
R20440 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t10 540.38
R20441 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t7 367.928
R20442 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n4 227.526
R20443 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t9 227.356
R20444 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n5 227.266
R20445 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n6 227.266
R20446 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t8 213.688
R20447 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n2 160.439
R20448 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n1 94.4341
R20449 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t0 42.7944
R20450 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t5 30.379
R20451 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t6 30.379
R20452 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t2 30.379
R20453 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t4 30.379
R20454 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t1 30.379
R20455 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.t3 30.379
R20456 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n0 13.4358
R20457 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B.n3 0.821842
R20458 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n9 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t8 540.38
R20459 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t12 491.64
R20460 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t17 491.64
R20461 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t16 491.64
R20462 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t7 491.64
R20463 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t10 367.928
R20464 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n1 227.526
R20465 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n8 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t15 227.356
R20466 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n2 227.266
R20467 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n3 227.266
R20468 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t11 213.688
R20469 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n6 162.852
R20470 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n9 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n8 160.439
R20471 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t13 139.78
R20472 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t18 139.78
R20473 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t9 139.78
R20474 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t14 139.78
R20475 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n8 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n7 94.4341
R20476 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t3 42.7831
R20477 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n5 38.6833
R20478 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t1 30.379
R20479 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t2 30.379
R20480 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t4 30.379
R20481 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t0 30.379
R20482 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t6 30.379
R20483 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t5 30.379
R20484 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n4 28.3986
R20485 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n0 18.8832
R20486 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n10 10.7052
R20487 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n10 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT 5.09176
R20488 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n10 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT 4.19292
R20489 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n9 0.794268
R20490 mux8_6.NAND4F_4.Y.n6 mux8_6.NAND4F_4.Y.t10 1032.02
R20491 mux8_6.NAND4F_4.Y.n6 mux8_6.NAND4F_4.Y.t11 336.962
R20492 mux8_6.NAND4F_4.Y.n6 mux8_6.NAND4F_4.Y.t9 326.154
R20493 mux8_6.NAND4F_4.Y.n0 mux8_6.NAND4F_4.Y.n1 187.373
R20494 mux8_6.NAND4F_4.Y.n0 mux8_6.NAND4F_4.Y.n2 187.192
R20495 mux8_6.NAND4F_4.Y.n0 mux8_6.NAND4F_4.Y.n3 187.192
R20496 mux8_6.NAND4F_4.Y.n5 mux8_6.NAND4F_4.Y.n4 187.192
R20497 mux8_6.NAND4F_4.Y mux8_6.NAND4F_4.Y.n6 162.942
R20498 mux8_6.NAND4F_4.Y.n7 mux8_6.NAND4F_4.Y 24.5377
R20499 mux8_6.NAND4F_4.Y.n7 mux8_6.NAND4F_4.Y.t4 22.6141
R20500 mux8_6.NAND4F_4.Y.n1 mux8_6.NAND4F_4.Y.t0 20.1899
R20501 mux8_6.NAND4F_4.Y.n1 mux8_6.NAND4F_4.Y.t1 20.1899
R20502 mux8_6.NAND4F_4.Y.n2 mux8_6.NAND4F_4.Y.t5 20.1899
R20503 mux8_6.NAND4F_4.Y.n2 mux8_6.NAND4F_4.Y.t6 20.1899
R20504 mux8_6.NAND4F_4.Y.n3 mux8_6.NAND4F_4.Y.t8 20.1899
R20505 mux8_6.NAND4F_4.Y.n3 mux8_6.NAND4F_4.Y.t7 20.1899
R20506 mux8_6.NAND4F_4.Y.n4 mux8_6.NAND4F_4.Y.t2 20.1899
R20507 mux8_6.NAND4F_4.Y.n4 mux8_6.NAND4F_4.Y.t3 20.1899
R20508 mux8_6.NAND4F_4.Y mux8_6.NAND4F_4.Y.n7 0.894894
R20509 mux8_6.NAND4F_4.Y mux8_6.NAND4F_4.Y.n5 0.452586
R20510 mux8_6.NAND4F_4.Y.n5 mux8_6.NAND4F_4.Y.n0 0.358709
R20511 mux8_6.NAND4F_8.Y.n1 mux8_6.NAND4F_8.Y.t14 379.173
R20512 mux8_6.NAND4F_8.Y.n2 mux8_6.NAND4F_8.Y.t13 312.599
R20513 mux8_6.NAND4F_8.Y.n1 mux8_6.NAND4F_8.Y.t9 247.428
R20514 mux8_6.NAND4F_8.Y.n4 mux8_6.NAND4F_8.Y.t10 247.428
R20515 mux8_6.NAND4F_8.Y.n3 mux8_6.NAND4F_8.Y.t12 247.428
R20516 mux8_6.NAND4F_8.Y.n2 mux8_6.NAND4F_8.Y.t11 247.428
R20517 mux8_6.NAND4F_8.Y.n0 mux8_6.NAND4F_8.Y.n6 187.373
R20518 mux8_6.NAND4F_8.Y.n0 mux8_6.NAND4F_8.Y.n7 187.192
R20519 mux8_6.NAND4F_8.Y.n0 mux8_6.NAND4F_8.Y.n8 187.192
R20520 mux8_6.NAND4F_8.Y.n10 mux8_6.NAND4F_8.Y.n9 187.192
R20521 mux8_6.NAND4F_8.Y mux8_6.NAND4F_8.Y.n5 162.139
R20522 mux8_6.NAND4F_8.Y.n4 mux8_6.NAND4F_8.Y.n3 65.1723
R20523 mux8_6.NAND4F_8.Y.n3 mux8_6.NAND4F_8.Y.n2 65.1723
R20524 mux8_6.NAND4F_8.Y.n5 mux8_6.NAND4F_8.Y.n4 33.2653
R20525 mux8_6.NAND4F_8.Y.n5 mux8_6.NAND4F_8.Y.n1 31.9075
R20526 mux8_6.NAND4F_8.Y mux8_6.NAND4F_8.Y.t2 22.6141
R20527 mux8_6.NAND4F_8.Y.n6 mux8_6.NAND4F_8.Y.t1 20.1899
R20528 mux8_6.NAND4F_8.Y.n6 mux8_6.NAND4F_8.Y.t0 20.1899
R20529 mux8_6.NAND4F_8.Y.n7 mux8_6.NAND4F_8.Y.t5 20.1899
R20530 mux8_6.NAND4F_8.Y.n7 mux8_6.NAND4F_8.Y.t6 20.1899
R20531 mux8_6.NAND4F_8.Y.n8 mux8_6.NAND4F_8.Y.t7 20.1899
R20532 mux8_6.NAND4F_8.Y.n8 mux8_6.NAND4F_8.Y.t8 20.1899
R20533 mux8_6.NAND4F_8.Y.n9 mux8_6.NAND4F_8.Y.t3 20.1899
R20534 mux8_6.NAND4F_8.Y.n9 mux8_6.NAND4F_8.Y.t4 20.1899
R20535 mux8_6.NAND4F_8.Y mux8_6.NAND4F_8.Y.n10 0.452586
R20536 mux8_6.NAND4F_8.Y.n10 mux8_6.NAND4F_8.Y.n0 0.358709
R20537 V_FLAG_0.XOR2_2.B.n0 V_FLAG_0.XOR2_2.B.t17 491.64
R20538 V_FLAG_0.XOR2_2.B.n0 V_FLAG_0.XOR2_2.B.t15 491.64
R20539 V_FLAG_0.XOR2_2.B.n0 V_FLAG_0.XOR2_2.B.t13 491.64
R20540 V_FLAG_0.XOR2_2.B.n0 V_FLAG_0.XOR2_2.B.t16 491.64
R20541 V_FLAG_0.XOR2_2.B V_FLAG_0.XOR2_2.B.n2 162.924
R20542 V_FLAG_0.XOR2_2.B.n1 V_FLAG_0.XOR2_2.B.t18 139.78
R20543 V_FLAG_0.XOR2_2.B.n1 V_FLAG_0.XOR2_2.B.t12 139.78
R20544 V_FLAG_0.XOR2_2.B.n1 V_FLAG_0.XOR2_2.B.t14 139.78
R20545 V_FLAG_0.XOR2_2.B.n1 V_FLAG_0.XOR2_2.B.t19 139.78
R20546 V_FLAG_0.XOR2_2.B.n5 V_FLAG_0.XOR2_2.B.n4 120.999
R20547 V_FLAG_0.XOR2_2.B.n5 V_FLAG_0.XOR2_2.B.n3 120.999
R20548 V_FLAG_0.XOR2_2.B.n17 V_FLAG_0.XOR2_2.B.n16 104.489
R20549 V_FLAG_0.XOR2_2.B.n7 V_FLAG_0.XOR2_2.B.n6 92.5005
R20550 V_FLAG_0.XOR2_2.B.n14 V_FLAG_0.XOR2_2.B.n12 86.2638
R20551 V_FLAG_0.XOR2_2.B.n12 V_FLAG_0.XOR2_2.B.n11 85.8873
R20552 V_FLAG_0.XOR2_2.B.n12 V_FLAG_0.XOR2_2.B.n9 85.724
R20553 V_FLAG_0.XOR2_2.B V_FLAG_0.XOR2_2.B.n17 84.0552
R20554 V_FLAG_0.XOR2_2.B.n15 V_FLAG_0.XOR2_2.B.n11 75.0672
R20555 V_FLAG_0.XOR2_2.B.n15 V_FLAG_0.XOR2_2.B.n14 75.0672
R20556 V_FLAG_0.XOR2_2.B.n9 V_FLAG_0.XOR2_2.B.n8 73.1255
R20557 V_FLAG_0.XOR2_2.B.n11 V_FLAG_0.XOR2_2.B.n10 73.1255
R20558 V_FLAG_0.XOR2_2.B.n14 V_FLAG_0.XOR2_2.B.n13 73.1255
R20559 V_FLAG_0.XOR2_2.B.n16 V_FLAG_0.XOR2_2.B.n9 68.8946
R20560 V_FLAG_0.XOR2_2.B.n17 V_FLAG_0.XOR2_2.B.n7 41.9827
R20561 V_FLAG_0.XOR2_2.B.n2 V_FLAG_0.XOR2_2.B.n1 38.6833
R20562 V_FLAG_0.XOR2_2.B.n6 V_FLAG_0.XOR2_2.B.t2 30.462
R20563 V_FLAG_0.XOR2_2.B.n6 V_FLAG_0.XOR2_2.B.t4 30.462
R20564 V_FLAG_0.XOR2_2.B.n4 V_FLAG_0.XOR2_2.B.t6 30.462
R20565 V_FLAG_0.XOR2_2.B.n4 V_FLAG_0.XOR2_2.B.t11 30.462
R20566 V_FLAG_0.XOR2_2.B.n3 V_FLAG_0.XOR2_2.B.t3 30.462
R20567 V_FLAG_0.XOR2_2.B.n3 V_FLAG_0.XOR2_2.B.t1 30.462
R20568 V_FLAG_0.XOR2_2.B.n2 V_FLAG_0.XOR2_2.B.n0 28.3986
R20569 V_FLAG_0.XOR2_2.B.n7 V_FLAG_0.XOR2_2.B.n5 28.124
R20570 V_FLAG_0.XOR2_2.B.n10 V_FLAG_0.XOR2_2.B.t8 11.8205
R20571 V_FLAG_0.XOR2_2.B.n10 V_FLAG_0.XOR2_2.B.t9 11.8205
R20572 V_FLAG_0.XOR2_2.B.n8 V_FLAG_0.XOR2_2.B.t10 11.8205
R20573 V_FLAG_0.XOR2_2.B.n8 V_FLAG_0.XOR2_2.B.t5 11.8205
R20574 V_FLAG_0.XOR2_2.B.n13 V_FLAG_0.XOR2_2.B.t7 11.8205
R20575 V_FLAG_0.XOR2_2.B.n13 V_FLAG_0.XOR2_2.B.t0 11.8205
R20576 V_FLAG_0.XOR2_2.B.n16 V_FLAG_0.XOR2_2.B.n15 9.3005
R20577 mux8_0.NAND4F_2.D.n4 mux8_0.NAND4F_2.D.t13 1388.16
R20578 mux8_0.NAND4F_2.D.n7 mux8_0.NAND4F_2.D.t5 1388.16
R20579 mux8_0.NAND4F_2.D.n10 mux8_0.NAND4F_2.D.t9 1388.16
R20580 mux8_0.NAND4F_2.D.n1 mux8_0.NAND4F_2.D.t7 1388.16
R20581 mux8_0.NAND4F_2.D.n4 mux8_0.NAND4F_2.D.t12 350.839
R20582 mux8_0.NAND4F_2.D.n7 mux8_0.NAND4F_2.D.t11 350.839
R20583 mux8_0.NAND4F_2.D.n10 mux8_0.NAND4F_2.D.t10 350.839
R20584 mux8_0.NAND4F_2.D.n1 mux8_0.NAND4F_2.D.t6 350.839
R20585 mux8_0.NAND4F_2.D.n5 mux8_0.NAND4F_2.D.t4 308.481
R20586 mux8_0.NAND4F_2.D.n8 mux8_0.NAND4F_2.D.t15 308.481
R20587 mux8_0.NAND4F_2.D.n11 mux8_0.NAND4F_2.D.t14 308.481
R20588 mux8_0.NAND4F_2.D.n2 mux8_0.NAND4F_2.D.t8 308.481
R20589 mux8_0.NAND4F_2.D.n0 mux8_0.NAND4F_2.D.t1 256.514
R20590 mux8_0.NAND4F_2.D.n0 mux8_0.NAND4F_2.D.n3 226.258
R20591 mux8_0.NAND4F_2.D mux8_0.NAND4F_2.D.n5 161.458
R20592 mux8_0.NAND4F_2.D mux8_0.NAND4F_2.D.n11 161.435
R20593 mux8_0.NAND4F_2.D mux8_0.NAND4F_2.D.n2 161.435
R20594 mux8_0.NAND4F_2.D mux8_0.NAND4F_2.D.n8 161.429
R20595 mux8_0.NAND4F_2.D.n0 mux8_0.NAND4F_2.D.t0 83.7172
R20596 mux8_0.NAND4F_2.D.n3 mux8_0.NAND4F_2.D.t2 30.379
R20597 mux8_0.NAND4F_2.D.n3 mux8_0.NAND4F_2.D.t3 30.379
R20598 mux8_0.NAND4F_2.D.n5 mux8_0.NAND4F_2.D.n4 27.752
R20599 mux8_0.NAND4F_2.D.n8 mux8_0.NAND4F_2.D.n7 27.752
R20600 mux8_0.NAND4F_2.D.n11 mux8_0.NAND4F_2.D.n10 27.752
R20601 mux8_0.NAND4F_2.D.n2 mux8_0.NAND4F_2.D.n1 27.752
R20602 mux8_0.NAND4F_2.D.n6 mux8_0.NAND4F_2.D.n0 12.759
R20603 mux8_0.NAND4F_2.D mux8_0.NAND4F_2.D.n12 10.6871
R20604 mux8_0.NAND4F_2.D.n6 mux8_0.NAND4F_2.D 9.0005
R20605 mux8_0.NAND4F_2.D.n12 mux8_0.NAND4F_2.D 9.0005
R20606 mux8_0.NAND4F_2.D.n9 mux8_0.NAND4F_2.D 9.0005
R20607 mux8_0.NAND4F_2.D.n9 mux8_0.NAND4F_2.D.n6 1.74507
R20608 mux8_0.NAND4F_2.D.n12 mux8_0.NAND4F_2.D.n9 1.69072
R20609 mux8_2.NAND4F_4.Y.n6 mux8_2.NAND4F_4.Y.t11 1032.02
R20610 mux8_2.NAND4F_4.Y.n6 mux8_2.NAND4F_4.Y.t10 336.962
R20611 mux8_2.NAND4F_4.Y.n6 mux8_2.NAND4F_4.Y.t9 326.154
R20612 mux8_2.NAND4F_4.Y.n0 mux8_2.NAND4F_4.Y.n1 187.373
R20613 mux8_2.NAND4F_4.Y.n0 mux8_2.NAND4F_4.Y.n2 187.192
R20614 mux8_2.NAND4F_4.Y.n0 mux8_2.NAND4F_4.Y.n3 187.192
R20615 mux8_2.NAND4F_4.Y.n5 mux8_2.NAND4F_4.Y.n4 187.192
R20616 mux8_2.NAND4F_4.Y mux8_2.NAND4F_4.Y.n6 162.942
R20617 mux8_2.NAND4F_4.Y.n7 mux8_2.NAND4F_4.Y 24.5377
R20618 mux8_2.NAND4F_4.Y.n7 mux8_2.NAND4F_4.Y.t0 22.6141
R20619 mux8_2.NAND4F_4.Y.n1 mux8_2.NAND4F_4.Y.t6 20.1899
R20620 mux8_2.NAND4F_4.Y.n1 mux8_2.NAND4F_4.Y.t5 20.1899
R20621 mux8_2.NAND4F_4.Y.n2 mux8_2.NAND4F_4.Y.t4 20.1899
R20622 mux8_2.NAND4F_4.Y.n2 mux8_2.NAND4F_4.Y.t3 20.1899
R20623 mux8_2.NAND4F_4.Y.n3 mux8_2.NAND4F_4.Y.t8 20.1899
R20624 mux8_2.NAND4F_4.Y.n3 mux8_2.NAND4F_4.Y.t7 20.1899
R20625 mux8_2.NAND4F_4.Y.n4 mux8_2.NAND4F_4.Y.t2 20.1899
R20626 mux8_2.NAND4F_4.Y.n4 mux8_2.NAND4F_4.Y.t1 20.1899
R20627 mux8_2.NAND4F_4.Y mux8_2.NAND4F_4.Y.n7 0.894894
R20628 mux8_2.NAND4F_4.Y mux8_2.NAND4F_4.Y.n5 0.452586
R20629 mux8_2.NAND4F_4.Y.n5 mux8_2.NAND4F_4.Y.n0 0.358709
R20630 a_n17677_n18225.n0 a_n17677_n18225.n2 231.24
R20631 a_n17677_n18225.n6 a_n17677_n18225.n1 231.24
R20632 a_n17677_n18225.n0 a_n17677_n18225.n3 231.03
R20633 a_n17677_n18225.n1 a_n17677_n18225.n4 231.03
R20634 a_n17677_n18225.n1 a_n17677_n18225.n5 231.03
R20635 a_n17677_n18225.n2 a_n17677_n18225.t3 25.395
R20636 a_n17677_n18225.n2 a_n17677_n18225.t2 25.395
R20637 a_n17677_n18225.n3 a_n17677_n18225.t1 25.395
R20638 a_n17677_n18225.n3 a_n17677_n18225.t0 25.395
R20639 a_n17677_n18225.n4 a_n17677_n18225.t4 25.395
R20640 a_n17677_n18225.n4 a_n17677_n18225.t6 25.395
R20641 a_n17677_n18225.n5 a_n17677_n18225.t5 25.395
R20642 a_n17677_n18225.n5 a_n17677_n18225.t9 25.395
R20643 a_n17677_n18225.t8 a_n17677_n18225.n6 25.395
R20644 a_n17677_n18225.n6 a_n17677_n18225.t7 25.395
R20645 a_n17677_n18225.n1 a_n17677_n18225.n0 0.421553
R20646 A0.n19 A0.t27 540.38
R20647 A0.n5 A0.t22 540.38
R20648 A0.n29 A0.t13 540.375
R20649 A0.n6 A0.t19 491.64
R20650 A0.n6 A0.t36 491.64
R20651 A0.n6 A0.t45 491.64
R20652 A0.n6 A0.t32 491.64
R20653 A0.n1 A0.t5 491.64
R20654 A0.n1 A0.t16 491.64
R20655 A0.n1 A0.t4 491.64
R20656 A0.n1 A0.t21 491.64
R20657 A0.n16 A0.t8 485.221
R20658 A0.n13 A0.t20 485.221
R20659 A0.n24 A0.t33 485.221
R20660 A0.n14 A0.t34 367.928
R20661 A0.n11 A0.t43 367.928
R20662 A0.n22 A0.t39 367.928
R20663 A0.n17 A0.t38 367.928
R20664 A0.n3 A0.t26 367.928
R20665 A0.n27 A0.t28 343.827
R20666 A0.n32 A0.t0 312.599
R20667 A0.n35 A0.t37 247.428
R20668 A0.n34 A0.t18 247.428
R20669 A0.n33 A0.t15 247.428
R20670 A0.n32 A0.t2 247.428
R20671 A0.n27 A0.t40 237.787
R20672 A0.n36 A0.t35 229.754
R20673 A0.n28 A0.t6 227.356
R20674 A0.n18 A0.t10 227.356
R20675 A0.n4 A0.t24 227.356
R20676 A0.n15 A0.t7 224.478
R20677 A0.n12 A0.t14 224.478
R20678 A0.n23 A0.t17 224.478
R20679 A0.n14 A0.t3 213.688
R20680 A0.n11 A0.t11 213.688
R20681 A0.n22 A0.t23 213.688
R20682 A0.n17 A0.t42 213.688
R20683 A0.n3 A0.t25 213.688
R20684 A0 A0.n2 163.036
R20685 A0.n9 A0.n8 162.867
R20686 A0 A0.n36 162.409
R20687 A0.n19 A0.n18 160.439
R20688 A0.n5 A0.n4 160.439
R20689 A0.n29 A0.n28 160.433
R20690 A0.n7 A0.t30 139.78
R20691 A0.n7 A0.t9 139.78
R20692 A0.n7 A0.t1 139.78
R20693 A0.n7 A0.t12 139.78
R20694 A0.n0 A0.t29 139.78
R20695 A0.n0 A0.t44 139.78
R20696 A0.n0 A0.t31 139.78
R20697 A0.n0 A0.t41 139.78
R20698 A0.n18 A0.n17 94.4341
R20699 A0.n4 A0.n3 94.4341
R20700 A0.n36 A0.n35 91.5805
R20701 A0.n16 A0.n15 84.5046
R20702 A0.n13 A0.n12 84.5046
R20703 A0.n24 A0.n23 84.5046
R20704 A0.n15 A0.n14 72.3005
R20705 A0.n12 A0.n11 72.3005
R20706 A0.n23 A0.n22 72.3005
R20707 A0.n28 A0.n27 70.3341
R20708 A0.n33 A0.n32 65.1723
R20709 A0.n34 A0.n33 65.1723
R20710 A0.n35 A0.n34 65.1723
R20711 A0 A0.n16 61.0566
R20712 A0 A0.n13 61.0566
R20713 A0 A0.n24 61.0566
R20714 A0.n2 A0.n0 38.8368
R20715 A0.n8 A0.n7 38.6833
R20716 A0.n26 A0 33.5593
R20717 A0.n8 A0.n6 28.3986
R20718 A0.n2 A0.n1 28.2451
R20719 A0 A0.n10 18.1908
R20720 A0.n38 A0.n37 15.3483
R20721 A0.n26 A0.n25 13.1591
R20722 A0.n37 A0 12.5899
R20723 A0.n31 A0.n30 12.4105
R20724 A0.n10 A0.n9 9.00496
R20725 A0.n20 A0 6.24054
R20726 A0.n10 A0 3.87912
R20727 A0.n37 A0.n31 3.5777
R20728 A0 A0.n26 2.72912
R20729 A0.n21 A0 2.42219
R20730 A0.n25 A0.n21 2.42068
R20731 A0.n38 A0 1.65812
R20732 A0.n30 A0 1.32855
R20733 A0 A0.n29 0.905186
R20734 A0 A0.n19 0.900886
R20735 A0 A0.n5 0.89693
R20736 A0.n25 A0 0.282595
R20737 A0.n20 A0 0.244944
R20738 A0.n21 A0 0.244944
R20739 A0.n30 A0 0.0861742
R20740 A0.n39 A0.n38 0.063
R20741 A0.n9 A0 0.0590664
R20742 A0.n39 A0 0.0434293
R20743 A0 A0.n20 0.0373976
R20744 A0 A0.n39 0.0359167
R20745 A0.n31 A0 0.00999495
R20746 a_n17677_n15425.n0 a_n17677_n15425.n2 231.24
R20747 a_n17677_n15425.n1 a_n17677_n15425.n5 231.24
R20748 a_n17677_n15425.n0 a_n17677_n15425.n3 231.03
R20749 a_n17677_n15425.n1 a_n17677_n15425.n4 231.03
R20750 a_n17677_n15425.n6 a_n17677_n15425.n1 231.03
R20751 a_n17677_n15425.n2 a_n17677_n15425.t4 25.395
R20752 a_n17677_n15425.n2 a_n17677_n15425.t3 25.395
R20753 a_n17677_n15425.n3 a_n17677_n15425.t2 25.395
R20754 a_n17677_n15425.n3 a_n17677_n15425.t1 25.395
R20755 a_n17677_n15425.n4 a_n17677_n15425.t0 25.395
R20756 a_n17677_n15425.n4 a_n17677_n15425.t9 25.395
R20757 a_n17677_n15425.n5 a_n17677_n15425.t6 25.395
R20758 a_n17677_n15425.n5 a_n17677_n15425.t5 25.395
R20759 a_n17677_n15425.t8 a_n17677_n15425.n6 25.395
R20760 a_n17677_n15425.n6 a_n17677_n15425.t7 25.395
R20761 a_n17677_n15425.n1 a_n17677_n15425.n0 0.421553
R20762 OR8_0.NOT8_0.A0.n3 OR8_0.NOT8_0.A0.t7 394.37
R20763 OR8_0.NOT8_0.A0.n2 OR8_0.NOT8_0.A0.t10 291.829
R20764 OR8_0.NOT8_0.A0.n2 OR8_0.NOT8_0.A0.t8 291.829
R20765 OR8_0.NOT8_0.A0.n0 OR8_0.NOT8_0.A0.t4 256.425
R20766 OR8_0.NOT8_0.A0.n0 OR8_0.NOT8_0.A0.n5 231.24
R20767 OR8_0.NOT8_0.A0.n0 OR8_0.NOT8_0.A0.n6 231.03
R20768 OR8_0.NOT8_0.A0.n2 OR8_0.NOT8_0.A0.t9 221.72
R20769 OR8_0.NOT8_0.A0.n4 OR8_0.NOT8_0.A0.n1 66.4681
R20770 OR8_0.NOT8_0.A0.n3 OR8_0.NOT8_0.A0.n2 53.374
R20771 OR8_0.NOT8_0.A0.n4 OR8_0.NOT8_0.A0 28.3993
R20772 OR8_0.NOT8_0.A0.n6 OR8_0.NOT8_0.A0.t3 25.395
R20773 OR8_0.NOT8_0.A0.n6 OR8_0.NOT8_0.A0.t2 25.395
R20774 OR8_0.NOT8_0.A0.n5 OR8_0.NOT8_0.A0.t1 25.395
R20775 OR8_0.NOT8_0.A0.n5 OR8_0.NOT8_0.A0.t0 25.395
R20776 OR8_0.NOT8_0.A0.n1 OR8_0.NOT8_0.A0.t5 19.8005
R20777 OR8_0.NOT8_0.A0.n1 OR8_0.NOT8_0.A0.t6 19.8005
R20778 OR8_0.NOT8_0.A0 OR8_0.NOT8_0.A0.n3 1.27931
R20779 OR8_0.NOT8_0.A0 OR8_0.NOT8_0.A0.n0 0.355237
R20780 OR8_0.NOT8_0.A0 OR8_0.NOT8_0.A0.n4 0.293873
R20781 a_n17446_n8419.n0 a_n17446_n8419.t5 539.788
R20782 a_n17446_n8419.n1 a_n17446_n8419.t7 531.496
R20783 a_n17446_n8419.n0 a_n17446_n8419.t6 490.034
R20784 a_n17446_n8419.n5 a_n17446_n8419.t0 283.788
R20785 a_n17446_n8419.t1 a_n17446_n8419.n5 205.489
R20786 a_n17446_n8419.n2 a_n17446_n8419.t2 182.625
R20787 a_n17446_n8419.n3 a_n17446_n8419.t4 179.054
R20788 a_n17446_n8419.n2 a_n17446_n8419.t3 139.78
R20789 a_n17446_n8419.n4 a_n17446_n8419.n3 101.368
R20790 a_n17446_n8419.n5 a_n17446_n8419.n4 77.9135
R20791 a_n17446_n8419.n4 a_n17446_n8419.n1 76.1557
R20792 a_n17446_n8419.n1 a_n17446_n8419.n0 8.29297
R20793 a_n17446_n8419.n3 a_n17446_n8419.n2 3.57087
R20794 a_n17266_n8419.n2 a_n17266_n8419.n1 121.353
R20795 a_n17266_n8419.n3 a_n17266_n8419.n2 121.001
R20796 a_n17266_n8419.n2 a_n17266_n8419.n0 120.977
R20797 a_n17266_n8419.n1 a_n17266_n8419.t1 30.462
R20798 a_n17266_n8419.n1 a_n17266_n8419.t0 30.462
R20799 a_n17266_n8419.n0 a_n17266_n8419.t5 30.462
R20800 a_n17266_n8419.n0 a_n17266_n8419.t4 30.462
R20801 a_n17266_n8419.n3 a_n17266_n8419.t3 30.462
R20802 a_n17266_n8419.t2 a_n17266_n8419.n3 30.462
R20803 OR8_0.NOT8_0.A3.n2 OR8_0.NOT8_0.A3.t8 394.37
R20804 OR8_0.NOT8_0.A3.n1 OR8_0.NOT8_0.A3.t7 291.829
R20805 OR8_0.NOT8_0.A3.n1 OR8_0.NOT8_0.A3.t9 291.829
R20806 OR8_0.NOT8_0.A3.n0 OR8_0.NOT8_0.A3.t4 256.425
R20807 OR8_0.NOT8_0.A3.n0 OR8_0.NOT8_0.A3.n4 231.24
R20808 OR8_0.NOT8_0.A3.n0 OR8_0.NOT8_0.A3.n5 231.03
R20809 OR8_0.NOT8_0.A3.n1 OR8_0.NOT8_0.A3.t10 221.72
R20810 OR8_0.NOT8_0.A3.n0 OR8_0.NOT8_0.A3.n3 66.4895
R20811 OR8_0.NOT8_0.A3.n2 OR8_0.NOT8_0.A3.n1 53.374
R20812 OR8_0.NOT8_0.A3.n5 OR8_0.NOT8_0.A3.t3 25.395
R20813 OR8_0.NOT8_0.A3.n5 OR8_0.NOT8_0.A3.t2 25.395
R20814 OR8_0.NOT8_0.A3.n4 OR8_0.NOT8_0.A3.t1 25.395
R20815 OR8_0.NOT8_0.A3.n4 OR8_0.NOT8_0.A3.t5 25.395
R20816 OR8_0.NOT8_0.A3.n3 OR8_0.NOT8_0.A3.t6 19.8005
R20817 OR8_0.NOT8_0.A3.n3 OR8_0.NOT8_0.A3.t0 19.8005
R20818 OR8_0.NOT8_0.A3.n0 OR8_0.NOT8_0.A3 11.3387
R20819 OR8_0.NOT8_0.A3 OR8_0.NOT8_0.A3.n2 1.23583
R20820 right_shifter_0.S0.n1 right_shifter_0.S0.t5 1032.02
R20821 right_shifter_0.S0.n1 right_shifter_0.S0.t4 336.962
R20822 right_shifter_0.S0.n1 right_shifter_0.S0.t6 326.154
R20823 right_shifter_0.S0.n0 right_shifter_0.S0.t3 256.514
R20824 right_shifter_0.S0.n0 right_shifter_0.S0.n2 226.258
R20825 mux8_1.NAND4F_6.A right_shifter_0.S0.n1 162.952
R20826 right_shifter_0.S0.n0 right_shifter_0.S0.t0 83.7172
R20827 mux8_1.A7 right_shifter_0.S0.n0 55.0298
R20828 right_shifter_0.S0.n2 right_shifter_0.S0.t1 30.379
R20829 right_shifter_0.S0.n2 right_shifter_0.S0.t2 30.379
R20830 mux8_1.A7 mux8_1.NAND4F_6.A 13.4456
R20831 Y3.n2 Y3.t4 960.788
R20832 Y3.n0 Y3.t7 883.668
R20833 Y3.n1 Y3.t6 740.381
R20834 Y3.n0 Y3.t5 729.428
R20835 Y3.n4 Y3.t0 256.514
R20836 Y3.n5 Y3.n3 226.251
R20837 Y3 Y3.n2 162.025
R20838 Y3.n4 Y3.t1 83.7599
R20839 Y3.n1 Y3.n0 72.3005
R20840 Y3.n3 Y3.t2 30.379
R20841 Y3.n3 Y3.t3 30.379
R20842 Y3.n2 Y3.n1 16.7975
R20843 Y3.n5 Y3.n4 0.0323878
R20844 Y3.n5 Y3 0.0262937
R20845 Y3 Y3.n5 0.0126173
R20846 ZFLAG_0.nor4_0.Y.n6 ZFLAG_0.nor4_0.Y.t9 485.221
R20847 ZFLAG_0.nor4_0.Y.n4 ZFLAG_0.nor4_0.Y.t10 367.928
R20848 ZFLAG_0.nor4_0.Y.n5 ZFLAG_0.nor4_0.Y.t8 224.478
R20849 ZFLAG_0.nor4_0.Y.n4 ZFLAG_0.nor4_0.Y.t7 213.688
R20850 ZFLAG_0.nor4_0.Y ZFLAG_0.nor4_0.Y.t0 148.181
R20851 ZFLAG_0.nor4_0.Y ZFLAG_0.nor4_0.Y.n3 140.613
R20852 ZFLAG_0.nor4_0.Y.n6 ZFLAG_0.nor4_0.Y.n5 84.5046
R20853 ZFLAG_0.nor4_0.Y.n5 ZFLAG_0.nor4_0.Y.n4 72.3005
R20854 ZFLAG_0.nor4_0.Y.n2 ZFLAG_0.nor4_0.Y.n0 66.4372
R20855 ZFLAG_0.nor4_0.Y.n2 ZFLAG_0.nor4_0.Y.n1 66.3172
R20856 ZFLAG_0.nor4_0.Y ZFLAG_0.nor4_0.Y.n6 61.0566
R20857 ZFLAG_0.nor4_0.Y.n0 ZFLAG_0.nor4_0.Y.t6 19.8005
R20858 ZFLAG_0.nor4_0.Y.n0 ZFLAG_0.nor4_0.Y.t4 19.8005
R20859 ZFLAG_0.nor4_0.Y.n1 ZFLAG_0.nor4_0.Y.t3 19.8005
R20860 ZFLAG_0.nor4_0.Y.n1 ZFLAG_0.nor4_0.Y.t5 19.8005
R20861 ZFLAG_0.nor4_0.Y.n3 ZFLAG_0.nor4_0.Y.t1 7.59513
R20862 ZFLAG_0.nor4_0.Y.n3 ZFLAG_0.nor4_0.Y.t2 7.59513
R20863 ZFLAG_0.nor4_0.Y ZFLAG_0.nor4_0.Y.n2 0.61307
R20864 B5.n6 B5.t27 491.64
R20865 B5.n5 B5.t21 491.64
R20866 B5.n4 B5.t2 491.64
R20867 B5.n3 B5.t33 491.64
R20868 B5.n23 B5.t7 491.64
R20869 B5.n22 B5.t22 491.64
R20870 B5.n21 B5.t4 491.64
R20871 B5.n20 B5.t32 491.64
R20872 B5.n10 B5.t6 485.443
R20873 B5.n27 B5.t16 394.37
R20874 B5.n31 B5.t28 394.37
R20875 B5.n1 B5.t3 394.37
R20876 B5.n13 B5.t13 379.173
R20877 B5.n8 B5.t15 343.827
R20878 B5.n14 B5.t5 312.599
R20879 B5.n26 B5.t25 291.829
R20880 B5.n26 B5.t24 291.829
R20881 B5.n30 B5.t10 291.829
R20882 B5.n30 B5.t30 291.829
R20883 B5.n0 B5.t18 291.829
R20884 B5.n0 B5.t14 291.829
R20885 B5.n7 B5.t23 255.588
R20886 B5.n24 B5.t26 255.588
R20887 B5.n14 B5.t34 247.428
R20888 B5.n15 B5.t31 247.428
R20889 B5.n16 B5.t20 247.428
R20890 B5.n13 B5.t17 247.428
R20891 B5.n8 B5.t29 237.787
R20892 B5.n9 B5.t1 224.478
R20893 B5.n26 B5.t0 221.72
R20894 B5.n30 B5.t12 221.72
R20895 B5.n0 B5.t11 221.72
R20896 B5.n20 B5.n19 209.407
R20897 B5.n3 B5.n2 209.19
R20898 B5 B5.n17 162.139
R20899 B5.n2 B5.t19 139.78
R20900 B5.n2 B5.t9 139.78
R20901 B5.n2 B5.t36 139.78
R20902 B5.n19 B5.t37 139.78
R20903 B5.n19 B5.t8 139.78
R20904 B5.n19 B5.t35 139.78
R20905 B5.n10 B5.n9 83.8438
R20906 B5.n16 B5.n15 65.1723
R20907 B5.n15 B5.n14 65.1723
R20908 B5 B5.n10 61.0461
R20909 B5.n27 B5.n26 53.374
R20910 B5.n31 B5.n30 53.374
R20911 B5.n1 B5.n0 53.374
R20912 B5.n9 B5.n8 48.2005
R20913 B5.n12 B5 41.7905
R20914 B5.n17 B5.n16 33.2653
R20915 B5.n17 B5.n13 31.9075
R20916 B5 B5.n24 27.4136
R20917 B5.n5 B5.n4 17.8661
R20918 B5.n4 B5.n3 17.8661
R20919 B5.n21 B5.n20 17.8661
R20920 B5.n22 B5.n21 17.8661
R20921 B5.n6 B5.n5 17.1217
R20922 B5.n23 B5.n22 17.1217
R20923 B5.n34 B5.n33 14.1808
R20924 B5.n18 B5 12.5696
R20925 B5.n25 B5 12.5587
R20926 B5.n29 B5.n28 12.5047
R20927 B5.n12 B5.n11 12.4162
R20928 B5.n33 B5.n32 12.4105
R20929 B5 B5.n7 11.1665
R20930 B5.n29 B5.n25 10.0354
R20931 B5.n25 B5.n18 7.8666
R20932 B5.n18 B5 5.13276
R20933 B5.n33 B5.n29 2.5871
R20934 B5.n7 B5.n6 1.8615
R20935 B5.n24 B5.n23 1.8615
R20936 B5.n11 B5 1.31161
R20937 B5.n28 B5.n27 1.23221
R20938 B5.n34 B5.n1 0.762507
R20939 B5.n32 B5.n31 0.759495
R20940 B5.n32 B5 0.0592349
R20941 B5.n11 B5 0.0577917
R20942 B5 B5.n34 0.0562229
R20943 B5.n28 B5 0.0476014
R20944 B5 B5.n12 0.00311111
R20945 a_7548_n16422.t0 a_7548_n16422.t1 9.9005
R20946 a_7644_n16422.t0 a_7644_n16422.t1 9.9005
R20947 B3.n32 B3.t31 540.38
R20948 B3.n39 B3.t17 540.38
R20949 B3.n28 B3.t15 491.64
R20950 B3.n27 B3.t47 491.64
R20951 B3.n26 B3.t38 491.64
R20952 B3.n25 B3.t26 491.64
R20953 B3.n20 B3.t13 491.64
R20954 B3.n19 B3.t35 491.64
R20955 B3.n18 B3.t12 491.64
R20956 B3.n17 B3.t49 491.64
R20957 B3.n47 B3.t7 485.443
R20958 B3.n35 B3.t48 485.221
R20959 B3.n42 B3.t41 485.221
R20960 B3.n13 B3.t27 394.37
R20961 B3.n9 B3.t45 394.37
R20962 B3.n6 B3.t6 394.37
R20963 B3.n0 B3.t16 379.173
R20964 B3.n30 B3.t30 367.928
R20965 B3.n33 B3.t5 367.928
R20966 B3.n40 B3.t52 367.928
R20967 B3.n37 B3.t51 367.928
R20968 B3.n45 B3.t18 343.827
R20969 B3.n1 B3.t8 312.599
R20970 B3.n12 B3.t39 291.829
R20971 B3.n12 B3.t37 291.829
R20972 B3.n8 B3.t9 291.829
R20973 B3.n8 B3.t36 291.829
R20974 B3.n5 B3.t24 291.829
R20975 B3.n5 B3.t23 291.829
R20976 B3.n29 B3.t11 255.588
R20977 B3.n21 B3.t40 255.588
R20978 B3.n1 B3.t46 247.428
R20979 B3.n2 B3.t42 247.428
R20980 B3.n3 B3.t25 247.428
R20981 B3.n0 B3.t21 247.428
R20982 B3.n45 B3.t22 237.787
R20983 B3.n31 B3.t4 227.356
R20984 B3.n38 B3.t50 227.356
R20985 B3.n46 B3.t44 224.478
R20986 B3.n34 B3.t43 224.478
R20987 B3.n41 B3.t29 224.478
R20988 B3.n12 B3.t1 221.72
R20989 B3.n8 B3.t10 221.72
R20990 B3.n5 B3.t19 221.72
R20991 B3.n30 B3.t28 213.688
R20992 B3.n33 B3.t2 213.688
R20993 B3.n40 B3.t33 213.688
R20994 B3.n37 B3.t32 213.688
R20995 B3.n17 B3.n16 209.407
R20996 B3.n25 B3.n24 209.19
R20997 B3 B3.n4 162.139
R20998 B3.n32 B3.n31 160.439
R20999 B3.n39 B3.n38 160.439
R21000 B3.n24 B3.t0 139.78
R21001 B3.n24 B3.t14 139.78
R21002 B3.n24 B3.t34 139.78
R21003 B3.n16 B3.t3 139.78
R21004 B3.n16 B3.t20 139.78
R21005 B3.n16 B3.t53 139.78
R21006 B3.n31 B3.n30 94.4341
R21007 B3.n38 B3.n37 94.4341
R21008 B3.n35 B3.n34 84.5046
R21009 B3.n42 B3.n41 84.5046
R21010 B3.n47 B3.n46 83.8438
R21011 B3.n34 B3.n33 72.3005
R21012 B3.n41 B3.n40 72.3005
R21013 B3.n3 B3.n2 65.1723
R21014 B3.n2 B3.n1 65.1723
R21015 B3 B3.n35 61.0566
R21016 B3 B3.n42 61.0566
R21017 B3 B3.n47 61.0461
R21018 B3.n13 B3.n12 53.374
R21019 B3.n9 B3.n8 53.374
R21020 B3.n6 B3.n5 53.374
R21021 B3.n46 B3.n45 48.2005
R21022 B3.n44 B3 36.3623
R21023 B3.n4 B3.n3 33.2653
R21024 B3.n4 B3.n0 31.9075
R21025 B3 B3.n21 27.4136
R21026 B3.n27 B3.n26 17.8661
R21027 B3.n26 B3.n25 17.8661
R21028 B3.n18 B3.n17 17.8661
R21029 B3.n19 B3.n18 17.8661
R21030 B3.n28 B3.n27 17.1217
R21031 B3.n20 B3.n19 17.1217
R21032 B3.n11 B3.n7 14.4293
R21033 B3.n23 B3 12.8136
R21034 B3.n15 B3.n14 12.5652
R21035 B3.n22 B3 12.4808
R21036 B3.n49 B3.n48 12.4105
R21037 B3.n11 B3.n10 12.4105
R21038 B3 B3.n29 11.1665
R21039 B3.n22 B3.n15 8.05642
R21040 B3.n23 B3.n22 7.04771
R21041 B3.n44 B3.n43 6.01478
R21042 B3 B3.n44 5.72519
R21043 B3.n50 B3.n23 5.15688
R21044 B3.n36 B3 3.59317
R21045 B3.n43 B3 3.54887
R21046 B3.n36 B3 3.32934
R21047 B3.n43 B3 3.3031
R21048 B3.n15 B3.n11 2.77827
R21049 B3.n29 B3.n28 1.8615
R21050 B3.n21 B3.n20 1.8615
R21051 B3 B3.n36 1.2542
R21052 B3.n14 B3.n13 1.22315
R21053 B3.n48 B3 1.16057
R21054 B3 B3.n32 0.900886
R21055 B3 B3.n39 0.900886
R21056 B3.n7 B3.n6 0.764013
R21057 B3.n10 B3.n9 0.758742
R21058 B3.n43 B3 0.178278
R21059 B3.n48 B3 0.151542
R21060 B3.n14 B3 0.0602826
R21061 B3.n10 B3 0.059988
R21062 B3.n7 B3 0.0547169
R21063 B3 B3.n50 0.0311806
R21064 B3.n50 B3.n49 0.024
R21065 B3.n49 B3 0.00393902
R21066 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t19 491.64
R21067 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t14 491.64
R21068 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t22 491.64
R21069 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t20 491.64
R21070 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t15 485.221
R21071 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t18 367.928
R21072 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t13 255.588
R21073 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t16 224.478
R21074 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t17 213.688
R21075 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n18 209.19
R21076 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t12 139.78
R21077 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t21 139.78
R21078 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t23 139.78
R21079 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n1 120.999
R21080 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n0 120.999
R21081 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n13 104.489
R21082 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 103.258
R21083 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n3 92.5005
R21084 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n8 86.2638
R21085 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n9 85.8873
R21086 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n6 85.724
R21087 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n16 84.5046
R21088 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n14 84.0545
R21089 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n11 75.0672
R21090 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n8 75.0672
R21091 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n10 73.1255
R21092 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n6 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n5 73.1255
R21093 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n8 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n7 73.1255
R21094 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n15 72.3005
R21095 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n6 68.8946
R21096 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n17 60.9816
R21097 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n4 41.9827
R21098 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t3 30.462
R21099 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t10 30.462
R21100 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t9 30.462
R21101 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t8 30.462
R21102 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t1 30.462
R21103 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t5 30.462
R21104 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n2 28.124
R21105 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n19 17.8661
R21106 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n20 17.8661
R21107 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n21 17.1217
R21108 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n23 15.6329
R21109 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t4 11.8205
R21110 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t7 11.8205
R21111 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t6 11.8205
R21112 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t11 11.8205
R21113 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t2 11.8205
R21114 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t0 11.8205
R21115 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 10.8165
R21116 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n12 9.3005
R21117 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n24 2.50602
R21118 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n22 1.8615
R21119 a_n10786_3190.n2 a_n10786_3190.n1 121.353
R21120 a_n10786_3190.n2 a_n10786_3190.n0 121.353
R21121 a_n10786_3190.n3 a_n10786_3190.n2 121.001
R21122 a_n10786_3190.n1 a_n10786_3190.t0 30.462
R21123 a_n10786_3190.n1 a_n10786_3190.t1 30.462
R21124 a_n10786_3190.n0 a_n10786_3190.t4 30.462
R21125 a_n10786_3190.n0 a_n10786_3190.t5 30.462
R21126 a_n10786_3190.n3 a_n10786_3190.t3 30.462
R21127 a_n10786_3190.t2 a_n10786_3190.n3 30.462
R21128 mux8_7.NAND4F_0.C.n6 mux8_7.NAND4F_0.C.t15 978.795
R21129 mux8_7.NAND4F_0.C.n4 mux8_7.NAND4F_0.C.t11 978.795
R21130 mux8_7.NAND4F_0.C.n11 mux8_7.NAND4F_0.C.t8 978.795
R21131 mux8_7.NAND4F_0.C.n2 mux8_7.NAND4F_0.C.t12 978.795
R21132 mux8_7.NAND4F_0.C.n5 mux8_7.NAND4F_0.C.t10 308.481
R21133 mux8_7.NAND4F_0.C.n5 mux8_7.NAND4F_0.C.t9 308.481
R21134 mux8_7.NAND4F_0.C.n3 mux8_7.NAND4F_0.C.t14 308.481
R21135 mux8_7.NAND4F_0.C.n3 mux8_7.NAND4F_0.C.t13 308.481
R21136 mux8_7.NAND4F_0.C.n10 mux8_7.NAND4F_0.C.t4 308.481
R21137 mux8_7.NAND4F_0.C.n10 mux8_7.NAND4F_0.C.t5 308.481
R21138 mux8_7.NAND4F_0.C.n1 mux8_7.NAND4F_0.C.t6 308.481
R21139 mux8_7.NAND4F_0.C.n1 mux8_7.NAND4F_0.C.t7 308.481
R21140 mux8_7.NAND4F_0.C.n0 mux8_7.NAND4F_0.C.t1 256.514
R21141 mux8_7.NAND4F_0.C.n0 mux8_7.NAND4F_0.C.n8 226.258
R21142 mux8_7.NAND4F_0.C mux8_7.NAND4F_0.C.n6 161.856
R21143 mux8_7.NAND4F_0.C mux8_7.NAND4F_0.C.n4 161.847
R21144 mux8_7.NAND4F_0.C mux8_7.NAND4F_0.C.n11 161.84
R21145 mux8_7.NAND4F_0.C mux8_7.NAND4F_0.C.n2 161.831
R21146 mux8_7.NAND4F_0.C.n0 mux8_7.NAND4F_0.C.t0 83.7172
R21147 mux8_7.NAND4F_0.C.n8 mux8_7.NAND4F_0.C.t3 30.379
R21148 mux8_7.NAND4F_0.C.n8 mux8_7.NAND4F_0.C.t2 30.379
R21149 mux8_7.NAND4F_0.C.n9 mux8_7.NAND4F_0.C.n0 13.5186
R21150 mux8_7.NAND4F_0.C mux8_7.NAND4F_0.C.n12 13.0862
R21151 mux8_7.NAND4F_0.C.n7 mux8_7.NAND4F_0.C 13.0435
R21152 mux8_7.NAND4F_0.C.n12 mux8_7.NAND4F_0.C 12.4135
R21153 mux8_7.NAND4F_0.C.n7 mux8_7.NAND4F_0.C 12.4105
R21154 mux8_7.NAND4F_0.C.n6 mux8_7.NAND4F_0.C.n5 11.0463
R21155 mux8_7.NAND4F_0.C.n4 mux8_7.NAND4F_0.C.n3 11.0463
R21156 mux8_7.NAND4F_0.C.n11 mux8_7.NAND4F_0.C.n10 11.0463
R21157 mux8_7.NAND4F_0.C.n2 mux8_7.NAND4F_0.C.n1 11.0463
R21158 mux8_7.NAND4F_0.C.n12 mux8_7.NAND4F_0.C.n9 3.46056
R21159 mux8_7.NAND4F_0.C.n9 mux8_7.NAND4F_0.C.n7 1.8134
R21160 mux8_7.NAND4F_1.Y.n2 mux8_7.NAND4F_1.Y.t11 978.795
R21161 mux8_7.NAND4F_1.Y.n1 mux8_7.NAND4F_1.Y.t9 308.481
R21162 mux8_7.NAND4F_1.Y.n1 mux8_7.NAND4F_1.Y.t10 308.481
R21163 mux8_7.NAND4F_1.Y.n0 mux8_7.NAND4F_1.Y.n3 187.373
R21164 mux8_7.NAND4F_1.Y.n0 mux8_7.NAND4F_1.Y.n4 187.192
R21165 mux8_7.NAND4F_1.Y.n0 mux8_7.NAND4F_1.Y.n5 187.192
R21166 mux8_7.NAND4F_1.Y.n7 mux8_7.NAND4F_1.Y.n6 187.192
R21167 mux8_7.NAND4F_1.Y mux8_7.NAND4F_1.Y.n2 161.84
R21168 mux8_7.NAND4F_1.Y mux8_7.NAND4F_1.Y.t6 23.4335
R21169 mux8_7.NAND4F_1.Y.n3 mux8_7.NAND4F_1.Y.t1 20.1899
R21170 mux8_7.NAND4F_1.Y.n3 mux8_7.NAND4F_1.Y.t0 20.1899
R21171 mux8_7.NAND4F_1.Y.n4 mux8_7.NAND4F_1.Y.t3 20.1899
R21172 mux8_7.NAND4F_1.Y.n4 mux8_7.NAND4F_1.Y.t2 20.1899
R21173 mux8_7.NAND4F_1.Y.n5 mux8_7.NAND4F_1.Y.t8 20.1899
R21174 mux8_7.NAND4F_1.Y.n5 mux8_7.NAND4F_1.Y.t7 20.1899
R21175 mux8_7.NAND4F_1.Y.n6 mux8_7.NAND4F_1.Y.t4 20.1899
R21176 mux8_7.NAND4F_1.Y.n6 mux8_7.NAND4F_1.Y.t5 20.1899
R21177 mux8_7.NAND4F_1.Y.n2 mux8_7.NAND4F_1.Y.n1 11.0463
R21178 mux8_7.NAND4F_1.Y mux8_7.NAND4F_1.Y.n7 0.527586
R21179 mux8_7.NAND4F_1.Y.n7 mux8_7.NAND4F_1.Y.n0 0.358709
R21180 MULT_0.4bit_ADDER_0.B2.t1 MULT_0.4bit_ADDER_0.B2.n0 83.7599
R21181 MULT_0.4bit_ADDER_0.B2.n0 MULT_0.4bit_ADDER_0.B2.n2 0.0323878
R21182 MULT_0.4bit_ADDER_0.B2.n2 MULT_0.4bit_ADDER_0.B2 8.92851
R21183 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_0.B2.n14 0.0198089
R21184 MULT_0.4bit_ADDER_0.B2.n14 MULT_0.4bit_ADDER_0.B2 0.0116789
R21185 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_0.B2.n14 0.0213333
R21186 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_0.B2.n9 0.840348
R21187 MULT_0.4bit_ADDER_0.B2.n13 MULT_0.4bit_ADDER_0.B2.n9 10.8165
R21188 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_0.B2.n13 0.0755
R21189 MULT_0.4bit_ADDER_0.B2.n10 MULT_0.4bit_ADDER_0.B2.n13 60.9816
R21190 MULT_0.4bit_ADDER_0.B2.n10 MULT_0.4bit_ADDER_0.B2.n12 84.5046
R21191 MULT_0.4bit_ADDER_0.B2.n12 MULT_0.4bit_ADDER_0.B2.t5 224.478
R21192 MULT_0.4bit_ADDER_0.B2.n12 MULT_0.4bit_ADDER_0.B2.n11 72.3005
R21193 MULT_0.4bit_ADDER_0.B2.n11 MULT_0.4bit_ADDER_0.B2.t11 213.688
R21194 MULT_0.4bit_ADDER_0.B2.n11 MULT_0.4bit_ADDER_0.B2.t12 367.928
R21195 MULT_0.4bit_ADDER_0.B2.n10 MULT_0.4bit_ADDER_0.B2.t7 485.221
R21196 MULT_0.4bit_ADDER_0.B2.n9 MULT_0.4bit_ADDER_0.B2 103.258
R21197 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_0.B2.n8 15.6329
R21198 MULT_0.4bit_ADDER_0.B2.n8 MULT_0.4bit_ADDER_0.B2.n7 1.8615
R21199 MULT_0.4bit_ADDER_0.B2.n7 MULT_0.4bit_ADDER_0.B2.n6 17.1217
R21200 MULT_0.4bit_ADDER_0.B2.n6 MULT_0.4bit_ADDER_0.B2.n5 17.8661
R21201 MULT_0.4bit_ADDER_0.B2.n5 MULT_0.4bit_ADDER_0.B2.n4 17.8661
R21202 MULT_0.4bit_ADDER_0.B2.t6 MULT_0.4bit_ADDER_0.B2.n8 255.588
R21203 MULT_0.4bit_ADDER_0.B2.n7 MULT_0.4bit_ADDER_0.B2.t8 491.64
R21204 MULT_0.4bit_ADDER_0.B2.n6 MULT_0.4bit_ADDER_0.B2.t15 491.64
R21205 MULT_0.4bit_ADDER_0.B2.n5 MULT_0.4bit_ADDER_0.B2.t14 491.64
R21206 MULT_0.4bit_ADDER_0.B2.n4 MULT_0.4bit_ADDER_0.B2.t13 491.64
R21207 MULT_0.4bit_ADDER_0.B2.n3 MULT_0.4bit_ADDER_0.B2.n4 209.19
R21208 MULT_0.4bit_ADDER_0.B2.t4 MULT_0.4bit_ADDER_0.B2.n3 139.78
R21209 MULT_0.4bit_ADDER_0.B2.t9 MULT_0.4bit_ADDER_0.B2.n3 139.78
R21210 MULT_0.4bit_ADDER_0.B2.t10 MULT_0.4bit_ADDER_0.B2.n3 139.78
R21211 MULT_0.4bit_ADDER_0.B2.n1 MULT_0.4bit_ADDER_0.B2.n2 226.251
R21212 MULT_0.4bit_ADDER_0.B2.t3 MULT_0.4bit_ADDER_0.B2.n1 30.379
R21213 MULT_0.4bit_ADDER_0.B2.n1 MULT_0.4bit_ADDER_0.B2.t2 30.379
R21214 MULT_0.4bit_ADDER_0.B2.n0 MULT_0.4bit_ADDER_0.B2.t0 256.514
R21215 a_n16822_3164.n0 a_n16822_3164.t7 539.788
R21216 a_n16822_3164.n1 a_n16822_3164.t5 531.496
R21217 a_n16822_3164.n0 a_n16822_3164.t3 490.034
R21218 a_n16822_3164.n5 a_n16822_3164.t0 283.788
R21219 a_n16822_3164.t1 a_n16822_3164.n5 205.489
R21220 a_n16822_3164.n2 a_n16822_3164.t6 182.625
R21221 a_n16822_3164.n3 a_n16822_3164.t4 179.054
R21222 a_n16822_3164.n2 a_n16822_3164.t2 139.78
R21223 a_n16822_3164.n4 a_n16822_3164.n3 101.368
R21224 a_n16822_3164.n5 a_n16822_3164.n4 77.9135
R21225 a_n16822_3164.n4 a_n16822_3164.n1 76.1557
R21226 a_n16822_3164.n1 a_n16822_3164.n0 8.29297
R21227 a_n16822_3164.n3 a_n16822_3164.n2 3.57087
R21228 a_n16792_3190.n2 a_n16792_3190.n0 121.353
R21229 a_n16792_3190.n2 a_n16792_3190.n1 121.001
R21230 a_n16792_3190.n3 a_n16792_3190.n2 120.977
R21231 a_n16792_3190.n1 a_n16792_3190.t3 30.462
R21232 a_n16792_3190.n1 a_n16792_3190.t1 30.462
R21233 a_n16792_3190.n0 a_n16792_3190.t5 30.462
R21234 a_n16792_3190.n0 a_n16792_3190.t4 30.462
R21235 a_n16792_3190.n3 a_n16792_3190.t2 30.462
R21236 a_n16792_3190.t0 a_n16792_3190.n3 30.462
R21237 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t14 491.64
R21238 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t12 491.64
R21239 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t13 491.64
R21240 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t22 491.64
R21241 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t18 485.221
R21242 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t19 367.928
R21243 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t16 255.588
R21244 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t20 224.478
R21245 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t21 213.688
R21246 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n18 209.19
R21247 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t17 139.78
R21248 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t23 139.78
R21249 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t15 139.78
R21250 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n1 120.999
R21251 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n0 120.999
R21252 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n13 104.489
R21253 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 103.258
R21254 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n3 92.5005
R21255 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n8 86.2638
R21256 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n9 85.8873
R21257 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n6 85.724
R21258 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n16 84.5046
R21259 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n14 84.0545
R21260 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n11 75.0672
R21261 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n8 75.0672
R21262 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n10 73.1255
R21263 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n8 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n7 73.1255
R21264 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n6 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n5 73.1255
R21265 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n15 72.3005
R21266 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n6 68.8946
R21267 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n17 60.9816
R21268 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n4 41.9827
R21269 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t0 30.462
R21270 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t8 30.462
R21271 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t7 30.462
R21272 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t6 30.462
R21273 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t1 30.462
R21274 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t2 30.462
R21275 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n2 28.124
R21276 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n19 17.8661
R21277 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n20 17.8661
R21278 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n21 17.1217
R21279 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n23 15.6329
R21280 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t4 11.8205
R21281 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t5 11.8205
R21282 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t10 11.8205
R21283 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t11 11.8205
R21284 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t3 11.8205
R21285 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t9 11.8205
R21286 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 10.8165
R21287 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n12 9.3005
R21288 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n24 2.50602
R21289 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n22 1.8615
R21290 a_n13372_1406.n0 a_n13372_1406.t3 539.788
R21291 a_n13372_1406.n1 a_n13372_1406.t5 531.496
R21292 a_n13372_1406.n0 a_n13372_1406.t6 490.034
R21293 a_n13372_1406.n5 a_n13372_1406.t0 283.788
R21294 a_n13372_1406.t1 a_n13372_1406.n5 205.489
R21295 a_n13372_1406.n2 a_n13372_1406.t7 182.625
R21296 a_n13372_1406.n3 a_n13372_1406.t2 179.054
R21297 a_n13372_1406.n2 a_n13372_1406.t4 139.78
R21298 a_n13372_1406.n4 a_n13372_1406.n3 101.368
R21299 a_n13372_1406.n5 a_n13372_1406.n4 77.9135
R21300 a_n13372_1406.n4 a_n13372_1406.n1 76.1557
R21301 a_n13372_1406.n1 a_n13372_1406.n0 8.29297
R21302 a_n13372_1406.n3 a_n13372_1406.n2 3.57087
R21303 a_7452_n20950.t0 a_7452_n20950.t1 9.9005
R21304 a_7548_n20950.t0 a_7548_n20950.t1 9.9005
R21305 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t10 540.38
R21306 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t9 367.928
R21307 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n5 227.526
R21308 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t8 227.356
R21309 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n6 227.266
R21310 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n4 227.266
R21311 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t7 213.688
R21312 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n2 160.439
R21313 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n1 94.4341
R21314 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t5 42.7944
R21315 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t3 30.379
R21316 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t0 30.379
R21317 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t6 30.379
R21318 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t4 30.379
R21319 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t1 30.379
R21320 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.t2 30.379
R21321 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n0 13.4358
R21322 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B.n3 0.821842
R21323 mux8_0.NAND4F_4.Y.n6 mux8_0.NAND4F_4.Y.t11 1032.02
R21324 mux8_0.NAND4F_4.Y.n6 mux8_0.NAND4F_4.Y.t9 336.962
R21325 mux8_0.NAND4F_4.Y.n6 mux8_0.NAND4F_4.Y.t10 326.154
R21326 mux8_0.NAND4F_4.Y.n0 mux8_0.NAND4F_4.Y.n1 187.373
R21327 mux8_0.NAND4F_4.Y.n0 mux8_0.NAND4F_4.Y.n2 187.192
R21328 mux8_0.NAND4F_4.Y.n0 mux8_0.NAND4F_4.Y.n3 187.192
R21329 mux8_0.NAND4F_4.Y.n5 mux8_0.NAND4F_4.Y.n4 187.192
R21330 mux8_0.NAND4F_4.Y mux8_0.NAND4F_4.Y.n6 162.942
R21331 mux8_0.NAND4F_4.Y.n7 mux8_0.NAND4F_4.Y 24.5377
R21332 mux8_0.NAND4F_4.Y.n7 mux8_0.NAND4F_4.Y.t6 22.6141
R21333 mux8_0.NAND4F_4.Y.n1 mux8_0.NAND4F_4.Y.t2 20.1899
R21334 mux8_0.NAND4F_4.Y.n1 mux8_0.NAND4F_4.Y.t3 20.1899
R21335 mux8_0.NAND4F_4.Y.n2 mux8_0.NAND4F_4.Y.t8 20.1899
R21336 mux8_0.NAND4F_4.Y.n2 mux8_0.NAND4F_4.Y.t7 20.1899
R21337 mux8_0.NAND4F_4.Y.n3 mux8_0.NAND4F_4.Y.t0 20.1899
R21338 mux8_0.NAND4F_4.Y.n3 mux8_0.NAND4F_4.Y.t1 20.1899
R21339 mux8_0.NAND4F_4.Y.n4 mux8_0.NAND4F_4.Y.t4 20.1899
R21340 mux8_0.NAND4F_4.Y.n4 mux8_0.NAND4F_4.Y.t5 20.1899
R21341 mux8_0.NAND4F_4.Y mux8_0.NAND4F_4.Y.n7 0.894894
R21342 mux8_0.NAND4F_4.Y mux8_0.NAND4F_4.Y.n5 0.452586
R21343 mux8_0.NAND4F_4.Y.n5 mux8_0.NAND4F_4.Y.n0 0.358709
R21344 a_n14751_2026.n1 a_n14751_2026.n5 81.2978
R21345 a_n14751_2026.n1 a_n14751_2026.n6 81.1637
R21346 a_n14751_2026.n0 a_n14751_2026.n4 81.1637
R21347 a_n14751_2026.n0 a_n14751_2026.n3 81.1637
R21348 a_n14751_2026.n7 a_n14751_2026.n1 81.1637
R21349 a_n14751_2026.n0 a_n14751_2026.n2 80.9213
R21350 a_n14751_2026.n5 a_n14751_2026.t7 11.8205
R21351 a_n14751_2026.n5 a_n14751_2026.t8 11.8205
R21352 a_n14751_2026.n6 a_n14751_2026.t3 11.8205
R21353 a_n14751_2026.n6 a_n14751_2026.t6 11.8205
R21354 a_n14751_2026.n4 a_n14751_2026.t2 11.8205
R21355 a_n14751_2026.n4 a_n14751_2026.t1 11.8205
R21356 a_n14751_2026.n3 a_n14751_2026.t9 11.8205
R21357 a_n14751_2026.n3 a_n14751_2026.t0 11.8205
R21358 a_n14751_2026.n2 a_n14751_2026.t11 11.8205
R21359 a_n14751_2026.n2 a_n14751_2026.t10 11.8205
R21360 a_n14751_2026.n7 a_n14751_2026.t4 11.8205
R21361 a_n14751_2026.t5 a_n14751_2026.n7 11.8205
R21362 a_n14751_2026.n1 a_n14751_2026.n0 0.402735
R21363 mux8_2.NAND4F_7.Y.n2 mux8_2.NAND4F_7.Y.t10 1388.16
R21364 mux8_2.NAND4F_7.Y.n2 mux8_2.NAND4F_7.Y.t9 350.839
R21365 mux8_2.NAND4F_7.Y.n3 mux8_2.NAND4F_7.Y.t11 308.481
R21366 mux8_2.NAND4F_7.Y.n1 mux8_2.NAND4F_7.Y.n4 187.373
R21367 mux8_2.NAND4F_7.Y.n1 mux8_2.NAND4F_7.Y.n5 187.192
R21368 mux8_2.NAND4F_7.Y.n1 mux8_2.NAND4F_7.Y.n6 187.192
R21369 mux8_2.NAND4F_7.Y.n0 mux8_2.NAND4F_7.Y.n7 187.192
R21370 mux8_2.NAND4F_7.Y mux8_2.NAND4F_7.Y.n3 161.492
R21371 mux8_2.NAND4F_7.Y.n3 mux8_2.NAND4F_7.Y.n2 27.752
R21372 mux8_2.NAND4F_7.Y mux8_2.NAND4F_7.Y.t3 23.5642
R21373 mux8_2.NAND4F_7.Y.n4 mux8_2.NAND4F_7.Y.t0 20.1899
R21374 mux8_2.NAND4F_7.Y.n4 mux8_2.NAND4F_7.Y.t1 20.1899
R21375 mux8_2.NAND4F_7.Y.n5 mux8_2.NAND4F_7.Y.t8 20.1899
R21376 mux8_2.NAND4F_7.Y.n5 mux8_2.NAND4F_7.Y.t7 20.1899
R21377 mux8_2.NAND4F_7.Y.n6 mux8_2.NAND4F_7.Y.t5 20.1899
R21378 mux8_2.NAND4F_7.Y.n6 mux8_2.NAND4F_7.Y.t6 20.1899
R21379 mux8_2.NAND4F_7.Y.n7 mux8_2.NAND4F_7.Y.t2 20.1899
R21380 mux8_2.NAND4F_7.Y.n7 mux8_2.NAND4F_7.Y.t4 20.1899
R21381 mux8_2.NAND4F_7.Y mux8_2.NAND4F_7.Y.n0 0.472662
R21382 mux8_2.NAND4F_7.Y.n0 mux8_2.NAND4F_7.Y.n1 0.358709
R21383 mux8_2.NAND4F_9.Y.n1 mux8_2.NAND4F_9.Y.t12 312.599
R21384 mux8_2.NAND4F_9.Y.n4 mux8_2.NAND4F_9.Y.t13 247.428
R21385 mux8_2.NAND4F_9.Y.n1 mux8_2.NAND4F_9.Y.t11 247.428
R21386 mux8_2.NAND4F_9.Y.n2 mux8_2.NAND4F_9.Y.t10 247.428
R21387 mux8_2.NAND4F_9.Y.n3 mux8_2.NAND4F_9.Y.t9 247.428
R21388 mux8_2.NAND4F_9.Y.n5 mux8_2.NAND4F_9.Y.t14 229.754
R21389 mux8_2.NAND4F_9.Y.n0 mux8_2.NAND4F_9.Y.n6 187.373
R21390 mux8_2.NAND4F_9.Y.n0 mux8_2.NAND4F_9.Y.n7 187.192
R21391 mux8_2.NAND4F_9.Y.n0 mux8_2.NAND4F_9.Y.n8 187.192
R21392 mux8_2.NAND4F_9.Y.n10 mux8_2.NAND4F_9.Y.n9 187.192
R21393 mux8_2.NAND4F_9.Y mux8_2.NAND4F_9.Y.n5 162.275
R21394 mux8_2.NAND4F_9.Y.n5 mux8_2.NAND4F_9.Y.n4 91.5805
R21395 mux8_2.NAND4F_9.Y.n2 mux8_2.NAND4F_9.Y.n1 65.1723
R21396 mux8_2.NAND4F_9.Y.n3 mux8_2.NAND4F_9.Y.n2 65.1723
R21397 mux8_2.NAND4F_9.Y.n4 mux8_2.NAND4F_9.Y.n3 65.1723
R21398 mux8_2.NAND4F_9.Y mux8_2.NAND4F_9.Y.t5 22.6141
R21399 mux8_2.NAND4F_9.Y.n6 mux8_2.NAND4F_9.Y.t1 20.1899
R21400 mux8_2.NAND4F_9.Y.n6 mux8_2.NAND4F_9.Y.t0 20.1899
R21401 mux8_2.NAND4F_9.Y.n7 mux8_2.NAND4F_9.Y.t3 20.1899
R21402 mux8_2.NAND4F_9.Y.n7 mux8_2.NAND4F_9.Y.t4 20.1899
R21403 mux8_2.NAND4F_9.Y.n8 mux8_2.NAND4F_9.Y.t2 20.1899
R21404 mux8_2.NAND4F_9.Y.n8 mux8_2.NAND4F_9.Y.t8 20.1899
R21405 mux8_2.NAND4F_9.Y.n9 mux8_2.NAND4F_9.Y.t6 20.1899
R21406 mux8_2.NAND4F_9.Y.n9 mux8_2.NAND4F_9.Y.t7 20.1899
R21407 mux8_2.NAND4F_9.Y mux8_2.NAND4F_9.Y.n10 0.396904
R21408 mux8_2.NAND4F_9.Y.n10 mux8_2.NAND4F_9.Y.n0 0.358709
R21409 a_n12345_n23105.n2 a_n12345_n23105.t7 541.395
R21410 a_n12345_n23105.n3 a_n12345_n23105.t4 527.402
R21411 a_n12345_n23105.n2 a_n12345_n23105.t5 491.64
R21412 a_n12345_n23105.n5 a_n12345_n23105.t0 281.906
R21413 a_n12345_n23105.t1 a_n12345_n23105.n5 204.359
R21414 a_n12345_n23105.n0 a_n12345_n23105.t3 180.73
R21415 a_n12345_n23105.n1 a_n12345_n23105.t2 179.45
R21416 a_n12345_n23105.n0 a_n12345_n23105.t6 139.78
R21417 a_n12345_n23105.n4 a_n12345_n23105.n1 105.635
R21418 a_n12345_n23105.n4 a_n12345_n23105.n3 76.0005
R21419 a_n12345_n23105.n5 a_n12345_n23105.n4 67.9685
R21420 a_n12345_n23105.n3 a_n12345_n23105.n2 13.994
R21421 a_n12345_n23105.n1 a_n12345_n23105.n0 1.28015
R21422 a_n6920_3190.n2 a_n6920_3190.n0 121.353
R21423 a_n6920_3190.n3 a_n6920_3190.n2 121.001
R21424 a_n6920_3190.n2 a_n6920_3190.n1 120.977
R21425 a_n6920_3190.n1 a_n6920_3190.t5 30.462
R21426 a_n6920_3190.n1 a_n6920_3190.t3 30.462
R21427 a_n6920_3190.n0 a_n6920_3190.t0 30.462
R21428 a_n6920_3190.n0 a_n6920_3190.t1 30.462
R21429 a_n6920_3190.t2 a_n6920_3190.n3 30.462
R21430 a_n6920_3190.n3 a_n6920_3190.t4 30.462
R21431 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n9 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t13 540.38
R21432 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t7 491.64
R21433 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t9 491.64
R21434 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t14 491.64
R21435 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t11 491.64
R21436 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n7 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t15 367.928
R21437 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n2 227.526
R21438 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n8 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t16 227.356
R21439 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n3 227.266
R21440 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n1 227.266
R21441 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n7 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t17 213.688
R21442 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n6 162.852
R21443 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n9 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n8 160.439
R21444 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t10 139.78
R21445 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t8 139.78
R21446 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t12 139.78
R21447 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t18 139.78
R21448 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n8 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n7 94.4341
R21449 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t0 42.7831
R21450 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n6 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n5 38.6833
R21451 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n3 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t5 30.379
R21452 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n3 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t2 30.379
R21453 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n1 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t1 30.379
R21454 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n1 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t6 30.379
R21455 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n2 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t3 30.379
R21456 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n2 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t4 30.379
R21457 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n6 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n4 28.3986
R21458 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n0 18.8832
R21459 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n10 10.7052
R21460 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n10 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 5.09176
R21461 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n10 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 4.19292
R21462 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n9 0.794268
R21463 a_n16483_2026.n0 a_n16483_2026.n2 81.2978
R21464 a_n16483_2026.n0 a_n16483_2026.n3 81.1637
R21465 a_n16483_2026.n0 a_n16483_2026.n4 81.1637
R21466 a_n16483_2026.n1 a_n16483_2026.n5 81.1637
R21467 a_n16483_2026.n1 a_n16483_2026.n6 81.1637
R21468 a_n16483_2026.n7 a_n16483_2026.n1 80.9213
R21469 a_n16483_2026.n2 a_n16483_2026.t11 11.8205
R21470 a_n16483_2026.n2 a_n16483_2026.t9 11.8205
R21471 a_n16483_2026.n3 a_n16483_2026.t2 11.8205
R21472 a_n16483_2026.n3 a_n16483_2026.t10 11.8205
R21473 a_n16483_2026.n4 a_n16483_2026.t1 11.8205
R21474 a_n16483_2026.n4 a_n16483_2026.t0 11.8205
R21475 a_n16483_2026.n5 a_n16483_2026.t8 11.8205
R21476 a_n16483_2026.n5 a_n16483_2026.t7 11.8205
R21477 a_n16483_2026.n6 a_n16483_2026.t4 11.8205
R21478 a_n16483_2026.n6 a_n16483_2026.t6 11.8205
R21479 a_n16483_2026.t5 a_n16483_2026.n7 11.8205
R21480 a_n16483_2026.n7 a_n16483_2026.t3 11.8205
R21481 a_n16483_2026.n1 a_n16483_2026.n0 0.402735
R21482 a_n22489_1406.n2 a_n22489_1406.n1 121.353
R21483 a_n22489_1406.n2 a_n22489_1406.n0 121.353
R21484 a_n22489_1406.n3 a_n22489_1406.n2 121.001
R21485 a_n22489_1406.n1 a_n22489_1406.t2 30.462
R21486 a_n22489_1406.n1 a_n22489_1406.t3 30.462
R21487 a_n22489_1406.n0 a_n22489_1406.t1 30.462
R21488 a_n22489_1406.n0 a_n22489_1406.t0 30.462
R21489 a_n22489_1406.n3 a_n22489_1406.t5 30.462
R21490 a_n22489_1406.t4 a_n22489_1406.n3 30.462
R21491 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t13 540.38
R21492 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t10 491.64
R21493 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t8 491.64
R21494 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t9 491.64
R21495 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t14 491.64
R21496 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t16 367.928
R21497 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n2 227.526
R21498 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t11 227.356
R21499 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n1 227.266
R21500 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n3 227.266
R21501 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n7 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t15 213.688
R21502 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n6 162.852
R21503 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n8 160.439
R21504 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t18 139.78
R21505 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t12 139.78
R21506 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t7 139.78
R21507 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t17 139.78
R21508 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n7 94.4341
R21509 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t5 42.7831
R21510 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n5 38.6833
R21511 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t0 30.379
R21512 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t1 30.379
R21513 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t6 30.379
R21514 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t4 30.379
R21515 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t3 30.379
R21516 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t2 30.379
R21517 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n4 28.3986
R21518 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n0 18.8832
R21519 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n10 10.7052
R21520 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT 5.09176
R21521 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT 4.19292
R21522 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n9 0.794268
R21523 a_n11840_n11683.n2 a_n11840_n11683.n0 121.353
R21524 a_n11840_n11683.n3 a_n11840_n11683.n2 121.353
R21525 a_n11840_n11683.n2 a_n11840_n11683.n1 121.001
R21526 a_n11840_n11683.n1 a_n11840_n11683.t4 30.462
R21527 a_n11840_n11683.n1 a_n11840_n11683.t0 30.462
R21528 a_n11840_n11683.n0 a_n11840_n11683.t5 30.462
R21529 a_n11840_n11683.n0 a_n11840_n11683.t3 30.462
R21530 a_n11840_n11683.n3 a_n11840_n11683.t1 30.462
R21531 a_n11840_n11683.t2 a_n11840_n11683.n3 30.462
R21532 a_n12345_n31403.n2 a_n12345_n31403.t3 539.788
R21533 a_n12345_n31403.n3 a_n12345_n31403.t5 531.496
R21534 a_n12345_n31403.n2 a_n12345_n31403.t4 490.034
R21535 a_n12345_n31403.n5 a_n12345_n31403.t0 283.788
R21536 a_n12345_n31403.t1 a_n12345_n31403.n5 205.489
R21537 a_n12345_n31403.n0 a_n12345_n31403.t6 182.625
R21538 a_n12345_n31403.n1 a_n12345_n31403.t2 179.054
R21539 a_n12345_n31403.n0 a_n12345_n31403.t7 139.78
R21540 a_n12345_n31403.n4 a_n12345_n31403.n1 101.368
R21541 a_n12345_n31403.n5 a_n12345_n31403.n4 77.9135
R21542 a_n12345_n31403.n4 a_n12345_n31403.n3 76.1557
R21543 a_n12345_n31403.n3 a_n12345_n31403.n2 8.29297
R21544 a_n12345_n31403.n1 a_n12345_n31403.n0 3.57087
R21545 a_n11274_n31661.n2 a_n11274_n31661.n1 121.353
R21546 a_n11274_n31661.n3 a_n11274_n31661.n2 121.001
R21547 a_n11274_n31661.n2 a_n11274_n31661.n0 120.977
R21548 a_n11274_n31661.n0 a_n11274_n31661.t1 30.462
R21549 a_n11274_n31661.n0 a_n11274_n31661.t0 30.462
R21550 a_n11274_n31661.n1 a_n11274_n31661.t4 30.462
R21551 a_n11274_n31661.n1 a_n11274_n31661.t5 30.462
R21552 a_n11274_n31661.t2 a_n11274_n31661.n3 30.462
R21553 a_n11274_n31661.n3 a_n11274_n31661.t3 30.462
R21554 a_n20659_3810.n0 a_n20659_3810.n2 81.2978
R21555 a_n20659_3810.n1 a_n20659_3810.n5 81.1637
R21556 a_n20659_3810.n0 a_n20659_3810.n4 81.1637
R21557 a_n20659_3810.n0 a_n20659_3810.n3 81.1637
R21558 a_n20659_3810.n7 a_n20659_3810.n1 81.1637
R21559 a_n20659_3810.n1 a_n20659_3810.n6 80.9213
R21560 a_n20659_3810.n6 a_n20659_3810.t0 11.8205
R21561 a_n20659_3810.n6 a_n20659_3810.t1 11.8205
R21562 a_n20659_3810.n5 a_n20659_3810.t6 11.8205
R21563 a_n20659_3810.n5 a_n20659_3810.t7 11.8205
R21564 a_n20659_3810.n4 a_n20659_3810.t10 11.8205
R21565 a_n20659_3810.n4 a_n20659_3810.t11 11.8205
R21566 a_n20659_3810.n3 a_n20659_3810.t3 11.8205
R21567 a_n20659_3810.n3 a_n20659_3810.t9 11.8205
R21568 a_n20659_3810.n2 a_n20659_3810.t4 11.8205
R21569 a_n20659_3810.n2 a_n20659_3810.t5 11.8205
R21570 a_n20659_3810.n7 a_n20659_3810.t8 11.8205
R21571 a_n20659_3810.t2 a_n20659_3810.n7 11.8205
R21572 a_n20659_3810.n1 a_n20659_3810.n0 0.402735
R21573 A6.n5 A6.t21 540.38
R21574 A6.n13 A6.t19 540.375
R21575 A6.n6 A6.t8 491.64
R21576 A6.n6 A6.t23 491.64
R21577 A6.n6 A6.t29 491.64
R21578 A6.n6 A6.t20 491.64
R21579 A6.n1 A6.t5 491.64
R21580 A6.n1 A6.t4 491.64
R21581 A6.n1 A6.t22 491.64
R21582 A6.n1 A6.t6 491.64
R21583 A6.n3 A6.t0 367.928
R21584 A6.n11 A6.t27 343.827
R21585 A6.n16 A6.t1 312.599
R21586 A6.n19 A6.t26 247.428
R21587 A6.n18 A6.t14 247.428
R21588 A6.n17 A6.t13 247.428
R21589 A6.n16 A6.t7 247.428
R21590 A6.n11 A6.t28 237.787
R21591 A6.n20 A6.t24 229.754
R21592 A6.n12 A6.t9 227.356
R21593 A6.n4 A6.t2 227.356
R21594 A6.n3 A6.t3 213.688
R21595 A6 A6.n2 163.036
R21596 A6.n9 A6.n8 162.867
R21597 A6 A6.n20 162.409
R21598 A6.n5 A6.n4 160.439
R21599 A6.n13 A6.n12 160.433
R21600 A6.n7 A6.t18 139.78
R21601 A6.n7 A6.t11 139.78
R21602 A6.n7 A6.t25 139.78
R21603 A6.n7 A6.t12 139.78
R21604 A6.n0 A6.t10 139.78
R21605 A6.n0 A6.t17 139.78
R21606 A6.n0 A6.t16 139.78
R21607 A6.n0 A6.t15 139.78
R21608 A6.n4 A6.n3 94.4341
R21609 A6.n20 A6.n19 91.5805
R21610 A6.n12 A6.n11 70.3341
R21611 A6.n17 A6.n16 65.1723
R21612 A6.n18 A6.n17 65.1723
R21613 A6.n19 A6.n18 65.1723
R21614 A6.n2 A6.n0 38.8368
R21615 A6.n8 A6.n7 38.6833
R21616 A6.n8 A6.n6 28.3986
R21617 A6.n2 A6.n1 28.2451
R21618 A6 A6.n21 19.5453
R21619 A6 A6.n10 18.1908
R21620 A6.n21 A6 12.7976
R21621 A6.n15 A6.n14 12.4105
R21622 A6.n10 A6.n9 9.00496
R21623 A6.n21 A6.n15 4.19023
R21624 A6.n10 A6 3.87912
R21625 A6.n14 A6 1.41239
R21626 A6 A6.n13 0.905186
R21627 A6 A6.n5 0.89693
R21628 A6.n14 A6 0.0721292
R21629 A6.n9 A6 0.0590664
R21630 A6.n15 A6 0.0109444
R21631 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t7 540.38
R21632 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t8 367.928
R21633 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n4 227.526
R21634 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t9 227.356
R21635 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n5 227.266
R21636 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n6 227.266
R21637 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t10 213.688
R21638 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n2 160.439
R21639 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n1 94.4341
R21640 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t0 42.7944
R21641 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t6 30.379
R21642 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t5 30.379
R21643 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t2 30.379
R21644 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t4 30.379
R21645 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t3 30.379
R21646 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.t1 30.379
R21647 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n0 13.4358
R21648 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B.n3 0.821842
R21649 a_n19028_n8445.n2 a_n19028_n8445.t2 541.395
R21650 a_n19028_n8445.n3 a_n19028_n8445.t5 527.402
R21651 a_n19028_n8445.n2 a_n19028_n8445.t7 491.64
R21652 a_n19028_n8445.n5 a_n19028_n8445.t0 281.906
R21653 a_n19028_n8445.t1 a_n19028_n8445.n5 204.359
R21654 a_n19028_n8445.n0 a_n19028_n8445.t3 180.73
R21655 a_n19028_n8445.n1 a_n19028_n8445.t6 179.45
R21656 a_n19028_n8445.n0 a_n19028_n8445.t4 139.78
R21657 a_n19028_n8445.n4 a_n19028_n8445.n1 105.635
R21658 a_n19028_n8445.n4 a_n19028_n8445.n3 76.0005
R21659 a_n19028_n8445.n5 a_n19028_n8445.n4 67.9685
R21660 a_n19028_n8445.n3 a_n19028_n8445.n2 13.994
R21661 a_n19028_n8445.n1 a_n19028_n8445.n0 1.28015
R21662 a_n18998_n7799.n7 a_n18998_n7799.n1 81.2978
R21663 a_n18998_n7799.n1 a_n18998_n7799.n6 81.1637
R21664 a_n18998_n7799.n1 a_n18998_n7799.n5 81.1637
R21665 a_n18998_n7799.n0 a_n18998_n7799.n4 81.1637
R21666 a_n18998_n7799.n0 a_n18998_n7799.n3 81.1637
R21667 a_n18998_n7799.n0 a_n18998_n7799.n2 80.9213
R21668 a_n18998_n7799.n6 a_n18998_n7799.t2 11.8205
R21669 a_n18998_n7799.n6 a_n18998_n7799.t3 11.8205
R21670 a_n18998_n7799.n5 a_n18998_n7799.t0 11.8205
R21671 a_n18998_n7799.n5 a_n18998_n7799.t1 11.8205
R21672 a_n18998_n7799.n4 a_n18998_n7799.t6 11.8205
R21673 a_n18998_n7799.n4 a_n18998_n7799.t8 11.8205
R21674 a_n18998_n7799.n3 a_n18998_n7799.t9 11.8205
R21675 a_n18998_n7799.n3 a_n18998_n7799.t7 11.8205
R21676 a_n18998_n7799.n2 a_n18998_n7799.t11 11.8205
R21677 a_n18998_n7799.n2 a_n18998_n7799.t10 11.8205
R21678 a_n18998_n7799.t5 a_n18998_n7799.n7 11.8205
R21679 a_n18998_n7799.n7 a_n18998_n7799.t4 11.8205
R21680 a_n18998_n7799.n1 a_n18998_n7799.n0 0.402735
R21681 a_11386_n35462.t0 a_11386_n35462.t1 9.9005
R21682 mux8_6.NAND4F_9.Y.n1 mux8_6.NAND4F_9.Y.t11 312.599
R21683 mux8_6.NAND4F_9.Y.n4 mux8_6.NAND4F_9.Y.t10 247.428
R21684 mux8_6.NAND4F_9.Y.n1 mux8_6.NAND4F_9.Y.t12 247.428
R21685 mux8_6.NAND4F_9.Y.n2 mux8_6.NAND4F_9.Y.t13 247.428
R21686 mux8_6.NAND4F_9.Y.n3 mux8_6.NAND4F_9.Y.t9 247.428
R21687 mux8_6.NAND4F_9.Y.n5 mux8_6.NAND4F_9.Y.t14 229.754
R21688 mux8_6.NAND4F_9.Y.n0 mux8_6.NAND4F_9.Y.n6 187.373
R21689 mux8_6.NAND4F_9.Y.n0 mux8_6.NAND4F_9.Y.n7 187.192
R21690 mux8_6.NAND4F_9.Y.n0 mux8_6.NAND4F_9.Y.n8 187.192
R21691 mux8_6.NAND4F_9.Y.n10 mux8_6.NAND4F_9.Y.n9 187.192
R21692 mux8_6.NAND4F_9.Y mux8_6.NAND4F_9.Y.n5 162.275
R21693 mux8_6.NAND4F_9.Y.n5 mux8_6.NAND4F_9.Y.n4 91.5805
R21694 mux8_6.NAND4F_9.Y.n2 mux8_6.NAND4F_9.Y.n1 65.1723
R21695 mux8_6.NAND4F_9.Y.n3 mux8_6.NAND4F_9.Y.n2 65.1723
R21696 mux8_6.NAND4F_9.Y.n4 mux8_6.NAND4F_9.Y.n3 65.1723
R21697 mux8_6.NAND4F_9.Y mux8_6.NAND4F_9.Y.t2 22.6141
R21698 mux8_6.NAND4F_9.Y.n6 mux8_6.NAND4F_9.Y.t7 20.1899
R21699 mux8_6.NAND4F_9.Y.n6 mux8_6.NAND4F_9.Y.t8 20.1899
R21700 mux8_6.NAND4F_9.Y.n7 mux8_6.NAND4F_9.Y.t5 20.1899
R21701 mux8_6.NAND4F_9.Y.n7 mux8_6.NAND4F_9.Y.t6 20.1899
R21702 mux8_6.NAND4F_9.Y.n8 mux8_6.NAND4F_9.Y.t0 20.1899
R21703 mux8_6.NAND4F_9.Y.n8 mux8_6.NAND4F_9.Y.t1 20.1899
R21704 mux8_6.NAND4F_9.Y.n9 mux8_6.NAND4F_9.Y.t4 20.1899
R21705 mux8_6.NAND4F_9.Y.n9 mux8_6.NAND4F_9.Y.t3 20.1899
R21706 mux8_6.NAND4F_9.Y mux8_6.NAND4F_9.Y.n10 0.396904
R21707 mux8_6.NAND4F_9.Y.n10 mux8_6.NAND4F_9.Y.n0 0.358709
R21708 a_n8200_1380.n2 a_n8200_1380.t7 541.395
R21709 a_n8200_1380.n3 a_n8200_1380.t6 527.402
R21710 a_n8200_1380.n2 a_n8200_1380.t3 491.64
R21711 a_n8200_1380.n5 a_n8200_1380.t0 281.906
R21712 a_n8200_1380.t1 a_n8200_1380.n5 204.359
R21713 a_n8200_1380.n0 a_n8200_1380.t5 180.73
R21714 a_n8200_1380.n1 a_n8200_1380.t2 179.45
R21715 a_n8200_1380.n0 a_n8200_1380.t4 139.78
R21716 a_n8200_1380.n4 a_n8200_1380.n1 105.635
R21717 a_n8200_1380.n4 a_n8200_1380.n3 76.0005
R21718 a_n8200_1380.n5 a_n8200_1380.n4 67.9685
R21719 a_n8200_1380.n3 a_n8200_1380.n2 13.994
R21720 a_n8200_1380.n1 a_n8200_1380.n0 1.28015
R21721 a_n15707_n11063.n0 a_n15707_n11063.n2 81.2978
R21722 a_n15707_n11063.n0 a_n15707_n11063.n3 81.1637
R21723 a_n15707_n11063.n0 a_n15707_n11063.n4 81.1637
R21724 a_n15707_n11063.n1 a_n15707_n11063.n5 81.1637
R21725 a_n15707_n11063.n1 a_n15707_n11063.n6 81.1637
R21726 a_n15707_n11063.n7 a_n15707_n11063.n1 80.9213
R21727 a_n15707_n11063.n2 a_n15707_n11063.t8 11.8205
R21728 a_n15707_n11063.n2 a_n15707_n11063.t7 11.8205
R21729 a_n15707_n11063.n3 a_n15707_n11063.t11 11.8205
R21730 a_n15707_n11063.n3 a_n15707_n11063.t9 11.8205
R21731 a_n15707_n11063.n4 a_n15707_n11063.t10 11.8205
R21732 a_n15707_n11063.n4 a_n15707_n11063.t6 11.8205
R21733 a_n15707_n11063.n5 a_n15707_n11063.t1 11.8205
R21734 a_n15707_n11063.n5 a_n15707_n11063.t0 11.8205
R21735 a_n15707_n11063.n6 a_n15707_n11063.t4 11.8205
R21736 a_n15707_n11063.n6 a_n15707_n11063.t2 11.8205
R21737 a_n15707_n11063.t5 a_n15707_n11063.n7 11.8205
R21738 a_n15707_n11063.n7 a_n15707_n11063.t3 11.8205
R21739 a_n15707_n11063.n1 a_n15707_n11063.n0 0.402735
R21740 a_n9305_n5154.n0 a_n9305_n5154.t3 539.788
R21741 a_n9305_n5154.n1 a_n9305_n5154.t6 531.496
R21742 a_n9305_n5154.n0 a_n9305_n5154.t4 490.034
R21743 a_n9305_n5154.n5 a_n9305_n5154.t0 283.788
R21744 a_n9305_n5154.t1 a_n9305_n5154.n5 205.489
R21745 a_n9305_n5154.n2 a_n9305_n5154.t7 182.625
R21746 a_n9305_n5154.n3 a_n9305_n5154.t5 179.054
R21747 a_n9305_n5154.n2 a_n9305_n5154.t2 139.78
R21748 a_n9305_n5154.n4 a_n9305_n5154.n3 101.368
R21749 a_n9305_n5154.n5 a_n9305_n5154.n4 77.9135
R21750 a_n9305_n5154.n4 a_n9305_n5154.n1 76.1557
R21751 a_n9305_n5154.n1 a_n9305_n5154.n0 8.29297
R21752 a_n9305_n5154.n3 a_n9305_n5154.n2 3.57087
R21753 MULT_0.S1.n0 MULT_0.S1.t14 1032.02
R21754 MULT_0.S1.n0 MULT_0.S1.t13 336.962
R21755 MULT_0.S1.n0 MULT_0.S1.t12 326.154
R21756 mux8_2.NAND4F_0.A MULT_0.S1.n0 162.952
R21757 MULT_0.S1.n3 MULT_0.S1.n2 120.999
R21758 MULT_0.S1.n3 MULT_0.S1.n1 120.999
R21759 MULT_0.S1.n15 MULT_0.S1.n14 104.489
R21760 MULT_0.S1.n5 MULT_0.S1.n4 92.5005
R21761 MULT_0.S1.n12 MULT_0.S1.n10 86.2638
R21762 MULT_0.S1.n10 MULT_0.S1.n9 85.8873
R21763 MULT_0.S1.n10 MULT_0.S1.n7 85.724
R21764 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.Y MULT_0.S1.n15 83.8907
R21765 MULT_0.S1.n13 MULT_0.S1.n12 75.0672
R21766 MULT_0.S1.n13 MULT_0.S1.n9 75.0672
R21767 MULT_0.S1.n12 MULT_0.S1.n11 73.1255
R21768 MULT_0.S1.n9 MULT_0.S1.n8 73.1255
R21769 MULT_0.S1.n7 MULT_0.S1.n6 73.1255
R21770 MULT_0.S1.n14 MULT_0.S1.n7 68.8946
R21771 MULT_0.4bit_ADDER_0.S0 mux8_2.A1 44.2371
R21772 MULT_0.S1.n15 MULT_0.S1.n5 41.9827
R21773 MULT_0.S1.n4 MULT_0.S1.t5 30.462
R21774 MULT_0.S1.n4 MULT_0.S1.t8 30.462
R21775 MULT_0.S1.n2 MULT_0.S1.t6 30.462
R21776 MULT_0.S1.n2 MULT_0.S1.t7 30.462
R21777 MULT_0.S1.n1 MULT_0.S1.t3 30.462
R21778 MULT_0.S1.n1 MULT_0.S1.t4 30.462
R21779 MULT_0.S1.n5 MULT_0.S1.n3 28.124
R21780 mux8_2.A1 mux8_2.NAND4F_0.A 17.2107
R21781 MULT_0.S1.n8 MULT_0.S1.t1 11.8205
R21782 MULT_0.S1.n8 MULT_0.S1.t2 11.8205
R21783 MULT_0.S1.n11 MULT_0.S1.t10 11.8205
R21784 MULT_0.S1.n11 MULT_0.S1.t9 11.8205
R21785 MULT_0.S1.n6 MULT_0.S1.t0 11.8205
R21786 MULT_0.S1.n6 MULT_0.S1.t11 11.8205
R21787 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.Y MULT_0.4bit_ADDER_0.S0 10.5465
R21788 MULT_0.S1.n14 MULT_0.S1.n13 9.3005
R21789 a_n9125_n5154.n2 a_n9125_n5154.n1 121.353
R21790 a_n9125_n5154.n3 a_n9125_n5154.n2 121.001
R21791 a_n9125_n5154.n2 a_n9125_n5154.n0 120.977
R21792 a_n9125_n5154.n1 a_n9125_n5154.t1 30.462
R21793 a_n9125_n5154.n1 a_n9125_n5154.t2 30.462
R21794 a_n9125_n5154.n0 a_n9125_n5154.t3 30.462
R21795 a_n9125_n5154.n0 a_n9125_n5154.t5 30.462
R21796 a_n9125_n5154.t4 a_n9125_n5154.n3 30.462
R21797 a_n9125_n5154.n3 a_n9125_n5154.t0 30.462
R21798 MULT_0.4bit_ADDER_0.A3.n3 MULT_0.4bit_ADDER_0.A3.t15 540.38
R21799 MULT_0.4bit_ADDER_0.A3.n4 MULT_0.4bit_ADDER_0.A3.t10 491.64
R21800 MULT_0.4bit_ADDER_0.A3.n4 MULT_0.4bit_ADDER_0.A3.t4 491.64
R21801 MULT_0.4bit_ADDER_0.A3.n4 MULT_0.4bit_ADDER_0.A3.t14 491.64
R21802 MULT_0.4bit_ADDER_0.A3.n4 MULT_0.4bit_ADDER_0.A3.t7 491.64
R21803 MULT_0.4bit_ADDER_0.A3.n1 MULT_0.4bit_ADDER_0.A3.t12 367.928
R21804 MULT_0.inv_11.Y MULT_0.4bit_ADDER_0.A3.t3 256.514
R21805 MULT_0.4bit_ADDER_0.A3.n2 MULT_0.4bit_ADDER_0.A3.t9 227.356
R21806 MULT_0.inv_11.Y MULT_0.4bit_ADDER_0.A3.n7 226.248
R21807 MULT_0.4bit_ADDER_0.A3.n1 MULT_0.4bit_ADDER_0.A3.t6 213.688
R21808 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_0.B MULT_0.4bit_ADDER_0.A3.n6 162.867
R21809 MULT_0.4bit_ADDER_0.A3.n3 MULT_0.4bit_ADDER_0.A3.n2 160.439
R21810 MULT_0.4bit_ADDER_0.A3.n5 MULT_0.4bit_ADDER_0.A3.t11 139.78
R21811 MULT_0.4bit_ADDER_0.A3.n5 MULT_0.4bit_ADDER_0.A3.t5 139.78
R21812 MULT_0.4bit_ADDER_0.A3.n5 MULT_0.4bit_ADDER_0.A3.t8 139.78
R21813 MULT_0.4bit_ADDER_0.A3.n5 MULT_0.4bit_ADDER_0.A3.t13 139.78
R21814 MULT_0.4bit_ADDER_0.A3.n2 MULT_0.4bit_ADDER_0.A3.n1 94.4341
R21815 MULT_0.inv_11.Y MULT_0.4bit_ADDER_0.A3.t0 83.8155
R21816 MULT_0.4bit_ADDER_0.A3.n6 MULT_0.4bit_ADDER_0.A3.n5 38.6833
R21817 MULT_0.4bit_ADDER_0.A3.n7 MULT_0.4bit_ADDER_0.A3.t2 30.379
R21818 MULT_0.4bit_ADDER_0.A3.n7 MULT_0.4bit_ADDER_0.A3.t1 30.379
R21819 MULT_0.4bit_ADDER_0.A3.n6 MULT_0.4bit_ADDER_0.A3.n4 28.3986
R21820 MULT_0.4bit_ADDER_0.A3.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_0.B 9.00496
R21821 MULT_0.4bit_ADDER_0.A3.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_0.B 3.87912
R21822 MULT_0.inv_11.Y MULT_0.4bit_ADDER_0.A3.n0 2.57842
R21823 MULT_0.4bit_ADDER_0.A3.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.A 1.47848
R21824 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_0.B MULT_0.4bit_ADDER_0.A3.n3 0.89693
R21825 a_n20557_n4534.n0 a_n20557_n4534.n3 81.2978
R21826 a_n20557_n4534.n0 a_n20557_n4534.n4 81.1637
R21827 a_n20557_n4534.n0 a_n20557_n4534.n5 81.1637
R21828 a_n20557_n4534.n1 a_n20557_n4534.n6 81.1637
R21829 a_n20557_n4534.n7 a_n20557_n4534.n1 81.1637
R21830 a_n20557_n4534.n1 a_n20557_n4534.n2 80.9213
R21831 a_n20557_n4534.n3 a_n20557_n4534.t7 11.8205
R21832 a_n20557_n4534.n3 a_n20557_n4534.t6 11.8205
R21833 a_n20557_n4534.n4 a_n20557_n4534.t5 11.8205
R21834 a_n20557_n4534.n4 a_n20557_n4534.t8 11.8205
R21835 a_n20557_n4534.n5 a_n20557_n4534.t3 11.8205
R21836 a_n20557_n4534.n5 a_n20557_n4534.t4 11.8205
R21837 a_n20557_n4534.n6 a_n20557_n4534.t10 11.8205
R21838 a_n20557_n4534.n6 a_n20557_n4534.t11 11.8205
R21839 a_n20557_n4534.n2 a_n20557_n4534.t1 11.8205
R21840 a_n20557_n4534.n2 a_n20557_n4534.t0 11.8205
R21841 a_n20557_n4534.t2 a_n20557_n4534.n7 11.8205
R21842 a_n20557_n4534.n7 a_n20557_n4534.t9 11.8205
R21843 a_n20557_n4534.n1 a_n20557_n4534.n0 0.402735
R21844 a_n19178_n8419.n0 a_n19178_n8419.t3 539.788
R21845 a_n19178_n8419.n1 a_n19178_n8419.t6 531.496
R21846 a_n19178_n8419.n0 a_n19178_n8419.t5 490.034
R21847 a_n19178_n8419.n5 a_n19178_n8419.t0 283.788
R21848 a_n19178_n8419.t1 a_n19178_n8419.n5 205.489
R21849 a_n19178_n8419.n2 a_n19178_n8419.t7 182.625
R21850 a_n19178_n8419.n3 a_n19178_n8419.t4 179.054
R21851 a_n19178_n8419.n2 a_n19178_n8419.t2 139.78
R21852 a_n19178_n8419.n4 a_n19178_n8419.n3 101.368
R21853 a_n19178_n8419.n5 a_n19178_n8419.n4 77.9135
R21854 a_n19178_n8419.n4 a_n19178_n8419.n1 76.1557
R21855 a_n19178_n8419.n1 a_n19178_n8419.n0 8.29297
R21856 a_n19178_n8419.n3 a_n19178_n8419.n2 3.57087
R21857 a_n18998_n8419.n2 a_n18998_n8419.n0 121.353
R21858 a_n18998_n8419.n2 a_n18998_n8419.n1 121.001
R21859 a_n18998_n8419.n3 a_n18998_n8419.n2 120.977
R21860 a_n18998_n8419.n0 a_n18998_n8419.t4 30.462
R21861 a_n18998_n8419.n0 a_n18998_n8419.t3 30.462
R21862 a_n18998_n8419.n1 a_n18998_n8419.t1 30.462
R21863 a_n18998_n8419.n1 a_n18998_n8419.t5 30.462
R21864 a_n18998_n8419.n3 a_n18998_n8419.t0 30.462
R21865 a_n18998_n8419.t2 a_n18998_n8419.n3 30.462
R21866 mux8_2.inv_0.A.n3 mux8_2.inv_0.A.t9 291.829
R21867 mux8_2.inv_0.A.n3 mux8_2.inv_0.A.t7 291.829
R21868 mux8_2.inv_0.A.n0 mux8_2.inv_0.A.t2 256.425
R21869 mux8_2.inv_0.A.n0 mux8_2.inv_0.A.n4 231.24
R21870 mux8_2.inv_0.A.n0 mux8_2.inv_0.A.n5 231.03
R21871 mux8_2.inv_0.A.n3 mux8_2.inv_0.A.t10 221.72
R21872 mux8_2.inv_0.A.t8 mux8_2.inv_0.A.n2 393.959
R21873 mux8_2.inv_0.A.n6 mux8_2.inv_0.A.n1 66.6316
R21874 mux8_2.inv_0.A.n2 mux8_2.inv_0.A.n3 53.4611
R21875 mux8_2.inv_0.A.n5 mux8_2.inv_0.A.t3 25.395
R21876 mux8_2.inv_0.A.n5 mux8_2.inv_0.A.t4 25.395
R21877 mux8_2.inv_0.A.n4 mux8_2.inv_0.A.t5 25.395
R21878 mux8_2.inv_0.A.n4 mux8_2.inv_0.A.t1 25.395
R21879 mux8_2.inv_0.A.n6 mux8_2.inv_0.A.t6 19.8005
R21880 mux8_2.inv_0.A.n6 mux8_2.inv_0.A.t0 19.8005
R21881 mux8_2.inv_0.A.n1 mux8_2.inv_0.A.n0 0.38953
R21882 mux8_2.inv_0.A.n1 mux8_2.inv_0.A.n2 0.294762
R21883 a_n10864_n11683.n0 a_n10864_n11683.t2 539.788
R21884 a_n10864_n11683.n1 a_n10864_n11683.t5 531.496
R21885 a_n10864_n11683.n0 a_n10864_n11683.t6 490.034
R21886 a_n10864_n11683.n5 a_n10864_n11683.t1 283.788
R21887 a_n10864_n11683.t0 a_n10864_n11683.n5 205.489
R21888 a_n10864_n11683.n2 a_n10864_n11683.t7 182.625
R21889 a_n10864_n11683.n3 a_n10864_n11683.t3 179.054
R21890 a_n10864_n11683.n2 a_n10864_n11683.t4 139.78
R21891 a_n10864_n11683.n4 a_n10864_n11683.n3 101.368
R21892 a_n10864_n11683.n5 a_n10864_n11683.n4 77.9135
R21893 a_n10864_n11683.n4 a_n10864_n11683.n1 76.1557
R21894 a_n10864_n11683.n1 a_n10864_n11683.n0 8.29297
R21895 a_n10864_n11683.n3 a_n10864_n11683.n2 3.57087
R21896 a_n13399_n11683.n2 a_n13399_n11683.n1 121.353
R21897 a_n13399_n11683.n2 a_n13399_n11683.n0 121.353
R21898 a_n13399_n11683.n3 a_n13399_n11683.n2 121.001
R21899 a_n13399_n11683.n1 a_n13399_n11683.t4 30.462
R21900 a_n13399_n11683.n1 a_n13399_n11683.t3 30.462
R21901 a_n13399_n11683.n0 a_n13399_n11683.t0 30.462
R21902 a_n13399_n11683.n0 a_n13399_n11683.t1 30.462
R21903 a_n13399_n11683.t2 a_n13399_n11683.n3 30.462
R21904 a_n13399_n11683.n3 a_n13399_n11683.t5 30.462
R21905 a_n19178_n5154.n0 a_n19178_n5154.t4 539.788
R21906 a_n19178_n5154.n1 a_n19178_n5154.t7 531.496
R21907 a_n19178_n5154.n0 a_n19178_n5154.t5 490.034
R21908 a_n19178_n5154.n5 a_n19178_n5154.t0 283.788
R21909 a_n19178_n5154.t1 a_n19178_n5154.n5 205.489
R21910 a_n19178_n5154.n2 a_n19178_n5154.t2 182.625
R21911 a_n19178_n5154.n3 a_n19178_n5154.t6 179.054
R21912 a_n19178_n5154.n2 a_n19178_n5154.t3 139.78
R21913 a_n19178_n5154.n4 a_n19178_n5154.n3 101.368
R21914 a_n19178_n5154.n5 a_n19178_n5154.n4 77.9135
R21915 a_n19178_n5154.n4 a_n19178_n5154.n1 76.1557
R21916 a_n19178_n5154.n1 a_n19178_n5154.n0 8.29297
R21917 a_n19178_n5154.n3 a_n19178_n5154.n2 3.57087
R21918 a_n18998_n5154.n2 a_n18998_n5154.n0 121.353
R21919 a_n18998_n5154.n2 a_n18998_n5154.n1 121.001
R21920 a_n18998_n5154.n3 a_n18998_n5154.n2 120.977
R21921 a_n18998_n5154.n0 a_n18998_n5154.t4 30.462
R21922 a_n18998_n5154.n0 a_n18998_n5154.t5 30.462
R21923 a_n18998_n5154.n1 a_n18998_n5154.t0 30.462
R21924 a_n18998_n5154.n1 a_n18998_n5154.t3 30.462
R21925 a_n18998_n5154.t2 a_n18998_n5154.n3 30.462
R21926 a_n18998_n5154.n3 a_n18998_n5154.t1 30.462
R21927 AND8_0.NOT8_0.A4.n2 AND8_0.NOT8_0.A4.t7 394.37
R21928 AND8_0.NOT8_0.A4.n1 AND8_0.NOT8_0.A4.t10 291.829
R21929 AND8_0.NOT8_0.A4.n1 AND8_0.NOT8_0.A4.t8 291.829
R21930 AND8_0.NOT8_0.A4.n0 AND8_0.NOT8_0.A4.n4 227.526
R21931 AND8_0.NOT8_0.A4.n0 AND8_0.NOT8_0.A4.n5 227.266
R21932 AND8_0.NOT8_0.A4.n0 AND8_0.NOT8_0.A4.n3 227.266
R21933 AND8_0.NOT8_0.A4.n1 AND8_0.NOT8_0.A4.t9 221.72
R21934 AND8_0.NOT8_0.A4.n2 AND8_0.NOT8_0.A4.n1 53.374
R21935 AND8_0.NOT8_0.A4.n0 AND8_0.NOT8_0.A4.t4 42.7663
R21936 AND8_0.NOT8_0.A4.n5 AND8_0.NOT8_0.A4.t6 30.379
R21937 AND8_0.NOT8_0.A4.n5 AND8_0.NOT8_0.A4.t1 30.379
R21938 AND8_0.NOT8_0.A4.n3 AND8_0.NOT8_0.A4.t3 30.379
R21939 AND8_0.NOT8_0.A4.n3 AND8_0.NOT8_0.A4.t5 30.379
R21940 AND8_0.NOT8_0.A4.n4 AND8_0.NOT8_0.A4.t0 30.379
R21941 AND8_0.NOT8_0.A4.n4 AND8_0.NOT8_0.A4.t2 30.379
R21942 AND8_0.NOT8_0.A4 AND8_0.NOT8_0.A4.n0 2.07191
R21943 AND8_0.NOT8_0.A4 AND8_0.NOT8_0.A4.n2 1.28112
R21944 AND8_0.S4.n1 AND8_0.S4.t6 1032.02
R21945 AND8_0.S4.n1 AND8_0.S4.t4 336.962
R21946 AND8_0.S4.n1 AND8_0.S4.t5 326.154
R21947 AND8_0.S4.n0 AND8_0.S4.t1 256.514
R21948 AND8_0.S4.n0 AND8_0.S4.n2 226.258
R21949 AND8_0.S4 AND8_0.S4.n1 162.945
R21950 AND8_0.S4.n0 AND8_0.S4.t0 83.7172
R21951 AND8_0.S4.n2 AND8_0.S4.t2 30.379
R21952 AND8_0.S4.n2 AND8_0.S4.t3 30.379
R21953 AND8_0.S4 AND8_0.S4.n0 1.93382
R21954 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t23 491.64
R21955 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t18 491.64
R21956 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t15 491.64
R21957 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t13 491.64
R21958 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t12 485.221
R21959 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t22 367.928
R21960 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t21 255.588
R21961 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t17 224.478
R21962 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t20 213.688
R21963 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n18 209.19
R21964 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t19 139.78
R21965 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t14 139.78
R21966 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t16 139.78
R21967 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n1 120.999
R21968 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n0 120.999
R21969 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n13 104.489
R21970 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 103.258
R21971 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n3 92.5005
R21972 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n8 86.2638
R21973 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n9 85.8873
R21974 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n6 85.724
R21975 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n16 84.5046
R21976 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n14 84.0545
R21977 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n8 75.0672
R21978 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n11 75.0672
R21979 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n6 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n5 73.1255
R21980 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n8 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n7 73.1255
R21981 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n10 73.1255
R21982 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n15 72.3005
R21983 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n6 68.8946
R21984 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n17 60.9816
R21985 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n4 41.9827
R21986 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t6 30.462
R21987 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t9 30.462
R21988 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t10 30.462
R21989 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t11 30.462
R21990 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t7 30.462
R21991 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t8 30.462
R21992 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n2 28.124
R21993 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n19 17.8661
R21994 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n20 17.8661
R21995 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n21 17.1217
R21996 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n23 15.6329
R21997 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t4 11.8205
R21998 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t5 11.8205
R21999 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t3 11.8205
R22000 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t2 11.8205
R22001 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t0 11.8205
R22002 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t1 11.8205
R22003 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 10.8165
R22004 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n12 9.3005
R22005 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n24 2.50602
R22006 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n22 1.8615
R22007 a_n7909_373.t0 a_n7909_373.t1 19.8005
R22008 a_n19187_n9452.t0 a_n19187_n9452.t1 19.8005
R22009 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t18 491.64
R22010 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t17 491.64
R22011 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t12 491.64
R22012 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t22 491.64
R22013 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t15 485.221
R22014 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t21 367.928
R22015 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t16 255.588
R22016 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t20 224.478
R22017 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t19 213.688
R22018 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n0 209.19
R22019 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t14 139.78
R22020 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t23 139.78
R22021 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t13 139.78
R22022 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n11 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n10 120.999
R22023 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n11 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n9 120.999
R22024 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n23 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n22 104.489
R22025 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n13 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n12 92.5005
R22026 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n20 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n18 86.2638
R22027 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n18 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n17 85.8873
R22028 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n18 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n15 85.724
R22029 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n8 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n7 84.5046
R22030 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n23 83.8907
R22031 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n21 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n20 75.0672
R22032 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n21 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n17 75.0672
R22033 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n20 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n19 73.1255
R22034 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n17 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n16 73.1255
R22035 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n15 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n14 73.1255
R22036 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n7 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n6 72.3005
R22037 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n22 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n15 68.8946
R22038 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n8 60.9797
R22039 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n23 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n13 41.9827
R22040 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n12 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t1 30.462
R22041 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n12 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t8 30.462
R22042 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t7 30.462
R22043 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n10 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t3 30.462
R22044 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t2 30.462
R22045 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t0 30.462
R22046 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n13 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n11 28.124
R22047 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n5 19.963
R22048 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n1 17.8661
R22049 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n2 17.8661
R22050 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n3 17.1217
R22051 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n16 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t10 11.8205
R22052 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n16 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t9 11.8205
R22053 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n19 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t6 11.8205
R22054 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n19 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t5 11.8205
R22055 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n14 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t11 11.8205
R22056 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n14 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t4 11.8205
R22057 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n22 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n21 9.3005
R22058 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n4 1.8615
R22059 a_n16690_n11683.n2 a_n16690_n11683.n1 121.353
R22060 a_n16690_n11683.n2 a_n16690_n11683.n0 121.353
R22061 a_n16690_n11683.n3 a_n16690_n11683.n2 121.001
R22062 a_n16690_n11683.n1 a_n16690_n11683.t0 30.462
R22063 a_n16690_n11683.n1 a_n16690_n11683.t1 30.462
R22064 a_n16690_n11683.n0 a_n16690_n11683.t3 30.462
R22065 a_n16690_n11683.n0 a_n16690_n11683.t4 30.462
R22066 a_n16690_n11683.n3 a_n16690_n11683.t5 30.462
R22067 a_n16690_n11683.t2 a_n16690_n11683.n3 30.462
R22068 a_n23374_3190.n2 a_n23374_3190.n0 121.353
R22069 a_n23374_3190.n3 a_n23374_3190.n2 121.001
R22070 a_n23374_3190.n2 a_n23374_3190.n1 120.977
R22071 a_n23374_3190.n1 a_n23374_3190.t4 30.462
R22072 a_n23374_3190.n1 a_n23374_3190.t0 30.462
R22073 a_n23374_3190.n0 a_n23374_3190.t1 30.462
R22074 a_n23374_3190.n0 a_n23374_3190.t2 30.462
R22075 a_n23374_3190.t3 a_n23374_3190.n3 30.462
R22076 a_n23374_3190.n3 a_n23374_3190.t5 30.462
R22077 MULT_0.NAND2_15.Y.n5 MULT_0.NAND2_15.Y.t7 291.829
R22078 MULT_0.NAND2_15.Y.n5 MULT_0.NAND2_15.Y.t9 291.829
R22079 MULT_0.NAND2_15.Y.n0 MULT_0.NAND2_15.Y.n3 227.526
R22080 MULT_0.NAND2_15.Y.n0 MULT_0.NAND2_15.Y.n2 227.266
R22081 MULT_0.NAND2_15.Y.n0 MULT_0.NAND2_15.Y.n4 227.266
R22082 MULT_0.NAND2_15.Y.n5 MULT_0.NAND2_15.Y.t8 221.72
R22083 MULT_0.NAND2_15.Y.t10 MULT_0.NAND2_15.Y.n1 393.897
R22084 MULT_0.NAND2_15.Y.n0 MULT_0.NAND2_15.Y.t0 42.7333
R22085 MULT_0.NAND2_15.Y.n3 MULT_0.NAND2_15.Y.t6 30.379
R22086 MULT_0.NAND2_15.Y.n3 MULT_0.NAND2_15.Y.t4 30.379
R22087 MULT_0.NAND2_15.Y.n2 MULT_0.NAND2_15.Y.t1 30.379
R22088 MULT_0.NAND2_15.Y.n2 MULT_0.NAND2_15.Y.t2 30.379
R22089 MULT_0.NAND2_15.Y.n4 MULT_0.NAND2_15.Y.t3 30.379
R22090 MULT_0.NAND2_15.Y.n4 MULT_0.NAND2_15.Y.t5 30.379
R22091 MULT_0.NAND2_15.Y.n5 MULT_0.NAND2_15.Y.n1 53.4915
R22092 MULT_0.NAND2_15.Y.n0 MULT_0.NAND2_15.Y.n1 0.622976
R22093 AND8_0.NOT8_0.A5.n2 AND8_0.NOT8_0.A5.t10 394.37
R22094 AND8_0.NOT8_0.A5.n1 AND8_0.NOT8_0.A5.t9 291.829
R22095 AND8_0.NOT8_0.A5.n1 AND8_0.NOT8_0.A5.t7 291.829
R22096 AND8_0.NOT8_0.A5.n0 AND8_0.NOT8_0.A5.n4 227.526
R22097 AND8_0.NOT8_0.A5.n0 AND8_0.NOT8_0.A5.n5 227.266
R22098 AND8_0.NOT8_0.A5.n0 AND8_0.NOT8_0.A5.n3 227.266
R22099 AND8_0.NOT8_0.A5.n1 AND8_0.NOT8_0.A5.t8 221.72
R22100 AND8_0.NOT8_0.A5.n2 AND8_0.NOT8_0.A5.n1 53.374
R22101 AND8_0.NOT8_0.A5.n0 AND8_0.NOT8_0.A5.t3 42.7768
R22102 AND8_0.NOT8_0.A5.n5 AND8_0.NOT8_0.A5.t5 30.379
R22103 AND8_0.NOT8_0.A5.n5 AND8_0.NOT8_0.A5.t1 30.379
R22104 AND8_0.NOT8_0.A5.n3 AND8_0.NOT8_0.A5.t4 30.379
R22105 AND8_0.NOT8_0.A5.n3 AND8_0.NOT8_0.A5.t6 30.379
R22106 AND8_0.NOT8_0.A5.n4 AND8_0.NOT8_0.A5.t0 30.379
R22107 AND8_0.NOT8_0.A5.n4 AND8_0.NOT8_0.A5.t2 30.379
R22108 AND8_0.NOT8_0.A5 AND8_0.NOT8_0.A5.n0 2.03413
R22109 AND8_0.NOT8_0.A5 AND8_0.NOT8_0.A5.n2 1.27931
R22110 a_n11490_1380.n2 a_n11490_1380.t3 541.395
R22111 a_n11490_1380.n3 a_n11490_1380.t7 527.402
R22112 a_n11490_1380.n2 a_n11490_1380.t5 491.64
R22113 a_n11490_1380.n5 a_n11490_1380.t0 281.906
R22114 a_n11490_1380.t1 a_n11490_1380.n5 204.359
R22115 a_n11490_1380.n0 a_n11490_1380.t2 180.73
R22116 a_n11490_1380.n1 a_n11490_1380.t4 179.45
R22117 a_n11490_1380.n0 a_n11490_1380.t6 139.78
R22118 a_n11490_1380.n4 a_n11490_1380.n1 105.635
R22119 a_n11490_1380.n4 a_n11490_1380.n3 76.0005
R22120 a_n11490_1380.n5 a_n11490_1380.n4 67.9685
R22121 a_n11490_1380.n3 a_n11490_1380.n2 13.994
R22122 a_n11490_1380.n1 a_n11490_1380.n0 1.28015
R22123 a_n11460_1406.n2 a_n11460_1406.n1 121.353
R22124 a_n11460_1406.n3 a_n11460_1406.n2 121.001
R22125 a_n11460_1406.n2 a_n11460_1406.n0 120.977
R22126 a_n11460_1406.n1 a_n11460_1406.t0 30.462
R22127 a_n11460_1406.n1 a_n11460_1406.t1 30.462
R22128 a_n11460_1406.n0 a_n11460_1406.t5 30.462
R22129 a_n11460_1406.n0 a_n11460_1406.t4 30.462
R22130 a_n11460_1406.n3 a_n11460_1406.t3 30.462
R22131 a_n11460_1406.t2 a_n11460_1406.n3 30.462
R22132 mux8_6.inv_0.A.n1 mux8_6.inv_0.A.t7 291.829
R22133 mux8_6.inv_0.A.n1 mux8_6.inv_0.A.t9 291.829
R22134 mux8_6.inv_0.A.n0 mux8_6.inv_0.A.t5 256.425
R22135 mux8_6.inv_0.A.n0 mux8_6.inv_0.A.n2 231.24
R22136 mux8_6.inv_0.A.n0 mux8_6.inv_0.A.n3 231.03
R22137 mux8_6.inv_0.A.n1 mux8_6.inv_0.A.t8 221.72
R22138 mux8_6.inv_0.A.t10 mux8_6.inv_0.A.n0 393.959
R22139 mux8_6.inv_0.A.n4 mux8_6.inv_0.A.n0 66.6316
R22140 mux8_6.inv_0.A.n0 mux8_6.inv_0.A.n1 54.1444
R22141 mux8_6.inv_0.A.n3 mux8_6.inv_0.A.t4 25.395
R22142 mux8_6.inv_0.A.n3 mux8_6.inv_0.A.t3 25.395
R22143 mux8_6.inv_0.A.n2 mux8_6.inv_0.A.t2 25.395
R22144 mux8_6.inv_0.A.n2 mux8_6.inv_0.A.t1 25.395
R22145 mux8_6.inv_0.A.n4 mux8_6.inv_0.A.t6 19.8005
R22146 mux8_6.inv_0.A.n4 mux8_6.inv_0.A.t0 19.8005
R22147 a_11865_n34471.n1 a_11865_n34471.n4 231.24
R22148 a_11865_n34471.n0 a_11865_n34471.n2 231.24
R22149 a_11865_n34471.n1 a_11865_n34471.n5 231.03
R22150 a_11865_n34471.n0 a_11865_n34471.n3 231.03
R22151 a_11865_n34471.n6 a_11865_n34471.n1 231.03
R22152 a_11865_n34471.n4 a_11865_n34471.t2 25.395
R22153 a_11865_n34471.n4 a_11865_n34471.t0 25.395
R22154 a_11865_n34471.n5 a_11865_n34471.t3 25.395
R22155 a_11865_n34471.n5 a_11865_n34471.t1 25.395
R22156 a_11865_n34471.n3 a_11865_n34471.t5 25.395
R22157 a_11865_n34471.n3 a_11865_n34471.t9 25.395
R22158 a_11865_n34471.n2 a_11865_n34471.t7 25.395
R22159 a_11865_n34471.n2 a_11865_n34471.t6 25.395
R22160 a_11865_n34471.n6 a_11865_n34471.t8 25.395
R22161 a_11865_n34471.t4 a_11865_n34471.n6 25.395
R22162 a_11865_n34471.n1 a_11865_n34471.n0 0.421553
R22163 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t12 491.64
R22164 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t17 491.64
R22165 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t14 491.64
R22166 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t22 491.64
R22167 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t18 485.221
R22168 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t19 367.928
R22169 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t16 255.588
R22170 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t20 224.478
R22171 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t21 213.688
R22172 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n18 209.19
R22173 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t23 139.78
R22174 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t13 139.78
R22175 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t15 139.78
R22176 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n1 120.999
R22177 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n0 120.999
R22178 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n13 104.489
R22179 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 103.258
R22180 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n3 92.5005
R22181 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n8 86.2638
R22182 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n9 85.8873
R22183 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n6 85.724
R22184 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n16 84.5046
R22185 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n14 84.0545
R22186 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n8 75.0672
R22187 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n11 75.0672
R22188 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n6 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n5 73.1255
R22189 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n8 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n7 73.1255
R22190 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n10 73.1255
R22191 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n15 72.3005
R22192 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n6 68.8946
R22193 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n17 60.9816
R22194 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n4 41.9827
R22195 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t11 30.462
R22196 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t2 30.462
R22197 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t1 30.462
R22198 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t0 30.462
R22199 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t9 30.462
R22200 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t10 30.462
R22201 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n2 28.124
R22202 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n19 17.8661
R22203 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n20 17.8661
R22204 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n21 17.1217
R22205 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n23 15.6329
R22206 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t6 11.8205
R22207 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t7 11.8205
R22208 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t8 11.8205
R22209 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t3 11.8205
R22210 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t4 11.8205
R22211 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t5 11.8205
R22212 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 10.8165
R22213 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n12 9.3005
R22214 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n24 2.50602
R22215 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n22 1.8615
R22216 a_n21333_2026.n1 a_n21333_2026.n6 81.2978
R22217 a_n21333_2026.n1 a_n21333_2026.n5 81.1637
R22218 a_n21333_2026.n0 a_n21333_2026.n4 81.1637
R22219 a_n21333_2026.n0 a_n21333_2026.n3 81.1637
R22220 a_n21333_2026.n7 a_n21333_2026.n1 81.1637
R22221 a_n21333_2026.n0 a_n21333_2026.n2 80.9213
R22222 a_n21333_2026.n6 a_n21333_2026.t1 11.8205
R22223 a_n21333_2026.n6 a_n21333_2026.t2 11.8205
R22224 a_n21333_2026.n5 a_n21333_2026.t8 11.8205
R22225 a_n21333_2026.n5 a_n21333_2026.t0 11.8205
R22226 a_n21333_2026.n4 a_n21333_2026.t9 11.8205
R22227 a_n21333_2026.n4 a_n21333_2026.t11 11.8205
R22228 a_n21333_2026.n3 a_n21333_2026.t5 11.8205
R22229 a_n21333_2026.n3 a_n21333_2026.t10 11.8205
R22230 a_n21333_2026.n2 a_n21333_2026.t6 11.8205
R22231 a_n21333_2026.n2 a_n21333_2026.t4 11.8205
R22232 a_n21333_2026.n7 a_n21333_2026.t7 11.8205
R22233 a_n21333_2026.t3 a_n21333_2026.n7 11.8205
R22234 a_n21333_2026.n1 a_n21333_2026.n0 0.402735
R22235 a_n12596_n11683.n0 a_n12596_n11683.t5 539.788
R22236 a_n12596_n11683.n1 a_n12596_n11683.t4 531.496
R22237 a_n12596_n11683.n0 a_n12596_n11683.t7 490.034
R22238 a_n12596_n11683.n5 a_n12596_n11683.t0 283.788
R22239 a_n12596_n11683.t1 a_n12596_n11683.n5 205.489
R22240 a_n12596_n11683.n2 a_n12596_n11683.t3 182.625
R22241 a_n12596_n11683.n3 a_n12596_n11683.t2 179.054
R22242 a_n12596_n11683.n2 a_n12596_n11683.t6 139.78
R22243 a_n12596_n11683.n4 a_n12596_n11683.n3 101.368
R22244 a_n12596_n11683.n5 a_n12596_n11683.n4 77.9135
R22245 a_n12596_n11683.n4 a_n12596_n11683.n1 76.1557
R22246 a_n12596_n11683.n1 a_n12596_n11683.n0 8.29297
R22247 a_n12596_n11683.n3 a_n12596_n11683.n2 3.57087
R22248 a_n1618_1380.n2 a_n1618_1380.t7 541.395
R22249 a_n1618_1380.n3 a_n1618_1380.t4 527.402
R22250 a_n1618_1380.n2 a_n1618_1380.t2 491.64
R22251 a_n1618_1380.n5 a_n1618_1380.t0 281.906
R22252 a_n1618_1380.t1 a_n1618_1380.n5 204.359
R22253 a_n1618_1380.n0 a_n1618_1380.t3 180.73
R22254 a_n1618_1380.n1 a_n1618_1380.t5 179.45
R22255 a_n1618_1380.n0 a_n1618_1380.t6 139.78
R22256 a_n1618_1380.n4 a_n1618_1380.n1 105.635
R22257 a_n1618_1380.n4 a_n1618_1380.n3 76.0005
R22258 a_n1618_1380.n5 a_n1618_1380.n4 67.9685
R22259 a_n1618_1380.n3 a_n1618_1380.n2 13.994
R22260 a_n1618_1380.n1 a_n1618_1380.n0 1.28015
R22261 a_n1588_2026.n0 a_n1588_2026.n2 81.2978
R22262 a_n1588_2026.n0 a_n1588_2026.n3 81.1637
R22263 a_n1588_2026.n0 a_n1588_2026.n4 81.1637
R22264 a_n1588_2026.n1 a_n1588_2026.n5 81.1637
R22265 a_n1588_2026.n1 a_n1588_2026.n6 81.1637
R22266 a_n1588_2026.n7 a_n1588_2026.n1 80.9213
R22267 a_n1588_2026.n2 a_n1588_2026.t9 11.8205
R22268 a_n1588_2026.n2 a_n1588_2026.t11 11.8205
R22269 a_n1588_2026.n3 a_n1588_2026.t3 11.8205
R22270 a_n1588_2026.n3 a_n1588_2026.t10 11.8205
R22271 a_n1588_2026.n4 a_n1588_2026.t4 11.8205
R22272 a_n1588_2026.n4 a_n1588_2026.t5 11.8205
R22273 a_n1588_2026.n5 a_n1588_2026.t8 11.8205
R22274 a_n1588_2026.n5 a_n1588_2026.t6 11.8205
R22275 a_n1588_2026.n6 a_n1588_2026.t1 11.8205
R22276 a_n1588_2026.n6 a_n1588_2026.t7 11.8205
R22277 a_n1588_2026.t2 a_n1588_2026.n7 11.8205
R22278 a_n1588_2026.n7 a_n1588_2026.t0 11.8205
R22279 a_n1588_2026.n1 a_n1588_2026.n0 0.402735
R22280 mux8_1.NAND4F_2.D.n4 mux8_1.NAND4F_2.D.t12 1388.16
R22281 mux8_1.NAND4F_2.D.n7 mux8_1.NAND4F_2.D.t9 1388.16
R22282 mux8_1.NAND4F_2.D.n10 mux8_1.NAND4F_2.D.t4 1388.16
R22283 mux8_1.NAND4F_2.D.n1 mux8_1.NAND4F_2.D.t10 1388.16
R22284 mux8_1.NAND4F_2.D.n4 mux8_1.NAND4F_2.D.t7 350.839
R22285 mux8_1.NAND4F_2.D.n7 mux8_1.NAND4F_2.D.t15 350.839
R22286 mux8_1.NAND4F_2.D.n10 mux8_1.NAND4F_2.D.t8 350.839
R22287 mux8_1.NAND4F_2.D.n1 mux8_1.NAND4F_2.D.t13 350.839
R22288 mux8_1.NAND4F_2.D.n5 mux8_1.NAND4F_2.D.t6 308.481
R22289 mux8_1.NAND4F_2.D.n8 mux8_1.NAND4F_2.D.t14 308.481
R22290 mux8_1.NAND4F_2.D.n11 mux8_1.NAND4F_2.D.t5 308.481
R22291 mux8_1.NAND4F_2.D.n2 mux8_1.NAND4F_2.D.t11 308.481
R22292 mux8_1.NAND4F_2.D.n0 mux8_1.NAND4F_2.D.t1 256.514
R22293 mux8_1.NAND4F_2.D.n0 mux8_1.NAND4F_2.D.n3 226.258
R22294 mux8_1.NAND4F_2.D mux8_1.NAND4F_2.D.n5 161.458
R22295 mux8_1.NAND4F_2.D mux8_1.NAND4F_2.D.n11 161.435
R22296 mux8_1.NAND4F_2.D mux8_1.NAND4F_2.D.n2 161.435
R22297 mux8_1.NAND4F_2.D mux8_1.NAND4F_2.D.n8 161.429
R22298 mux8_1.NAND4F_2.D.n0 mux8_1.NAND4F_2.D.t0 83.7172
R22299 mux8_1.NAND4F_2.D.n3 mux8_1.NAND4F_2.D.t3 30.379
R22300 mux8_1.NAND4F_2.D.n3 mux8_1.NAND4F_2.D.t2 30.379
R22301 mux8_1.NAND4F_2.D.n5 mux8_1.NAND4F_2.D.n4 27.752
R22302 mux8_1.NAND4F_2.D.n8 mux8_1.NAND4F_2.D.n7 27.752
R22303 mux8_1.NAND4F_2.D.n11 mux8_1.NAND4F_2.D.n10 27.752
R22304 mux8_1.NAND4F_2.D.n2 mux8_1.NAND4F_2.D.n1 27.752
R22305 mux8_1.NAND4F_2.D.n6 mux8_1.NAND4F_2.D.n0 12.759
R22306 mux8_1.NAND4F_2.D mux8_1.NAND4F_2.D.n12 10.6871
R22307 mux8_1.NAND4F_2.D.n6 mux8_1.NAND4F_2.D 9.0005
R22308 mux8_1.NAND4F_2.D.n12 mux8_1.NAND4F_2.D 9.0005
R22309 mux8_1.NAND4F_2.D.n9 mux8_1.NAND4F_2.D 9.0005
R22310 mux8_1.NAND4F_2.D.n9 mux8_1.NAND4F_2.D.n6 1.74507
R22311 mux8_1.NAND4F_2.D.n12 mux8_1.NAND4F_2.D.n9 1.69072
R22312 a_9336_n2838.t0 a_9336_n2838.t1 9.9005
R22313 a_n8350_1406.n0 a_n8350_1406.t5 539.788
R22314 a_n8350_1406.n1 a_n8350_1406.t2 531.496
R22315 a_n8350_1406.n0 a_n8350_1406.t4 490.034
R22316 a_n8350_1406.n5 a_n8350_1406.t0 283.788
R22317 a_n8350_1406.t1 a_n8350_1406.n5 205.489
R22318 a_n8350_1406.n2 a_n8350_1406.t3 182.625
R22319 a_n8350_1406.n3 a_n8350_1406.t6 179.054
R22320 a_n8350_1406.n2 a_n8350_1406.t7 139.78
R22321 a_n8350_1406.n4 a_n8350_1406.n3 101.368
R22322 a_n8350_1406.n5 a_n8350_1406.n4 77.9135
R22323 a_n8350_1406.n4 a_n8350_1406.n1 76.1557
R22324 a_n8350_1406.n1 a_n8350_1406.n0 8.29297
R22325 a_n8350_1406.n3 a_n8350_1406.n2 3.57087
R22326 a_n8170_2026.n7 a_n8170_2026.n1 81.2978
R22327 a_n8170_2026.n1 a_n8170_2026.n6 81.1637
R22328 a_n8170_2026.n1 a_n8170_2026.n5 81.1637
R22329 a_n8170_2026.n0 a_n8170_2026.n4 81.1637
R22330 a_n8170_2026.n0 a_n8170_2026.n3 81.1637
R22331 a_n8170_2026.n0 a_n8170_2026.n2 80.9213
R22332 a_n8170_2026.n6 a_n8170_2026.t8 11.8205
R22333 a_n8170_2026.n6 a_n8170_2026.t0 11.8205
R22334 a_n8170_2026.n5 a_n8170_2026.t6 11.8205
R22335 a_n8170_2026.n5 a_n8170_2026.t7 11.8205
R22336 a_n8170_2026.n4 a_n8170_2026.t11 11.8205
R22337 a_n8170_2026.n4 a_n8170_2026.t9 11.8205
R22338 a_n8170_2026.n3 a_n8170_2026.t3 11.8205
R22339 a_n8170_2026.n3 a_n8170_2026.t10 11.8205
R22340 a_n8170_2026.n2 a_n8170_2026.t4 11.8205
R22341 a_n8170_2026.n2 a_n8170_2026.t5 11.8205
R22342 a_n8170_2026.n7 a_n8170_2026.t1 11.8205
R22343 a_n8170_2026.t2 a_n8170_2026.n7 11.8205
R22344 a_n8170_2026.n1 a_n8170_2026.n0 0.402735
R22345 MULT_0.NAND2_1.Y.n5 MULT_0.NAND2_1.Y.t7 291.829
R22346 MULT_0.NAND2_1.Y.n5 MULT_0.NAND2_1.Y.t9 291.829
R22347 MULT_0.NAND2_1.Y.n0 MULT_0.NAND2_1.Y.n2 227.526
R22348 MULT_0.NAND2_1.Y.n0 MULT_0.NAND2_1.Y.n3 227.266
R22349 MULT_0.NAND2_1.Y.n0 MULT_0.NAND2_1.Y.n4 227.266
R22350 MULT_0.NAND2_1.Y.n5 MULT_0.NAND2_1.Y.t8 221.72
R22351 MULT_0.NAND2_1.Y.t10 MULT_0.NAND2_1.Y.n1 393.897
R22352 MULT_0.NAND2_1.Y.n0 MULT_0.NAND2_1.Y.t0 42.7333
R22353 MULT_0.NAND2_1.Y.n2 MULT_0.NAND2_1.Y.t5 30.379
R22354 MULT_0.NAND2_1.Y.n2 MULT_0.NAND2_1.Y.t4 30.379
R22355 MULT_0.NAND2_1.Y.n3 MULT_0.NAND2_1.Y.t2 30.379
R22356 MULT_0.NAND2_1.Y.n3 MULT_0.NAND2_1.Y.t6 30.379
R22357 MULT_0.NAND2_1.Y.n4 MULT_0.NAND2_1.Y.t1 30.379
R22358 MULT_0.NAND2_1.Y.n4 MULT_0.NAND2_1.Y.t3 30.379
R22359 MULT_0.NAND2_1.Y.n5 MULT_0.NAND2_1.Y.n1 53.4917
R22360 MULT_0.NAND2_1.Y.n0 MULT_0.NAND2_1.Y.n1 0.623962
R22361 MULT_0.4bit_ADDER_0.B1.n6 MULT_0.4bit_ADDER_0.B1.t6 491.64
R22362 MULT_0.4bit_ADDER_0.B1.n7 MULT_0.4bit_ADDER_0.B1.t12 491.64
R22363 MULT_0.4bit_ADDER_0.B1.n8 MULT_0.4bit_ADDER_0.B1.t11 491.64
R22364 MULT_0.4bit_ADDER_0.B1.n9 MULT_0.4bit_ADDER_0.B1.t14 491.64
R22365 MULT_0.4bit_ADDER_0.B1.n4 MULT_0.4bit_ADDER_0.B1.t13 485.221
R22366 MULT_0.4bit_ADDER_0.B1.n2 MULT_0.4bit_ADDER_0.B1.t5 367.928
R22367 MULT_0.4bit_ADDER_0.B1.n0 MULT_0.4bit_ADDER_0.B1.t1 256.514
R22368 MULT_0.4bit_ADDER_0.B1.n10 MULT_0.4bit_ADDER_0.B1.t10 255.588
R22369 MULT_0.4bit_ADDER_0.B1.n0 MULT_0.4bit_ADDER_0.B1.n1 226.251
R22370 MULT_0.4bit_ADDER_0.B1.n3 MULT_0.4bit_ADDER_0.B1.t9 224.478
R22371 MULT_0.4bit_ADDER_0.B1.n2 MULT_0.4bit_ADDER_0.B1.t8 213.688
R22372 MULT_0.4bit_ADDER_0.B1.n6 MULT_0.4bit_ADDER_0.B1.n5 209.19
R22373 MULT_0.4bit_ADDER_0.B1.n5 MULT_0.4bit_ADDER_0.B1.t4 139.78
R22374 MULT_0.4bit_ADDER_0.B1.n5 MULT_0.4bit_ADDER_0.B1.t15 139.78
R22375 MULT_0.4bit_ADDER_0.B1.n5 MULT_0.4bit_ADDER_0.B1.t7 139.78
R22376 MULT_0.4bit_ADDER_0.B1.n11 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_0.A 103.258
R22377 MULT_0.4bit_ADDER_0.B1.n4 MULT_0.4bit_ADDER_0.B1.n3 84.5046
R22378 MULT_0.4bit_ADDER_0.B1.n0 MULT_0.4bit_ADDER_0.B1.t0 83.7599
R22379 MULT_0.4bit_ADDER_0.B1.n3 MULT_0.4bit_ADDER_0.B1.n2 72.3005
R22380 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_0.A MULT_0.4bit_ADDER_0.B1.n4 60.9816
R22381 MULT_0.4bit_ADDER_0.B1.n1 MULT_0.4bit_ADDER_0.B1.t3 30.379
R22382 MULT_0.4bit_ADDER_0.B1.n1 MULT_0.4bit_ADDER_0.B1.t2 30.379
R22383 MULT_0.4bit_ADDER_0.B1.n7 MULT_0.4bit_ADDER_0.B1.n6 17.8661
R22384 MULT_0.4bit_ADDER_0.B1.n8 MULT_0.4bit_ADDER_0.B1.n7 17.8661
R22385 MULT_0.4bit_ADDER_0.FULL_ADDER_2.B MULT_0.4bit_ADDER_0.B1.n0 17.8223
R22386 MULT_0.4bit_ADDER_0.B1.n9 MULT_0.4bit_ADDER_0.B1.n8 17.1217
R22387 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_0.A MULT_0.4bit_ADDER_0.B1.n10 15.6329
R22388 MULT_0.4bit_ADDER_0.B1.n11 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_0.A 10.8165
R22389 MULT_0.4bit_ADDER_0.B1.n10 MULT_0.4bit_ADDER_0.B1.n9 1.8615
R22390 MULT_0.4bit_ADDER_0.FULL_ADDER_2.B MULT_0.4bit_ADDER_0.B1.n11 0.868086
R22391 a_n10714_n5180.n2 a_n10714_n5180.t2 541.395
R22392 a_n10714_n5180.n3 a_n10714_n5180.t3 527.402
R22393 a_n10714_n5180.n2 a_n10714_n5180.t5 491.64
R22394 a_n10714_n5180.n5 a_n10714_n5180.t1 281.906
R22395 a_n10714_n5180.t0 a_n10714_n5180.n5 204.359
R22396 a_n10714_n5180.n0 a_n10714_n5180.t4 180.73
R22397 a_n10714_n5180.n1 a_n10714_n5180.t7 179.45
R22398 a_n10714_n5180.n0 a_n10714_n5180.t6 139.78
R22399 a_n10714_n5180.n4 a_n10714_n5180.n1 105.635
R22400 a_n10714_n5180.n4 a_n10714_n5180.n3 76.0005
R22401 a_n10714_n5180.n5 a_n10714_n5180.n4 67.9685
R22402 a_n10714_n5180.n3 a_n10714_n5180.n2 13.994
R22403 a_n10714_n5180.n1 a_n10714_n5180.n0 1.28015
R22404 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t20 491.64
R22405 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t23 491.64
R22406 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t12 491.64
R22407 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t18 491.64
R22408 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n8 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t22 485.221
R22409 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t13 367.928
R22410 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t15 255.588
R22411 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t19 224.478
R22412 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t17 213.688
R22413 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n0 209.19
R22414 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t16 139.78
R22415 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t14 139.78
R22416 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t21 139.78
R22417 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n11 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n10 120.999
R22418 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n11 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n9 120.999
R22419 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n23 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n22 104.489
R22420 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n13 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n12 92.5005
R22421 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n20 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n18 86.2638
R22422 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n18 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n17 85.8873
R22423 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n18 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n15 85.724
R22424 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n8 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n7 84.5046
R22425 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n23 83.8907
R22426 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n21 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n20 75.0672
R22427 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n21 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n17 75.0672
R22428 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n20 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n19 73.1255
R22429 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n15 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n14 73.1255
R22430 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n17 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n16 73.1255
R22431 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n6 72.3005
R22432 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n22 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n15 68.8946
R22433 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n8 60.9797
R22434 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n23 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n13 41.9827
R22435 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n12 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t6 30.462
R22436 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n12 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t0 30.462
R22437 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n10 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t1 30.462
R22438 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n10 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t2 30.462
R22439 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n9 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t8 30.462
R22440 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n9 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t7 30.462
R22441 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n13 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n11 28.124
R22442 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n5 19.963
R22443 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n1 17.8661
R22444 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n2 17.8661
R22445 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n3 17.1217
R22446 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n14 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t5 11.8205
R22447 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n14 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t9 11.8205
R22448 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n19 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t10 11.8205
R22449 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n19 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t11 11.8205
R22450 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n16 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t4 11.8205
R22451 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n16 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t3 11.8205
R22452 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n22 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n21 9.3005
R22453 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n4 1.8615
R22454 a_n10684_n4534.n0 a_n10684_n4534.n4 81.2978
R22455 a_n10684_n4534.n0 a_n10684_n4534.n5 81.1637
R22456 a_n10684_n4534.n0 a_n10684_n4534.n6 81.1637
R22457 a_n10684_n4534.n1 a_n10684_n4534.n3 81.1637
R22458 a_n10684_n4534.n7 a_n10684_n4534.n1 81.1637
R22459 a_n10684_n4534.n1 a_n10684_n4534.n2 80.9213
R22460 a_n10684_n4534.n4 a_n10684_n4534.t8 11.8205
R22461 a_n10684_n4534.n4 a_n10684_n4534.t7 11.8205
R22462 a_n10684_n4534.n5 a_n10684_n4534.t11 11.8205
R22463 a_n10684_n4534.n5 a_n10684_n4534.t6 11.8205
R22464 a_n10684_n4534.n6 a_n10684_n4534.t9 11.8205
R22465 a_n10684_n4534.n6 a_n10684_n4534.t10 11.8205
R22466 a_n10684_n4534.n3 a_n10684_n4534.t3 11.8205
R22467 a_n10684_n4534.n3 a_n10684_n4534.t1 11.8205
R22468 a_n10684_n4534.n2 a_n10684_n4534.t4 11.8205
R22469 a_n10684_n4534.n2 a_n10684_n4534.t5 11.8205
R22470 a_n10684_n4534.n7 a_n10684_n4534.t0 11.8205
R22471 a_n10684_n4534.t2 a_n10684_n4534.n7 11.8205
R22472 a_n10684_n4534.n1 a_n10684_n4534.n0 0.402735
R22473 a_n9155_n5180.n2 a_n9155_n5180.t2 541.395
R22474 a_n9155_n5180.n3 a_n9155_n5180.t4 527.402
R22475 a_n9155_n5180.n2 a_n9155_n5180.t5 491.64
R22476 a_n9155_n5180.n5 a_n9155_n5180.t0 281.906
R22477 a_n9155_n5180.t1 a_n9155_n5180.n5 204.359
R22478 a_n9155_n5180.n0 a_n9155_n5180.t3 180.73
R22479 a_n9155_n5180.n1 a_n9155_n5180.t7 179.45
R22480 a_n9155_n5180.n0 a_n9155_n5180.t6 139.78
R22481 a_n9155_n5180.n4 a_n9155_n5180.n1 105.635
R22482 a_n9155_n5180.n4 a_n9155_n5180.n3 76.0005
R22483 a_n9155_n5180.n5 a_n9155_n5180.n4 67.9685
R22484 a_n9155_n5180.n3 a_n9155_n5180.n2 13.994
R22485 a_n9155_n5180.n1 a_n9155_n5180.n0 1.28015
R22486 a_n17677_n23825.n0 a_n17677_n23825.n2 231.24
R22487 a_n17677_n23825.n1 a_n17677_n23825.n5 231.24
R22488 a_n17677_n23825.n0 a_n17677_n23825.n3 231.03
R22489 a_n17677_n23825.n1 a_n17677_n23825.n4 231.03
R22490 a_n17677_n23825.n6 a_n17677_n23825.n1 231.03
R22491 a_n17677_n23825.n2 a_n17677_n23825.t1 25.395
R22492 a_n17677_n23825.n2 a_n17677_n23825.t0 25.395
R22493 a_n17677_n23825.n3 a_n17677_n23825.t4 25.395
R22494 a_n17677_n23825.n3 a_n17677_n23825.t3 25.395
R22495 a_n17677_n23825.n4 a_n17677_n23825.t2 25.395
R22496 a_n17677_n23825.n4 a_n17677_n23825.t9 25.395
R22497 a_n17677_n23825.n5 a_n17677_n23825.t6 25.395
R22498 a_n17677_n23825.n5 a_n17677_n23825.t5 25.395
R22499 a_n17677_n23825.t8 a_n17677_n23825.n6 25.395
R22500 a_n17677_n23825.n6 a_n17677_n23825.t7 25.395
R22501 a_n17677_n23825.n1 a_n17677_n23825.n0 0.421553
R22502 OR8_0.NOT8_0.A6.n3 OR8_0.NOT8_0.A6.t10 394.37
R22503 OR8_0.NOT8_0.A6.n2 OR8_0.NOT8_0.A6.t8 291.829
R22504 OR8_0.NOT8_0.A6.n2 OR8_0.NOT8_0.A6.t9 291.829
R22505 OR8_0.NOT8_0.A6.n0 OR8_0.NOT8_0.A6.t4 256.425
R22506 OR8_0.NOT8_0.A6.n0 OR8_0.NOT8_0.A6.n5 231.24
R22507 OR8_0.NOT8_0.A6.n0 OR8_0.NOT8_0.A6.n6 231.03
R22508 OR8_0.NOT8_0.A6.n2 OR8_0.NOT8_0.A6.t7 221.72
R22509 OR8_0.NOT8_0.A6.n4 OR8_0.NOT8_0.A6.n1 66.4681
R22510 OR8_0.NOT8_0.A6.n3 OR8_0.NOT8_0.A6.n2 53.374
R22511 OR8_0.NOT8_0.A6.n4 OR8_0.NOT8_0.A6 26.6429
R22512 OR8_0.NOT8_0.A6.n6 OR8_0.NOT8_0.A6.t3 25.395
R22513 OR8_0.NOT8_0.A6.n6 OR8_0.NOT8_0.A6.t2 25.395
R22514 OR8_0.NOT8_0.A6.n5 OR8_0.NOT8_0.A6.t1 25.395
R22515 OR8_0.NOT8_0.A6.n5 OR8_0.NOT8_0.A6.t0 25.395
R22516 OR8_0.NOT8_0.A6.n1 OR8_0.NOT8_0.A6.t5 19.8005
R22517 OR8_0.NOT8_0.A6.n1 OR8_0.NOT8_0.A6.t6 19.8005
R22518 OR8_0.NOT8_0.A6 OR8_0.NOT8_0.A6.n3 1.25939
R22519 OR8_0.NOT8_0.A6 OR8_0.NOT8_0.A6.n0 0.355237
R22520 OR8_0.NOT8_0.A6 OR8_0.NOT8_0.A6.n4 0.293873
R22521 mux8_6.NAND4F_0.C.n6 mux8_6.NAND4F_0.C.t11 978.795
R22522 mux8_6.NAND4F_0.C.n4 mux8_6.NAND4F_0.C.t6 978.795
R22523 mux8_6.NAND4F_0.C.n11 mux8_6.NAND4F_0.C.t8 978.795
R22524 mux8_6.NAND4F_0.C.n2 mux8_6.NAND4F_0.C.t10 978.795
R22525 mux8_6.NAND4F_0.C.n5 mux8_6.NAND4F_0.C.t13 308.481
R22526 mux8_6.NAND4F_0.C.n5 mux8_6.NAND4F_0.C.t12 308.481
R22527 mux8_6.NAND4F_0.C.n3 mux8_6.NAND4F_0.C.t9 308.481
R22528 mux8_6.NAND4F_0.C.n3 mux8_6.NAND4F_0.C.t7 308.481
R22529 mux8_6.NAND4F_0.C.n10 mux8_6.NAND4F_0.C.t4 308.481
R22530 mux8_6.NAND4F_0.C.n10 mux8_6.NAND4F_0.C.t5 308.481
R22531 mux8_6.NAND4F_0.C.n1 mux8_6.NAND4F_0.C.t14 308.481
R22532 mux8_6.NAND4F_0.C.n1 mux8_6.NAND4F_0.C.t15 308.481
R22533 mux8_6.NAND4F_0.C.n0 mux8_6.NAND4F_0.C.t1 256.514
R22534 mux8_6.NAND4F_0.C.n0 mux8_6.NAND4F_0.C.n8 226.258
R22535 mux8_6.NAND4F_0.C mux8_6.NAND4F_0.C.n6 161.856
R22536 mux8_6.NAND4F_0.C mux8_6.NAND4F_0.C.n4 161.847
R22537 mux8_6.NAND4F_0.C mux8_6.NAND4F_0.C.n11 161.84
R22538 mux8_6.NAND4F_0.C mux8_6.NAND4F_0.C.n2 161.831
R22539 mux8_6.NAND4F_0.C.n0 mux8_6.NAND4F_0.C.t0 83.7172
R22540 mux8_6.NAND4F_0.C.n8 mux8_6.NAND4F_0.C.t3 30.379
R22541 mux8_6.NAND4F_0.C.n8 mux8_6.NAND4F_0.C.t2 30.379
R22542 mux8_6.NAND4F_0.C.n9 mux8_6.NAND4F_0.C.n0 13.5186
R22543 mux8_6.NAND4F_0.C mux8_6.NAND4F_0.C.n12 13.0862
R22544 mux8_6.NAND4F_0.C.n7 mux8_6.NAND4F_0.C 13.0435
R22545 mux8_6.NAND4F_0.C.n12 mux8_6.NAND4F_0.C 12.4135
R22546 mux8_6.NAND4F_0.C.n7 mux8_6.NAND4F_0.C 12.4105
R22547 mux8_6.NAND4F_0.C.n6 mux8_6.NAND4F_0.C.n5 11.0463
R22548 mux8_6.NAND4F_0.C.n4 mux8_6.NAND4F_0.C.n3 11.0463
R22549 mux8_6.NAND4F_0.C.n11 mux8_6.NAND4F_0.C.n10 11.0463
R22550 mux8_6.NAND4F_0.C.n2 mux8_6.NAND4F_0.C.n1 11.0463
R22551 mux8_6.NAND4F_0.C.n12 mux8_6.NAND4F_0.C.n9 3.46056
R22552 mux8_6.NAND4F_0.C.n9 mux8_6.NAND4F_0.C.n7 1.8134
R22553 mux8_6.NAND4F_1.Y.n2 mux8_6.NAND4F_1.Y.t11 978.795
R22554 mux8_6.NAND4F_1.Y.n1 mux8_6.NAND4F_1.Y.t9 308.481
R22555 mux8_6.NAND4F_1.Y.n1 mux8_6.NAND4F_1.Y.t10 308.481
R22556 mux8_6.NAND4F_1.Y.n0 mux8_6.NAND4F_1.Y.n3 187.373
R22557 mux8_6.NAND4F_1.Y.n0 mux8_6.NAND4F_1.Y.n4 187.192
R22558 mux8_6.NAND4F_1.Y.n0 mux8_6.NAND4F_1.Y.n5 187.192
R22559 mux8_6.NAND4F_1.Y.n7 mux8_6.NAND4F_1.Y.n6 187.192
R22560 mux8_6.NAND4F_1.Y mux8_6.NAND4F_1.Y.n2 161.84
R22561 mux8_6.NAND4F_1.Y mux8_6.NAND4F_1.Y.t8 23.4335
R22562 mux8_6.NAND4F_1.Y.n3 mux8_6.NAND4F_1.Y.t1 20.1899
R22563 mux8_6.NAND4F_1.Y.n3 mux8_6.NAND4F_1.Y.t0 20.1899
R22564 mux8_6.NAND4F_1.Y.n4 mux8_6.NAND4F_1.Y.t3 20.1899
R22565 mux8_6.NAND4F_1.Y.n4 mux8_6.NAND4F_1.Y.t2 20.1899
R22566 mux8_6.NAND4F_1.Y.n5 mux8_6.NAND4F_1.Y.t5 20.1899
R22567 mux8_6.NAND4F_1.Y.n5 mux8_6.NAND4F_1.Y.t4 20.1899
R22568 mux8_6.NAND4F_1.Y.n6 mux8_6.NAND4F_1.Y.t6 20.1899
R22569 mux8_6.NAND4F_1.Y.n6 mux8_6.NAND4F_1.Y.t7 20.1899
R22570 mux8_6.NAND4F_1.Y.n2 mux8_6.NAND4F_1.Y.n1 11.0463
R22571 mux8_6.NAND4F_1.Y mux8_6.NAND4F_1.Y.n7 0.527586
R22572 mux8_6.NAND4F_1.Y.n7 mux8_6.NAND4F_1.Y.n0 0.358709
R22573 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t9 540.38
R22574 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t8 367.928
R22575 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n5 227.526
R22576 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t10 227.356
R22577 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n6 227.266
R22578 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n4 227.266
R22579 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t7 213.688
R22580 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n2 160.439
R22581 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n1 94.4341
R22582 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t3 42.7944
R22583 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t6 30.379
R22584 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t1 30.379
R22585 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t4 30.379
R22586 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t5 30.379
R22587 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t0 30.379
R22588 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.t2 30.379
R22589 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n0 13.4358
R22590 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B.n3 0.821842
R22591 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t9 485.221
R22592 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t8 367.928
R22593 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n5 227.526
R22594 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n4 227.266
R22595 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n6 227.266
R22596 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t7 224.478
R22597 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t10 213.688
R22598 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n2 84.5046
R22599 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n1 72.3005
R22600 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n3 61.0566
R22601 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t3 42.7747
R22602 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t1 30.379
R22603 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t0 30.379
R22604 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t4 30.379
R22605 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t6 30.379
R22606 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t5 30.379
R22607 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.t2 30.379
R22608 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A.n0 0.583137
R22609 mux8_3.NAND4F_5.Y.n1 mux8_3.NAND4F_5.Y.t11 1032.02
R22610 mux8_3.NAND4F_5.Y.n1 mux8_3.NAND4F_5.Y.t9 336.962
R22611 mux8_3.NAND4F_5.Y.n1 mux8_3.NAND4F_5.Y.t10 326.154
R22612 mux8_3.NAND4F_5.Y.n0 mux8_3.NAND4F_5.Y.n3 187.373
R22613 mux8_3.NAND4F_5.Y.n0 mux8_3.NAND4F_5.Y.n4 187.192
R22614 mux8_3.NAND4F_5.Y.n0 mux8_3.NAND4F_5.Y.n5 187.192
R22615 mux8_3.NAND4F_5.Y.n7 mux8_3.NAND4F_5.Y.n6 187.192
R22616 mux8_3.NAND4F_5.Y mux8_3.NAND4F_5.Y.n1 162.94
R22617 mux8_3.NAND4F_5.Y.n2 mux8_3.NAND4F_5.Y 24.4721
R22618 mux8_3.NAND4F_5.Y.n2 mux8_3.NAND4F_5.Y.t8 22.6141
R22619 mux8_3.NAND4F_5.Y.n3 mux8_3.NAND4F_5.Y.t1 20.1899
R22620 mux8_3.NAND4F_5.Y.n3 mux8_3.NAND4F_5.Y.t0 20.1899
R22621 mux8_3.NAND4F_5.Y.n4 mux8_3.NAND4F_5.Y.t2 20.1899
R22622 mux8_3.NAND4F_5.Y.n4 mux8_3.NAND4F_5.Y.t3 20.1899
R22623 mux8_3.NAND4F_5.Y.n5 mux8_3.NAND4F_5.Y.t4 20.1899
R22624 mux8_3.NAND4F_5.Y.n5 mux8_3.NAND4F_5.Y.t5 20.1899
R22625 mux8_3.NAND4F_5.Y.n6 mux8_3.NAND4F_5.Y.t6 20.1899
R22626 mux8_3.NAND4F_5.Y.n6 mux8_3.NAND4F_5.Y.t7 20.1899
R22627 mux8_3.NAND4F_5.Y mux8_3.NAND4F_5.Y.n2 0.950576
R22628 mux8_3.NAND4F_5.Y mux8_3.NAND4F_5.Y.n7 0.396904
R22629 mux8_3.NAND4F_5.Y.n7 mux8_3.NAND4F_5.Y.n0 0.358709
R22630 a_n9901_1406.n2 a_n9901_1406.n0 121.353
R22631 a_n9901_1406.n2 a_n9901_1406.n1 121.001
R22632 a_n9901_1406.n3 a_n9901_1406.n2 120.977
R22633 a_n9901_1406.n0 a_n9901_1406.t4 30.462
R22634 a_n9901_1406.n0 a_n9901_1406.t3 30.462
R22635 a_n9901_1406.n1 a_n9901_1406.t2 30.462
R22636 a_n9901_1406.n1 a_n9901_1406.t5 30.462
R22637 a_n9901_1406.t0 a_n9901_1406.n3 30.462
R22638 a_n9901_1406.n3 a_n9901_1406.t1 30.462
R22639 mux8_4.A0.n0 mux8_4.A0.t13 1032.02
R22640 mux8_4.A0.n0 mux8_4.A0.t12 336.962
R22641 mux8_4.A0.n0 mux8_4.A0.t14 326.154
R22642 mux8_4.A0 mux8_4.A0.n0 162.952
R22643 mux8_4.A0.n3 mux8_4.A0.n2 120.999
R22644 mux8_4.A0.n3 mux8_4.A0.n1 120.999
R22645 mux8_4.A0.n15 mux8_4.A0.n14 104.489
R22646 mux8_4.A0.n5 mux8_4.A0.n4 92.5005
R22647 mux8_4.A0.n12 mux8_4.A0.n10 86.2638
R22648 mux8_4.A0.n10 mux8_4.A0.n9 85.8873
R22649 mux8_4.A0.n10 mux8_4.A0.n7 85.724
R22650 mux8_4.A0 mux8_4.A0.n15 83.8907
R22651 mux8_4.A0.n13 mux8_4.A0.n12 75.0672
R22652 mux8_4.A0.n13 mux8_4.A0.n9 75.0672
R22653 mux8_4.A0.n12 mux8_4.A0.n11 73.1255
R22654 mux8_4.A0.n7 mux8_4.A0.n6 73.1255
R22655 mux8_4.A0.n9 mux8_4.A0.n8 73.1255
R22656 mux8_4.A0.n14 mux8_4.A0.n7 68.8946
R22657 mux8_4.A0.n15 mux8_4.A0.n5 41.9827
R22658 mux8_4.A0.n4 mux8_4.A0.t1 30.462
R22659 mux8_4.A0.n4 mux8_4.A0.t4 30.462
R22660 mux8_4.A0.n2 mux8_4.A0.t5 30.462
R22661 mux8_4.A0.n2 mux8_4.A0.t6 30.462
R22662 mux8_4.A0.n1 mux8_4.A0.t2 30.462
R22663 mux8_4.A0.n1 mux8_4.A0.t3 30.462
R22664 mux8_4.A0.n5 mux8_4.A0.n3 28.124
R22665 mux8_4.A0.n6 mux8_4.A0.t11 11.8205
R22666 mux8_4.A0.n6 mux8_4.A0.t9 11.8205
R22667 mux8_4.A0.n11 mux8_4.A0.t7 11.8205
R22668 mux8_4.A0.n11 mux8_4.A0.t8 11.8205
R22669 mux8_4.A0.n8 mux8_4.A0.t10 11.8205
R22670 mux8_4.A0.n8 mux8_4.A0.t0 11.8205
R22671 mux8_4.A0.n14 mux8_4.A0.n13 9.3005
R22672 AND8_0.S1.n2 AND8_0.S1.t4 1032.02
R22673 AND8_0.S1.n2 AND8_0.S1.t6 336.962
R22674 AND8_0.S1.n2 AND8_0.S1.t5 326.154
R22675 AND8_0.S1.n0 AND8_0.S1.t1 256.514
R22676 AND8_0.S1.n0 AND8_0.S1.n1 226.258
R22677 AND8_0.S1 AND8_0.S1.n2 162.945
R22678 AND8_0.S1.n0 AND8_0.S1.t0 83.7172
R22679 AND8_0.S1.n1 AND8_0.S1.t2 30.379
R22680 AND8_0.S1.n1 AND8_0.S1.t3 30.379
R22681 AND8_0.S1 AND8_0.S1.n0 1.91499
R22682 right_shifter_0.S5.n1 right_shifter_0.S5.t4 1032.02
R22683 right_shifter_0.S5.n1 right_shifter_0.S5.t5 336.962
R22684 right_shifter_0.S5.n1 right_shifter_0.S5.t6 326.154
R22685 right_shifter_0.S5.n0 right_shifter_0.S5.t1 256.514
R22686 right_shifter_0.S5.n0 right_shifter_0.S5.n2 226.258
R22687 mux8_7.NAND4F_6.A right_shifter_0.S5.n1 162.952
R22688 right_shifter_0.S5.n0 right_shifter_0.S5.t0 83.7172
R22689 mux8_7.A7 right_shifter_0.S5.n0 33.1497
R22690 right_shifter_0.S5.n2 right_shifter_0.S5.t3 30.379
R22691 right_shifter_0.S5.n2 right_shifter_0.S5.t2 30.379
R22692 mux8_7.A7 mux8_7.NAND4F_6.A 13.4456
R22693 a_8592_n26406.t0 a_8592_n26406.t1 9.9005
R22694 mux8_7.NAND4F_6.Y.n1 mux8_7.NAND4F_6.Y.t9 933.563
R22695 mux8_7.NAND4F_6.Y.n1 mux8_7.NAND4F_6.Y.t10 367.635
R22696 mux8_7.NAND4F_6.Y.n2 mux8_7.NAND4F_6.Y.t11 308.481
R22697 mux8_7.NAND4F_6.Y.n0 mux8_7.NAND4F_6.Y.n4 187.373
R22698 mux8_7.NAND4F_6.Y.n0 mux8_7.NAND4F_6.Y.n5 187.192
R22699 mux8_7.NAND4F_6.Y.n0 mux8_7.NAND4F_6.Y.n6 187.192
R22700 mux8_7.NAND4F_6.Y.n8 mux8_7.NAND4F_6.Y.n7 187.192
R22701 mux8_7.NAND4F_6.Y mux8_7.NAND4F_6.Y.n2 162.047
R22702 mux8_7.NAND4F_6.Y.n3 mux8_7.NAND4F_6.Y.t2 22.7831
R22703 mux8_7.NAND4F_6.Y.n3 mux8_7.NAND4F_6.Y 22.171
R22704 mux8_7.NAND4F_6.Y.n4 mux8_7.NAND4F_6.Y.t1 20.1899
R22705 mux8_7.NAND4F_6.Y.n4 mux8_7.NAND4F_6.Y.t0 20.1899
R22706 mux8_7.NAND4F_6.Y.n5 mux8_7.NAND4F_6.Y.t6 20.1899
R22707 mux8_7.NAND4F_6.Y.n5 mux8_7.NAND4F_6.Y.t5 20.1899
R22708 mux8_7.NAND4F_6.Y.n6 mux8_7.NAND4F_6.Y.t7 20.1899
R22709 mux8_7.NAND4F_6.Y.n6 mux8_7.NAND4F_6.Y.t8 20.1899
R22710 mux8_7.NAND4F_6.Y.n7 mux8_7.NAND4F_6.Y.t4 20.1899
R22711 mux8_7.NAND4F_6.Y.n7 mux8_7.NAND4F_6.Y.t3 20.1899
R22712 mux8_7.NAND4F_6.Y.n2 mux8_7.NAND4F_6.Y.n1 10.955
R22713 mux8_7.NAND4F_6.Y mux8_7.NAND4F_6.Y.n3 0.781576
R22714 mux8_7.NAND4F_6.Y mux8_7.NAND4F_6.Y.n8 0.396904
R22715 mux8_7.NAND4F_6.Y.n8 mux8_7.NAND4F_6.Y.n0 0.358709
R22716 a_n1012_1406.n2 a_n1012_1406.n0 121.353
R22717 a_n1012_1406.n3 a_n1012_1406.n2 121.353
R22718 a_n1012_1406.n2 a_n1012_1406.n1 121.001
R22719 a_n1012_1406.n0 a_n1012_1406.t4 30.462
R22720 a_n1012_1406.n0 a_n1012_1406.t3 30.462
R22721 a_n1012_1406.n1 a_n1012_1406.t1 30.462
R22722 a_n1012_1406.n1 a_n1012_1406.t5 30.462
R22723 a_n1012_1406.t2 a_n1012_1406.n3 30.462
R22724 a_n1012_1406.n3 a_n1012_1406.t0 30.462
R22725 a_10363_n26405.t0 a_10363_n26405.t1 9.9005
R22726 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t7 485.221
R22727 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t9 367.928
R22728 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n5 227.526
R22729 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n4 227.266
R22730 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n6 227.266
R22731 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t8 224.478
R22732 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t10 213.688
R22733 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n2 84.5046
R22734 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n1 72.3005
R22735 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n3 61.0566
R22736 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t0 42.7747
R22737 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t6 30.379
R22738 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t4 30.379
R22739 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t1 30.379
R22740 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t2 30.379
R22741 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t3 30.379
R22742 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.t5 30.379
R22743 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A.n0 0.583137
R22744 a_n10240_3164.n0 a_n10240_3164.t6 539.788
R22745 a_n10240_3164.n1 a_n10240_3164.t4 531.496
R22746 a_n10240_3164.n0 a_n10240_3164.t2 490.034
R22747 a_n10240_3164.n5 a_n10240_3164.t0 283.788
R22748 a_n10240_3164.t1 a_n10240_3164.n5 205.489
R22749 a_n10240_3164.n2 a_n10240_3164.t5 182.625
R22750 a_n10240_3164.n3 a_n10240_3164.t3 179.054
R22751 a_n10240_3164.n2 a_n10240_3164.t7 139.78
R22752 a_n10240_3164.n4 a_n10240_3164.n3 101.368
R22753 a_n10240_3164.n5 a_n10240_3164.n4 77.9135
R22754 a_n10240_3164.n4 a_n10240_3164.n1 76.1557
R22755 a_n10240_3164.n1 a_n10240_3164.n0 8.29297
R22756 a_n10240_3164.n3 a_n10240_3164.n2 3.57087
R22757 a_n10786_3810.n0 a_n10786_3810.n2 81.2978
R22758 a_n10786_3810.n1 a_n10786_3810.n5 81.1637
R22759 a_n10786_3810.n0 a_n10786_3810.n4 81.1637
R22760 a_n10786_3810.n0 a_n10786_3810.n3 81.1637
R22761 a_n10786_3810.n7 a_n10786_3810.n1 81.1637
R22762 a_n10786_3810.n1 a_n10786_3810.n6 80.9213
R22763 a_n10786_3810.n6 a_n10786_3810.t0 11.8205
R22764 a_n10786_3810.n6 a_n10786_3810.t1 11.8205
R22765 a_n10786_3810.n5 a_n10786_3810.t7 11.8205
R22766 a_n10786_3810.n5 a_n10786_3810.t6 11.8205
R22767 a_n10786_3810.n4 a_n10786_3810.t5 11.8205
R22768 a_n10786_3810.n4 a_n10786_3810.t3 11.8205
R22769 a_n10786_3810.n3 a_n10786_3810.t10 11.8205
R22770 a_n10786_3810.n3 a_n10786_3810.t4 11.8205
R22771 a_n10786_3810.n2 a_n10786_3810.t8 11.8205
R22772 a_n10786_3810.n2 a_n10786_3810.t9 11.8205
R22773 a_n10786_3810.n7 a_n10786_3810.t11 11.8205
R22774 a_n10786_3810.t2 a_n10786_3810.n7 11.8205
R22775 a_n10786_3810.n1 a_n10786_3810.n0 0.402735
R22776 a_n20587_n5180.n2 a_n20587_n5180.t7 541.395
R22777 a_n20587_n5180.n3 a_n20587_n5180.t4 527.402
R22778 a_n20587_n5180.n2 a_n20587_n5180.t5 491.64
R22779 a_n20587_n5180.n5 a_n20587_n5180.t0 281.906
R22780 a_n20587_n5180.t1 a_n20587_n5180.n5 204.359
R22781 a_n20587_n5180.n0 a_n20587_n5180.t2 180.73
R22782 a_n20587_n5180.n1 a_n20587_n5180.t6 179.45
R22783 a_n20587_n5180.n0 a_n20587_n5180.t3 139.78
R22784 a_n20587_n5180.n4 a_n20587_n5180.n1 105.635
R22785 a_n20587_n5180.n4 a_n20587_n5180.n3 76.0005
R22786 a_n20587_n5180.n5 a_n20587_n5180.n4 67.9685
R22787 a_n20587_n5180.n3 a_n20587_n5180.n2 13.994
R22788 a_n20587_n5180.n1 a_n20587_n5180.n0 1.28015
R22789 right_shifter_0.buffer_5.inv_1.A.n0 right_shifter_0.buffer_5.inv_1.A.t4 393.921
R22790 right_shifter_0.buffer_5.inv_1.A.n2 right_shifter_0.buffer_5.inv_1.A.t7 291.829
R22791 right_shifter_0.buffer_5.inv_1.A.n2 right_shifter_0.buffer_5.inv_1.A.t6 291.829
R22792 right_shifter_0.buffer_5.inv_1.A.n0 right_shifter_0.buffer_5.inv_1.A.t1 256.514
R22793 right_shifter_0.buffer_5.inv_1.A.n0 right_shifter_0.buffer_5.inv_1.A.n1 226.162
R22794 right_shifter_0.buffer_5.inv_1.A.n2 right_shifter_0.buffer_5.inv_1.A.t5 221.72
R22795 right_shifter_0.buffer_5.inv_1.A.n0 right_shifter_0.buffer_5.inv_1.A.t0 83.795
R22796 right_shifter_0.buffer_5.inv_1.A.n0 right_shifter_0.buffer_5.inv_1.A.n2 53.7938
R22797 right_shifter_0.buffer_5.inv_1.A.n1 right_shifter_0.buffer_5.inv_1.A.t3 30.379
R22798 right_shifter_0.buffer_5.inv_1.A.n1 right_shifter_0.buffer_5.inv_1.A.t2 30.379
R22799 right_shifter_0.S2.n1 right_shifter_0.S2.t6 1032.02
R22800 right_shifter_0.S2.n1 right_shifter_0.S2.t4 336.962
R22801 right_shifter_0.S2.n1 right_shifter_0.S2.t5 326.154
R22802 right_shifter_0.S2.n0 right_shifter_0.S2.t1 256.514
R22803 right_shifter_0.S2.n0 right_shifter_0.S2.n2 226.258
R22804 mux8_3.NAND4F_6.A right_shifter_0.S2.n1 162.952
R22805 right_shifter_0.S2.n0 right_shifter_0.S2.t0 83.7172
R22806 right_shifter_0.S2.n2 right_shifter_0.S2.t3 30.379
R22807 right_shifter_0.S2.n2 right_shifter_0.S2.t2 30.379
R22808 mux8_3.A7 right_shifter_0.S2.n0 25.5824
R22809 mux8_3.A7 mux8_3.NAND4F_6.A 13.4205
R22810 a_n17368_3810.n0 a_n17368_3810.n2 81.2978
R22811 a_n17368_3810.n1 a_n17368_3810.n6 81.1637
R22812 a_n17368_3810.n1 a_n17368_3810.n5 81.1637
R22813 a_n17368_3810.n0 a_n17368_3810.n4 81.1637
R22814 a_n17368_3810.n0 a_n17368_3810.n3 81.1637
R22815 a_n17368_3810.n7 a_n17368_3810.n1 80.9213
R22816 a_n17368_3810.n6 a_n17368_3810.t11 11.8205
R22817 a_n17368_3810.n6 a_n17368_3810.t0 11.8205
R22818 a_n17368_3810.n5 a_n17368_3810.t9 11.8205
R22819 a_n17368_3810.n5 a_n17368_3810.t10 11.8205
R22820 a_n17368_3810.n4 a_n17368_3810.t5 11.8205
R22821 a_n17368_3810.n4 a_n17368_3810.t3 11.8205
R22822 a_n17368_3810.n3 a_n17368_3810.t6 11.8205
R22823 a_n17368_3810.n3 a_n17368_3810.t4 11.8205
R22824 a_n17368_3810.n2 a_n17368_3810.t7 11.8205
R22825 a_n17368_3810.n2 a_n17368_3810.t8 11.8205
R22826 a_n17368_3810.n7 a_n17368_3810.t1 11.8205
R22827 a_n17368_3810.t2 a_n17368_3810.n7 11.8205
R22828 a_n17368_3810.n1 a_n17368_3810.n0 0.402735
R22829 a_n15131_n8419.n2 a_n15131_n8419.n0 121.353
R22830 a_n15131_n8419.n3 a_n15131_n8419.n2 121.353
R22831 a_n15131_n8419.n2 a_n15131_n8419.n1 121.001
R22832 a_n15131_n8419.n0 a_n15131_n8419.t2 30.462
R22833 a_n15131_n8419.n0 a_n15131_n8419.t0 30.462
R22834 a_n15131_n8419.n1 a_n15131_n8419.t3 30.462
R22835 a_n15131_n8419.n1 a_n15131_n8419.t1 30.462
R22836 a_n15131_n8419.n3 a_n15131_n8419.t5 30.462
R22837 a_n15131_n8419.t4 a_n15131_n8419.n3 30.462
R22838 a_n6641_1380.n2 a_n6641_1380.t3 541.395
R22839 a_n6641_1380.n3 a_n6641_1380.t5 527.402
R22840 a_n6641_1380.n2 a_n6641_1380.t7 491.64
R22841 a_n6641_1380.n5 a_n6641_1380.t0 281.906
R22842 a_n6641_1380.t1 a_n6641_1380.n5 204.359
R22843 a_n6641_1380.n0 a_n6641_1380.t4 180.73
R22844 a_n6641_1380.n1 a_n6641_1380.t6 179.45
R22845 a_n6641_1380.n0 a_n6641_1380.t2 139.78
R22846 a_n6641_1380.n4 a_n6641_1380.n1 105.635
R22847 a_n6641_1380.n4 a_n6641_1380.n3 76.0005
R22848 a_n6641_1380.n5 a_n6641_1380.n4 67.9685
R22849 a_n6641_1380.n3 a_n6641_1380.n2 13.994
R22850 a_n6641_1380.n1 a_n6641_1380.n0 1.28015
R22851 a_n6611_1406.n3 a_n6611_1406.n2 121.353
R22852 a_n6611_1406.n2 a_n6611_1406.n1 121.001
R22853 a_n6611_1406.n2 a_n6611_1406.n0 120.977
R22854 a_n6611_1406.n1 a_n6611_1406.t4 30.462
R22855 a_n6611_1406.n1 a_n6611_1406.t2 30.462
R22856 a_n6611_1406.n0 a_n6611_1406.t5 30.462
R22857 a_n6611_1406.n0 a_n6611_1406.t0 30.462
R22858 a_n6611_1406.t3 a_n6611_1406.n3 30.462
R22859 a_n6611_1406.n3 a_n6611_1406.t1 30.462
R22860 a_n4879_1406.n2 a_n4879_1406.n0 121.353
R22861 a_n4879_1406.n2 a_n4879_1406.n1 121.001
R22862 a_n4879_1406.n3 a_n4879_1406.n2 120.977
R22863 a_n4879_1406.n0 a_n4879_1406.t5 30.462
R22864 a_n4879_1406.n0 a_n4879_1406.t3 30.462
R22865 a_n4879_1406.n1 a_n4879_1406.t1 30.462
R22866 a_n4879_1406.n1 a_n4879_1406.t4 30.462
R22867 a_n4879_1406.t2 a_n4879_1406.n3 30.462
R22868 a_n4879_1406.n3 a_n4879_1406.t0 30.462
R22869 mux8_0.NAND4F_6.Y.n1 mux8_0.NAND4F_6.Y.t9 933.563
R22870 mux8_0.NAND4F_6.Y.n1 mux8_0.NAND4F_6.Y.t10 367.635
R22871 mux8_0.NAND4F_6.Y.n2 mux8_0.NAND4F_6.Y.t11 308.481
R22872 mux8_0.NAND4F_6.Y.n0 mux8_0.NAND4F_6.Y.n4 187.373
R22873 mux8_0.NAND4F_6.Y.n0 mux8_0.NAND4F_6.Y.n5 187.192
R22874 mux8_0.NAND4F_6.Y.n0 mux8_0.NAND4F_6.Y.n6 187.192
R22875 mux8_0.NAND4F_6.Y.n8 mux8_0.NAND4F_6.Y.n7 187.192
R22876 mux8_0.NAND4F_6.Y mux8_0.NAND4F_6.Y.n2 162.047
R22877 mux8_0.NAND4F_6.Y.n3 mux8_0.NAND4F_6.Y.t6 22.7831
R22878 mux8_0.NAND4F_6.Y.n3 mux8_0.NAND4F_6.Y 22.171
R22879 mux8_0.NAND4F_6.Y.n4 mux8_0.NAND4F_6.Y.t1 20.1899
R22880 mux8_0.NAND4F_6.Y.n4 mux8_0.NAND4F_6.Y.t0 20.1899
R22881 mux8_0.NAND4F_6.Y.n5 mux8_0.NAND4F_6.Y.t3 20.1899
R22882 mux8_0.NAND4F_6.Y.n5 mux8_0.NAND4F_6.Y.t2 20.1899
R22883 mux8_0.NAND4F_6.Y.n6 mux8_0.NAND4F_6.Y.t8 20.1899
R22884 mux8_0.NAND4F_6.Y.n6 mux8_0.NAND4F_6.Y.t7 20.1899
R22885 mux8_0.NAND4F_6.Y.n7 mux8_0.NAND4F_6.Y.t4 20.1899
R22886 mux8_0.NAND4F_6.Y.n7 mux8_0.NAND4F_6.Y.t5 20.1899
R22887 mux8_0.NAND4F_6.Y.n2 mux8_0.NAND4F_6.Y.n1 10.955
R22888 mux8_0.NAND4F_6.Y mux8_0.NAND4F_6.Y.n3 0.781576
R22889 mux8_0.NAND4F_6.Y mux8_0.NAND4F_6.Y.n8 0.396904
R22890 mux8_0.NAND4F_6.Y.n8 mux8_0.NAND4F_6.Y.n0 0.358709
R22891 a_7173_4939.t0 a_7173_4939.t1 19.8005
R22892 a_n17677_n22425.n0 a_n17677_n22425.n2 231.24
R22893 a_n17677_n22425.n6 a_n17677_n22425.n1 231.24
R22894 a_n17677_n22425.n0 a_n17677_n22425.n3 231.03
R22895 a_n17677_n22425.n1 a_n17677_n22425.n4 231.03
R22896 a_n17677_n22425.n1 a_n17677_n22425.n5 231.03
R22897 a_n17677_n22425.n2 a_n17677_n22425.t8 25.395
R22898 a_n17677_n22425.n2 a_n17677_n22425.t7 25.395
R22899 a_n17677_n22425.n3 a_n17677_n22425.t6 25.395
R22900 a_n17677_n22425.n3 a_n17677_n22425.t5 25.395
R22901 a_n17677_n22425.n4 a_n17677_n22425.t9 25.395
R22902 a_n17677_n22425.n4 a_n17677_n22425.t3 25.395
R22903 a_n17677_n22425.n5 a_n17677_n22425.t2 25.395
R22904 a_n17677_n22425.n5 a_n17677_n22425.t1 25.395
R22905 a_n17677_n22425.n6 a_n17677_n22425.t0 25.395
R22906 a_n17677_n22425.t4 a_n17677_n22425.n6 25.395
R22907 a_n17677_n22425.n1 a_n17677_n22425.n0 0.421553
R22908 a_n20587_n8445.n2 a_n20587_n8445.t2 541.395
R22909 a_n20587_n8445.n3 a_n20587_n8445.t5 527.402
R22910 a_n20587_n8445.n2 a_n20587_n8445.t6 491.64
R22911 a_n20587_n8445.n5 a_n20587_n8445.t0 281.906
R22912 a_n20587_n8445.t1 a_n20587_n8445.n5 204.359
R22913 a_n20587_n8445.n0 a_n20587_n8445.t3 180.73
R22914 a_n20587_n8445.n1 a_n20587_n8445.t7 179.45
R22915 a_n20587_n8445.n0 a_n20587_n8445.t4 139.78
R22916 a_n20587_n8445.n4 a_n20587_n8445.n1 105.635
R22917 a_n20587_n8445.n4 a_n20587_n8445.n3 76.0005
R22918 a_n20587_n8445.n5 a_n20587_n8445.n4 67.9685
R22919 a_n20587_n8445.n3 a_n20587_n8445.n2 13.994
R22920 a_n20587_n8445.n1 a_n20587_n8445.n0 1.28015
R22921 a_n20557_n7799.n0 a_n20557_n7799.n4 81.2978
R22922 a_n20557_n7799.n0 a_n20557_n7799.n5 81.1637
R22923 a_n20557_n7799.n0 a_n20557_n7799.n6 81.1637
R22924 a_n20557_n7799.n1 a_n20557_n7799.n3 81.1637
R22925 a_n20557_n7799.n7 a_n20557_n7799.n1 81.1637
R22926 a_n20557_n7799.n1 a_n20557_n7799.n2 80.9213
R22927 a_n20557_n7799.n4 a_n20557_n7799.t3 11.8205
R22928 a_n20557_n7799.n4 a_n20557_n7799.t5 11.8205
R22929 a_n20557_n7799.n5 a_n20557_n7799.t11 11.8205
R22930 a_n20557_n7799.n5 a_n20557_n7799.t4 11.8205
R22931 a_n20557_n7799.n6 a_n20557_n7799.t9 11.8205
R22932 a_n20557_n7799.n6 a_n20557_n7799.t10 11.8205
R22933 a_n20557_n7799.n3 a_n20557_n7799.t7 11.8205
R22934 a_n20557_n7799.n3 a_n20557_n7799.t1 11.8205
R22935 a_n20557_n7799.n2 a_n20557_n7799.t6 11.8205
R22936 a_n20557_n7799.n2 a_n20557_n7799.t8 11.8205
R22937 a_n20557_n7799.n7 a_n20557_n7799.t0 11.8205
R22938 a_n20557_n7799.t2 a_n20557_n7799.n7 11.8205
R22939 a_n20557_n7799.n1 a_n20557_n7799.n0 0.402735
R22940 mux8_1.NAND4F_3.Y.n7 mux8_1.NAND4F_3.Y.t11 978.795
R22941 mux8_1.NAND4F_3.Y.n6 mux8_1.NAND4F_3.Y.t9 308.481
R22942 mux8_1.NAND4F_3.Y.n6 mux8_1.NAND4F_3.Y.t10 308.481
R22943 mux8_1.NAND4F_3.Y.n0 mux8_1.NAND4F_3.Y.n1 187.373
R22944 mux8_1.NAND4F_3.Y.n0 mux8_1.NAND4F_3.Y.n2 187.192
R22945 mux8_1.NAND4F_3.Y.n0 mux8_1.NAND4F_3.Y.n3 187.192
R22946 mux8_1.NAND4F_3.Y.n5 mux8_1.NAND4F_3.Y.n4 187.192
R22947 mux8_1.NAND4F_3.Y mux8_1.NAND4F_3.Y.n7 161.839
R22948 mux8_1.NAND4F_3.Y mux8_1.NAND4F_3.Y.t2 23.4426
R22949 mux8_1.NAND4F_3.Y.n1 mux8_1.NAND4F_3.Y.t5 20.1899
R22950 mux8_1.NAND4F_3.Y.n1 mux8_1.NAND4F_3.Y.t6 20.1899
R22951 mux8_1.NAND4F_3.Y.n2 mux8_1.NAND4F_3.Y.t1 20.1899
R22952 mux8_1.NAND4F_3.Y.n2 mux8_1.NAND4F_3.Y.t0 20.1899
R22953 mux8_1.NAND4F_3.Y.n3 mux8_1.NAND4F_3.Y.t8 20.1899
R22954 mux8_1.NAND4F_3.Y.n3 mux8_1.NAND4F_3.Y.t7 20.1899
R22955 mux8_1.NAND4F_3.Y.n4 mux8_1.NAND4F_3.Y.t3 20.1899
R22956 mux8_1.NAND4F_3.Y.n4 mux8_1.NAND4F_3.Y.t4 20.1899
R22957 mux8_1.NAND4F_3.Y.n7 mux8_1.NAND4F_3.Y.n6 11.0463
R22958 mux8_1.NAND4F_3.Y mux8_1.NAND4F_3.Y.n5 0.518495
R22959 mux8_1.NAND4F_3.Y.n5 mux8_1.NAND4F_3.Y.n0 0.358709
R22960 OR8_0.S1.n1 OR8_0.S1.t4 1032.02
R22961 OR8_0.S1.n1 OR8_0.S1.t6 336.962
R22962 OR8_0.S1.n1 OR8_0.S1.t5 326.154
R22963 OR8_0.S1.n0 OR8_0.S1.t2 256.514
R22964 OR8_0.S1.n0 OR8_0.S1.n2 226.258
R22965 OR8_0.S1 OR8_0.S1.n1 162.952
R22966 OR8_0.S1.n0 OR8_0.S1.t3 83.7172
R22967 OR8_0.S1.n2 OR8_0.S1.t1 30.379
R22968 OR8_0.S1.n2 OR8_0.S1.t0 30.379
R22969 OR8_0.S1 OR8_0.S1.n0 1.9208
R22970 a_8592_n7266.t0 a_8592_n7266.t1 9.9005
R22971 mux8_2.NAND4F_2.Y.n6 mux8_2.NAND4F_2.Y.t9 933.563
R22972 mux8_2.NAND4F_2.Y.n6 mux8_2.NAND4F_2.Y.t11 367.635
R22973 mux8_2.NAND4F_2.Y.n7 mux8_2.NAND4F_2.Y.t10 308.481
R22974 mux8_2.NAND4F_2.Y.n0 mux8_2.NAND4F_2.Y.n1 187.373
R22975 mux8_2.NAND4F_2.Y.n0 mux8_2.NAND4F_2.Y.n2 187.192
R22976 mux8_2.NAND4F_2.Y.n0 mux8_2.NAND4F_2.Y.n3 187.192
R22977 mux8_2.NAND4F_2.Y.n5 mux8_2.NAND4F_2.Y.n4 187.192
R22978 mux8_2.NAND4F_2.Y mux8_2.NAND4F_2.Y.n7 162.102
R22979 mux8_2.NAND4F_2.Y.n8 mux8_2.NAND4F_2.Y.t6 22.7096
R22980 mux8_2.NAND4F_2.Y.n8 mux8_2.NAND4F_2.Y 22.4285
R22981 mux8_2.NAND4F_2.Y.n1 mux8_2.NAND4F_2.Y.t5 20.1899
R22982 mux8_2.NAND4F_2.Y.n1 mux8_2.NAND4F_2.Y.t4 20.1899
R22983 mux8_2.NAND4F_2.Y.n2 mux8_2.NAND4F_2.Y.t1 20.1899
R22984 mux8_2.NAND4F_2.Y.n2 mux8_2.NAND4F_2.Y.t0 20.1899
R22985 mux8_2.NAND4F_2.Y.n3 mux8_2.NAND4F_2.Y.t2 20.1899
R22986 mux8_2.NAND4F_2.Y.n3 mux8_2.NAND4F_2.Y.t3 20.1899
R22987 mux8_2.NAND4F_2.Y.n4 mux8_2.NAND4F_2.Y.t7 20.1899
R22988 mux8_2.NAND4F_2.Y.n4 mux8_2.NAND4F_2.Y.t8 20.1899
R22989 mux8_2.NAND4F_2.Y.n7 mux8_2.NAND4F_2.Y.n6 10.955
R22990 mux8_2.NAND4F_2.Y mux8_2.NAND4F_2.Y.n8 0.799394
R22991 mux8_2.NAND4F_2.Y mux8_2.NAND4F_2.Y.n5 0.452586
R22992 mux8_2.NAND4F_2.Y.n5 mux8_2.NAND4F_2.Y.n0 0.358709
R22993 a_11290_n7266.t0 a_11290_n7266.t1 9.9005
R22994 a_11386_n7266.t0 a_11386_n7266.t1 9.9005
R22995 a_3313_4914.n0 a_3313_4914.t4 539.788
R22996 a_3313_4914.n1 a_3313_4914.t2 531.496
R22997 a_3313_4914.n0 a_3313_4914.t5 490.034
R22998 a_3313_4914.n5 a_3313_4914.t0 283.788
R22999 a_3313_4914.t1 a_3313_4914.n5 205.489
R23000 a_3313_4914.n2 a_3313_4914.t7 182.625
R23001 a_3313_4914.n3 a_3313_4914.t6 179.054
R23002 a_3313_4914.n2 a_3313_4914.t3 139.78
R23003 a_3313_4914.n4 a_3313_4914.n3 101.368
R23004 a_3313_4914.n5 a_3313_4914.n4 77.9135
R23005 a_3313_4914.n4 a_3313_4914.n1 76.1557
R23006 a_3313_4914.n1 a_3313_4914.n0 8.29297
R23007 a_3313_4914.n3 a_3313_4914.n2 3.57087
R23008 a_n20737_n8419.n0 a_n20737_n8419.t4 539.788
R23009 a_n20737_n8419.n1 a_n20737_n8419.t6 531.496
R23010 a_n20737_n8419.n0 a_n20737_n8419.t5 490.034
R23011 a_n20737_n8419.n5 a_n20737_n8419.t0 283.788
R23012 a_n20737_n8419.t1 a_n20737_n8419.n5 205.489
R23013 a_n20737_n8419.n2 a_n20737_n8419.t7 182.625
R23014 a_n20737_n8419.n3 a_n20737_n8419.t3 179.054
R23015 a_n20737_n8419.n2 a_n20737_n8419.t2 139.78
R23016 a_n20737_n8419.n4 a_n20737_n8419.n3 101.368
R23017 a_n20737_n8419.n5 a_n20737_n8419.n4 77.9135
R23018 a_n20737_n8419.n4 a_n20737_n8419.n1 76.1557
R23019 a_n20737_n8419.n1 a_n20737_n8419.n0 8.29297
R23020 a_n20737_n8419.n3 a_n20737_n8419.n2 3.57087
R23021 a_n20557_n8419.n2 a_n20557_n8419.n1 121.353
R23022 a_n20557_n8419.n3 a_n20557_n8419.n2 121.001
R23023 a_n20557_n8419.n2 a_n20557_n8419.n0 120.977
R23024 a_n20557_n8419.n1 a_n20557_n8419.t1 30.462
R23025 a_n20557_n8419.n1 a_n20557_n8419.t0 30.462
R23026 a_n20557_n8419.n0 a_n20557_n8419.t3 30.462
R23027 a_n20557_n8419.n0 a_n20557_n8419.t5 30.462
R23028 a_n20557_n8419.n3 a_n20557_n8419.t4 30.462
R23029 a_n20557_n8419.t2 a_n20557_n8419.n3 30.462
R23030 a_n368_3164.n0 a_n368_3164.t3 539.788
R23031 a_n368_3164.n1 a_n368_3164.t7 531.496
R23032 a_n368_3164.n0 a_n368_3164.t5 490.034
R23033 a_n368_3164.n5 a_n368_3164.t0 283.788
R23034 a_n368_3164.t1 a_n368_3164.n5 205.489
R23035 a_n368_3164.n2 a_n368_3164.t2 182.625
R23036 a_n368_3164.n3 a_n368_3164.t6 179.054
R23037 a_n368_3164.n2 a_n368_3164.t4 139.78
R23038 a_n368_3164.n4 a_n368_3164.n3 101.368
R23039 a_n368_3164.n5 a_n368_3164.n4 77.9135
R23040 a_n368_3164.n4 a_n368_3164.n1 76.1557
R23041 a_n368_3164.n1 a_n368_3164.n0 8.29297
R23042 a_n368_3164.n3 a_n368_3164.n2 3.57087
R23043 a_8400_n25478.t0 a_8400_n25478.t1 9.9005
R23044 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t16 491.64
R23045 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t12 491.64
R23046 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t21 491.64
R23047 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t14 491.64
R23048 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t15 485.221
R23049 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t19 367.928
R23050 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t23 255.588
R23051 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t13 224.478
R23052 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n15 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t18 213.688
R23053 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n19 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n18 209.19
R23054 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t20 139.78
R23055 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t22 139.78
R23056 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n18 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t17 139.78
R23057 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n1 120.999
R23058 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n2 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n0 120.999
R23059 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n13 104.489
R23060 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 103.258
R23061 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n3 92.5005
R23062 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n8 86.2638
R23063 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n9 85.8873
R23064 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n9 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n6 85.724
R23065 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n17 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n16 84.5046
R23066 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n14 84.0545
R23067 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n11 75.0672
R23068 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n12 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n8 75.0672
R23069 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n11 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n10 73.1255
R23070 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n8 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n7 73.1255
R23071 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n6 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n5 73.1255
R23072 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n16 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n15 72.3005
R23073 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n6 68.8946
R23074 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n17 60.9816
R23075 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n14 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n4 41.9827
R23076 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t5 30.462
R23077 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n3 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t9 30.462
R23078 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t10 30.462
R23079 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n1 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t11 30.462
R23080 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t3 30.462
R23081 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t4 30.462
R23082 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n4 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n2 28.124
R23083 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n20 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n19 17.8661
R23084 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n21 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n20 17.8661
R23085 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n22 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n21 17.1217
R23086 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n23 15.6329
R23087 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t6 11.8205
R23088 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n7 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t7 11.8205
R23089 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t1 11.8205
R23090 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n10 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t0 11.8205
R23091 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t8 11.8205
R23092 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n5 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t2 11.8205
R23093 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n24 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 10.8165
R23094 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n13 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n12 9.3005
R23095 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n24 2.50602
R23096 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n23 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n22 1.8615
R23097 a_n338_3190.n2 a_n338_3190.n0 121.353
R23098 a_n338_3190.n2 a_n338_3190.n1 121.001
R23099 a_n338_3190.n3 a_n338_3190.n2 120.977
R23100 a_n338_3190.n1 a_n338_3190.t2 30.462
R23101 a_n338_3190.n1 a_n338_3190.t3 30.462
R23102 a_n338_3190.n0 a_n338_3190.t1 30.462
R23103 a_n338_3190.n0 a_n338_3190.t0 30.462
R23104 a_n338_3190.t4 a_n338_3190.n3 30.462
R23105 a_n338_3190.n3 a_n338_3190.t5 30.462
R23106 a_n9931_1380.n2 a_n9931_1380.t5 541.395
R23107 a_n9931_1380.n3 a_n9931_1380.t2 527.402
R23108 a_n9931_1380.n2 a_n9931_1380.t7 491.64
R23109 a_n9931_1380.n5 a_n9931_1380.t0 281.906
R23110 a_n9931_1380.t1 a_n9931_1380.n5 204.359
R23111 a_n9931_1380.n0 a_n9931_1380.t6 180.73
R23112 a_n9931_1380.n1 a_n9931_1380.t3 179.45
R23113 a_n9931_1380.n0 a_n9931_1380.t4 139.78
R23114 a_n9931_1380.n4 a_n9931_1380.n1 105.635
R23115 a_n9931_1380.n4 a_n9931_1380.n3 76.0005
R23116 a_n9931_1380.n5 a_n9931_1380.n4 67.9685
R23117 a_n9931_1380.n3 a_n9931_1380.n2 13.994
R23118 a_n9931_1380.n1 a_n9931_1380.n0 1.28015
R23119 a_n9901_2026.n0 a_n9901_2026.n3 81.2978
R23120 a_n9901_2026.n0 a_n9901_2026.n4 81.1637
R23121 a_n9901_2026.n0 a_n9901_2026.n5 81.1637
R23122 a_n9901_2026.n1 a_n9901_2026.n6 81.1637
R23123 a_n9901_2026.n7 a_n9901_2026.n1 81.1637
R23124 a_n9901_2026.n1 a_n9901_2026.n2 80.9213
R23125 a_n9901_2026.n3 a_n9901_2026.t7 11.8205
R23126 a_n9901_2026.n3 a_n9901_2026.t8 11.8205
R23127 a_n9901_2026.n4 a_n9901_2026.t10 11.8205
R23128 a_n9901_2026.n4 a_n9901_2026.t6 11.8205
R23129 a_n9901_2026.n5 a_n9901_2026.t11 11.8205
R23130 a_n9901_2026.n5 a_n9901_2026.t9 11.8205
R23131 a_n9901_2026.n6 a_n9901_2026.t0 11.8205
R23132 a_n9901_2026.n6 a_n9901_2026.t1 11.8205
R23133 a_n9901_2026.n2 a_n9901_2026.t3 11.8205
R23134 a_n9901_2026.n2 a_n9901_2026.t4 11.8205
R23135 a_n9901_2026.n7 a_n9901_2026.t5 11.8205
R23136 a_n9901_2026.t2 a_n9901_2026.n7 11.8205
R23137 a_n9901_2026.n1 a_n9901_2026.n0 0.402735
R23138 a_n20737_n5154.n0 a_n20737_n5154.t5 539.788
R23139 a_n20737_n5154.n1 a_n20737_n5154.t7 531.496
R23140 a_n20737_n5154.n0 a_n20737_n5154.t6 490.034
R23141 a_n20737_n5154.n5 a_n20737_n5154.t0 283.788
R23142 a_n20737_n5154.t1 a_n20737_n5154.n5 205.489
R23143 a_n20737_n5154.n2 a_n20737_n5154.t2 182.625
R23144 a_n20737_n5154.n3 a_n20737_n5154.t4 179.054
R23145 a_n20737_n5154.n2 a_n20737_n5154.t3 139.78
R23146 a_n20737_n5154.n4 a_n20737_n5154.n3 101.368
R23147 a_n20737_n5154.n5 a_n20737_n5154.n4 77.9135
R23148 a_n20737_n5154.n4 a_n20737_n5154.n1 76.1557
R23149 a_n20737_n5154.n1 a_n20737_n5154.n0 8.29297
R23150 a_n20737_n5154.n3 a_n20737_n5154.n2 3.57087
R23151 a_n20557_n5154.n3 a_n20557_n5154.n2 121.353
R23152 a_n20557_n5154.n2 a_n20557_n5154.n1 121.001
R23153 a_n20557_n5154.n2 a_n20557_n5154.n0 120.977
R23154 a_n20557_n5154.n1 a_n20557_n5154.t0 30.462
R23155 a_n20557_n5154.n1 a_n20557_n5154.t5 30.462
R23156 a_n20557_n5154.n0 a_n20557_n5154.t2 30.462
R23157 a_n20557_n5154.n0 a_n20557_n5154.t1 30.462
R23158 a_n20557_n5154.t4 a_n20557_n5154.n3 30.462
R23159 a_n20557_n5154.n3 a_n20557_n5154.t3 30.462
R23160 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t22 491.64
R23161 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t23 491.64
R23162 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t12 491.64
R23163 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t20 491.64
R23164 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n8 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t18 485.221
R23165 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t13 367.928
R23166 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t16 255.588
R23167 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t21 224.478
R23168 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t14 213.688
R23169 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n0 209.19
R23170 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t17 139.78
R23171 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t15 139.78
R23172 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t19 139.78
R23173 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n11 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n10 120.999
R23174 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n11 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n9 120.999
R23175 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n23 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n22 104.489
R23176 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n13 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n12 92.5005
R23177 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n20 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n18 86.2638
R23178 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n18 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n17 85.8873
R23179 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n18 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n15 85.724
R23180 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n8 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n7 84.5046
R23181 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n23 83.8907
R23182 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n21 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n20 75.0672
R23183 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n21 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n17 75.0672
R23184 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n20 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n19 73.1255
R23185 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n17 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n16 73.1255
R23186 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n15 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n14 73.1255
R23187 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n6 72.3005
R23188 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n22 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n15 68.8946
R23189 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n8 60.9797
R23190 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n23 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n13 41.9827
R23191 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n12 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t9 30.462
R23192 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n12 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t2 30.462
R23193 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n10 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t1 30.462
R23194 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n10 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t0 30.462
R23195 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n9 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t11 30.462
R23196 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n9 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t10 30.462
R23197 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n13 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n11 28.124
R23198 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n5 19.963
R23199 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n1 17.8661
R23200 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n2 17.8661
R23201 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n3 17.1217
R23202 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n16 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t8 11.8205
R23203 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n16 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t7 11.8205
R23204 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n19 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t4 11.8205
R23205 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n19 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t3 11.8205
R23206 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n14 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t6 11.8205
R23207 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n14 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t5 11.8205
R23208 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n22 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n21 9.3005
R23209 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n4 1.8615
R23210 a_n11274_n23075.n2 a_n11274_n23075.n0 121.353
R23211 a_n11274_n23075.n3 a_n11274_n23075.n2 121.353
R23212 a_n11274_n23075.n2 a_n11274_n23075.n1 121.001
R23213 a_n11274_n23075.n1 a_n11274_n23075.t0 30.462
R23214 a_n11274_n23075.n1 a_n11274_n23075.t3 30.462
R23215 a_n11274_n23075.n0 a_n11274_n23075.t5 30.462
R23216 a_n11274_n23075.n0 a_n11274_n23075.t4 30.462
R23217 a_n11274_n23075.t2 a_n11274_n23075.n3 30.462
R23218 a_n11274_n23075.n3 a_n11274_n23075.t1 30.462
R23219 AND8_0.S3.n1 AND8_0.S3.t6 1032.02
R23220 AND8_0.S3.n1 AND8_0.S3.t4 336.962
R23221 AND8_0.S3.n1 AND8_0.S3.t5 326.154
R23222 AND8_0.S3.n0 AND8_0.S3.t3 256.514
R23223 AND8_0.S3.n0 AND8_0.S3.n2 226.258
R23224 AND8_0.S3 AND8_0.S3.n1 162.945
R23225 AND8_0.S3.n0 AND8_0.S3.t0 83.7172
R23226 AND8_0.S3.n2 AND8_0.S3.t1 30.379
R23227 AND8_0.S3.n2 AND8_0.S3.t2 30.379
R23228 AND8_0.S3 AND8_0.S3.n0 1.92801
R23229 a_n13222_1380.n2 a_n13222_1380.t3 541.395
R23230 a_n13222_1380.n3 a_n13222_1380.t2 527.402
R23231 a_n13222_1380.n2 a_n13222_1380.t5 491.64
R23232 a_n13222_1380.n5 a_n13222_1380.t0 281.906
R23233 a_n13222_1380.t1 a_n13222_1380.n5 204.359
R23234 a_n13222_1380.n0 a_n13222_1380.t7 180.73
R23235 a_n13222_1380.n1 a_n13222_1380.t4 179.45
R23236 a_n13222_1380.n0 a_n13222_1380.t6 139.78
R23237 a_n13222_1380.n4 a_n13222_1380.n1 105.635
R23238 a_n13222_1380.n4 a_n13222_1380.n3 76.0005
R23239 a_n13222_1380.n5 a_n13222_1380.n4 67.9685
R23240 a_n13222_1380.n3 a_n13222_1380.n2 13.994
R23241 a_n13222_1380.n1 a_n13222_1380.n0 1.28015
R23242 mux8_1.NAND4F_4.Y.n6 mux8_1.NAND4F_4.Y.t9 1032.02
R23243 mux8_1.NAND4F_4.Y.n6 mux8_1.NAND4F_4.Y.t11 336.962
R23244 mux8_1.NAND4F_4.Y.n6 mux8_1.NAND4F_4.Y.t10 326.154
R23245 mux8_1.NAND4F_4.Y.n0 mux8_1.NAND4F_4.Y.n1 187.373
R23246 mux8_1.NAND4F_4.Y.n0 mux8_1.NAND4F_4.Y.n2 187.192
R23247 mux8_1.NAND4F_4.Y.n0 mux8_1.NAND4F_4.Y.n3 187.192
R23248 mux8_1.NAND4F_4.Y.n5 mux8_1.NAND4F_4.Y.n4 187.192
R23249 mux8_1.NAND4F_4.Y mux8_1.NAND4F_4.Y.n6 162.942
R23250 mux8_1.NAND4F_4.Y.n7 mux8_1.NAND4F_4.Y 24.5377
R23251 mux8_1.NAND4F_4.Y.n7 mux8_1.NAND4F_4.Y.t0 22.6141
R23252 mux8_1.NAND4F_4.Y.n1 mux8_1.NAND4F_4.Y.t3 20.1899
R23253 mux8_1.NAND4F_4.Y.n1 mux8_1.NAND4F_4.Y.t4 20.1899
R23254 mux8_1.NAND4F_4.Y.n2 mux8_1.NAND4F_4.Y.t5 20.1899
R23255 mux8_1.NAND4F_4.Y.n2 mux8_1.NAND4F_4.Y.t6 20.1899
R23256 mux8_1.NAND4F_4.Y.n3 mux8_1.NAND4F_4.Y.t7 20.1899
R23257 mux8_1.NAND4F_4.Y.n3 mux8_1.NAND4F_4.Y.t8 20.1899
R23258 mux8_1.NAND4F_4.Y.n4 mux8_1.NAND4F_4.Y.t1 20.1899
R23259 mux8_1.NAND4F_4.Y.n4 mux8_1.NAND4F_4.Y.t2 20.1899
R23260 mux8_1.NAND4F_4.Y mux8_1.NAND4F_4.Y.n7 0.894894
R23261 mux8_1.NAND4F_4.Y mux8_1.NAND4F_4.Y.n5 0.452586
R23262 mux8_1.NAND4F_4.Y.n5 mux8_1.NAND4F_4.Y.n0 0.358709
R23263 a_n7496_3190.n2 a_n7496_3190.n1 121.353
R23264 a_n7496_3190.n2 a_n7496_3190.n0 121.353
R23265 a_n7496_3190.n3 a_n7496_3190.n2 121.001
R23266 a_n7496_3190.n1 a_n7496_3190.t0 30.462
R23267 a_n7496_3190.n1 a_n7496_3190.t1 30.462
R23268 a_n7496_3190.n0 a_n7496_3190.t3 30.462
R23269 a_n7496_3190.n0 a_n7496_3190.t4 30.462
R23270 a_n7496_3190.n3 a_n7496_3190.t5 30.462
R23271 a_n7496_3190.t2 a_n7496_3190.n3 30.462
R23272 a_n16663_1406.n0 a_n16663_1406.t5 539.788
R23273 a_n16663_1406.n1 a_n16663_1406.t7 531.496
R23274 a_n16663_1406.n0 a_n16663_1406.t2 490.034
R23275 a_n16663_1406.n5 a_n16663_1406.t0 283.788
R23276 a_n16663_1406.t1 a_n16663_1406.n5 205.489
R23277 a_n16663_1406.n2 a_n16663_1406.t3 182.625
R23278 a_n16663_1406.n3 a_n16663_1406.t4 179.054
R23279 a_n16663_1406.n2 a_n16663_1406.t6 139.78
R23280 a_n16663_1406.n4 a_n16663_1406.n3 101.368
R23281 a_n16663_1406.n5 a_n16663_1406.n4 77.9135
R23282 a_n16663_1406.n4 a_n16663_1406.n1 76.1557
R23283 a_n16663_1406.n1 a_n16663_1406.n0 8.29297
R23284 a_n16663_1406.n3 a_n16663_1406.n2 3.57087
R23285 a_n17677_n19625.n0 a_n17677_n19625.n2 231.24
R23286 a_n17677_n19625.n1 a_n17677_n19625.n4 231.24
R23287 a_n17677_n19625.n0 a_n17677_n19625.n3 231.03
R23288 a_n17677_n19625.n1 a_n17677_n19625.n5 231.03
R23289 a_n17677_n19625.n6 a_n17677_n19625.n1 231.03
R23290 a_n17677_n19625.n2 a_n17677_n19625.t3 25.395
R23291 a_n17677_n19625.n2 a_n17677_n19625.t2 25.395
R23292 a_n17677_n19625.n3 a_n17677_n19625.t1 25.395
R23293 a_n17677_n19625.n3 a_n17677_n19625.t0 25.395
R23294 a_n17677_n19625.n5 a_n17677_n19625.t7 25.395
R23295 a_n17677_n19625.n5 a_n17677_n19625.t6 25.395
R23296 a_n17677_n19625.n4 a_n17677_n19625.t5 25.395
R23297 a_n17677_n19625.n4 a_n17677_n19625.t9 25.395
R23298 a_n17677_n19625.t4 a_n17677_n19625.n6 25.395
R23299 a_n17677_n19625.n6 a_n17677_n19625.t8 25.395
R23300 a_n17677_n19625.n1 a_n17677_n19625.n0 0.421553
R23301 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t7 540.38
R23302 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t10 367.928
R23303 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n5 227.526
R23304 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t8 227.356
R23305 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n6 227.266
R23306 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n4 227.266
R23307 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t9 213.688
R23308 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n2 160.439
R23309 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n1 94.4341
R23310 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t3 42.7944
R23311 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t6 30.379
R23312 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t1 30.379
R23313 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t4 30.379
R23314 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t5 30.379
R23315 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t2 30.379
R23316 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.t0 30.379
R23317 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n0 13.4358
R23318 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B.n3 0.821842
R23319 A4.n5 A4.t0 540.38
R23320 A4.n13 A4.t7 540.375
R23321 A4.n6 A4.t26 491.64
R23322 A4.n6 A4.t6 491.64
R23323 A4.n6 A4.t20 491.64
R23324 A4.n6 A4.t14 491.64
R23325 A4.n1 A4.t23 491.64
R23326 A4.n1 A4.t25 491.64
R23327 A4.n1 A4.t21 491.64
R23328 A4.n1 A4.t4 491.64
R23329 A4.n3 A4.t1 367.928
R23330 A4.n11 A4.t5 343.827
R23331 A4.n16 A4.t17 312.599
R23332 A4.n19 A4.t12 247.428
R23333 A4.n18 A4.t29 247.428
R23334 A4.n17 A4.t27 247.428
R23335 A4.n16 A4.t18 247.428
R23336 A4.n11 A4.t15 237.787
R23337 A4.n20 A4.t10 229.754
R23338 A4.n12 A4.t24 227.356
R23339 A4.n4 A4.t2 227.356
R23340 A4.n3 A4.t3 213.688
R23341 A4 A4.n2 163.036
R23342 A4.n9 A4.n8 162.867
R23343 A4 A4.n20 162.409
R23344 A4.n5 A4.n4 160.439
R23345 A4.n13 A4.n12 160.433
R23346 A4.n7 A4.t9 139.78
R23347 A4.n7 A4.t28 139.78
R23348 A4.n7 A4.t16 139.78
R23349 A4.n7 A4.t22 139.78
R23350 A4.n0 A4.t8 139.78
R23351 A4.n0 A4.t19 139.78
R23352 A4.n0 A4.t11 139.78
R23353 A4.n0 A4.t13 139.78
R23354 A4.n4 A4.n3 94.4341
R23355 A4.n20 A4.n19 91.5805
R23356 A4.n12 A4.n11 70.3341
R23357 A4.n17 A4.n16 65.1723
R23358 A4.n18 A4.n17 65.1723
R23359 A4.n19 A4.n18 65.1723
R23360 A4.n2 A4.n0 38.8368
R23361 A4.n8 A4.n7 38.6833
R23362 A4.n8 A4.n6 28.3986
R23363 A4.n2 A4.n1 28.2451
R23364 A4 A4.n22 20.476
R23365 A4 A4.n10 18.1908
R23366 A4.n15 A4.n14 12.4105
R23367 A4.n22 A4.n21 12.4105
R23368 A4.n10 A4.n9 9.00496
R23369 A4.n22 A4.n15 4.17016
R23370 A4.n10 A4 3.87912
R23371 A4.n21 A4 1.49721
R23372 A4.n14 A4 1.34555
R23373 A4 A4.n13 0.905186
R23374 A4 A4.n5 0.89693
R23375 A4.n14 A4 0.0770306
R23376 A4.n9 A4 0.0590664
R23377 A4.n15 A4 0.0133182
R23378 A4.n21 A4 0.0115294
R23379 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t7 540.38
R23380 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t8 367.928
R23381 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n4 227.526
R23382 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t9 227.356
R23383 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n5 227.266
R23384 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n6 227.266
R23385 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t10 213.688
R23386 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n2 160.439
R23387 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n1 94.4341
R23388 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t0 42.7944
R23389 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t5 30.379
R23390 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t6 30.379
R23391 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t2 30.379
R23392 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t4 30.379
R23393 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t3 30.379
R23394 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.t1 30.379
R23395 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n0 13.4358
R23396 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B.n3 0.821842
R23397 a_n12446_n5180.n2 a_n12446_n5180.t2 541.395
R23398 a_n12446_n5180.n3 a_n12446_n5180.t4 527.402
R23399 a_n12446_n5180.n2 a_n12446_n5180.t5 491.64
R23400 a_n12446_n5180.n5 a_n12446_n5180.t0 281.906
R23401 a_n12446_n5180.t1 a_n12446_n5180.n5 204.359
R23402 a_n12446_n5180.n0 a_n12446_n5180.t3 180.73
R23403 a_n12446_n5180.n1 a_n12446_n5180.t7 179.45
R23404 a_n12446_n5180.n0 a_n12446_n5180.t6 139.78
R23405 a_n12446_n5180.n4 a_n12446_n5180.n1 105.635
R23406 a_n12446_n5180.n4 a_n12446_n5180.n3 76.0005
R23407 a_n12446_n5180.n5 a_n12446_n5180.n4 67.9685
R23408 a_n12446_n5180.n3 a_n12446_n5180.n2 13.994
R23409 a_n12446_n5180.n1 a_n12446_n5180.n0 1.28015
R23410 MULT_0.4bit_ADDER_1.B0.n4 MULT_0.4bit_ADDER_1.B0.t21 491.64
R23411 MULT_0.4bit_ADDER_1.B0.n5 MULT_0.4bit_ADDER_1.B0.t14 491.64
R23412 MULT_0.4bit_ADDER_1.B0.n6 MULT_0.4bit_ADDER_1.B0.t16 491.64
R23413 MULT_0.4bit_ADDER_1.B0.n7 MULT_0.4bit_ADDER_1.B0.t22 491.64
R23414 MULT_0.4bit_ADDER_1.B0.n2 MULT_0.4bit_ADDER_1.B0.t19 485.221
R23415 MULT_0.4bit_ADDER_1.B0.n0 MULT_0.4bit_ADDER_1.B0.t12 367.928
R23416 MULT_0.4bit_ADDER_1.B0.n8 MULT_0.4bit_ADDER_1.B0.t18 255.588
R23417 MULT_0.4bit_ADDER_1.B0.n1 MULT_0.4bit_ADDER_1.B0.t15 224.478
R23418 MULT_0.4bit_ADDER_1.B0.n0 MULT_0.4bit_ADDER_1.B0.t13 213.688
R23419 MULT_0.4bit_ADDER_1.B0.n4 MULT_0.4bit_ADDER_1.B0.n3 209.19
R23420 MULT_0.4bit_ADDER_1.B0.n3 MULT_0.4bit_ADDER_1.B0.t17 139.78
R23421 MULT_0.4bit_ADDER_1.B0.n3 MULT_0.4bit_ADDER_1.B0.t23 139.78
R23422 MULT_0.4bit_ADDER_1.B0.n3 MULT_0.4bit_ADDER_1.B0.t20 139.78
R23423 MULT_0.4bit_ADDER_1.B0.n12 MULT_0.4bit_ADDER_1.B0.n11 120.999
R23424 MULT_0.4bit_ADDER_1.B0.n12 MULT_0.4bit_ADDER_1.B0.n10 120.999
R23425 MULT_0.4bit_ADDER_1.B0.n24 MULT_0.4bit_ADDER_1.B0.n23 104.489
R23426 MULT_0.4bit_ADDER_1.B0.n9 MULT_0.4bit_ADDER_1.B0 103.258
R23427 MULT_0.4bit_ADDER_1.B0.n14 MULT_0.4bit_ADDER_1.B0.n13 92.5005
R23428 MULT_0.4bit_ADDER_1.B0.n21 MULT_0.4bit_ADDER_1.B0.n19 86.2638
R23429 MULT_0.4bit_ADDER_1.B0.n19 MULT_0.4bit_ADDER_1.B0.n18 85.8873
R23430 MULT_0.4bit_ADDER_1.B0.n19 MULT_0.4bit_ADDER_1.B0.n16 85.724
R23431 MULT_0.4bit_ADDER_1.B0.n2 MULT_0.4bit_ADDER_1.B0.n1 84.5046
R23432 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_1.B0.n24 83.8907
R23433 MULT_0.4bit_ADDER_1.B0.n22 MULT_0.4bit_ADDER_1.B0.n21 75.0672
R23434 MULT_0.4bit_ADDER_1.B0.n22 MULT_0.4bit_ADDER_1.B0.n18 75.0672
R23435 MULT_0.4bit_ADDER_1.B0.n21 MULT_0.4bit_ADDER_1.B0.n20 73.1255
R23436 MULT_0.4bit_ADDER_1.B0.n18 MULT_0.4bit_ADDER_1.B0.n17 73.1255
R23437 MULT_0.4bit_ADDER_1.B0.n16 MULT_0.4bit_ADDER_1.B0.n15 73.1255
R23438 MULT_0.4bit_ADDER_1.B0.n1 MULT_0.4bit_ADDER_1.B0.n0 72.3005
R23439 MULT_0.4bit_ADDER_1.B0.n23 MULT_0.4bit_ADDER_1.B0.n16 68.8946
R23440 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_1.B0.n2 60.9816
R23441 MULT_0.4bit_ADDER_1.B0.n24 MULT_0.4bit_ADDER_1.B0.n14 41.9827
R23442 MULT_0.4bit_ADDER_1.B0.n13 MULT_0.4bit_ADDER_1.B0.t9 30.462
R23443 MULT_0.4bit_ADDER_1.B0.n13 MULT_0.4bit_ADDER_1.B0.t2 30.462
R23444 MULT_0.4bit_ADDER_1.B0.n11 MULT_0.4bit_ADDER_1.B0.t1 30.462
R23445 MULT_0.4bit_ADDER_1.B0.n11 MULT_0.4bit_ADDER_1.B0.t8 30.462
R23446 MULT_0.4bit_ADDER_1.B0.n10 MULT_0.4bit_ADDER_1.B0.t11 30.462
R23447 MULT_0.4bit_ADDER_1.B0.n10 MULT_0.4bit_ADDER_1.B0.t10 30.462
R23448 MULT_0.4bit_ADDER_1.B0.n14 MULT_0.4bit_ADDER_1.B0.n12 28.124
R23449 MULT_0.4bit_ADDER_1.B0.n5 MULT_0.4bit_ADDER_1.B0.n4 17.8661
R23450 MULT_0.4bit_ADDER_1.B0.n6 MULT_0.4bit_ADDER_1.B0.n5 17.8661
R23451 MULT_0.4bit_ADDER_1.B0.n7 MULT_0.4bit_ADDER_1.B0.n6 17.1217
R23452 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_1.B0.n8 15.6329
R23453 MULT_0.4bit_ADDER_1.B0.n17 MULT_0.4bit_ADDER_1.B0.t4 11.8205
R23454 MULT_0.4bit_ADDER_1.B0.n17 MULT_0.4bit_ADDER_1.B0.t3 11.8205
R23455 MULT_0.4bit_ADDER_1.B0.n20 MULT_0.4bit_ADDER_1.B0.t6 11.8205
R23456 MULT_0.4bit_ADDER_1.B0.n20 MULT_0.4bit_ADDER_1.B0.t0 11.8205
R23457 MULT_0.4bit_ADDER_1.B0.n15 MULT_0.4bit_ADDER_1.B0.t5 11.8205
R23458 MULT_0.4bit_ADDER_1.B0.n15 MULT_0.4bit_ADDER_1.B0.t7 11.8205
R23459 MULT_0.4bit_ADDER_1.B0.n9 MULT_0.4bit_ADDER_1.B0 10.8165
R23460 MULT_0.4bit_ADDER_1.B0.n23 MULT_0.4bit_ADDER_1.B0.n22 9.3005
R23461 MULT_0.4bit_ADDER_1.B0.n8 MULT_0.4bit_ADDER_1.B0.n7 1.8615
R23462 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_1.B0.n9 0.855699
R23463 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t10 485.221
R23464 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t7 367.928
R23465 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n5 227.526
R23466 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n4 227.266
R23467 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n6 227.266
R23468 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t9 224.478
R23469 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t8 213.688
R23470 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n2 84.5046
R23471 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n1 72.3005
R23472 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n3 61.0566
R23473 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t6 42.7747
R23474 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t1 30.379
R23475 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t0 30.379
R23476 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t5 30.379
R23477 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t4 30.379
R23478 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t3 30.379
R23479 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.t2 30.379
R23480 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A.n0 0.583137
R23481 mux8_0.NAND4F_4.B.n10 mux8_0.NAND4F_4.B.t11 933.563
R23482 mux8_0.NAND4F_4.B.n5 mux8_0.NAND4F_4.B.t5 933.563
R23483 mux8_0.NAND4F_4.B.n3 mux8_0.NAND4F_4.B.t7 933.563
R23484 mux8_0.NAND4F_4.B.n1 mux8_0.NAND4F_4.B.t13 933.563
R23485 mux8_0.NAND4F_4.B.n10 mux8_0.NAND4F_4.B.t6 367.635
R23486 mux8_0.NAND4F_4.B.n5 mux8_0.NAND4F_4.B.t9 367.635
R23487 mux8_0.NAND4F_4.B.n3 mux8_0.NAND4F_4.B.t12 367.635
R23488 mux8_0.NAND4F_4.B.n1 mux8_0.NAND4F_4.B.t15 367.635
R23489 mux8_0.NAND4F_4.B.n11 mux8_0.NAND4F_4.B.t8 308.481
R23490 mux8_0.NAND4F_4.B.n6 mux8_0.NAND4F_4.B.t10 308.481
R23491 mux8_0.NAND4F_4.B.n4 mux8_0.NAND4F_4.B.t14 308.481
R23492 mux8_0.NAND4F_4.B.n2 mux8_0.NAND4F_4.B.t4 308.481
R23493 mux8_0.NAND4F_4.B.n0 mux8_0.NAND4F_4.B.t2 256.514
R23494 mux8_0.NAND4F_4.B.n0 mux8_0.NAND4F_4.B.n8 226.258
R23495 mux8_0.NAND4F_4.B mux8_0.NAND4F_4.B.n2 162.173
R23496 mux8_0.NAND4F_4.B mux8_0.NAND4F_4.B.n6 162.137
R23497 mux8_0.NAND4F_4.B mux8_0.NAND4F_4.B.n11 162.117
R23498 mux8_0.NAND4F_4.B.n7 mux8_0.NAND4F_4.B.n4 161.703
R23499 mux8_0.NAND4F_4.B.n0 mux8_0.NAND4F_4.B.t0 83.7172
R23500 mux8_0.NAND4F_4.B.n8 mux8_0.NAND4F_4.B.t3 30.379
R23501 mux8_0.NAND4F_4.B.n8 mux8_0.NAND4F_4.B.t1 30.379
R23502 mux8_0.NAND4F_4.B.n12 mux8_0.NAND4F_4.B 24.8912
R23503 mux8_0.NAND4F_4.B.n7 mux8_0.NAND4F_4.B 21.6618
R23504 mux8_0.NAND4F_4.B.n11 mux8_0.NAND4F_4.B.n10 10.955
R23505 mux8_0.NAND4F_4.B.n6 mux8_0.NAND4F_4.B.n5 10.955
R23506 mux8_0.NAND4F_4.B.n4 mux8_0.NAND4F_4.B.n3 10.955
R23507 mux8_0.NAND4F_4.B.n2 mux8_0.NAND4F_4.B.n1 10.955
R23508 mux8_0.NAND4F_4.B.n12 mux8_0.NAND4F_4.B.n9 3.67985
R23509 mux8_0.NAND4F_4.B.n9 mux8_0.NAND4F_4.B.n0 1.46835
R23510 mux8_0.NAND4F_4.B mux8_0.NAND4F_4.B.n12 0.502677
R23511 mux8_0.NAND4F_4.B.n9 mux8_0.NAND4F_4.B 0.498606
R23512 mux8_0.NAND4F_4.B mux8_0.NAND4F_4.B.n7 0.470197
R23513 mux8_0.NAND4F_5.Y.n1 mux8_0.NAND4F_5.Y.t9 1032.02
R23514 mux8_0.NAND4F_5.Y.n1 mux8_0.NAND4F_5.Y.t10 336.962
R23515 mux8_0.NAND4F_5.Y.n1 mux8_0.NAND4F_5.Y.t11 326.154
R23516 mux8_0.NAND4F_5.Y.n0 mux8_0.NAND4F_5.Y.n3 187.373
R23517 mux8_0.NAND4F_5.Y.n0 mux8_0.NAND4F_5.Y.n4 187.192
R23518 mux8_0.NAND4F_5.Y.n0 mux8_0.NAND4F_5.Y.n5 187.192
R23519 mux8_0.NAND4F_5.Y.n7 mux8_0.NAND4F_5.Y.n6 187.192
R23520 mux8_0.NAND4F_5.Y mux8_0.NAND4F_5.Y.n1 162.94
R23521 mux8_0.NAND4F_5.Y.n2 mux8_0.NAND4F_5.Y 24.4721
R23522 mux8_0.NAND4F_5.Y.n2 mux8_0.NAND4F_5.Y.t6 22.6141
R23523 mux8_0.NAND4F_5.Y.n3 mux8_0.NAND4F_5.Y.t0 20.1899
R23524 mux8_0.NAND4F_5.Y.n3 mux8_0.NAND4F_5.Y.t1 20.1899
R23525 mux8_0.NAND4F_5.Y.n4 mux8_0.NAND4F_5.Y.t8 20.1899
R23526 mux8_0.NAND4F_5.Y.n4 mux8_0.NAND4F_5.Y.t7 20.1899
R23527 mux8_0.NAND4F_5.Y.n5 mux8_0.NAND4F_5.Y.t2 20.1899
R23528 mux8_0.NAND4F_5.Y.n5 mux8_0.NAND4F_5.Y.t3 20.1899
R23529 mux8_0.NAND4F_5.Y.n6 mux8_0.NAND4F_5.Y.t4 20.1899
R23530 mux8_0.NAND4F_5.Y.n6 mux8_0.NAND4F_5.Y.t5 20.1899
R23531 mux8_0.NAND4F_5.Y mux8_0.NAND4F_5.Y.n2 0.950576
R23532 mux8_0.NAND4F_5.Y mux8_0.NAND4F_5.Y.n7 0.396904
R23533 mux8_0.NAND4F_5.Y.n7 mux8_0.NAND4F_5.Y.n0 0.358709
R23534 a_n6611_2026.n7 a_n6611_2026.n1 81.2978
R23535 a_n6611_2026.n1 a_n6611_2026.n6 81.1637
R23536 a_n6611_2026.n1 a_n6611_2026.n5 81.1637
R23537 a_n6611_2026.n0 a_n6611_2026.n4 81.1637
R23538 a_n6611_2026.n0 a_n6611_2026.n3 81.1637
R23539 a_n6611_2026.n0 a_n6611_2026.n2 80.9213
R23540 a_n6611_2026.n6 a_n6611_2026.t6 11.8205
R23541 a_n6611_2026.n6 a_n6611_2026.t3 11.8205
R23542 a_n6611_2026.n5 a_n6611_2026.t7 11.8205
R23543 a_n6611_2026.n5 a_n6611_2026.t11 11.8205
R23544 a_n6611_2026.n4 a_n6611_2026.t8 11.8205
R23545 a_n6611_2026.n4 a_n6611_2026.t10 11.8205
R23546 a_n6611_2026.n3 a_n6611_2026.t2 11.8205
R23547 a_n6611_2026.n3 a_n6611_2026.t9 11.8205
R23548 a_n6611_2026.n2 a_n6611_2026.t1 11.8205
R23549 a_n6611_2026.n2 a_n6611_2026.t0 11.8205
R23550 a_n6611_2026.n7 a_n6611_2026.t4 11.8205
R23551 a_n6611_2026.t5 a_n6611_2026.n7 11.8205
R23552 a_n6611_2026.n1 a_n6611_2026.n0 0.402735
R23553 mux8_4.NAND4F_0.C.n6 mux8_4.NAND4F_0.C.t4 978.795
R23554 mux8_4.NAND4F_0.C.n4 mux8_4.NAND4F_0.C.t12 978.795
R23555 mux8_4.NAND4F_0.C.n11 mux8_4.NAND4F_0.C.t11 978.795
R23556 mux8_4.NAND4F_0.C.n2 mux8_4.NAND4F_0.C.t13 978.795
R23557 mux8_4.NAND4F_0.C.n5 mux8_4.NAND4F_0.C.t7 308.481
R23558 mux8_4.NAND4F_0.C.n5 mux8_4.NAND4F_0.C.t5 308.481
R23559 mux8_4.NAND4F_0.C.n3 mux8_4.NAND4F_0.C.t15 308.481
R23560 mux8_4.NAND4F_0.C.n3 mux8_4.NAND4F_0.C.t14 308.481
R23561 mux8_4.NAND4F_0.C.n10 mux8_4.NAND4F_0.C.t6 308.481
R23562 mux8_4.NAND4F_0.C.n10 mux8_4.NAND4F_0.C.t8 308.481
R23563 mux8_4.NAND4F_0.C.n1 mux8_4.NAND4F_0.C.t9 308.481
R23564 mux8_4.NAND4F_0.C.n1 mux8_4.NAND4F_0.C.t10 308.481
R23565 mux8_4.NAND4F_0.C.n0 mux8_4.NAND4F_0.C.t1 256.514
R23566 mux8_4.NAND4F_0.C.n0 mux8_4.NAND4F_0.C.n8 226.258
R23567 mux8_4.NAND4F_0.C mux8_4.NAND4F_0.C.n6 161.856
R23568 mux8_4.NAND4F_0.C mux8_4.NAND4F_0.C.n4 161.847
R23569 mux8_4.NAND4F_0.C mux8_4.NAND4F_0.C.n11 161.84
R23570 mux8_4.NAND4F_0.C mux8_4.NAND4F_0.C.n2 161.831
R23571 mux8_4.NAND4F_0.C.n0 mux8_4.NAND4F_0.C.t0 83.7172
R23572 mux8_4.NAND4F_0.C.n8 mux8_4.NAND4F_0.C.t3 30.379
R23573 mux8_4.NAND4F_0.C.n8 mux8_4.NAND4F_0.C.t2 30.379
R23574 mux8_4.NAND4F_0.C.n9 mux8_4.NAND4F_0.C.n0 13.5186
R23575 mux8_4.NAND4F_0.C mux8_4.NAND4F_0.C.n12 13.0862
R23576 mux8_4.NAND4F_0.C.n7 mux8_4.NAND4F_0.C 13.0435
R23577 mux8_4.NAND4F_0.C.n12 mux8_4.NAND4F_0.C 12.4135
R23578 mux8_4.NAND4F_0.C.n7 mux8_4.NAND4F_0.C 12.4105
R23579 mux8_4.NAND4F_0.C.n6 mux8_4.NAND4F_0.C.n5 11.0463
R23580 mux8_4.NAND4F_0.C.n4 mux8_4.NAND4F_0.C.n3 11.0463
R23581 mux8_4.NAND4F_0.C.n11 mux8_4.NAND4F_0.C.n10 11.0463
R23582 mux8_4.NAND4F_0.C.n2 mux8_4.NAND4F_0.C.n1 11.0463
R23583 mux8_4.NAND4F_0.C.n12 mux8_4.NAND4F_0.C.n9 3.46056
R23584 mux8_4.NAND4F_0.C.n9 mux8_4.NAND4F_0.C.n7 1.8134
R23585 a_9336_n16422.t0 a_9336_n16422.t1 9.9005
R23586 a_9432_n16422.t0 a_9432_n16422.t1 9.9005
R23587 mux8_5.NAND4F_2.Y.n6 mux8_5.NAND4F_2.Y.t11 933.563
R23588 mux8_5.NAND4F_2.Y.n6 mux8_5.NAND4F_2.Y.t9 367.635
R23589 mux8_5.NAND4F_2.Y.n7 mux8_5.NAND4F_2.Y.t10 308.481
R23590 mux8_5.NAND4F_2.Y.n0 mux8_5.NAND4F_2.Y.n1 187.373
R23591 mux8_5.NAND4F_2.Y.n0 mux8_5.NAND4F_2.Y.n2 187.192
R23592 mux8_5.NAND4F_2.Y.n0 mux8_5.NAND4F_2.Y.n3 187.192
R23593 mux8_5.NAND4F_2.Y.n5 mux8_5.NAND4F_2.Y.n4 187.192
R23594 mux8_5.NAND4F_2.Y mux8_5.NAND4F_2.Y.n7 162.102
R23595 mux8_5.NAND4F_2.Y.n8 mux8_5.NAND4F_2.Y.t4 22.7096
R23596 mux8_5.NAND4F_2.Y.n8 mux8_5.NAND4F_2.Y 22.4285
R23597 mux8_5.NAND4F_2.Y.n1 mux8_5.NAND4F_2.Y.t0 20.1899
R23598 mux8_5.NAND4F_2.Y.n1 mux8_5.NAND4F_2.Y.t1 20.1899
R23599 mux8_5.NAND4F_2.Y.n2 mux8_5.NAND4F_2.Y.t6 20.1899
R23600 mux8_5.NAND4F_2.Y.n2 mux8_5.NAND4F_2.Y.t5 20.1899
R23601 mux8_5.NAND4F_2.Y.n3 mux8_5.NAND4F_2.Y.t7 20.1899
R23602 mux8_5.NAND4F_2.Y.n3 mux8_5.NAND4F_2.Y.t8 20.1899
R23603 mux8_5.NAND4F_2.Y.n4 mux8_5.NAND4F_2.Y.t2 20.1899
R23604 mux8_5.NAND4F_2.Y.n4 mux8_5.NAND4F_2.Y.t3 20.1899
R23605 mux8_5.NAND4F_2.Y.n7 mux8_5.NAND4F_2.Y.n6 10.955
R23606 mux8_5.NAND4F_2.Y mux8_5.NAND4F_2.Y.n8 0.799394
R23607 mux8_5.NAND4F_2.Y mux8_5.NAND4F_2.Y.n5 0.452586
R23608 mux8_5.NAND4F_2.Y.n5 mux8_5.NAND4F_2.Y.n0 0.358709
R23609 B7.n4 B7.t40 491.64
R23610 B7.n3 B7.t19 491.64
R23611 B7.n2 B7.t14 491.64
R23612 B7.n1 B7.t1 491.64
R23613 B7.n7 B7.t15 491.64
R23614 B7.n7 B7.t0 491.64
R23615 B7.n7 B7.t21 491.64
R23616 B7.n7 B7.t6 491.64
R23617 B7.n27 B7.t44 491.64
R23618 B7.n26 B7.t9 491.64
R23619 B7.n25 B7.t41 491.64
R23620 B7.n24 B7.t22 491.64
R23621 B7.n13 B7.t16 485.443
R23622 B7.n32 B7.t24 394.37
R23623 B7.n36 B7.t20 394.37
R23624 B7.n39 B7.t37 394.37
R23625 B7.n16 B7.t31 379.173
R23626 B7.n11 B7.t23 343.827
R23627 B7.n17 B7.t27 312.599
R23628 B7.n31 B7.t33 291.829
R23629 B7.n31 B7.t32 291.829
R23630 B7.n35 B7.t28 291.829
R23631 B7.n35 B7.t8 291.829
R23632 B7.n38 B7.t5 291.829
R23633 B7.n38 B7.t4 291.829
R23634 B7.n5 B7.t30 255.588
R23635 B7.n28 B7.t17 255.588
R23636 B7.n17 B7.t12 247.428
R23637 B7.n18 B7.t11 247.428
R23638 B7.n19 B7.t38 247.428
R23639 B7.n16 B7.t36 247.428
R23640 B7.n11 B7.t42 237.787
R23641 B7.n12 B7.t13 224.478
R23642 B7.n31 B7.t7 221.72
R23643 B7.n35 B7.t34 221.72
R23644 B7.n38 B7.t2 221.72
R23645 B7.n24 B7.n23 209.407
R23646 B7.n1 B7.n0 209.19
R23647 B7.n29 B7 206.742
R23648 B7 B7.n9 162.924
R23649 B7 B7.n20 162.139
R23650 B7.n0 B7.t26 139.78
R23651 B7.n0 B7.t35 139.78
R23652 B7.n0 B7.t18 139.78
R23653 B7.n8 B7.t3 139.78
R23654 B7.n8 B7.t29 139.78
R23655 B7.n8 B7.t43 139.78
R23656 B7.n8 B7.t25 139.78
R23657 B7.n23 B7.t45 139.78
R23658 B7.n23 B7.t10 139.78
R23659 B7.n23 B7.t39 139.78
R23660 B7.n13 B7.n12 83.8438
R23661 B7.n19 B7.n18 65.1723
R23662 B7.n18 B7.n17 65.1723
R23663 B7 B7.n13 61.0461
R23664 B7.n32 B7.n31 53.374
R23665 B7.n36 B7.n35 53.374
R23666 B7.n39 B7.n38 53.374
R23667 B7.n12 B7.n11 48.2005
R23668 B7.n9 B7.n8 38.6833
R23669 B7.n10 B7 37.3234
R23670 B7.n20 B7.n19 33.2653
R23671 B7.n20 B7.n16 31.9075
R23672 B7.n9 B7.n7 28.3986
R23673 B7 B7.n10 28.3317
R23674 B7 B7.n28 27.4136
R23675 B7.n3 B7.n2 17.8661
R23676 B7.n2 B7.n1 17.8661
R23677 B7.n25 B7.n24 17.8661
R23678 B7.n26 B7.n25 17.8661
R23679 B7.n4 B7.n3 17.1217
R23680 B7.n27 B7.n26 17.1217
R23681 B7.n40 B7.n37 14.3915
R23682 B7.n10 B7.n6 13.2852
R23683 B7.n37 B7 12.7234
R23684 B7.n34 B7.n30 12.62
R23685 B7.n34 B7 12.5598
R23686 B7.n15 B7.n14 12.4179
R23687 B7.n22 B7.n21 12.4105
R23688 B7.n30 B7.n29 12.4105
R23689 B7 B7.n5 11.1665
R23690 B7.n30 B7.n22 9.43705
R23691 B7.n22 B7.n15 5.31737
R23692 B7.n37 B7.n34 2.81006
R23693 B7.n5 B7.n4 1.8615
R23694 B7.n28 B7.n27 1.8615
R23695 B7.n14 B7 1.31242
R23696 B7.n33 B7.n32 1.19598
R23697 B7.n21 B7 1.08194
R23698 B7 B7.n36 0.81823
R23699 B7.n40 B7.n39 0.816926
R23700 B7.n15 B7 0.108208
R23701 B7.n29 B7 0.0769706
R23702 B7.n33 B7 0.067529
R23703 B7.n14 B7 0.0612639
R23704 B7 B7.n33 0.0456389
R23705 B7.n21 B7 0.0421667
R23706 B7.n6 B7 0.00999367
R23707 B7.n6 B7 0.00287342
R23708 B7 B7.n40 0.00272209
R23709 a_1887_5534.n1 a_1887_5534.n6 81.2978
R23710 a_1887_5534.n1 a_1887_5534.n5 81.1637
R23711 a_1887_5534.n0 a_1887_5534.n4 81.1637
R23712 a_1887_5534.n0 a_1887_5534.n3 81.1637
R23713 a_1887_5534.n7 a_1887_5534.n1 81.1637
R23714 a_1887_5534.n0 a_1887_5534.n2 80.9213
R23715 a_1887_5534.n6 a_1887_5534.t2 11.8205
R23716 a_1887_5534.n6 a_1887_5534.t1 11.8205
R23717 a_1887_5534.n5 a_1887_5534.t4 11.8205
R23718 a_1887_5534.n5 a_1887_5534.t5 11.8205
R23719 a_1887_5534.n4 a_1887_5534.t10 11.8205
R23720 a_1887_5534.n4 a_1887_5534.t11 11.8205
R23721 a_1887_5534.n3 a_1887_5534.t8 11.8205
R23722 a_1887_5534.n3 a_1887_5534.t9 11.8205
R23723 a_1887_5534.n2 a_1887_5534.t7 11.8205
R23724 a_1887_5534.n2 a_1887_5534.t6 11.8205
R23725 a_1887_5534.n7 a_1887_5534.t0 11.8205
R23726 a_1887_5534.t3 a_1887_5534.n7 11.8205
R23727 a_1887_5534.n1 a_1887_5534.n0 0.402735
R23728 mux8_5.inv_0.A.n3 mux8_5.inv_0.A.t8 291.829
R23729 mux8_5.inv_0.A.n3 mux8_5.inv_0.A.t7 291.829
R23730 mux8_5.inv_0.A.n0 mux8_5.inv_0.A.t1 256.425
R23731 mux8_5.inv_0.A.n0 mux8_5.inv_0.A.n4 231.24
R23732 mux8_5.inv_0.A.n0 mux8_5.inv_0.A.n5 231.03
R23733 mux8_5.inv_0.A.n3 mux8_5.inv_0.A.t10 221.72
R23734 mux8_5.inv_0.A.t9 mux8_5.inv_0.A.n2 393.959
R23735 mux8_5.inv_0.A.n6 mux8_5.inv_0.A.n1 66.6316
R23736 mux8_5.inv_0.A.n2 mux8_5.inv_0.A.n3 53.4611
R23737 mux8_5.inv_0.A.n4 mux8_5.inv_0.A.t3 25.395
R23738 mux8_5.inv_0.A.n4 mux8_5.inv_0.A.t2 25.395
R23739 mux8_5.inv_0.A.n5 mux8_5.inv_0.A.t5 25.395
R23740 mux8_5.inv_0.A.n5 mux8_5.inv_0.A.t4 25.395
R23741 mux8_5.inv_0.A.n6 mux8_5.inv_0.A.t6 19.8005
R23742 mux8_5.inv_0.A.n6 mux8_5.inv_0.A.t0 19.8005
R23743 mux8_5.inv_0.A.n1 mux8_5.inv_0.A.n0 0.38953
R23744 mux8_5.inv_0.A.n1 mux8_5.inv_0.A.n2 0.294762
R23745 mux8_5.NAND4F_2.D.n4 mux8_5.NAND4F_2.D.t7 1388.16
R23746 mux8_5.NAND4F_2.D.n7 mux8_5.NAND4F_2.D.t12 1388.16
R23747 mux8_5.NAND4F_2.D.n10 mux8_5.NAND4F_2.D.t4 1388.16
R23748 mux8_5.NAND4F_2.D.n1 mux8_5.NAND4F_2.D.t11 1388.16
R23749 mux8_5.NAND4F_2.D.n4 mux8_5.NAND4F_2.D.t6 350.839
R23750 mux8_5.NAND4F_2.D.n7 mux8_5.NAND4F_2.D.t9 350.839
R23751 mux8_5.NAND4F_2.D.n10 mux8_5.NAND4F_2.D.t5 350.839
R23752 mux8_5.NAND4F_2.D.n1 mux8_5.NAND4F_2.D.t14 350.839
R23753 mux8_5.NAND4F_2.D.n5 mux8_5.NAND4F_2.D.t13 308.481
R23754 mux8_5.NAND4F_2.D.n8 mux8_5.NAND4F_2.D.t10 308.481
R23755 mux8_5.NAND4F_2.D.n11 mux8_5.NAND4F_2.D.t8 308.481
R23756 mux8_5.NAND4F_2.D.n2 mux8_5.NAND4F_2.D.t15 308.481
R23757 mux8_5.NAND4F_2.D.n0 mux8_5.NAND4F_2.D.t2 256.514
R23758 mux8_5.NAND4F_2.D.n0 mux8_5.NAND4F_2.D.n3 226.258
R23759 mux8_5.NAND4F_2.D mux8_5.NAND4F_2.D.n5 161.458
R23760 mux8_5.NAND4F_2.D mux8_5.NAND4F_2.D.n11 161.435
R23761 mux8_5.NAND4F_2.D mux8_5.NAND4F_2.D.n2 161.435
R23762 mux8_5.NAND4F_2.D mux8_5.NAND4F_2.D.n8 161.429
R23763 mux8_5.NAND4F_2.D.n0 mux8_5.NAND4F_2.D.t0 83.7172
R23764 mux8_5.NAND4F_2.D.n3 mux8_5.NAND4F_2.D.t1 30.379
R23765 mux8_5.NAND4F_2.D.n3 mux8_5.NAND4F_2.D.t3 30.379
R23766 mux8_5.NAND4F_2.D.n5 mux8_5.NAND4F_2.D.n4 27.752
R23767 mux8_5.NAND4F_2.D.n8 mux8_5.NAND4F_2.D.n7 27.752
R23768 mux8_5.NAND4F_2.D.n11 mux8_5.NAND4F_2.D.n10 27.752
R23769 mux8_5.NAND4F_2.D.n2 mux8_5.NAND4F_2.D.n1 27.752
R23770 mux8_5.NAND4F_2.D.n6 mux8_5.NAND4F_2.D.n0 12.759
R23771 mux8_5.NAND4F_2.D mux8_5.NAND4F_2.D.n12 10.6871
R23772 mux8_5.NAND4F_2.D.n6 mux8_5.NAND4F_2.D 9.0005
R23773 mux8_5.NAND4F_2.D.n12 mux8_5.NAND4F_2.D 9.0005
R23774 mux8_5.NAND4F_2.D.n9 mux8_5.NAND4F_2.D 9.0005
R23775 mux8_5.NAND4F_2.D.n9 mux8_5.NAND4F_2.D.n6 1.74507
R23776 mux8_5.NAND4F_2.D.n12 mux8_5.NAND4F_2.D.n9 1.69072
R23777 a_n20446_n2915.t0 a_n20446_n2915.t1 19.8005
R23778 a_n12347_n34023.n2 a_n12347_n34023.t3 539.788
R23779 a_n12347_n34023.n3 a_n12347_n34023.t5 531.496
R23780 a_n12347_n34023.n2 a_n12347_n34023.t4 490.034
R23781 a_n12347_n34023.n5 a_n12347_n34023.t0 283.788
R23782 a_n12347_n34023.t1 a_n12347_n34023.n5 205.489
R23783 a_n12347_n34023.n0 a_n12347_n34023.t6 182.625
R23784 a_n12347_n34023.n1 a_n12347_n34023.t2 179.054
R23785 a_n12347_n34023.n0 a_n12347_n34023.t7 139.78
R23786 a_n12347_n34023.n4 a_n12347_n34023.n1 101.368
R23787 a_n12347_n34023.n5 a_n12347_n34023.n4 77.9135
R23788 a_n12347_n34023.n4 a_n12347_n34023.n3 76.1557
R23789 a_n12347_n34023.n3 a_n12347_n34023.n2 8.29297
R23790 a_n12347_n34023.n1 a_n12347_n34023.n0 3.57087
R23791 a_n11276_n34281.n2 a_n11276_n34281.n1 121.353
R23792 a_n11276_n34281.n3 a_n11276_n34281.n2 121.001
R23793 a_n11276_n34281.n2 a_n11276_n34281.n0 120.977
R23794 a_n11276_n34281.n0 a_n11276_n34281.t4 30.462
R23795 a_n11276_n34281.n0 a_n11276_n34281.t3 30.462
R23796 a_n11276_n34281.n1 a_n11276_n34281.t1 30.462
R23797 a_n11276_n34281.n1 a_n11276_n34281.t2 30.462
R23798 a_n11276_n34281.n3 a_n11276_n34281.t5 30.462
R23799 a_n11276_n34281.t0 a_n11276_n34281.n3 30.462
R23800 XOR8_0.S7.n0 XOR8_0.S7.t14 1032.02
R23801 XOR8_0.S7.n0 XOR8_0.S7.t12 336.962
R23802 XOR8_0.S7.n0 XOR8_0.S7.t13 326.154
R23803 XOR8_0.S7 XOR8_0.S7.n0 162.946
R23804 XOR8_0.S7.n3 XOR8_0.S7.n1 120.999
R23805 XOR8_0.S7.n3 XOR8_0.S7.n2 120.999
R23806 XOR8_0.S7.n15 XOR8_0.S7.n14 104.865
R23807 XOR8_0.S7.n5 XOR8_0.S7.n4 92.5005
R23808 XOR8_0.S7.n12 XOR8_0.S7.n10 86.2638
R23809 XOR8_0.S7.n10 XOR8_0.S7.n9 85.8873
R23810 XOR8_0.S7.n10 XOR8_0.S7.n7 85.724
R23811 XOR8_0.S7 XOR8_0.S7.n15 83.8907
R23812 XOR8_0.S7.n13 XOR8_0.S7.n12 75.0672
R23813 XOR8_0.S7.n13 XOR8_0.S7.n9 75.0672
R23814 XOR8_0.S7.n7 XOR8_0.S7.n6 73.1255
R23815 XOR8_0.S7.n12 XOR8_0.S7.n11 73.1255
R23816 XOR8_0.S7.n9 XOR8_0.S7.n8 73.1255
R23817 XOR8_0.S7.n14 XOR8_0.S7.n7 68.5181
R23818 XOR8_0.S7.n15 XOR8_0.S7.n5 41.9827
R23819 XOR8_0.S7.n4 XOR8_0.S7.t11 30.462
R23820 XOR8_0.S7.n4 XOR8_0.S7.t7 30.462
R23821 XOR8_0.S7.n1 XOR8_0.S7.t10 30.462
R23822 XOR8_0.S7.n1 XOR8_0.S7.t9 30.462
R23823 XOR8_0.S7.n2 XOR8_0.S7.t6 30.462
R23824 XOR8_0.S7.n2 XOR8_0.S7.t8 30.462
R23825 XOR8_0.S7.n5 XOR8_0.S7.n3 28.124
R23826 XOR8_0.S7.n11 XOR8_0.S7.t4 11.8205
R23827 XOR8_0.S7.n11 XOR8_0.S7.t3 11.8205
R23828 XOR8_0.S7.n6 XOR8_0.S7.t2 11.8205
R23829 XOR8_0.S7.n6 XOR8_0.S7.t5 11.8205
R23830 XOR8_0.S7.n8 XOR8_0.S7.t0 11.8205
R23831 XOR8_0.S7.n8 XOR8_0.S7.t1 11.8205
R23832 XOR8_0.S7.n14 XOR8_0.S7.n13 9.3005
R23833 mux8_6.A1.n1 mux8_6.A1.t8 1032.02
R23834 mux8_6.A1.n1 mux8_6.A1.t7 336.962
R23835 mux8_6.A1.n1 mux8_6.A1.t9 326.154
R23836 mux8_6.A1.n0 mux8_6.A1.n2 227.526
R23837 mux8_6.A1.n0 mux8_6.A1.n3 227.266
R23838 mux8_6.A1.n0 mux8_6.A1.n4 227.266
R23839 mux8_6.A1 mux8_6.A1.n1 162.952
R23840 mux8_6.A1.n0 mux8_6.A1.t0 42.7831
R23841 mux8_6.A1.n2 mux8_6.A1.t5 30.379
R23842 mux8_6.A1.n2 mux8_6.A1.t6 30.379
R23843 mux8_6.A1.n3 mux8_6.A1.t2 30.379
R23844 mux8_6.A1.n3 mux8_6.A1.t4 30.379
R23845 mux8_6.A1.n4 mux8_6.A1.t1 30.379
R23846 mux8_6.A1.n4 mux8_6.A1.t3 30.379
R23847 mux8_6.A1 mux8_6.A1.n0 18.8681
R23848 right_shifter_0.S7.n1 right_shifter_0.S7.t4 1032.02
R23849 right_shifter_0.S7.n1 right_shifter_0.S7.t5 336.962
R23850 right_shifter_0.S7.n1 right_shifter_0.S7.t6 326.154
R23851 right_shifter_0.S7.n0 right_shifter_0.S7.t1 256.514
R23852 right_shifter_0.S7.n0 right_shifter_0.S7.n2 226.258
R23853 mux8_6.NAND4F_6.A right_shifter_0.S7.n1 162.952
R23854 right_shifter_0.S7.n0 right_shifter_0.S7.t0 83.7172
R23855 mux8_6.A7 right_shifter_0.S7.n0 44.354
R23856 right_shifter_0.S7.n2 right_shifter_0.S7.t3 30.379
R23857 right_shifter_0.S7.n2 right_shifter_0.S7.t2 30.379
R23858 mux8_6.A7 mux8_6.NAND4F_6.A 13.4456
R23859 a_8592_n35462.t0 a_8592_n35462.t1 9.9005
R23860 mux8_6.NAND4F_6.Y.n1 mux8_6.NAND4F_6.Y.t9 933.563
R23861 mux8_6.NAND4F_6.Y.n1 mux8_6.NAND4F_6.Y.t10 367.635
R23862 mux8_6.NAND4F_6.Y.n2 mux8_6.NAND4F_6.Y.t11 308.481
R23863 mux8_6.NAND4F_6.Y.n0 mux8_6.NAND4F_6.Y.n4 187.373
R23864 mux8_6.NAND4F_6.Y.n0 mux8_6.NAND4F_6.Y.n5 187.192
R23865 mux8_6.NAND4F_6.Y.n0 mux8_6.NAND4F_6.Y.n6 187.192
R23866 mux8_6.NAND4F_6.Y.n8 mux8_6.NAND4F_6.Y.n7 187.192
R23867 mux8_6.NAND4F_6.Y mux8_6.NAND4F_6.Y.n2 162.047
R23868 mux8_6.NAND4F_6.Y.n3 mux8_6.NAND4F_6.Y.t2 22.7831
R23869 mux8_6.NAND4F_6.Y.n3 mux8_6.NAND4F_6.Y 22.171
R23870 mux8_6.NAND4F_6.Y.n4 mux8_6.NAND4F_6.Y.t1 20.1899
R23871 mux8_6.NAND4F_6.Y.n4 mux8_6.NAND4F_6.Y.t0 20.1899
R23872 mux8_6.NAND4F_6.Y.n5 mux8_6.NAND4F_6.Y.t6 20.1899
R23873 mux8_6.NAND4F_6.Y.n5 mux8_6.NAND4F_6.Y.t5 20.1899
R23874 mux8_6.NAND4F_6.Y.n6 mux8_6.NAND4F_6.Y.t7 20.1899
R23875 mux8_6.NAND4F_6.Y.n6 mux8_6.NAND4F_6.Y.t8 20.1899
R23876 mux8_6.NAND4F_6.Y.n7 mux8_6.NAND4F_6.Y.t4 20.1899
R23877 mux8_6.NAND4F_6.Y.n7 mux8_6.NAND4F_6.Y.t3 20.1899
R23878 mux8_6.NAND4F_6.Y.n2 mux8_6.NAND4F_6.Y.n1 10.955
R23879 mux8_6.NAND4F_6.Y mux8_6.NAND4F_6.Y.n3 0.781576
R23880 mux8_6.NAND4F_6.Y mux8_6.NAND4F_6.Y.n8 0.396904
R23881 mux8_6.NAND4F_6.Y.n8 mux8_6.NAND4F_6.Y.n0 0.358709
R23882 right_shifter_0.C.n1 right_shifter_0.C.t6 1032.02
R23883 right_shifter_0.C.n1 right_shifter_0.C.t4 336.962
R23884 right_shifter_0.C.n1 right_shifter_0.C.t5 326.154
R23885 right_shifter_0.C.n0 right_shifter_0.C.t3 256.514
R23886 right_shifter_0.C.n0 right_shifter_0.C.n2 226.258
R23887 mux8_0.NAND4F_6.A right_shifter_0.C.n1 162.952
R23888 right_shifter_0.C.n0 right_shifter_0.C.t0 83.7172
R23889 mux8_0.A7 right_shifter_0.C.n0 60.0185
R23890 right_shifter_0.C.n2 right_shifter_0.C.t1 30.379
R23891 right_shifter_0.C.n2 right_shifter_0.C.t2 30.379
R23892 mux8_0.A7 mux8_0.NAND4F_6.A 13.4456
R23893 mux8_3.NAND4F_4.B.n10 mux8_3.NAND4F_4.B.t12 933.563
R23894 mux8_3.NAND4F_4.B.n5 mux8_3.NAND4F_4.B.t4 933.563
R23895 mux8_3.NAND4F_4.B.n3 mux8_3.NAND4F_4.B.t9 933.563
R23896 mux8_3.NAND4F_4.B.n1 mux8_3.NAND4F_4.B.t15 933.563
R23897 mux8_3.NAND4F_4.B.n10 mux8_3.NAND4F_4.B.t7 367.635
R23898 mux8_3.NAND4F_4.B.n5 mux8_3.NAND4F_4.B.t5 367.635
R23899 mux8_3.NAND4F_4.B.n3 mux8_3.NAND4F_4.B.t10 367.635
R23900 mux8_3.NAND4F_4.B.n1 mux8_3.NAND4F_4.B.t13 367.635
R23901 mux8_3.NAND4F_4.B.n11 mux8_3.NAND4F_4.B.t8 308.481
R23902 mux8_3.NAND4F_4.B.n6 mux8_3.NAND4F_4.B.t6 308.481
R23903 mux8_3.NAND4F_4.B.n4 mux8_3.NAND4F_4.B.t11 308.481
R23904 mux8_3.NAND4F_4.B.n2 mux8_3.NAND4F_4.B.t14 308.481
R23905 mux8_3.NAND4F_4.B.n0 mux8_3.NAND4F_4.B.t1 256.514
R23906 mux8_3.NAND4F_4.B.n0 mux8_3.NAND4F_4.B.n8 226.258
R23907 mux8_3.NAND4F_4.B mux8_3.NAND4F_4.B.n2 162.173
R23908 mux8_3.NAND4F_4.B mux8_3.NAND4F_4.B.n6 162.137
R23909 mux8_3.NAND4F_4.B mux8_3.NAND4F_4.B.n11 162.117
R23910 mux8_3.NAND4F_4.B.n7 mux8_3.NAND4F_4.B.n4 161.703
R23911 mux8_3.NAND4F_4.B.n0 mux8_3.NAND4F_4.B.t0 83.7172
R23912 mux8_3.NAND4F_4.B.n8 mux8_3.NAND4F_4.B.t3 30.379
R23913 mux8_3.NAND4F_4.B.n8 mux8_3.NAND4F_4.B.t2 30.379
R23914 mux8_3.NAND4F_4.B.n12 mux8_3.NAND4F_4.B 24.8912
R23915 mux8_3.NAND4F_4.B.n7 mux8_3.NAND4F_4.B 21.6618
R23916 mux8_3.NAND4F_4.B.n11 mux8_3.NAND4F_4.B.n10 10.955
R23917 mux8_3.NAND4F_4.B.n6 mux8_3.NAND4F_4.B.n5 10.955
R23918 mux8_3.NAND4F_4.B.n4 mux8_3.NAND4F_4.B.n3 10.955
R23919 mux8_3.NAND4F_4.B.n2 mux8_3.NAND4F_4.B.n1 10.955
R23920 mux8_3.NAND4F_4.B.n12 mux8_3.NAND4F_4.B.n9 3.67985
R23921 mux8_3.NAND4F_4.B.n9 mux8_3.NAND4F_4.B.n0 1.46835
R23922 mux8_3.NAND4F_4.B mux8_3.NAND4F_4.B.n12 0.502677
R23923 mux8_3.NAND4F_4.B.n9 mux8_3.NAND4F_4.B 0.498606
R23924 mux8_3.NAND4F_4.B mux8_3.NAND4F_4.B.n7 0.470197
R23925 a_8496_n30006.t0 a_8496_n30006.t1 9.9005
R23926 a_8592_n30006.t0 a_8592_n30006.t1 9.9005
R23927 a_10363_n35461.t0 a_10363_n35461.t1 9.9005
R23928 a_n24162_n7992.t0 a_n24162_n7992.t1 19.8005
R23929 MULT_0.inv_6.A.n5 MULT_0.inv_6.A.t8 291.829
R23930 MULT_0.inv_6.A.n5 MULT_0.inv_6.A.t10 291.829
R23931 MULT_0.inv_6.A.n0 MULT_0.inv_6.A.n2 227.526
R23932 MULT_0.inv_6.A.n0 MULT_0.inv_6.A.n3 227.266
R23933 MULT_0.inv_6.A.n0 MULT_0.inv_6.A.n4 227.266
R23934 MULT_0.inv_6.A.n5 MULT_0.inv_6.A.t9 221.72
R23935 MULT_0.inv_6.A.t7 MULT_0.inv_6.A.n1 393.897
R23936 MULT_0.inv_6.A.n0 MULT_0.inv_6.A.t3 42.7333
R23937 MULT_0.inv_6.A.n2 MULT_0.inv_6.A.t6 30.379
R23938 MULT_0.inv_6.A.n2 MULT_0.inv_6.A.t5 30.379
R23939 MULT_0.inv_6.A.n3 MULT_0.inv_6.A.t1 30.379
R23940 MULT_0.inv_6.A.n3 MULT_0.inv_6.A.t4 30.379
R23941 MULT_0.inv_6.A.n4 MULT_0.inv_6.A.t2 30.379
R23942 MULT_0.inv_6.A.n4 MULT_0.inv_6.A.t0 30.379
R23943 MULT_0.inv_6.A.n5 MULT_0.inv_6.A.n1 53.4911
R23944 MULT_0.inv_6.A.n0 MULT_0.inv_6.A.n1 0.620756
R23945 a_n10108_n5154.n2 a_n10108_n5154.n0 121.353
R23946 a_n10108_n5154.n3 a_n10108_n5154.n2 121.353
R23947 a_n10108_n5154.n2 a_n10108_n5154.n1 121.001
R23948 a_n10108_n5154.n1 a_n10108_n5154.t2 30.462
R23949 a_n10108_n5154.n1 a_n10108_n5154.t5 30.462
R23950 a_n10108_n5154.n0 a_n10108_n5154.t0 30.462
R23951 a_n10108_n5154.n0 a_n10108_n5154.t1 30.462
R23952 a_n10108_n5154.t4 a_n10108_n5154.n3 30.462
R23953 a_n10108_n5154.n3 a_n10108_n5154.t3 30.462
R23954 mux8_5.A0.n0 mux8_5.A0.t14 1032.02
R23955 mux8_5.A0.n0 mux8_5.A0.t12 336.962
R23956 mux8_5.A0.n0 mux8_5.A0.t13 326.154
R23957 mux8_5.A0 mux8_5.A0.n0 162.952
R23958 mux8_5.A0.n3 mux8_5.A0.n2 120.999
R23959 mux8_5.A0.n3 mux8_5.A0.n1 120.999
R23960 mux8_5.A0.n15 mux8_5.A0.n14 104.489
R23961 mux8_5.A0.n5 mux8_5.A0.n4 92.5005
R23962 mux8_5.A0.n12 mux8_5.A0.n10 86.2638
R23963 mux8_5.A0.n10 mux8_5.A0.n9 85.8873
R23964 mux8_5.A0.n10 mux8_5.A0.n7 85.724
R23965 mux8_5.A0 mux8_5.A0.n15 83.8907
R23966 mux8_5.A0.n13 mux8_5.A0.n12 75.0672
R23967 mux8_5.A0.n13 mux8_5.A0.n9 75.0672
R23968 mux8_5.A0.n12 mux8_5.A0.n11 73.1255
R23969 mux8_5.A0.n9 mux8_5.A0.n8 73.1255
R23970 mux8_5.A0.n7 mux8_5.A0.n6 73.1255
R23971 mux8_5.A0.n14 mux8_5.A0.n7 68.8946
R23972 mux8_5.A0.n15 mux8_5.A0.n5 41.9827
R23973 mux8_5.A0.n4 mux8_5.A0.t1 30.462
R23974 mux8_5.A0.n4 mux8_5.A0.t3 30.462
R23975 mux8_5.A0.n2 mux8_5.A0.t4 30.462
R23976 mux8_5.A0.n2 mux8_5.A0.t5 30.462
R23977 mux8_5.A0.n1 mux8_5.A0.t2 30.462
R23978 mux8_5.A0.n1 mux8_5.A0.t0 30.462
R23979 mux8_5.A0.n5 mux8_5.A0.n3 28.124
R23980 mux8_5.A0.n8 mux8_5.A0.t11 11.8205
R23981 mux8_5.A0.n8 mux8_5.A0.t9 11.8205
R23982 mux8_5.A0.n11 mux8_5.A0.t6 11.8205
R23983 mux8_5.A0.n11 mux8_5.A0.t7 11.8205
R23984 mux8_5.A0.n6 mux8_5.A0.t10 11.8205
R23985 mux8_5.A0.n6 mux8_5.A0.t8 11.8205
R23986 mux8_5.A0.n14 mux8_5.A0.n13 9.3005
R23987 a_n19981_n8419.n2 a_n19981_n8419.n1 121.353
R23988 a_n19981_n8419.n2 a_n19981_n8419.n0 121.353
R23989 a_n19981_n8419.n3 a_n19981_n8419.n2 121.001
R23990 a_n19981_n8419.n1 a_n19981_n8419.t1 30.462
R23991 a_n19981_n8419.n1 a_n19981_n8419.t0 30.462
R23992 a_n19981_n8419.n0 a_n19981_n8419.t5 30.462
R23993 a_n19981_n8419.n0 a_n19981_n8419.t4 30.462
R23994 a_n19981_n8419.n3 a_n19981_n8419.t3 30.462
R23995 a_n19981_n8419.t2 a_n19981_n8419.n3 30.462
R23996 a_7452_n2838.t0 a_7452_n2838.t1 9.9005
R23997 a_7548_n2838.t0 a_7548_n2838.t1 9.9005
R23998 a_n10884_1406.n2 a_n10884_1406.n0 121.353
R23999 a_n10884_1406.n3 a_n10884_1406.n2 121.353
R24000 a_n10884_1406.n2 a_n10884_1406.n1 121.001
R24001 a_n10884_1406.n0 a_n10884_1406.t5 30.462
R24002 a_n10884_1406.n0 a_n10884_1406.t3 30.462
R24003 a_n10884_1406.n1 a_n10884_1406.t1 30.462
R24004 a_n10884_1406.n1 a_n10884_1406.t4 30.462
R24005 a_n10884_1406.t2 a_n10884_1406.n3 30.462
R24006 a_n10884_1406.n3 a_n10884_1406.t0 30.462
R24007 a_n8170_1406.n2 a_n8170_1406.n0 121.353
R24008 a_n8170_1406.n2 a_n8170_1406.n1 121.001
R24009 a_n8170_1406.n3 a_n8170_1406.n2 120.977
R24010 a_n8170_1406.n0 a_n8170_1406.t4 30.462
R24011 a_n8170_1406.n0 a_n8170_1406.t5 30.462
R24012 a_n8170_1406.n1 a_n8170_1406.t1 30.462
R24013 a_n8170_1406.n1 a_n8170_1406.t3 30.462
R24014 a_n8170_1406.t2 a_n8170_1406.n3 30.462
R24015 a_n8170_1406.n3 a_n8170_1406.t0 30.462
R24016 MULT_0.inv_7.A.n5 MULT_0.inv_7.A.t10 291.829
R24017 MULT_0.inv_7.A.n5 MULT_0.inv_7.A.t8 291.829
R24018 MULT_0.inv_7.A.n0 MULT_0.inv_7.A.n3 227.526
R24019 MULT_0.inv_7.A.n0 MULT_0.inv_7.A.n2 227.266
R24020 MULT_0.inv_7.A.n0 MULT_0.inv_7.A.n4 227.266
R24021 MULT_0.inv_7.A.n5 MULT_0.inv_7.A.t7 221.72
R24022 MULT_0.inv_7.A.t9 MULT_0.inv_7.A.n1 393.897
R24023 MULT_0.inv_7.A.n0 MULT_0.inv_7.A.t3 42.7333
R24024 MULT_0.inv_7.A.n3 MULT_0.inv_7.A.t1 30.379
R24025 MULT_0.inv_7.A.n3 MULT_0.inv_7.A.t0 30.379
R24026 MULT_0.inv_7.A.n2 MULT_0.inv_7.A.t4 30.379
R24027 MULT_0.inv_7.A.n2 MULT_0.inv_7.A.t5 30.379
R24028 MULT_0.inv_7.A.n4 MULT_0.inv_7.A.t6 30.379
R24029 MULT_0.inv_7.A.n4 MULT_0.inv_7.A.t2 30.379
R24030 MULT_0.inv_7.A.n5 MULT_0.inv_7.A.n1 53.4911
R24031 MULT_0.inv_7.A.n0 MULT_0.inv_7.A.n1 0.620447
R24032 a_n12345_n31115.n2 a_n12345_n31115.t6 541.395
R24033 a_n12345_n31115.n3 a_n12345_n31115.t3 527.402
R24034 a_n12345_n31115.n2 a_n12345_n31115.t4 491.64
R24035 a_n12345_n31115.n5 a_n12345_n31115.t0 281.906
R24036 a_n12345_n31115.t1 a_n12345_n31115.n5 204.359
R24037 a_n12345_n31115.n0 a_n12345_n31115.t2 180.73
R24038 a_n12345_n31115.n1 a_n12345_n31115.t7 179.45
R24039 a_n12345_n31115.n0 a_n12345_n31115.t5 139.78
R24040 a_n12345_n31115.n4 a_n12345_n31115.n1 105.635
R24041 a_n12345_n31115.n4 a_n12345_n31115.n3 76.0005
R24042 a_n12345_n31115.n5 a_n12345_n31115.n4 67.9685
R24043 a_n12345_n31115.n3 a_n12345_n31115.n2 13.994
R24044 a_n12345_n31115.n1 a_n12345_n31115.n0 1.28015
R24045 a_n13192_1406.n2 a_n13192_1406.n1 121.353
R24046 a_n13192_1406.n3 a_n13192_1406.n2 121.001
R24047 a_n13192_1406.n2 a_n13192_1406.n0 120.977
R24048 a_n13192_1406.n1 a_n13192_1406.t4 30.462
R24049 a_n13192_1406.n1 a_n13192_1406.t5 30.462
R24050 a_n13192_1406.n0 a_n13192_1406.t0 30.462
R24051 a_n13192_1406.n0 a_n13192_1406.t1 30.462
R24052 a_n13192_1406.t2 a_n13192_1406.n3 30.462
R24053 a_n13192_1406.n3 a_n13192_1406.t3 30.462
R24054 a_11865_n11831.n1 a_11865_n11831.n5 231.24
R24055 a_11865_n11831.n0 a_11865_n11831.n2 231.24
R24056 a_11865_n11831.n1 a_11865_n11831.n4 231.03
R24057 a_11865_n11831.n0 a_11865_n11831.n3 231.03
R24058 a_11865_n11831.n6 a_11865_n11831.n1 231.03
R24059 a_11865_n11831.n5 a_11865_n11831.t3 25.395
R24060 a_11865_n11831.n5 a_11865_n11831.t1 25.395
R24061 a_11865_n11831.n4 a_11865_n11831.t5 25.395
R24062 a_11865_n11831.n4 a_11865_n11831.t0 25.395
R24063 a_11865_n11831.n3 a_11865_n11831.t7 25.395
R24064 a_11865_n11831.n3 a_11865_n11831.t6 25.395
R24065 a_11865_n11831.n2 a_11865_n11831.t9 25.395
R24066 a_11865_n11831.n2 a_11865_n11831.t8 25.395
R24067 a_11865_n11831.t4 a_11865_n11831.n6 25.395
R24068 a_11865_n11831.n6 a_11865_n11831.t2 25.395
R24069 a_11865_n11831.n1 a_11865_n11831.n0 0.421553
R24070 right_shifter_0.buffer_3.inv_1.A.n0 right_shifter_0.buffer_3.inv_1.A.t4 393.921
R24071 right_shifter_0.buffer_3.inv_1.A.n2 right_shifter_0.buffer_3.inv_1.A.t7 291.829
R24072 right_shifter_0.buffer_3.inv_1.A.n2 right_shifter_0.buffer_3.inv_1.A.t6 291.829
R24073 right_shifter_0.buffer_3.inv_1.A.n0 right_shifter_0.buffer_3.inv_1.A.t1 256.514
R24074 right_shifter_0.buffer_3.inv_1.A.n0 right_shifter_0.buffer_3.inv_1.A.n1 226.162
R24075 right_shifter_0.buffer_3.inv_1.A.n2 right_shifter_0.buffer_3.inv_1.A.t5 221.72
R24076 right_shifter_0.buffer_3.inv_1.A.n0 right_shifter_0.buffer_3.inv_1.A.t0 83.795
R24077 right_shifter_0.buffer_3.inv_1.A.n0 right_shifter_0.buffer_3.inv_1.A.n2 53.7938
R24078 right_shifter_0.buffer_3.inv_1.A.n1 right_shifter_0.buffer_3.inv_1.A.t3 30.379
R24079 right_shifter_0.buffer_3.inv_1.A.n1 right_shifter_0.buffer_3.inv_1.A.t2 30.379
R24080 right_shifter_0.S4.n1 right_shifter_0.S4.t4 1032.02
R24081 right_shifter_0.S4.n1 right_shifter_0.S4.t5 336.962
R24082 right_shifter_0.S4.n1 right_shifter_0.S4.t6 326.154
R24083 right_shifter_0.S4.n0 right_shifter_0.S4.t1 256.514
R24084 right_shifter_0.S4.n0 right_shifter_0.S4.n2 226.258
R24085 mux8_5.NAND4F_6.A right_shifter_0.S4.n1 162.952
R24086 right_shifter_0.S4.n0 right_shifter_0.S4.t0 83.7172
R24087 right_shifter_0.S4.n2 right_shifter_0.S4.t3 30.379
R24088 right_shifter_0.S4.n2 right_shifter_0.S4.t2 30.379
R24089 mux8_5.A7 right_shifter_0.S4.n0 25.8449
R24090 mux8_5.A7 mux8_5.NAND4F_6.A 13.3456
R24091 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n9 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t11 540.38
R24092 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t9 491.64
R24093 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t17 491.64
R24094 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t8 491.64
R24095 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t10 491.64
R24096 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n7 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t16 367.928
R24097 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n1 227.526
R24098 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n8 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t14 227.356
R24099 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n2 227.266
R24100 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n3 227.266
R24101 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n7 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t13 213.688
R24102 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n6 162.852
R24103 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n9 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n8 160.439
R24104 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t15 139.78
R24105 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t7 139.78
R24106 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t18 139.78
R24107 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t12 139.78
R24108 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n8 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n7 94.4341
R24109 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t0 42.7831
R24110 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n6 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n5 38.6833
R24111 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n1 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t6 30.379
R24112 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n1 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t5 30.379
R24113 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n2 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t2 30.379
R24114 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n2 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t4 30.379
R24115 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n3 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t3 30.379
R24116 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n3 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t1 30.379
R24117 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n6 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n4 28.3986
R24118 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n0 18.8832
R24119 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n10 10.7052
R24120 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n10 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 5.09176
R24121 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n10 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 4.19292
R24122 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n9 0.794268
R24123 a_n23095_1380.n2 a_n23095_1380.t6 541.395
R24124 a_n23095_1380.n3 a_n23095_1380.t5 527.402
R24125 a_n23095_1380.n2 a_n23095_1380.t4 491.64
R24126 a_n23095_1380.n5 a_n23095_1380.t0 281.906
R24127 a_n23095_1380.t1 a_n23095_1380.n5 204.359
R24128 a_n23095_1380.n0 a_n23095_1380.t3 180.73
R24129 a_n23095_1380.n1 a_n23095_1380.t2 179.45
R24130 a_n23095_1380.n0 a_n23095_1380.t7 139.78
R24131 a_n23095_1380.n4 a_n23095_1380.n1 105.635
R24132 a_n23095_1380.n4 a_n23095_1380.n3 76.0005
R24133 a_n23095_1380.n5 a_n23095_1380.n4 67.9685
R24134 a_n23095_1380.n3 a_n23095_1380.n2 13.994
R24135 a_n23095_1380.n1 a_n23095_1380.n0 1.28015
R24136 a_n9305_n11683.n0 a_n9305_n11683.t5 539.788
R24137 a_n9305_n11683.n1 a_n9305_n11683.t7 531.496
R24138 a_n9305_n11683.n0 a_n9305_n11683.t4 490.034
R24139 a_n9305_n11683.n5 a_n9305_n11683.t0 283.788
R24140 a_n9305_n11683.t1 a_n9305_n11683.n5 205.489
R24141 a_n9305_n11683.n2 a_n9305_n11683.t3 182.625
R24142 a_n9305_n11683.n3 a_n9305_n11683.t6 179.054
R24143 a_n9305_n11683.n2 a_n9305_n11683.t2 139.78
R24144 a_n9305_n11683.n4 a_n9305_n11683.n3 101.368
R24145 a_n9305_n11683.n5 a_n9305_n11683.n4 77.9135
R24146 a_n9305_n11683.n4 a_n9305_n11683.n1 76.1557
R24147 a_n9305_n11683.n1 a_n9305_n11683.n0 8.29297
R24148 a_n9305_n11683.n3 a_n9305_n11683.n2 3.57087
R24149 mux8_4.A1.n0 mux8_4.A1.t12 1032.02
R24150 mux8_4.A1.n0 mux8_4.A1.t14 336.962
R24151 mux8_4.A1.n0 mux8_4.A1.t13 326.154
R24152 mux8_4.A1 mux8_4.A1.n0 162.952
R24153 mux8_4.A1.n3 mux8_4.A1.n2 120.999
R24154 mux8_4.A1.n3 mux8_4.A1.n1 120.999
R24155 mux8_4.A1.n15 mux8_4.A1.n14 104.489
R24156 mux8_4.A1.n5 mux8_4.A1.n4 92.5005
R24157 mux8_4.A1.n12 mux8_4.A1.n10 86.2638
R24158 mux8_4.A1.n10 mux8_4.A1.n9 85.8873
R24159 mux8_4.A1.n10 mux8_4.A1.n7 85.724
R24160 mux8_4.A1 mux8_4.A1.n15 83.8907
R24161 mux8_4.A1.n13 mux8_4.A1.n12 75.0672
R24162 mux8_4.A1.n13 mux8_4.A1.n9 75.0672
R24163 mux8_4.A1.n12 mux8_4.A1.n11 73.1255
R24164 mux8_4.A1.n9 mux8_4.A1.n8 73.1255
R24165 mux8_4.A1.n7 mux8_4.A1.n6 73.1255
R24166 mux8_4.A1.n14 mux8_4.A1.n7 68.8946
R24167 mux8_4.A1.n15 mux8_4.A1.n5 41.9827
R24168 mux8_4.A1.n4 mux8_4.A1.t5 30.462
R24169 mux8_4.A1.n4 mux8_4.A1.t10 30.462
R24170 mux8_4.A1.n2 mux8_4.A1.t11 30.462
R24171 mux8_4.A1.n2 mux8_4.A1.t9 30.462
R24172 mux8_4.A1.n1 mux8_4.A1.t3 30.462
R24173 mux8_4.A1.n1 mux8_4.A1.t4 30.462
R24174 mux8_4.A1.n5 mux8_4.A1.n3 28.124
R24175 mux8_4.A1.n8 mux8_4.A1.t2 11.8205
R24176 mux8_4.A1.n8 mux8_4.A1.t1 11.8205
R24177 mux8_4.A1.n11 mux8_4.A1.t8 11.8205
R24178 mux8_4.A1.n11 mux8_4.A1.t6 11.8205
R24179 mux8_4.A1.n6 mux8_4.A1.t0 11.8205
R24180 mux8_4.A1.n6 mux8_4.A1.t7 11.8205
R24181 mux8_4.A1.n14 mux8_4.A1.n13 9.3005
R24182 a_n9125_n11683.n2 a_n9125_n11683.n0 121.353
R24183 a_n9125_n11683.n2 a_n9125_n11683.n1 121.001
R24184 a_n9125_n11683.n3 a_n9125_n11683.n2 120.977
R24185 a_n9125_n11683.n0 a_n9125_n11683.t2 30.462
R24186 a_n9125_n11683.n0 a_n9125_n11683.t0 30.462
R24187 a_n9125_n11683.n1 a_n9125_n11683.t3 30.462
R24188 a_n9125_n11683.n1 a_n9125_n11683.t1 30.462
R24189 a_n9125_n11683.t4 a_n9125_n11683.n3 30.462
R24190 a_n9125_n11683.n3 a_n9125_n11683.t5 30.462
R24191 a_11290_n26406.t0 a_11290_n26406.t1 9.9005
R24192 a_n13399_n5154.n2 a_n13399_n5154.n0 121.353
R24193 a_n13399_n5154.n3 a_n13399_n5154.n2 121.353
R24194 a_n13399_n5154.n2 a_n13399_n5154.n1 121.001
R24195 a_n13399_n5154.n0 a_n13399_n5154.t5 30.462
R24196 a_n13399_n5154.n0 a_n13399_n5154.t4 30.462
R24197 a_n13399_n5154.n1 a_n13399_n5154.t0 30.462
R24198 a_n13399_n5154.n1 a_n13399_n5154.t3 30.462
R24199 a_n13399_n5154.n3 a_n13399_n5154.t1 30.462
R24200 a_n13399_n5154.t2 a_n13399_n5154.n3 30.462
R24201 Y4.n2 Y4.t7 960.788
R24202 Y4.n0 Y4.t6 883.668
R24203 Y4.n1 Y4.t5 740.381
R24204 Y4.n0 Y4.t4 729.428
R24205 Y4.n4 Y4.t3 256.514
R24206 Y4.n5 Y4.n3 226.251
R24207 Y4 Y4.n2 162.037
R24208 Y4.n4 Y4.t0 83.7599
R24209 Y4.n1 Y4.n0 72.3005
R24210 Y4.n3 Y4.t2 30.379
R24211 Y4.n3 Y4.t1 30.379
R24212 Y4.n2 Y4.n1 16.7975
R24213 Y4.n5 Y4 0.0547328
R24214 Y4.n5 Y4.n4 0.0323878
R24215 Y4 Y4.n5 0.0126173
R24216 mux8_8.NAND4F_4.Y.n6 mux8_8.NAND4F_4.Y.t9 1032.02
R24217 mux8_8.NAND4F_4.Y.n6 mux8_8.NAND4F_4.Y.t10 336.962
R24218 mux8_8.NAND4F_4.Y.n6 mux8_8.NAND4F_4.Y.t11 326.154
R24219 mux8_8.NAND4F_4.Y.n0 mux8_8.NAND4F_4.Y.n1 187.373
R24220 mux8_8.NAND4F_4.Y.n0 mux8_8.NAND4F_4.Y.n2 187.192
R24221 mux8_8.NAND4F_4.Y.n0 mux8_8.NAND4F_4.Y.n3 187.192
R24222 mux8_8.NAND4F_4.Y.n5 mux8_8.NAND4F_4.Y.n4 187.192
R24223 mux8_8.NAND4F_4.Y mux8_8.NAND4F_4.Y.n6 162.942
R24224 mux8_8.NAND4F_4.Y.n7 mux8_8.NAND4F_4.Y 24.5377
R24225 mux8_8.NAND4F_4.Y.n7 mux8_8.NAND4F_4.Y.t2 22.6141
R24226 mux8_8.NAND4F_4.Y.n1 mux8_8.NAND4F_4.Y.t3 20.1899
R24227 mux8_8.NAND4F_4.Y.n1 mux8_8.NAND4F_4.Y.t4 20.1899
R24228 mux8_8.NAND4F_4.Y.n2 mux8_8.NAND4F_4.Y.t5 20.1899
R24229 mux8_8.NAND4F_4.Y.n2 mux8_8.NAND4F_4.Y.t6 20.1899
R24230 mux8_8.NAND4F_4.Y.n3 mux8_8.NAND4F_4.Y.t7 20.1899
R24231 mux8_8.NAND4F_4.Y.n3 mux8_8.NAND4F_4.Y.t8 20.1899
R24232 mux8_8.NAND4F_4.Y.n4 mux8_8.NAND4F_4.Y.t0 20.1899
R24233 mux8_8.NAND4F_4.Y.n4 mux8_8.NAND4F_4.Y.t1 20.1899
R24234 mux8_8.NAND4F_4.Y mux8_8.NAND4F_4.Y.n7 0.894894
R24235 mux8_8.NAND4F_4.Y mux8_8.NAND4F_4.Y.n5 0.452586
R24236 mux8_8.NAND4F_4.Y.n5 mux8_8.NAND4F_4.Y.n0 0.358709
R24237 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t7 540.38
R24238 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t10 367.928
R24239 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n5 227.526
R24240 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t8 227.356
R24241 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n6 227.266
R24242 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n4 227.266
R24243 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t9 213.688
R24244 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n2 160.439
R24245 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n1 94.4341
R24246 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t3 42.7944
R24247 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t5 30.379
R24248 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t0 30.379
R24249 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t6 30.379
R24250 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t4 30.379
R24251 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t1 30.379
R24252 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.t2 30.379
R24253 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n0 13.4358
R24254 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B.n3 0.821842
R24255 a_n12499_373.t0 a_n12499_373.t1 19.8005
R24256 MULT_0.NAND2_4.Y.n5 MULT_0.NAND2_4.Y.t8 291.829
R24257 MULT_0.NAND2_4.Y.n5 MULT_0.NAND2_4.Y.t10 291.829
R24258 MULT_0.NAND2_4.Y.n0 MULT_0.NAND2_4.Y.n2 227.526
R24259 MULT_0.NAND2_4.Y.n0 MULT_0.NAND2_4.Y.n3 227.266
R24260 MULT_0.NAND2_4.Y.n0 MULT_0.NAND2_4.Y.n4 227.266
R24261 MULT_0.NAND2_4.Y.n5 MULT_0.NAND2_4.Y.t9 221.72
R24262 MULT_0.NAND2_4.Y.t7 MULT_0.NAND2_4.Y.n1 393.897
R24263 MULT_0.NAND2_4.Y.n0 MULT_0.NAND2_4.Y.t0 42.7333
R24264 MULT_0.NAND2_4.Y.n2 MULT_0.NAND2_4.Y.t6 30.379
R24265 MULT_0.NAND2_4.Y.n2 MULT_0.NAND2_4.Y.t5 30.379
R24266 MULT_0.NAND2_4.Y.n3 MULT_0.NAND2_4.Y.t2 30.379
R24267 MULT_0.NAND2_4.Y.n3 MULT_0.NAND2_4.Y.t4 30.379
R24268 MULT_0.NAND2_4.Y.n4 MULT_0.NAND2_4.Y.t3 30.379
R24269 MULT_0.NAND2_4.Y.n4 MULT_0.NAND2_4.Y.t1 30.379
R24270 MULT_0.NAND2_4.Y.n5 MULT_0.NAND2_4.Y.n1 53.4911
R24271 MULT_0.NAND2_4.Y.n0 MULT_0.NAND2_4.Y.n1 0.620756
R24272 a_n17548_3190.n2 a_n17548_3190.t4 541.395
R24273 a_n17548_3190.n3 a_n17548_3190.t2 527.402
R24274 a_n17548_3190.n2 a_n17548_3190.t5 491.64
R24275 a_n17548_3190.n5 a_n17548_3190.t0 281.906
R24276 a_n17548_3190.t1 a_n17548_3190.n5 204.359
R24277 a_n17548_3190.n0 a_n17548_3190.t6 180.73
R24278 a_n17548_3190.n1 a_n17548_3190.t3 179.45
R24279 a_n17548_3190.n0 a_n17548_3190.t7 139.78
R24280 a_n17548_3190.n4 a_n17548_3190.n1 105.635
R24281 a_n17548_3190.n4 a_n17548_3190.n3 76.0005
R24282 a_n17548_3190.n5 a_n17548_3190.n4 67.9685
R24283 a_n17548_3190.n3 a_n17548_3190.n2 13.994
R24284 a_n17548_3190.n1 a_n17548_3190.n0 1.28015
R24285 a_8400_1690.t0 a_8400_1690.t1 9.9005
R24286 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n9 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t12 540.38
R24287 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t7 491.64
R24288 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t9 491.64
R24289 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t17 491.64
R24290 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t11 491.64
R24291 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n7 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t14 367.928
R24292 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n1 227.526
R24293 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n8 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t16 227.356
R24294 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n3 227.266
R24295 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n2 227.266
R24296 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n7 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t13 213.688
R24297 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n6 162.852
R24298 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n9 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n8 160.439
R24299 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t10 139.78
R24300 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t8 139.78
R24301 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t15 139.78
R24302 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t18 139.78
R24303 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n8 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n7 94.4341
R24304 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t3 42.7831
R24305 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n6 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n5 38.6833
R24306 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n3 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t4 30.379
R24307 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n3 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t6 30.379
R24308 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n1 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t1 30.379
R24309 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n1 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t0 30.379
R24310 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n2 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t5 30.379
R24311 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n2 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t2 30.379
R24312 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n6 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n4 28.3986
R24313 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n0 18.8832
R24314 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n10 11.2587
R24315 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n10 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 5.09176
R24316 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n10 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 4.19292
R24317 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n9 0.794268
R24318 a_n19774_2026.n0 a_n19774_2026.n2 81.2978
R24319 a_n19774_2026.n0 a_n19774_2026.n3 81.1637
R24320 a_n19774_2026.n0 a_n19774_2026.n4 81.1637
R24321 a_n19774_2026.n1 a_n19774_2026.n5 81.1637
R24322 a_n19774_2026.n1 a_n19774_2026.n6 81.1637
R24323 a_n19774_2026.n7 a_n19774_2026.n1 80.9213
R24324 a_n19774_2026.n2 a_n19774_2026.t0 11.8205
R24325 a_n19774_2026.n2 a_n19774_2026.t10 11.8205
R24326 a_n19774_2026.n3 a_n19774_2026.t7 11.8205
R24327 a_n19774_2026.n3 a_n19774_2026.t9 11.8205
R24328 a_n19774_2026.n4 a_n19774_2026.t11 11.8205
R24329 a_n19774_2026.n4 a_n19774_2026.t8 11.8205
R24330 a_n19774_2026.n5 a_n19774_2026.t4 11.8205
R24331 a_n19774_2026.n5 a_n19774_2026.t6 11.8205
R24332 a_n19774_2026.n6 a_n19774_2026.t2 11.8205
R24333 a_n19774_2026.n6 a_n19774_2026.t5 11.8205
R24334 a_n19774_2026.t3 a_n19774_2026.n7 11.8205
R24335 a_n19774_2026.n7 a_n19774_2026.t1 11.8205
R24336 a_n19774_2026.n1 a_n19774_2026.n0 0.402735
R24337 a_n7496_3810.n0 a_n7496_3810.n2 81.2978
R24338 a_n7496_3810.n1 a_n7496_3810.n5 81.1637
R24339 a_n7496_3810.n0 a_n7496_3810.n4 81.1637
R24340 a_n7496_3810.n0 a_n7496_3810.n3 81.1637
R24341 a_n7496_3810.n7 a_n7496_3810.n1 81.1637
R24342 a_n7496_3810.n1 a_n7496_3810.n6 80.9213
R24343 a_n7496_3810.n6 a_n7496_3810.t0 11.8205
R24344 a_n7496_3810.n6 a_n7496_3810.t1 11.8205
R24345 a_n7496_3810.n5 a_n7496_3810.t5 11.8205
R24346 a_n7496_3810.n5 a_n7496_3810.t3 11.8205
R24347 a_n7496_3810.n4 a_n7496_3810.t8 11.8205
R24348 a_n7496_3810.n4 a_n7496_3810.t6 11.8205
R24349 a_n7496_3810.n3 a_n7496_3810.t11 11.8205
R24350 a_n7496_3810.n3 a_n7496_3810.t7 11.8205
R24351 a_n7496_3810.n2 a_n7496_3810.t9 11.8205
R24352 a_n7496_3810.n2 a_n7496_3810.t10 11.8205
R24353 a_n7496_3810.n7 a_n7496_3810.t4 11.8205
R24354 a_n7496_3810.t2 a_n7496_3810.n7 11.8205
R24355 a_n7496_3810.n1 a_n7496_3810.n0 0.402735
R24356 a_n20296_n9452.t0 a_n20296_n9452.t1 19.8005
R24357 a_10363_n3765.t0 a_10363_n3765.t1 9.9005
R24358 a_10459_n3765.t0 a_10459_n3765.t1 9.9005
R24359 mux8_7.NAND4F_0.Y.n1 mux8_7.NAND4F_0.Y.t9 1388.16
R24360 mux8_7.NAND4F_0.Y.n1 mux8_7.NAND4F_0.Y.t11 350.839
R24361 mux8_7.NAND4F_0.Y.n2 mux8_7.NAND4F_0.Y.t10 308.481
R24362 mux8_7.NAND4F_0.Y.n0 mux8_7.NAND4F_0.Y.n3 187.373
R24363 mux8_7.NAND4F_0.Y.n0 mux8_7.NAND4F_0.Y.n4 187.192
R24364 mux8_7.NAND4F_0.Y.n0 mux8_7.NAND4F_0.Y.n5 187.192
R24365 mux8_7.NAND4F_0.Y mux8_7.NAND4F_0.Y.n6 187.192
R24366 mux8_7.NAND4F_0.Y mux8_7.NAND4F_0.Y.n2 161.492
R24367 mux8_7.NAND4F_0.Y.n2 mux8_7.NAND4F_0.Y.n1 27.752
R24368 mux8_7.NAND4F_0.Y mux8_7.NAND4F_0.Y.t3 23.5085
R24369 mux8_7.NAND4F_0.Y.n3 mux8_7.NAND4F_0.Y.t7 20.1899
R24370 mux8_7.NAND4F_0.Y.n3 mux8_7.NAND4F_0.Y.t8 20.1899
R24371 mux8_7.NAND4F_0.Y.n4 mux8_7.NAND4F_0.Y.t1 20.1899
R24372 mux8_7.NAND4F_0.Y.n4 mux8_7.NAND4F_0.Y.t0 20.1899
R24373 mux8_7.NAND4F_0.Y.n5 mux8_7.NAND4F_0.Y.t6 20.1899
R24374 mux8_7.NAND4F_0.Y.n5 mux8_7.NAND4F_0.Y.t5 20.1899
R24375 mux8_7.NAND4F_0.Y.n6 mux8_7.NAND4F_0.Y.t4 20.1899
R24376 mux8_7.NAND4F_0.Y.n6 mux8_7.NAND4F_0.Y.t2 20.1899
R24377 mux8_7.NAND4F_0.Y mux8_7.NAND4F_0.Y.n0 0.358709
R24378 a_n15131_n5154.n2 a_n15131_n5154.n0 121.353
R24379 a_n15131_n5154.n3 a_n15131_n5154.n2 121.353
R24380 a_n15131_n5154.n2 a_n15131_n5154.n1 121.001
R24381 a_n15131_n5154.n1 a_n15131_n5154.t3 30.462
R24382 a_n15131_n5154.n1 a_n15131_n5154.t0 30.462
R24383 a_n15131_n5154.n0 a_n15131_n5154.t5 30.462
R24384 a_n15131_n5154.n0 a_n15131_n5154.t4 30.462
R24385 a_n15131_n5154.n3 a_n15131_n5154.t1 30.462
R24386 a_n15131_n5154.t2 a_n15131_n5154.n3 30.462
R24387 a_n12314_n31661.n0 a_n12314_n31661.n2 81.2978
R24388 a_n12314_n31661.n1 a_n12314_n31661.n6 81.1637
R24389 a_n12314_n31661.n1 a_n12314_n31661.n5 81.1637
R24390 a_n12314_n31661.n0 a_n12314_n31661.n4 81.1637
R24391 a_n12314_n31661.n0 a_n12314_n31661.n3 81.1637
R24392 a_n12314_n31661.n7 a_n12314_n31661.n1 80.9213
R24393 a_n12314_n31661.n6 a_n12314_n31661.t1 11.8205
R24394 a_n12314_n31661.n6 a_n12314_n31661.t8 11.8205
R24395 a_n12314_n31661.n5 a_n12314_n31661.t7 11.8205
R24396 a_n12314_n31661.n5 a_n12314_n31661.t6 11.8205
R24397 a_n12314_n31661.n4 a_n12314_n31661.t11 11.8205
R24398 a_n12314_n31661.n4 a_n12314_n31661.t10 11.8205
R24399 a_n12314_n31661.n3 a_n12314_n31661.t9 11.8205
R24400 a_n12314_n31661.n3 a_n12314_n31661.t3 11.8205
R24401 a_n12314_n31661.n2 a_n12314_n31661.t5 11.8205
R24402 a_n12314_n31661.n2 a_n12314_n31661.t4 11.8205
R24403 a_n12314_n31661.n7 a_n12314_n31661.t0 11.8205
R24404 a_n12314_n31661.t2 a_n12314_n31661.n7 11.8205
R24405 a_n12314_n31661.n1 a_n12314_n31661.n0 0.402735
R24406 mux8_0.NAND4F_1.Y.n2 mux8_0.NAND4F_1.Y.t9 978.795
R24407 mux8_0.NAND4F_1.Y.n1 mux8_0.NAND4F_1.Y.t11 308.481
R24408 mux8_0.NAND4F_1.Y.n1 mux8_0.NAND4F_1.Y.t10 308.481
R24409 mux8_0.NAND4F_1.Y.n0 mux8_0.NAND4F_1.Y.n3 187.373
R24410 mux8_0.NAND4F_1.Y.n0 mux8_0.NAND4F_1.Y.n4 187.192
R24411 mux8_0.NAND4F_1.Y.n0 mux8_0.NAND4F_1.Y.n5 187.192
R24412 mux8_0.NAND4F_1.Y.n7 mux8_0.NAND4F_1.Y.n6 187.192
R24413 mux8_0.NAND4F_1.Y mux8_0.NAND4F_1.Y.n2 161.84
R24414 mux8_0.NAND4F_1.Y mux8_0.NAND4F_1.Y.t6 23.4335
R24415 mux8_0.NAND4F_1.Y.n3 mux8_0.NAND4F_1.Y.t1 20.1899
R24416 mux8_0.NAND4F_1.Y.n3 mux8_0.NAND4F_1.Y.t0 20.1899
R24417 mux8_0.NAND4F_1.Y.n4 mux8_0.NAND4F_1.Y.t5 20.1899
R24418 mux8_0.NAND4F_1.Y.n4 mux8_0.NAND4F_1.Y.t4 20.1899
R24419 mux8_0.NAND4F_1.Y.n5 mux8_0.NAND4F_1.Y.t3 20.1899
R24420 mux8_0.NAND4F_1.Y.n5 mux8_0.NAND4F_1.Y.t2 20.1899
R24421 mux8_0.NAND4F_1.Y.n6 mux8_0.NAND4F_1.Y.t8 20.1899
R24422 mux8_0.NAND4F_1.Y.n6 mux8_0.NAND4F_1.Y.t7 20.1899
R24423 mux8_0.NAND4F_1.Y.n2 mux8_0.NAND4F_1.Y.n1 11.0463
R24424 mux8_0.NAND4F_1.Y mux8_0.NAND4F_1.Y.n7 0.527586
R24425 mux8_0.NAND4F_1.Y.n7 mux8_0.NAND4F_1.Y.n0 0.358709
R24426 a_11194_762.t0 a_11194_762.t1 9.9005
R24427 a_11290_762.t0 a_11290_762.t1 9.9005
R24428 mux8_7.NAND4F_2.D.n4 mux8_7.NAND4F_2.D.t5 1388.16
R24429 mux8_7.NAND4F_2.D.n7 mux8_7.NAND4F_2.D.t8 1388.16
R24430 mux8_7.NAND4F_2.D.n10 mux8_7.NAND4F_2.D.t12 1388.16
R24431 mux8_7.NAND4F_2.D.n1 mux8_7.NAND4F_2.D.t7 1388.16
R24432 mux8_7.NAND4F_2.D.n4 mux8_7.NAND4F_2.D.t10 350.839
R24433 mux8_7.NAND4F_2.D.n7 mux8_7.NAND4F_2.D.t13 350.839
R24434 mux8_7.NAND4F_2.D.n10 mux8_7.NAND4F_2.D.t9 350.839
R24435 mux8_7.NAND4F_2.D.n1 mux8_7.NAND4F_2.D.t4 350.839
R24436 mux8_7.NAND4F_2.D.n5 mux8_7.NAND4F_2.D.t15 308.481
R24437 mux8_7.NAND4F_2.D.n8 mux8_7.NAND4F_2.D.t14 308.481
R24438 mux8_7.NAND4F_2.D.n11 mux8_7.NAND4F_2.D.t11 308.481
R24439 mux8_7.NAND4F_2.D.n2 mux8_7.NAND4F_2.D.t6 308.481
R24440 mux8_7.NAND4F_2.D.n0 mux8_7.NAND4F_2.D.t1 256.514
R24441 mux8_7.NAND4F_2.D.n0 mux8_7.NAND4F_2.D.n3 226.258
R24442 mux8_7.NAND4F_2.D mux8_7.NAND4F_2.D.n5 161.458
R24443 mux8_7.NAND4F_2.D mux8_7.NAND4F_2.D.n11 161.435
R24444 mux8_7.NAND4F_2.D mux8_7.NAND4F_2.D.n2 161.435
R24445 mux8_7.NAND4F_2.D mux8_7.NAND4F_2.D.n8 161.429
R24446 mux8_7.NAND4F_2.D.n0 mux8_7.NAND4F_2.D.t0 83.7172
R24447 mux8_7.NAND4F_2.D.n3 mux8_7.NAND4F_2.D.t3 30.379
R24448 mux8_7.NAND4F_2.D.n3 mux8_7.NAND4F_2.D.t2 30.379
R24449 mux8_7.NAND4F_2.D.n5 mux8_7.NAND4F_2.D.n4 27.752
R24450 mux8_7.NAND4F_2.D.n8 mux8_7.NAND4F_2.D.n7 27.752
R24451 mux8_7.NAND4F_2.D.n11 mux8_7.NAND4F_2.D.n10 27.752
R24452 mux8_7.NAND4F_2.D.n2 mux8_7.NAND4F_2.D.n1 27.752
R24453 mux8_7.NAND4F_2.D.n6 mux8_7.NAND4F_2.D.n0 12.759
R24454 mux8_7.NAND4F_2.D mux8_7.NAND4F_2.D.n12 10.6871
R24455 mux8_7.NAND4F_2.D.n6 mux8_7.NAND4F_2.D 9.0005
R24456 mux8_7.NAND4F_2.D.n12 mux8_7.NAND4F_2.D 9.0005
R24457 mux8_7.NAND4F_2.D.n9 mux8_7.NAND4F_2.D 9.0005
R24458 mux8_7.NAND4F_2.D.n9 mux8_7.NAND4F_2.D.n6 1.74507
R24459 mux8_7.NAND4F_2.D.n12 mux8_7.NAND4F_2.D.n9 1.69072
R24460 mux8_8.NAND4F_4.B.n10 mux8_8.NAND4F_4.B.t4 933.563
R24461 mux8_8.NAND4F_4.B.n5 mux8_8.NAND4F_4.B.t10 933.563
R24462 mux8_8.NAND4F_4.B.n3 mux8_8.NAND4F_4.B.t13 933.563
R24463 mux8_8.NAND4F_4.B.n1 mux8_8.NAND4F_4.B.t9 933.563
R24464 mux8_8.NAND4F_4.B.n10 mux8_8.NAND4F_4.B.t14 367.635
R24465 mux8_8.NAND4F_4.B.n5 mux8_8.NAND4F_4.B.t6 367.635
R24466 mux8_8.NAND4F_4.B.n3 mux8_8.NAND4F_4.B.t11 367.635
R24467 mux8_8.NAND4F_4.B.n1 mux8_8.NAND4F_4.B.t5 367.635
R24468 mux8_8.NAND4F_4.B.n11 mux8_8.NAND4F_4.B.t15 308.481
R24469 mux8_8.NAND4F_4.B.n6 mux8_8.NAND4F_4.B.t8 308.481
R24470 mux8_8.NAND4F_4.B.n4 mux8_8.NAND4F_4.B.t12 308.481
R24471 mux8_8.NAND4F_4.B.n2 mux8_8.NAND4F_4.B.t7 308.481
R24472 mux8_8.NAND4F_4.B.n0 mux8_8.NAND4F_4.B.t1 256.514
R24473 mux8_8.NAND4F_4.B.n0 mux8_8.NAND4F_4.B.n8 226.258
R24474 mux8_8.NAND4F_4.B mux8_8.NAND4F_4.B.n2 162.173
R24475 mux8_8.NAND4F_4.B mux8_8.NAND4F_4.B.n6 162.137
R24476 mux8_8.NAND4F_4.B mux8_8.NAND4F_4.B.n11 162.117
R24477 mux8_8.NAND4F_4.B.n7 mux8_8.NAND4F_4.B.n4 161.703
R24478 mux8_8.NAND4F_4.B.n0 mux8_8.NAND4F_4.B.t0 83.7172
R24479 mux8_8.NAND4F_4.B.n8 mux8_8.NAND4F_4.B.t3 30.379
R24480 mux8_8.NAND4F_4.B.n8 mux8_8.NAND4F_4.B.t2 30.379
R24481 mux8_8.NAND4F_4.B.n12 mux8_8.NAND4F_4.B 24.8912
R24482 mux8_8.NAND4F_4.B.n7 mux8_8.NAND4F_4.B 21.6618
R24483 mux8_8.NAND4F_4.B.n11 mux8_8.NAND4F_4.B.n10 10.955
R24484 mux8_8.NAND4F_4.B.n6 mux8_8.NAND4F_4.B.n5 10.955
R24485 mux8_8.NAND4F_4.B.n4 mux8_8.NAND4F_4.B.n3 10.955
R24486 mux8_8.NAND4F_4.B.n2 mux8_8.NAND4F_4.B.n1 10.955
R24487 mux8_8.NAND4F_4.B.n12 mux8_8.NAND4F_4.B.n9 3.67985
R24488 mux8_8.NAND4F_4.B.n9 mux8_8.NAND4F_4.B.n0 1.46835
R24489 mux8_8.NAND4F_4.B mux8_8.NAND4F_4.B.n12 0.502677
R24490 mux8_8.NAND4F_4.B.n9 mux8_8.NAND4F_4.B 0.498606
R24491 mux8_8.NAND4F_4.B mux8_8.NAND4F_4.B.n7 0.470197
R24492 mux8_0.NAND4F_9.Y.n1 mux8_0.NAND4F_9.Y.t12 312.599
R24493 mux8_0.NAND4F_9.Y.n4 mux8_0.NAND4F_9.Y.t13 247.428
R24494 mux8_0.NAND4F_9.Y.n1 mux8_0.NAND4F_9.Y.t14 247.428
R24495 mux8_0.NAND4F_9.Y.n2 mux8_0.NAND4F_9.Y.t9 247.428
R24496 mux8_0.NAND4F_9.Y.n3 mux8_0.NAND4F_9.Y.t11 247.428
R24497 mux8_0.NAND4F_9.Y.n5 mux8_0.NAND4F_9.Y.t10 229.754
R24498 mux8_0.NAND4F_9.Y.n0 mux8_0.NAND4F_9.Y.n6 187.373
R24499 mux8_0.NAND4F_9.Y.n0 mux8_0.NAND4F_9.Y.n7 187.192
R24500 mux8_0.NAND4F_9.Y.n0 mux8_0.NAND4F_9.Y.n8 187.192
R24501 mux8_0.NAND4F_9.Y.n10 mux8_0.NAND4F_9.Y.n9 187.192
R24502 mux8_0.NAND4F_9.Y mux8_0.NAND4F_9.Y.n5 162.275
R24503 mux8_0.NAND4F_9.Y.n5 mux8_0.NAND4F_9.Y.n4 91.5805
R24504 mux8_0.NAND4F_9.Y.n2 mux8_0.NAND4F_9.Y.n1 65.1723
R24505 mux8_0.NAND4F_9.Y.n3 mux8_0.NAND4F_9.Y.n2 65.1723
R24506 mux8_0.NAND4F_9.Y.n4 mux8_0.NAND4F_9.Y.n3 65.1723
R24507 mux8_0.NAND4F_9.Y mux8_0.NAND4F_9.Y.t0 22.6141
R24508 mux8_0.NAND4F_9.Y.n6 mux8_0.NAND4F_9.Y.t7 20.1899
R24509 mux8_0.NAND4F_9.Y.n6 mux8_0.NAND4F_9.Y.t8 20.1899
R24510 mux8_0.NAND4F_9.Y.n7 mux8_0.NAND4F_9.Y.t3 20.1899
R24511 mux8_0.NAND4F_9.Y.n7 mux8_0.NAND4F_9.Y.t4 20.1899
R24512 mux8_0.NAND4F_9.Y.n8 mux8_0.NAND4F_9.Y.t6 20.1899
R24513 mux8_0.NAND4F_9.Y.n8 mux8_0.NAND4F_9.Y.t5 20.1899
R24514 mux8_0.NAND4F_9.Y.n9 mux8_0.NAND4F_9.Y.t2 20.1899
R24515 mux8_0.NAND4F_9.Y.n9 mux8_0.NAND4F_9.Y.t1 20.1899
R24516 mux8_0.NAND4F_9.Y mux8_0.NAND4F_9.Y.n10 0.396904
R24517 mux8_0.NAND4F_9.Y.n10 mux8_0.NAND4F_9.Y.n0 0.358709
R24518 mux8_2.NAND4F_0.C.n6 mux8_2.NAND4F_0.C.t4 978.795
R24519 mux8_2.NAND4F_0.C.n4 mux8_2.NAND4F_0.C.t9 978.795
R24520 mux8_2.NAND4F_0.C.n11 mux8_2.NAND4F_0.C.t14 978.795
R24521 mux8_2.NAND4F_0.C.n2 mux8_2.NAND4F_0.C.t12 978.795
R24522 mux8_2.NAND4F_0.C.n5 mux8_2.NAND4F_0.C.t5 308.481
R24523 mux8_2.NAND4F_0.C.n5 mux8_2.NAND4F_0.C.t7 308.481
R24524 mux8_2.NAND4F_0.C.n3 mux8_2.NAND4F_0.C.t13 308.481
R24525 mux8_2.NAND4F_0.C.n3 mux8_2.NAND4F_0.C.t15 308.481
R24526 mux8_2.NAND4F_0.C.n10 mux8_2.NAND4F_0.C.t8 308.481
R24527 mux8_2.NAND4F_0.C.n10 mux8_2.NAND4F_0.C.t6 308.481
R24528 mux8_2.NAND4F_0.C.n1 mux8_2.NAND4F_0.C.t11 308.481
R24529 mux8_2.NAND4F_0.C.n1 mux8_2.NAND4F_0.C.t10 308.481
R24530 mux8_2.NAND4F_0.C.n0 mux8_2.NAND4F_0.C.t2 256.514
R24531 mux8_2.NAND4F_0.C.n0 mux8_2.NAND4F_0.C.n8 226.258
R24532 mux8_2.NAND4F_0.C mux8_2.NAND4F_0.C.n6 161.856
R24533 mux8_2.NAND4F_0.C mux8_2.NAND4F_0.C.n4 161.847
R24534 mux8_2.NAND4F_0.C mux8_2.NAND4F_0.C.n11 161.84
R24535 mux8_2.NAND4F_0.C mux8_2.NAND4F_0.C.n2 161.831
R24536 mux8_2.NAND4F_0.C.n0 mux8_2.NAND4F_0.C.t0 83.7172
R24537 mux8_2.NAND4F_0.C.n8 mux8_2.NAND4F_0.C.t1 30.379
R24538 mux8_2.NAND4F_0.C.n8 mux8_2.NAND4F_0.C.t3 30.379
R24539 mux8_2.NAND4F_0.C.n9 mux8_2.NAND4F_0.C.n0 13.5186
R24540 mux8_2.NAND4F_0.C mux8_2.NAND4F_0.C.n12 13.0862
R24541 mux8_2.NAND4F_0.C.n7 mux8_2.NAND4F_0.C 13.0435
R24542 mux8_2.NAND4F_0.C.n12 mux8_2.NAND4F_0.C 12.4135
R24543 mux8_2.NAND4F_0.C.n7 mux8_2.NAND4F_0.C 12.4105
R24544 mux8_2.NAND4F_0.C.n6 mux8_2.NAND4F_0.C.n5 11.0463
R24545 mux8_2.NAND4F_0.C.n4 mux8_2.NAND4F_0.C.n3 11.0463
R24546 mux8_2.NAND4F_0.C.n11 mux8_2.NAND4F_0.C.n10 11.0463
R24547 mux8_2.NAND4F_0.C.n2 mux8_2.NAND4F_0.C.n1 11.0463
R24548 mux8_2.NAND4F_0.C.n12 mux8_2.NAND4F_0.C.n9 3.46056
R24549 mux8_2.NAND4F_0.C.n9 mux8_2.NAND4F_0.C.n7 1.8134
R24550 a_n9314_n12716.t0 a_n9314_n12716.t1 19.8005
R24551 a_7452_n16422.t0 a_7452_n16422.t1 9.9005
R24552 mux8_1.inv_0.A.n3 mux8_1.inv_0.A.t9 291.829
R24553 mux8_1.inv_0.A.n3 mux8_1.inv_0.A.t8 291.829
R24554 mux8_1.inv_0.A.n0 mux8_1.inv_0.A.t1 256.425
R24555 mux8_1.inv_0.A.n0 mux8_1.inv_0.A.n4 231.24
R24556 mux8_1.inv_0.A.n0 mux8_1.inv_0.A.n5 231.03
R24557 mux8_1.inv_0.A.n3 mux8_1.inv_0.A.t7 221.72
R24558 mux8_1.inv_0.A.t10 mux8_1.inv_0.A.n2 393.959
R24559 mux8_1.inv_0.A.n6 mux8_1.inv_0.A.n1 66.6316
R24560 mux8_1.inv_0.A.n2 mux8_1.inv_0.A.n3 53.4611
R24561 mux8_1.inv_0.A.n5 mux8_1.inv_0.A.t2 25.395
R24562 mux8_1.inv_0.A.n5 mux8_1.inv_0.A.t3 25.395
R24563 mux8_1.inv_0.A.n4 mux8_1.inv_0.A.t4 25.395
R24564 mux8_1.inv_0.A.n4 mux8_1.inv_0.A.t5 25.395
R24565 mux8_1.inv_0.A.n6 mux8_1.inv_0.A.t6 19.8005
R24566 mux8_1.inv_0.A.n6 mux8_1.inv_0.A.t0 19.8005
R24567 mux8_1.inv_0.A.n1 mux8_1.inv_0.A.n0 0.38953
R24568 mux8_1.inv_0.A.n1 mux8_1.inv_0.A.n2 0.294762
R24569 Y0.n0 Y0.t4 883.668
R24570 Y0.n1 Y0.t6 729.428
R24571 Y0.n0 Y0.t5 729.428
R24572 Y0.n2 Y0.t7 462.137
R24573 Y0.n2 Y0.n1 437.014
R24574 Y0.n4 Y0.t2 256.514
R24575 Y0.n5 Y0.n3 226.251
R24576 Y0.n6 Y0.n2 163.262
R24577 Y0.n1 Y0.n0 154.24
R24578 Y0.n4 Y0.t0 83.7599
R24579 Y0.n6 Y0 31.6771
R24580 Y0.n3 Y0.t1 30.379
R24581 Y0.n3 Y0.t3 30.379
R24582 Y0 Y0.n6 0.0402727
R24583 Y0.n5 Y0.n4 0.0323878
R24584 Y0 Y0.n5 0.0189949
R24585 Y7.n0 Y7.t8 883.668
R24586 Y7.n1 Y7.t10 729.428
R24587 Y7.n0 Y7.t9 729.428
R24588 Y7.n2 Y7.t11 462.137
R24589 Y7.n2 Y7.n1 437.014
R24590 Y7.n9 Y7.t6 394.152
R24591 Y7.n8 Y7.t5 291.829
R24592 Y7.n8 Y7.t7 291.829
R24593 Y7.n6 Y7.t1 256.514
R24594 Y7.n5 Y7.n4 226.218
R24595 Y7.n8 Y7.t4 221.72
R24596 Y7.n3 Y7.n2 163.258
R24597 Y7.n1 Y7.n0 154.24
R24598 Y7.n7 Y7.t0 83.7172
R24599 Y7.n9 Y7.n8 53.4762
R24600 Y7.n5 Y7.n3 32.3263
R24601 Y7.n4 Y7.t3 30.379
R24602 Y7.n4 Y7.t2 30.379
R24603 Y7 Y7.n7 1.19779
R24604 Y7 Y7.n9 0.356178
R24605 Y7 Y7.n6 0.0469744
R24606 Y7.n3 Y7 0.0440606
R24607 Y7.n6 Y7.n5 0.0410411
R24608 Y7.n7 Y7 0.0189295
R24609 buffer_0.inv_1.A.n2 buffer_0.inv_1.A.t5 291.829
R24610 buffer_0.inv_1.A.n2 buffer_0.inv_1.A.t7 291.829
R24611 buffer_0.inv_1.A.n0 buffer_0.inv_1.A.t2 256.89
R24612 buffer_0.inv_1.A.n0 buffer_0.inv_1.A.n1 226.538
R24613 buffer_0.inv_1.A.n2 buffer_0.inv_1.A.t4 221.72
R24614 buffer_0.inv_1.A.t6 buffer_0.inv_1.A.n0 393.921
R24615 buffer_0.inv_1.A.n0 buffer_0.inv_1.A.t0 83.795
R24616 buffer_0.inv_1.A.n0 buffer_0.inv_1.A.n2 53.7938
R24617 buffer_0.inv_1.A.n1 buffer_0.inv_1.A.t1 30.379
R24618 buffer_0.inv_1.A.n1 buffer_0.inv_1.A.t3 30.379
R24619 a_n14781_1380.n2 a_n14781_1380.t4 541.395
R24620 a_n14781_1380.n3 a_n14781_1380.t3 527.402
R24621 a_n14781_1380.n2 a_n14781_1380.t6 491.64
R24622 a_n14781_1380.n5 a_n14781_1380.t0 281.906
R24623 a_n14781_1380.t1 a_n14781_1380.n5 204.359
R24624 a_n14781_1380.n0 a_n14781_1380.t2 180.73
R24625 a_n14781_1380.n1 a_n14781_1380.t5 179.45
R24626 a_n14781_1380.n0 a_n14781_1380.t7 139.78
R24627 a_n14781_1380.n4 a_n14781_1380.n1 105.635
R24628 a_n14781_1380.n4 a_n14781_1380.n3 76.0005
R24629 a_n14781_1380.n5 a_n14781_1380.n4 67.9685
R24630 a_n14781_1380.n3 a_n14781_1380.n2 13.994
R24631 a_n14781_1380.n1 a_n14781_1380.n0 1.28015
R24632 a_n15896_n6187.t0 a_n15896_n6187.t1 19.8005
R24633 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t9 485.221
R24634 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t10 367.928
R24635 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n5 227.526
R24636 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n6 227.266
R24637 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n4 227.266
R24638 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t8 224.478
R24639 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t7 213.688
R24640 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n2 84.5046
R24641 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n1 72.3005
R24642 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n3 61.0566
R24643 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t3 42.7747
R24644 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t4 30.379
R24645 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t1 30.379
R24646 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t6 30.379
R24647 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t5 30.379
R24648 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t0 30.379
R24649 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.t2 30.379
R24650 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A.n0 0.583137
R24651 mux8_2.NAND4F_4.B.n10 mux8_2.NAND4F_4.B.t14 933.563
R24652 mux8_2.NAND4F_4.B.n5 mux8_2.NAND4F_4.B.t4 933.563
R24653 mux8_2.NAND4F_4.B.n3 mux8_2.NAND4F_4.B.t5 933.563
R24654 mux8_2.NAND4F_4.B.n1 mux8_2.NAND4F_4.B.t15 933.563
R24655 mux8_2.NAND4F_4.B.n10 mux8_2.NAND4F_4.B.t13 367.635
R24656 mux8_2.NAND4F_4.B.n5 mux8_2.NAND4F_4.B.t12 367.635
R24657 mux8_2.NAND4F_4.B.n3 mux8_2.NAND4F_4.B.t8 367.635
R24658 mux8_2.NAND4F_4.B.n1 mux8_2.NAND4F_4.B.t9 367.635
R24659 mux8_2.NAND4F_4.B.n11 mux8_2.NAND4F_4.B.t11 308.481
R24660 mux8_2.NAND4F_4.B.n6 mux8_2.NAND4F_4.B.t10 308.481
R24661 mux8_2.NAND4F_4.B.n4 mux8_2.NAND4F_4.B.t6 308.481
R24662 mux8_2.NAND4F_4.B.n2 mux8_2.NAND4F_4.B.t7 308.481
R24663 mux8_2.NAND4F_4.B.n0 mux8_2.NAND4F_4.B.t2 256.514
R24664 mux8_2.NAND4F_4.B.n0 mux8_2.NAND4F_4.B.n8 226.258
R24665 mux8_2.NAND4F_4.B mux8_2.NAND4F_4.B.n2 162.173
R24666 mux8_2.NAND4F_4.B mux8_2.NAND4F_4.B.n6 162.137
R24667 mux8_2.NAND4F_4.B mux8_2.NAND4F_4.B.n11 162.117
R24668 mux8_2.NAND4F_4.B.n7 mux8_2.NAND4F_4.B.n4 161.703
R24669 mux8_2.NAND4F_4.B.n0 mux8_2.NAND4F_4.B.t0 83.7172
R24670 mux8_2.NAND4F_4.B.n8 mux8_2.NAND4F_4.B.t1 30.379
R24671 mux8_2.NAND4F_4.B.n8 mux8_2.NAND4F_4.B.t3 30.379
R24672 mux8_2.NAND4F_4.B.n12 mux8_2.NAND4F_4.B 24.8912
R24673 mux8_2.NAND4F_4.B.n7 mux8_2.NAND4F_4.B 21.6618
R24674 mux8_2.NAND4F_4.B.n11 mux8_2.NAND4F_4.B.n10 10.955
R24675 mux8_2.NAND4F_4.B.n6 mux8_2.NAND4F_4.B.n5 10.955
R24676 mux8_2.NAND4F_4.B.n4 mux8_2.NAND4F_4.B.n3 10.955
R24677 mux8_2.NAND4F_4.B.n2 mux8_2.NAND4F_4.B.n1 10.955
R24678 mux8_2.NAND4F_4.B.n12 mux8_2.NAND4F_4.B.n9 3.67985
R24679 mux8_2.NAND4F_4.B.n9 mux8_2.NAND4F_4.B.n0 1.46835
R24680 mux8_2.NAND4F_4.B mux8_2.NAND4F_4.B.n12 0.502677
R24681 mux8_2.NAND4F_4.B.n9 mux8_2.NAND4F_4.B 0.498606
R24682 mux8_2.NAND4F_4.B mux8_2.NAND4F_4.B.n7 0.470197
R24683 a_n11274_n26419.n2 a_n11274_n26419.n0 121.353
R24684 a_n11274_n26419.n2 a_n11274_n26419.n1 121.001
R24685 a_n11274_n26419.n3 a_n11274_n26419.n2 120.977
R24686 a_n11274_n26419.n1 a_n11274_n26419.t5 30.462
R24687 a_n11274_n26419.n1 a_n11274_n26419.t0 30.462
R24688 a_n11274_n26419.n0 a_n11274_n26419.t1 30.462
R24689 a_n11274_n26419.n0 a_n11274_n26419.t2 30.462
R24690 a_n11274_n26419.t4 a_n11274_n26419.n3 30.462
R24691 a_n11274_n26419.n3 a_n11274_n26419.t3 30.462
R24692 8bit_ADDER_0.C.n4 8bit_ADDER_0.C.t9 1032.02
R24693 8bit_ADDER_0.C.n4 8bit_ADDER_0.C.t8 336.962
R24694 8bit_ADDER_0.C.n4 8bit_ADDER_0.C.t7 326.154
R24695 8bit_ADDER_0.C.n0 8bit_ADDER_0.C.n1 227.526
R24696 8bit_ADDER_0.C.n0 8bit_ADDER_0.C.n3 227.266
R24697 8bit_ADDER_0.C.n0 8bit_ADDER_0.C.n2 227.266
R24698 8bit_ADDER_0.C 8bit_ADDER_0.C.n4 162.952
R24699 8bit_ADDER_0.C.n0 8bit_ADDER_0.C.t0 42.7831
R24700 8bit_ADDER_0.C.n3 8bit_ADDER_0.C.t1 30.379
R24701 8bit_ADDER_0.C.n3 8bit_ADDER_0.C.t3 30.379
R24702 8bit_ADDER_0.C.n1 8bit_ADDER_0.C.t6 30.379
R24703 8bit_ADDER_0.C.n1 8bit_ADDER_0.C.t5 30.379
R24704 8bit_ADDER_0.C.n2 8bit_ADDER_0.C.t2 30.379
R24705 8bit_ADDER_0.C.n2 8bit_ADDER_0.C.t4 30.379
R24706 8bit_ADDER_0.C 8bit_ADDER_0.C.n0 18.8873
R24707 a_1857_4888.n2 a_1857_4888.t7 541.395
R24708 a_1857_4888.n3 a_1857_4888.t3 527.402
R24709 a_1857_4888.n2 a_1857_4888.t4 491.64
R24710 a_1857_4888.n5 a_1857_4888.t0 281.906
R24711 a_1857_4888.t1 a_1857_4888.n5 204.359
R24712 a_1857_4888.n0 a_1857_4888.t5 180.73
R24713 a_1857_4888.n1 a_1857_4888.t2 179.45
R24714 a_1857_4888.n0 a_1857_4888.t6 139.78
R24715 a_1857_4888.n4 a_1857_4888.n1 105.635
R24716 a_1857_4888.n4 a_1857_4888.n3 76.0005
R24717 a_1857_4888.n5 a_1857_4888.n4 67.9685
R24718 a_1857_4888.n3 a_1857_4888.n2 13.994
R24719 a_1857_4888.n1 a_1857_4888.n0 1.28015
R24720 a_1887_4914.n3 a_1887_4914.n2 121.353
R24721 a_1887_4914.n2 a_1887_4914.n1 121.001
R24722 a_1887_4914.n2 a_1887_4914.n0 120.977
R24723 a_1887_4914.n1 a_1887_4914.t5 30.462
R24724 a_1887_4914.n1 a_1887_4914.t2 30.462
R24725 a_1887_4914.n0 a_1887_4914.t0 30.462
R24726 a_1887_4914.n0 a_1887_4914.t4 30.462
R24727 a_1887_4914.n3 a_1887_4914.t1 30.462
R24728 a_1887_4914.t3 a_1887_4914.n3 30.462
R24729 mux8_1.NAND4F_5.Y.n1 mux8_1.NAND4F_5.Y.t11 1032.02
R24730 mux8_1.NAND4F_5.Y.n1 mux8_1.NAND4F_5.Y.t10 336.962
R24731 mux8_1.NAND4F_5.Y.n1 mux8_1.NAND4F_5.Y.t9 326.154
R24732 mux8_1.NAND4F_5.Y.n0 mux8_1.NAND4F_5.Y.n3 187.373
R24733 mux8_1.NAND4F_5.Y.n0 mux8_1.NAND4F_5.Y.n4 187.192
R24734 mux8_1.NAND4F_5.Y.n0 mux8_1.NAND4F_5.Y.n5 187.192
R24735 mux8_1.NAND4F_5.Y.n7 mux8_1.NAND4F_5.Y.n6 187.192
R24736 mux8_1.NAND4F_5.Y mux8_1.NAND4F_5.Y.n1 162.94
R24737 mux8_1.NAND4F_5.Y.n2 mux8_1.NAND4F_5.Y 24.4721
R24738 mux8_1.NAND4F_5.Y.n2 mux8_1.NAND4F_5.Y.t2 22.6141
R24739 mux8_1.NAND4F_5.Y.n3 mux8_1.NAND4F_5.Y.t0 20.1899
R24740 mux8_1.NAND4F_5.Y.n3 mux8_1.NAND4F_5.Y.t1 20.1899
R24741 mux8_1.NAND4F_5.Y.n4 mux8_1.NAND4F_5.Y.t5 20.1899
R24742 mux8_1.NAND4F_5.Y.n4 mux8_1.NAND4F_5.Y.t6 20.1899
R24743 mux8_1.NAND4F_5.Y.n5 mux8_1.NAND4F_5.Y.t7 20.1899
R24744 mux8_1.NAND4F_5.Y.n5 mux8_1.NAND4F_5.Y.t8 20.1899
R24745 mux8_1.NAND4F_5.Y.n6 mux8_1.NAND4F_5.Y.t3 20.1899
R24746 mux8_1.NAND4F_5.Y.n6 mux8_1.NAND4F_5.Y.t4 20.1899
R24747 mux8_1.NAND4F_5.Y mux8_1.NAND4F_5.Y.n2 0.950576
R24748 mux8_1.NAND4F_5.Y mux8_1.NAND4F_5.Y.n7 0.396904
R24749 mux8_1.NAND4F_5.Y.n7 mux8_1.NAND4F_5.Y.n0 0.358709
R24750 a_11290_n35462.t0 a_11290_n35462.t1 9.9005
R24751 a_11386_n2838.t0 a_11386_n2838.t1 9.9005
R24752 mux8_8.NAND4F_3.Y.n7 mux8_8.NAND4F_3.Y.t9 978.795
R24753 mux8_8.NAND4F_3.Y.n6 mux8_8.NAND4F_3.Y.t11 308.481
R24754 mux8_8.NAND4F_3.Y.n6 mux8_8.NAND4F_3.Y.t10 308.481
R24755 mux8_8.NAND4F_3.Y.n0 mux8_8.NAND4F_3.Y.n1 187.373
R24756 mux8_8.NAND4F_3.Y.n0 mux8_8.NAND4F_3.Y.n2 187.192
R24757 mux8_8.NAND4F_3.Y.n0 mux8_8.NAND4F_3.Y.n3 187.192
R24758 mux8_8.NAND4F_3.Y.n5 mux8_8.NAND4F_3.Y.n4 187.192
R24759 mux8_8.NAND4F_3.Y mux8_8.NAND4F_3.Y.n7 161.839
R24760 mux8_8.NAND4F_3.Y mux8_8.NAND4F_3.Y.t4 23.4426
R24761 mux8_8.NAND4F_3.Y.n1 mux8_8.NAND4F_3.Y.t0 20.1899
R24762 mux8_8.NAND4F_3.Y.n1 mux8_8.NAND4F_3.Y.t6 20.1899
R24763 mux8_8.NAND4F_3.Y.n2 mux8_8.NAND4F_3.Y.t7 20.1899
R24764 mux8_8.NAND4F_3.Y.n2 mux8_8.NAND4F_3.Y.t8 20.1899
R24765 mux8_8.NAND4F_3.Y.n3 mux8_8.NAND4F_3.Y.t2 20.1899
R24766 mux8_8.NAND4F_3.Y.n3 mux8_8.NAND4F_3.Y.t1 20.1899
R24767 mux8_8.NAND4F_3.Y.n4 mux8_8.NAND4F_3.Y.t5 20.1899
R24768 mux8_8.NAND4F_3.Y.n4 mux8_8.NAND4F_3.Y.t3 20.1899
R24769 mux8_8.NAND4F_3.Y.n7 mux8_8.NAND4F_3.Y.n6 11.0463
R24770 mux8_8.NAND4F_3.Y mux8_8.NAND4F_3.Y.n5 0.518495
R24771 mux8_8.NAND4F_3.Y.n5 mux8_8.NAND4F_3.Y.n0 0.358709
R24772 a_11194_n30006.t0 a_11194_n30006.t1 9.9005
R24773 a_11290_n30006.t0 a_11290_n30006.t1 9.9005
R24774 Y6.n0 Y6.t5 883.668
R24775 Y6.n1 Y6.t7 740.381
R24776 Y6.n0 Y6.t6 729.428
R24777 Y6.n2 Y6.t4 700.508
R24778 Y6.n4 Y6.t3 256.514
R24779 Y6 Y6.n3 226.239
R24780 Y6 Y6.n2 162.989
R24781 Y6.n5 Y6.t0 83.7901
R24782 Y6.n1 Y6.n0 72.3005
R24783 Y6.n3 Y6.t2 30.379
R24784 Y6.n3 Y6.t1 30.379
R24785 Y6.n2 Y6.n1 16.7975
R24786 Y6.n5 Y6.n4 0.0574096
R24787 Y6 Y6.n5 0.0300905
R24788 Y6.n4 Y6 0.00182275
R24789 a_n12345_n17569.n2 a_n12345_n17569.t7 541.395
R24790 a_n12345_n17569.n3 a_n12345_n17569.t4 527.402
R24791 a_n12345_n17569.n2 a_n12345_n17569.t6 491.64
R24792 a_n12345_n17569.n5 a_n12345_n17569.t0 281.906
R24793 a_n12345_n17569.t1 a_n12345_n17569.n5 204.359
R24794 a_n12345_n17569.n0 a_n12345_n17569.t2 180.73
R24795 a_n12345_n17569.n1 a_n12345_n17569.t5 179.45
R24796 a_n12345_n17569.n0 a_n12345_n17569.t3 139.78
R24797 a_n12345_n17569.n4 a_n12345_n17569.n1 105.635
R24798 a_n12345_n17569.n4 a_n12345_n17569.n3 76.0005
R24799 a_n12345_n17569.n5 a_n12345_n17569.n4 67.9685
R24800 a_n12345_n17569.n3 a_n12345_n17569.n2 13.994
R24801 a_n12345_n17569.n1 a_n12345_n17569.n0 1.28015
R24802 a_n12316_n15299.n0 a_n12316_n15299.n2 81.2978
R24803 a_n12316_n15299.n1 a_n12316_n15299.n6 81.1637
R24804 a_n12316_n15299.n1 a_n12316_n15299.n5 81.1637
R24805 a_n12316_n15299.n0 a_n12316_n15299.n4 81.1637
R24806 a_n12316_n15299.n0 a_n12316_n15299.n3 81.1637
R24807 a_n12316_n15299.n7 a_n12316_n15299.n1 80.9213
R24808 a_n12316_n15299.n6 a_n12316_n15299.t0 11.8205
R24809 a_n12316_n15299.n6 a_n12316_n15299.t4 11.8205
R24810 a_n12316_n15299.n5 a_n12316_n15299.t5 11.8205
R24811 a_n12316_n15299.n5 a_n12316_n15299.t3 11.8205
R24812 a_n12316_n15299.n4 a_n12316_n15299.t8 11.8205
R24813 a_n12316_n15299.n4 a_n12316_n15299.t7 11.8205
R24814 a_n12316_n15299.n3 a_n12316_n15299.t6 11.8205
R24815 a_n12316_n15299.n3 a_n12316_n15299.t9 11.8205
R24816 a_n12316_n15299.n2 a_n12316_n15299.t11 11.8205
R24817 a_n12316_n15299.n2 a_n12316_n15299.t10 11.8205
R24818 a_n12316_n15299.t2 a_n12316_n15299.n7 11.8205
R24819 a_n12316_n15299.n7 a_n12316_n15299.t1 11.8205
R24820 a_n12316_n15299.n1 a_n12316_n15299.n0 0.402735
R24821 a_n10714_n11709.n2 a_n10714_n11709.t2 541.395
R24822 a_n10714_n11709.n3 a_n10714_n11709.t5 527.402
R24823 a_n10714_n11709.n2 a_n10714_n11709.t4 491.64
R24824 a_n10714_n11709.n5 a_n10714_n11709.t0 281.906
R24825 a_n10714_n11709.t1 a_n10714_n11709.n5 204.359
R24826 a_n10714_n11709.n0 a_n10714_n11709.t3 180.73
R24827 a_n10714_n11709.n1 a_n10714_n11709.t6 179.45
R24828 a_n10714_n11709.n0 a_n10714_n11709.t7 139.78
R24829 a_n10714_n11709.n4 a_n10714_n11709.n1 105.635
R24830 a_n10714_n11709.n4 a_n10714_n11709.n3 76.0005
R24831 a_n10714_n11709.n5 a_n10714_n11709.n4 67.9685
R24832 a_n10714_n11709.n3 a_n10714_n11709.n2 13.994
R24833 a_n10714_n11709.n1 a_n10714_n11709.n0 1.28015
R24834 a_n18305_n9452.t0 a_n18305_n9452.t1 19.8005
R24835 a_n23065_1406.n3 a_n23065_1406.n2 121.353
R24836 a_n23065_1406.n2 a_n23065_1406.n1 121.001
R24837 a_n23065_1406.n2 a_n23065_1406.n0 120.977
R24838 a_n23065_1406.n1 a_n23065_1406.t4 30.462
R24839 a_n23065_1406.n1 a_n23065_1406.t1 30.462
R24840 a_n23065_1406.n0 a_n23065_1406.t5 30.462
R24841 a_n23065_1406.n0 a_n23065_1406.t3 30.462
R24842 a_n23065_1406.n3 a_n23065_1406.t0 30.462
R24843 a_n23065_1406.t2 a_n23065_1406.n3 30.462
R24844 MULT_0.4bit_ADDER_0.A0.n3 MULT_0.4bit_ADDER_0.A0.t4 540.38
R24845 MULT_0.4bit_ADDER_0.A0.n4 MULT_0.4bit_ADDER_0.A0.t11 491.64
R24846 MULT_0.4bit_ADDER_0.A0.n4 MULT_0.4bit_ADDER_0.A0.t6 491.64
R24847 MULT_0.4bit_ADDER_0.A0.n4 MULT_0.4bit_ADDER_0.A0.t13 491.64
R24848 MULT_0.4bit_ADDER_0.A0.n4 MULT_0.4bit_ADDER_0.A0.t5 491.64
R24849 MULT_0.4bit_ADDER_0.A0.n1 MULT_0.4bit_ADDER_0.A0.t7 367.928
R24850 MULT_0.4bit_ADDER_0.A0.n0 MULT_0.4bit_ADDER_0.A0.t1 256.514
R24851 MULT_0.4bit_ADDER_0.A0.n2 MULT_0.4bit_ADDER_0.A0.t12 227.356
R24852 MULT_0.4bit_ADDER_0.A0.n0 MULT_0.4bit_ADDER_0.A0.n8 226.136
R24853 MULT_0.4bit_ADDER_0.A0.n1 MULT_0.4bit_ADDER_0.A0.t8 213.688
R24854 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_0.B MULT_0.4bit_ADDER_0.A0.n6 162.867
R24855 MULT_0.4bit_ADDER_0.A0.n3 MULT_0.4bit_ADDER_0.A0.n2 160.439
R24856 MULT_0.4bit_ADDER_0.A0.n5 MULT_0.4bit_ADDER_0.A0.t10 139.78
R24857 MULT_0.4bit_ADDER_0.A0.n5 MULT_0.4bit_ADDER_0.A0.t14 139.78
R24858 MULT_0.4bit_ADDER_0.A0.n5 MULT_0.4bit_ADDER_0.A0.t9 139.78
R24859 MULT_0.4bit_ADDER_0.A0.n5 MULT_0.4bit_ADDER_0.A0.t15 139.78
R24860 MULT_0.4bit_ADDER_0.A0.n2 MULT_0.4bit_ADDER_0.A0.n1 94.4341
R24861 MULT_0.4bit_ADDER_0.A0.n0 MULT_0.4bit_ADDER_0.A0.t0 83.8336
R24862 MULT_0.4bit_ADDER_0.A0.n6 MULT_0.4bit_ADDER_0.A0.n5 38.6833
R24863 MULT_0.4bit_ADDER_0.A0.n8 MULT_0.4bit_ADDER_0.A0.t3 30.379
R24864 MULT_0.4bit_ADDER_0.A0.n8 MULT_0.4bit_ADDER_0.A0.t2 30.379
R24865 MULT_0.4bit_ADDER_0.A0.n6 MULT_0.4bit_ADDER_0.A0.n4 28.3986
R24866 MULT_0.4bit_ADDER_0.A0.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.A 24.1898
R24867 MULT_0.4bit_ADDER_0.FULL_ADDER_3.A MULT_0.4bit_ADDER_0.A0.n7 16.8273
R24868 MULT_0.4bit_ADDER_0.A0.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_0.B 9.00496
R24869 MULT_0.4bit_ADDER_0.A0.n7 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_0.B 3.87912
R24870 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_0.B MULT_0.4bit_ADDER_0.A0.n3 0.89693
R24871 MULT_0.inv_15.Y.n3 MULT_0.inv_15.Y.t14 540.38
R24872 MULT_0.inv_15.Y.n4 MULT_0.inv_15.Y.t9 491.64
R24873 MULT_0.inv_15.Y.n4 MULT_0.inv_15.Y.t4 491.64
R24874 MULT_0.inv_15.Y.n4 MULT_0.inv_15.Y.t5 491.64
R24875 MULT_0.inv_15.Y.n4 MULT_0.inv_15.Y.t10 491.64
R24876 MULT_0.inv_15.Y.n1 MULT_0.inv_15.Y.t15 367.928
R24877 MULT_0.inv_15.Y MULT_0.inv_15.Y.t1 256.514
R24878 MULT_0.inv_15.Y.n2 MULT_0.inv_15.Y.t8 227.356
R24879 MULT_0.inv_15.Y MULT_0.inv_15.Y.n7 226.248
R24880 MULT_0.inv_15.Y.n1 MULT_0.inv_15.Y.t13 213.688
R24881 MULT_0.inv_15.Y MULT_0.inv_15.Y.n6 162.867
R24882 MULT_0.inv_15.Y.n3 MULT_0.inv_15.Y.n2 160.439
R24883 MULT_0.inv_15.Y.n5 MULT_0.inv_15.Y.t12 139.78
R24884 MULT_0.inv_15.Y.n5 MULT_0.inv_15.Y.t7 139.78
R24885 MULT_0.inv_15.Y.n5 MULT_0.inv_15.Y.t6 139.78
R24886 MULT_0.inv_15.Y.n5 MULT_0.inv_15.Y.t11 139.78
R24887 MULT_0.inv_15.Y.n2 MULT_0.inv_15.Y.n1 94.4341
R24888 MULT_0.inv_15.Y MULT_0.inv_15.Y.t0 83.8155
R24889 MULT_0.inv_15.Y.n6 MULT_0.inv_15.Y.n5 38.6833
R24890 MULT_0.inv_15.Y.n7 MULT_0.inv_15.Y.t3 30.379
R24891 MULT_0.inv_15.Y.n7 MULT_0.inv_15.Y.t2 30.379
R24892 MULT_0.inv_15.Y.n6 MULT_0.inv_15.Y.n4 28.3986
R24893 MULT_0.inv_15.Y.n0 MULT_0.inv_15.Y 9.00496
R24894 MULT_0.inv_15.Y.n0 MULT_0.inv_15.Y 3.87912
R24895 MULT_0.inv_15.Y MULT_0.inv_15.Y.n0 2.57951
R24896 MULT_0.inv_15.Y.n0 MULT_0.inv_15.Y 1.47848
R24897 MULT_0.inv_15.Y MULT_0.inv_15.Y.n3 0.89693
R24898 a_n20557_n11063.n7 a_n20557_n11063.n1 81.2978
R24899 a_n20557_n11063.n1 a_n20557_n11063.n6 81.1637
R24900 a_n20557_n11063.n1 a_n20557_n11063.n5 81.1637
R24901 a_n20557_n11063.n0 a_n20557_n11063.n4 81.1637
R24902 a_n20557_n11063.n0 a_n20557_n11063.n3 81.1637
R24903 a_n20557_n11063.n0 a_n20557_n11063.n2 80.9213
R24904 a_n20557_n11063.n6 a_n20557_n11063.t3 11.8205
R24905 a_n20557_n11063.n6 a_n20557_n11063.t0 11.8205
R24906 a_n20557_n11063.n5 a_n20557_n11063.t4 11.8205
R24907 a_n20557_n11063.n5 a_n20557_n11063.t5 11.8205
R24908 a_n20557_n11063.n4 a_n20557_n11063.t7 11.8205
R24909 a_n20557_n11063.n4 a_n20557_n11063.t6 11.8205
R24910 a_n20557_n11063.n3 a_n20557_n11063.t11 11.8205
R24911 a_n20557_n11063.n3 a_n20557_n11063.t8 11.8205
R24912 a_n20557_n11063.n2 a_n20557_n11063.t9 11.8205
R24913 a_n20557_n11063.n2 a_n20557_n11063.t10 11.8205
R24914 a_n20557_n11063.n7 a_n20557_n11063.t1 11.8205
R24915 a_n20557_n11063.t2 a_n20557_n11063.n7 11.8205
R24916 a_n20557_n11063.n1 a_n20557_n11063.n0 0.402735
R24917 mux8_0.NAND4F_7.Y.n2 mux8_0.NAND4F_7.Y.t9 1388.16
R24918 mux8_0.NAND4F_7.Y.n2 mux8_0.NAND4F_7.Y.t10 350.839
R24919 mux8_0.NAND4F_7.Y.n3 mux8_0.NAND4F_7.Y.t11 308.481
R24920 mux8_0.NAND4F_7.Y.n1 mux8_0.NAND4F_7.Y.n4 187.373
R24921 mux8_0.NAND4F_7.Y.n1 mux8_0.NAND4F_7.Y.n5 187.192
R24922 mux8_0.NAND4F_7.Y.n1 mux8_0.NAND4F_7.Y.n6 187.192
R24923 mux8_0.NAND4F_7.Y.n0 mux8_0.NAND4F_7.Y.n7 187.192
R24924 mux8_0.NAND4F_7.Y mux8_0.NAND4F_7.Y.n3 161.492
R24925 mux8_0.NAND4F_7.Y.n3 mux8_0.NAND4F_7.Y.n2 27.752
R24926 mux8_0.NAND4F_7.Y mux8_0.NAND4F_7.Y.t4 23.5642
R24927 mux8_0.NAND4F_7.Y.n4 mux8_0.NAND4F_7.Y.t1 20.1899
R24928 mux8_0.NAND4F_7.Y.n4 mux8_0.NAND4F_7.Y.t0 20.1899
R24929 mux8_0.NAND4F_7.Y.n5 mux8_0.NAND4F_7.Y.t3 20.1899
R24930 mux8_0.NAND4F_7.Y.n5 mux8_0.NAND4F_7.Y.t2 20.1899
R24931 mux8_0.NAND4F_7.Y.n6 mux8_0.NAND4F_7.Y.t7 20.1899
R24932 mux8_0.NAND4F_7.Y.n6 mux8_0.NAND4F_7.Y.t8 20.1899
R24933 mux8_0.NAND4F_7.Y.n7 mux8_0.NAND4F_7.Y.t6 20.1899
R24934 mux8_0.NAND4F_7.Y.n7 mux8_0.NAND4F_7.Y.t5 20.1899
R24935 mux8_0.NAND4F_7.Y mux8_0.NAND4F_7.Y.n0 0.472662
R24936 mux8_0.NAND4F_7.Y.n0 mux8_0.NAND4F_7.Y.n1 0.358709
R24937 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t7 485.221
R24938 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t10 367.928
R24939 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n5 227.526
R24940 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n6 227.266
R24941 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n4 227.266
R24942 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t8 224.478
R24943 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t9 213.688
R24944 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n2 84.5046
R24945 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n1 72.3005
R24946 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n3 61.0566
R24947 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t2 42.7747
R24948 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t0 30.379
R24949 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t4 30.379
R24950 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t3 30.379
R24951 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t1 30.379
R24952 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t5 30.379
R24953 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.t6 30.379
R24954 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A.n0 0.583137
R24955 a_n5918_373.t0 a_n5918_373.t1 19.8005
R24956 mux8_1.NAND4F_0.C.n6 mux8_1.NAND4F_0.C.t5 978.795
R24957 mux8_1.NAND4F_0.C.n4 mux8_1.NAND4F_0.C.t7 978.795
R24958 mux8_1.NAND4F_0.C.n11 mux8_1.NAND4F_0.C.t14 978.795
R24959 mux8_1.NAND4F_0.C.n2 mux8_1.NAND4F_0.C.t12 978.795
R24960 mux8_1.NAND4F_0.C.n5 mux8_1.NAND4F_0.C.t8 308.481
R24961 mux8_1.NAND4F_0.C.n5 mux8_1.NAND4F_0.C.t10 308.481
R24962 mux8_1.NAND4F_0.C.n3 mux8_1.NAND4F_0.C.t4 308.481
R24963 mux8_1.NAND4F_0.C.n3 mux8_1.NAND4F_0.C.t6 308.481
R24964 mux8_1.NAND4F_0.C.n10 mux8_1.NAND4F_0.C.t11 308.481
R24965 mux8_1.NAND4F_0.C.n10 mux8_1.NAND4F_0.C.t9 308.481
R24966 mux8_1.NAND4F_0.C.n1 mux8_1.NAND4F_0.C.t15 308.481
R24967 mux8_1.NAND4F_0.C.n1 mux8_1.NAND4F_0.C.t13 308.481
R24968 mux8_1.NAND4F_0.C.n0 mux8_1.NAND4F_0.C.t1 256.514
R24969 mux8_1.NAND4F_0.C.n0 mux8_1.NAND4F_0.C.n8 226.258
R24970 mux8_1.NAND4F_0.C mux8_1.NAND4F_0.C.n6 161.856
R24971 mux8_1.NAND4F_0.C mux8_1.NAND4F_0.C.n4 161.847
R24972 mux8_1.NAND4F_0.C mux8_1.NAND4F_0.C.n11 161.84
R24973 mux8_1.NAND4F_0.C mux8_1.NAND4F_0.C.n2 161.831
R24974 mux8_1.NAND4F_0.C.n0 mux8_1.NAND4F_0.C.t0 83.7172
R24975 mux8_1.NAND4F_0.C.n8 mux8_1.NAND4F_0.C.t3 30.379
R24976 mux8_1.NAND4F_0.C.n8 mux8_1.NAND4F_0.C.t2 30.379
R24977 mux8_1.NAND4F_0.C.n9 mux8_1.NAND4F_0.C.n0 13.5186
R24978 mux8_1.NAND4F_0.C mux8_1.NAND4F_0.C.n12 13.0862
R24979 mux8_1.NAND4F_0.C.n7 mux8_1.NAND4F_0.C 13.0435
R24980 mux8_1.NAND4F_0.C.n12 mux8_1.NAND4F_0.C 12.4135
R24981 mux8_1.NAND4F_0.C.n7 mux8_1.NAND4F_0.C 12.4105
R24982 mux8_1.NAND4F_0.C.n6 mux8_1.NAND4F_0.C.n5 11.0463
R24983 mux8_1.NAND4F_0.C.n4 mux8_1.NAND4F_0.C.n3 11.0463
R24984 mux8_1.NAND4F_0.C.n11 mux8_1.NAND4F_0.C.n10 11.0463
R24985 mux8_1.NAND4F_0.C.n2 mux8_1.NAND4F_0.C.n1 11.0463
R24986 mux8_1.NAND4F_0.C.n12 mux8_1.NAND4F_0.C.n9 3.46056
R24987 mux8_1.NAND4F_0.C.n9 mux8_1.NAND4F_0.C.n7 1.8134
R24988 mux8_1.NAND4F_0.Y.n1 mux8_1.NAND4F_0.Y.t10 1388.16
R24989 mux8_1.NAND4F_0.Y.n1 mux8_1.NAND4F_0.Y.t9 350.839
R24990 mux8_1.NAND4F_0.Y.n2 mux8_1.NAND4F_0.Y.t11 308.481
R24991 mux8_1.NAND4F_0.Y.n0 mux8_1.NAND4F_0.Y.n3 187.373
R24992 mux8_1.NAND4F_0.Y.n0 mux8_1.NAND4F_0.Y.n4 187.192
R24993 mux8_1.NAND4F_0.Y.n0 mux8_1.NAND4F_0.Y.n5 187.192
R24994 mux8_1.NAND4F_0.Y mux8_1.NAND4F_0.Y.n6 187.192
R24995 mux8_1.NAND4F_0.Y mux8_1.NAND4F_0.Y.n2 161.492
R24996 mux8_1.NAND4F_0.Y.n2 mux8_1.NAND4F_0.Y.n1 27.752
R24997 mux8_1.NAND4F_0.Y mux8_1.NAND4F_0.Y.t2 23.5085
R24998 mux8_1.NAND4F_0.Y.n3 mux8_1.NAND4F_0.Y.t5 20.1899
R24999 mux8_1.NAND4F_0.Y.n3 mux8_1.NAND4F_0.Y.t6 20.1899
R25000 mux8_1.NAND4F_0.Y.n4 mux8_1.NAND4F_0.Y.t3 20.1899
R25001 mux8_1.NAND4F_0.Y.n4 mux8_1.NAND4F_0.Y.t4 20.1899
R25002 mux8_1.NAND4F_0.Y.n5 mux8_1.NAND4F_0.Y.t7 20.1899
R25003 mux8_1.NAND4F_0.Y.n5 mux8_1.NAND4F_0.Y.t8 20.1899
R25004 mux8_1.NAND4F_0.Y.n6 mux8_1.NAND4F_0.Y.t1 20.1899
R25005 mux8_1.NAND4F_0.Y.n6 mux8_1.NAND4F_0.Y.t0 20.1899
R25006 mux8_1.NAND4F_0.Y mux8_1.NAND4F_0.Y.n0 0.358709
R25007 right_shifter_0.buffer_7.inv_1.A.n0 right_shifter_0.buffer_7.inv_1.A.t4 393.921
R25008 right_shifter_0.buffer_7.inv_1.A.n2 right_shifter_0.buffer_7.inv_1.A.t7 291.829
R25009 right_shifter_0.buffer_7.inv_1.A.n2 right_shifter_0.buffer_7.inv_1.A.t6 291.829
R25010 right_shifter_0.buffer_7.inv_1.A.n0 right_shifter_0.buffer_7.inv_1.A.t1 256.514
R25011 right_shifter_0.buffer_7.inv_1.A.n0 right_shifter_0.buffer_7.inv_1.A.n1 226.162
R25012 right_shifter_0.buffer_7.inv_1.A.n2 right_shifter_0.buffer_7.inv_1.A.t5 221.72
R25013 right_shifter_0.buffer_7.inv_1.A.n0 right_shifter_0.buffer_7.inv_1.A.t0 83.795
R25014 right_shifter_0.buffer_7.inv_1.A.n0 right_shifter_0.buffer_7.inv_1.A.n2 53.7938
R25015 right_shifter_0.buffer_7.inv_1.A.n1 right_shifter_0.buffer_7.inv_1.A.t3 30.379
R25016 right_shifter_0.buffer_7.inv_1.A.n1 right_shifter_0.buffer_7.inv_1.A.t2 30.379
R25017 a_11386_762.t0 a_11386_762.t1 9.9005
R25018 OR8_0.NOT8_0.A4.n3 OR8_0.NOT8_0.A4.t7 394.37
R25019 OR8_0.NOT8_0.A4.n2 OR8_0.NOT8_0.A4.t10 291.829
R25020 OR8_0.NOT8_0.A4.n2 OR8_0.NOT8_0.A4.t8 291.829
R25021 OR8_0.NOT8_0.A4.n1 OR8_0.NOT8_0.A4.t3 256.425
R25022 OR8_0.NOT8_0.A4.n1 OR8_0.NOT8_0.A4.n5 231.24
R25023 OR8_0.NOT8_0.A4.n1 OR8_0.NOT8_0.A4.n6 231.03
R25024 OR8_0.NOT8_0.A4.n2 OR8_0.NOT8_0.A4.t9 221.72
R25025 OR8_0.NOT8_0.A4.n0 OR8_0.NOT8_0.A4.n4 66.4895
R25026 OR8_0.NOT8_0.A4.n3 OR8_0.NOT8_0.A4.n2 53.374
R25027 OR8_0.NOT8_0.A4.n6 OR8_0.NOT8_0.A4.t2 25.395
R25028 OR8_0.NOT8_0.A4.n6 OR8_0.NOT8_0.A4.t1 25.395
R25029 OR8_0.NOT8_0.A4.n5 OR8_0.NOT8_0.A4.t0 25.395
R25030 OR8_0.NOT8_0.A4.n5 OR8_0.NOT8_0.A4.t4 25.395
R25031 OR8_0.NOT8_0.A4.n4 OR8_0.NOT8_0.A4.t5 19.8005
R25032 OR8_0.NOT8_0.A4.n4 OR8_0.NOT8_0.A4.t6 19.8005
R25033 OR8_0.NOT8_0.A4.n0 OR8_0.NOT8_0.A4 12.5431
R25034 OR8_0.NOT8_0.A4 OR8_0.NOT8_0.A4.n3 1.25033
R25035 OR8_0.NOT8_0.A4.n1 OR8_0.NOT8_0.A4.n0 0.566868
R25036 OR8_0.S4.n1 OR8_0.S4.t6 1032.02
R25037 OR8_0.S4.n1 OR8_0.S4.t4 336.962
R25038 OR8_0.S4.n1 OR8_0.S4.t5 326.154
R25039 OR8_0.S4.n0 OR8_0.S4.t1 256.514
R25040 OR8_0.S4.n0 OR8_0.S4.n2 226.258
R25041 mux8_5.NAND4F_2.A OR8_0.S4.n1 162.952
R25042 OR8_0.S4.n0 OR8_0.S4.t0 83.7172
R25043 OR8_0.NOT8_0.S4 mux8_5.A3 63.8509
R25044 OR8_0.S4.n2 OR8_0.S4.t2 30.379
R25045 OR8_0.S4.n2 OR8_0.S4.t3 30.379
R25046 mux8_5.A3 mux8_5.NAND4F_2.A 14.0763
R25047 OR8_0.NOT8_0.S4 OR8_0.S4.n0 1.9182
R25048 a_n15887_n11683.n0 a_n15887_n11683.t3 539.788
R25049 a_n15887_n11683.n1 a_n15887_n11683.t5 531.496
R25050 a_n15887_n11683.n0 a_n15887_n11683.t2 490.034
R25051 a_n15887_n11683.n5 a_n15887_n11683.t0 283.788
R25052 a_n15887_n11683.t1 a_n15887_n11683.n5 205.489
R25053 a_n15887_n11683.n2 a_n15887_n11683.t7 182.625
R25054 a_n15887_n11683.n3 a_n15887_n11683.t4 179.054
R25055 a_n15887_n11683.n2 a_n15887_n11683.t6 139.78
R25056 a_n15887_n11683.n4 a_n15887_n11683.n3 101.368
R25057 a_n15887_n11683.n5 a_n15887_n11683.n4 77.9135
R25058 a_n15887_n11683.n4 a_n15887_n11683.n1 76.1557
R25059 a_n15887_n11683.n1 a_n15887_n11683.n0 8.29297
R25060 a_n15887_n11683.n3 a_n15887_n11683.n2 3.57087
R25061 mux8_7.A1.n0 mux8_7.A1.t13 1032.02
R25062 mux8_7.A1.n0 mux8_7.A1.t14 336.962
R25063 mux8_7.A1.n0 mux8_7.A1.t12 326.154
R25064 mux8_7.A1 mux8_7.A1.n0 162.952
R25065 mux8_7.A1.n3 mux8_7.A1.n2 120.999
R25066 mux8_7.A1.n3 mux8_7.A1.n1 120.999
R25067 mux8_7.A1.n15 mux8_7.A1.n14 104.489
R25068 mux8_7.A1.n5 mux8_7.A1.n4 92.5005
R25069 mux8_7.A1.n12 mux8_7.A1.n10 86.2638
R25070 mux8_7.A1.n10 mux8_7.A1.n9 85.8873
R25071 mux8_7.A1.n10 mux8_7.A1.n7 85.724
R25072 mux8_7.A1 mux8_7.A1.n15 83.8907
R25073 mux8_7.A1.n13 mux8_7.A1.n9 75.0672
R25074 mux8_7.A1.n13 mux8_7.A1.n12 75.0672
R25075 mux8_7.A1.n7 mux8_7.A1.n6 73.1255
R25076 mux8_7.A1.n9 mux8_7.A1.n8 73.1255
R25077 mux8_7.A1.n12 mux8_7.A1.n11 73.1255
R25078 mux8_7.A1.n14 mux8_7.A1.n7 68.8946
R25079 mux8_7.A1.n15 mux8_7.A1.n5 41.9827
R25080 mux8_7.A1.n4 mux8_7.A1.t8 30.462
R25081 mux8_7.A1.n4 mux8_7.A1.t0 30.462
R25082 mux8_7.A1.n2 mux8_7.A1.t2 30.462
R25083 mux8_7.A1.n2 mux8_7.A1.t1 30.462
R25084 mux8_7.A1.n1 mux8_7.A1.t6 30.462
R25085 mux8_7.A1.n1 mux8_7.A1.t7 30.462
R25086 mux8_7.A1.n5 mux8_7.A1.n3 28.124
R25087 mux8_7.A1.n8 mux8_7.A1.t11 11.8205
R25088 mux8_7.A1.n8 mux8_7.A1.t10 11.8205
R25089 mux8_7.A1.n6 mux8_7.A1.t9 11.8205
R25090 mux8_7.A1.n6 mux8_7.A1.t4 11.8205
R25091 mux8_7.A1.n11 mux8_7.A1.t5 11.8205
R25092 mux8_7.A1.n11 mux8_7.A1.t3 11.8205
R25093 mux8_7.A1.n14 mux8_7.A1.n13 9.3005
R25094 mux8_6.NAND4F_2.D.n4 mux8_6.NAND4F_2.D.t15 1388.16
R25095 mux8_6.NAND4F_2.D.n7 mux8_6.NAND4F_2.D.t8 1388.16
R25096 mux8_6.NAND4F_2.D.n10 mux8_6.NAND4F_2.D.t12 1388.16
R25097 mux8_6.NAND4F_2.D.n1 mux8_6.NAND4F_2.D.t5 1388.16
R25098 mux8_6.NAND4F_2.D.n4 mux8_6.NAND4F_2.D.t6 350.839
R25099 mux8_6.NAND4F_2.D.n7 mux8_6.NAND4F_2.D.t9 350.839
R25100 mux8_6.NAND4F_2.D.n10 mux8_6.NAND4F_2.D.t4 350.839
R25101 mux8_6.NAND4F_2.D.n1 mux8_6.NAND4F_2.D.t13 350.839
R25102 mux8_6.NAND4F_2.D.n5 mux8_6.NAND4F_2.D.t11 308.481
R25103 mux8_6.NAND4F_2.D.n8 mux8_6.NAND4F_2.D.t10 308.481
R25104 mux8_6.NAND4F_2.D.n11 mux8_6.NAND4F_2.D.t7 308.481
R25105 mux8_6.NAND4F_2.D.n2 mux8_6.NAND4F_2.D.t14 308.481
R25106 mux8_6.NAND4F_2.D.n0 mux8_6.NAND4F_2.D.t1 256.514
R25107 mux8_6.NAND4F_2.D.n0 mux8_6.NAND4F_2.D.n3 226.258
R25108 mux8_6.NAND4F_2.D mux8_6.NAND4F_2.D.n5 161.458
R25109 mux8_6.NAND4F_2.D mux8_6.NAND4F_2.D.n11 161.435
R25110 mux8_6.NAND4F_2.D mux8_6.NAND4F_2.D.n2 161.435
R25111 mux8_6.NAND4F_2.D mux8_6.NAND4F_2.D.n8 161.429
R25112 mux8_6.NAND4F_2.D.n0 mux8_6.NAND4F_2.D.t0 83.7172
R25113 mux8_6.NAND4F_2.D.n3 mux8_6.NAND4F_2.D.t3 30.379
R25114 mux8_6.NAND4F_2.D.n3 mux8_6.NAND4F_2.D.t2 30.379
R25115 mux8_6.NAND4F_2.D.n5 mux8_6.NAND4F_2.D.n4 27.752
R25116 mux8_6.NAND4F_2.D.n8 mux8_6.NAND4F_2.D.n7 27.752
R25117 mux8_6.NAND4F_2.D.n11 mux8_6.NAND4F_2.D.n10 27.752
R25118 mux8_6.NAND4F_2.D.n2 mux8_6.NAND4F_2.D.n1 27.752
R25119 mux8_6.NAND4F_2.D.n6 mux8_6.NAND4F_2.D.n0 12.759
R25120 mux8_6.NAND4F_2.D mux8_6.NAND4F_2.D.n12 10.6871
R25121 mux8_6.NAND4F_2.D.n6 mux8_6.NAND4F_2.D 9.0005
R25122 mux8_6.NAND4F_2.D.n12 mux8_6.NAND4F_2.D 9.0005
R25123 mux8_6.NAND4F_2.D.n9 mux8_6.NAND4F_2.D 9.0005
R25124 mux8_6.NAND4F_2.D.n9 mux8_6.NAND4F_2.D.n6 1.74507
R25125 mux8_6.NAND4F_2.D.n12 mux8_6.NAND4F_2.D.n9 1.69072
R25126 a_n11723_n12716.t0 a_n11723_n12716.t1 19.8005
R25127 a_n12347_n33735.n2 a_n12347_n33735.t7 541.395
R25128 a_n12347_n33735.n3 a_n12347_n33735.t4 527.402
R25129 a_n12347_n33735.n2 a_n12347_n33735.t5 491.64
R25130 a_n12347_n33735.n5 a_n12347_n33735.t0 281.906
R25131 a_n12347_n33735.t1 a_n12347_n33735.n5 204.359
R25132 a_n12347_n33735.n0 a_n12347_n33735.t2 180.73
R25133 a_n12347_n33735.n1 a_n12347_n33735.t6 179.45
R25134 a_n12347_n33735.n0 a_n12347_n33735.t3 139.78
R25135 a_n12347_n33735.n4 a_n12347_n33735.n1 105.635
R25136 a_n12347_n33735.n4 a_n12347_n33735.n3 76.0005
R25137 a_n12347_n33735.n5 a_n12347_n33735.n4 67.9685
R25138 a_n12347_n33735.n3 a_n12347_n33735.n2 13.994
R25139 a_n12347_n33735.n1 a_n12347_n33735.n0 1.28015
R25140 a_n19178_n11683.n0 a_n19178_n11683.t6 539.788
R25141 a_n19178_n11683.n1 a_n19178_n11683.t2 531.496
R25142 a_n19178_n11683.n0 a_n19178_n11683.t5 490.034
R25143 a_n19178_n11683.n5 a_n19178_n11683.t0 283.788
R25144 a_n19178_n11683.t1 a_n19178_n11683.n5 205.489
R25145 a_n19178_n11683.n2 a_n19178_n11683.t4 182.625
R25146 a_n19178_n11683.n3 a_n19178_n11683.t7 179.054
R25147 a_n19178_n11683.n2 a_n19178_n11683.t3 139.78
R25148 a_n19178_n11683.n4 a_n19178_n11683.n3 101.368
R25149 a_n19178_n11683.n5 a_n19178_n11683.n4 77.9135
R25150 a_n19178_n11683.n4 a_n19178_n11683.n1 76.1557
R25151 a_n19178_n11683.n1 a_n19178_n11683.n0 8.29297
R25152 a_n19178_n11683.n3 a_n19178_n11683.n2 3.57087
R25153 a_7452_n21878.t0 a_7452_n21878.t1 9.9005
R25154 OR8_0.NOT8_0.A1.n3 OR8_0.NOT8_0.A1.t10 394.37
R25155 OR8_0.NOT8_0.A1.n2 OR8_0.NOT8_0.A1.t9 291.829
R25156 OR8_0.NOT8_0.A1.n2 OR8_0.NOT8_0.A1.t7 291.829
R25157 OR8_0.NOT8_0.A1.n0 OR8_0.NOT8_0.A1.t2 256.425
R25158 OR8_0.NOT8_0.A1.n0 OR8_0.NOT8_0.A1.n4 231.24
R25159 OR8_0.NOT8_0.A1.n0 OR8_0.NOT8_0.A1.n5 231.03
R25160 OR8_0.NOT8_0.A1.n2 OR8_0.NOT8_0.A1.t8 221.72
R25161 OR8_0.NOT8_0.A1.n0 OR8_0.NOT8_0.A1.n1 66.4724
R25162 OR8_0.NOT8_0.A1.n3 OR8_0.NOT8_0.A1.n2 53.374
R25163 OR8_0.NOT8_0.A1.n0 OR8_0.NOT8_0.A1 37.2016
R25164 OR8_0.NOT8_0.A1.n4 OR8_0.NOT8_0.A1.t4 25.395
R25165 OR8_0.NOT8_0.A1.n4 OR8_0.NOT8_0.A1.t3 25.395
R25166 OR8_0.NOT8_0.A1.n5 OR8_0.NOT8_0.A1.t1 25.395
R25167 OR8_0.NOT8_0.A1.n5 OR8_0.NOT8_0.A1.t5 25.395
R25168 OR8_0.NOT8_0.A1.n1 OR8_0.NOT8_0.A1.t6 19.8005
R25169 OR8_0.NOT8_0.A1.n1 OR8_0.NOT8_0.A1.t0 19.8005
R25170 OR8_0.NOT8_0.A1 OR8_0.NOT8_0.A1.n3 1.28475
R25171 a_9432_1690.t0 a_9432_1690.t1 9.9005
R25172 a_9528_1690.t0 a_9528_1690.t1 9.9005
R25173 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t22 491.64
R25174 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t12 491.64
R25175 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t13 491.64
R25176 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t20 491.64
R25177 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n8 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t15 485.221
R25178 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t18 367.928
R25179 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t16 255.588
R25180 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t23 224.478
R25181 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t21 213.688
R25182 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n0 209.19
R25183 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t17 139.78
R25184 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t14 139.78
R25185 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t19 139.78
R25186 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n11 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n10 120.999
R25187 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n11 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n9 120.999
R25188 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n23 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n22 104.489
R25189 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n13 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n12 92.5005
R25190 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n20 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n18 86.2638
R25191 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n18 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n17 85.8873
R25192 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n18 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n15 85.724
R25193 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n8 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n7 84.5046
R25194 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n23 83.8907
R25195 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n21 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n20 75.0672
R25196 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n21 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n17 75.0672
R25197 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n20 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n19 73.1255
R25198 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n17 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n16 73.1255
R25199 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n15 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n14 73.1255
R25200 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n7 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n6 72.3005
R25201 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n22 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n15 68.8946
R25202 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n8 60.9797
R25203 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n23 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n13 41.9827
R25204 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n12 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t3 30.462
R25205 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n12 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t11 30.462
R25206 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n10 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t0 30.462
R25207 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n10 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t8 30.462
R25208 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n9 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t2 30.462
R25209 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n9 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t4 30.462
R25210 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n13 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n11 28.124
R25211 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n5 19.963
R25212 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n1 17.8661
R25213 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n2 17.8661
R25214 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n3 17.1217
R25215 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n16 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t5 11.8205
R25216 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n16 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t6 11.8205
R25217 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n19 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t9 11.8205
R25218 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n19 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t10 11.8205
R25219 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n14 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t7 11.8205
R25220 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n14 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t1 11.8205
R25221 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n22 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n21 9.3005
R25222 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n4 1.8615
R25223 a_n9125_n7799.n7 a_n9125_n7799.n1 81.2978
R25224 a_n9125_n7799.n1 a_n9125_n7799.n6 81.1637
R25225 a_n9125_n7799.n1 a_n9125_n7799.n5 81.1637
R25226 a_n9125_n7799.n0 a_n9125_n7799.n4 81.1637
R25227 a_n9125_n7799.n0 a_n9125_n7799.n3 81.1637
R25228 a_n9125_n7799.n0 a_n9125_n7799.n2 80.9213
R25229 a_n9125_n7799.n6 a_n9125_n7799.t2 11.8205
R25230 a_n9125_n7799.n6 a_n9125_n7799.t3 11.8205
R25231 a_n9125_n7799.n5 a_n9125_n7799.t0 11.8205
R25232 a_n9125_n7799.n5 a_n9125_n7799.t1 11.8205
R25233 a_n9125_n7799.n4 a_n9125_n7799.t8 11.8205
R25234 a_n9125_n7799.n4 a_n9125_n7799.t6 11.8205
R25235 a_n9125_n7799.n3 a_n9125_n7799.t9 11.8205
R25236 a_n9125_n7799.n3 a_n9125_n7799.t7 11.8205
R25237 a_n9125_n7799.n2 a_n9125_n7799.t11 11.8205
R25238 a_n9125_n7799.n2 a_n9125_n7799.t10 11.8205
R25239 a_n9125_n7799.t5 a_n9125_n7799.n7 11.8205
R25240 a_n9125_n7799.n7 a_n9125_n7799.t4 11.8205
R25241 a_n9125_n7799.n1 a_n9125_n7799.n0 0.402735
R25242 a_n11640_1406.n0 a_n11640_1406.t2 539.788
R25243 a_n11640_1406.n1 a_n11640_1406.t5 531.496
R25244 a_n11640_1406.n0 a_n11640_1406.t7 490.034
R25245 a_n11640_1406.n5 a_n11640_1406.t0 283.788
R25246 a_n11640_1406.t1 a_n11640_1406.n5 205.489
R25247 a_n11640_1406.n2 a_n11640_1406.t6 182.625
R25248 a_n11640_1406.n3 a_n11640_1406.t3 179.054
R25249 a_n11640_1406.n2 a_n11640_1406.t4 139.78
R25250 a_n11640_1406.n4 a_n11640_1406.n3 101.368
R25251 a_n11640_1406.n5 a_n11640_1406.n4 77.9135
R25252 a_n11640_1406.n4 a_n11640_1406.n1 76.1557
R25253 a_n11640_1406.n1 a_n11640_1406.n0 8.29297
R25254 a_n11640_1406.n3 a_n11640_1406.n2 3.57087
R25255 a_n11460_2026.n0 a_n11460_2026.n4 81.2978
R25256 a_n11460_2026.n0 a_n11460_2026.n5 81.1637
R25257 a_n11460_2026.n0 a_n11460_2026.n6 81.1637
R25258 a_n11460_2026.n1 a_n11460_2026.n3 81.1637
R25259 a_n11460_2026.n7 a_n11460_2026.n1 81.1637
R25260 a_n11460_2026.n1 a_n11460_2026.n2 80.9213
R25261 a_n11460_2026.n4 a_n11460_2026.t8 11.8205
R25262 a_n11460_2026.n4 a_n11460_2026.t6 11.8205
R25263 a_n11460_2026.n5 a_n11460_2026.t10 11.8205
R25264 a_n11460_2026.n5 a_n11460_2026.t7 11.8205
R25265 a_n11460_2026.n6 a_n11460_2026.t11 11.8205
R25266 a_n11460_2026.n6 a_n11460_2026.t9 11.8205
R25267 a_n11460_2026.n3 a_n11460_2026.t5 11.8205
R25268 a_n11460_2026.n3 a_n11460_2026.t0 11.8205
R25269 a_n11460_2026.n2 a_n11460_2026.t3 11.8205
R25270 a_n11460_2026.n2 a_n11460_2026.t4 11.8205
R25271 a_n11460_2026.n7 a_n11460_2026.t1 11.8205
R25272 a_n11460_2026.t2 a_n11460_2026.n7 11.8205
R25273 a_n11460_2026.n1 a_n11460_2026.n0 0.402735
R25274 a_n16513_1380.n2 a_n16513_1380.t4 541.395
R25275 a_n16513_1380.n3 a_n16513_1380.t2 527.402
R25276 a_n16513_1380.n2 a_n16513_1380.t7 491.64
R25277 a_n16513_1380.n5 a_n16513_1380.t0 281.906
R25278 a_n16513_1380.t1 a_n16513_1380.n5 204.359
R25279 a_n16513_1380.n0 a_n16513_1380.t3 180.73
R25280 a_n16513_1380.n1 a_n16513_1380.t5 179.45
R25281 a_n16513_1380.n0 a_n16513_1380.t6 139.78
R25282 a_n16513_1380.n4 a_n16513_1380.n1 105.635
R25283 a_n16513_1380.n4 a_n16513_1380.n3 76.0005
R25284 a_n16513_1380.n5 a_n16513_1380.n4 67.9685
R25285 a_n16513_1380.n3 a_n16513_1380.n2 13.994
R25286 a_n16513_1380.n1 a_n16513_1380.n0 1.28015
R25287 Y5.n0 Y5.t4 883.668
R25288 Y5.n1 Y5.t6 740.381
R25289 Y5.n0 Y5.t7 729.428
R25290 Y5.n2 Y5.t5 700.508
R25291 Y5.n4 Y5.t1 256.514
R25292 Y5 Y5.n3 226.236
R25293 Y5 Y5.n2 162.625
R25294 Y5.n5 Y5.t0 83.7901
R25295 Y5.n1 Y5.n0 72.3005
R25296 Y5.n3 Y5.t3 30.379
R25297 Y5.n3 Y5.t2 30.379
R25298 Y5.n2 Y5.n1 16.7975
R25299 Y5.n5 Y5 0.0349228
R25300 Y5 Y5.n5 0.0300905
R25301 Y5.n4 Y5 0.0276164
R25302 Y5 Y5.n4 0.0229868
R25303 a_15855_n19505.n2 a_15855_n19505.n1 140.274
R25304 a_15855_n19505.n2 a_15855_n19505.n0 140.274
R25305 a_15855_n19505.n3 a_15855_n19505.n2 140.21
R25306 a_15855_n19505.n1 a_15855_n19505.t5 7.59513
R25307 a_15855_n19505.n1 a_15855_n19505.t3 7.59513
R25308 a_15855_n19505.n0 a_15855_n19505.t1 7.59513
R25309 a_15855_n19505.n0 a_15855_n19505.t0 7.59513
R25310 a_15855_n19505.n3 a_15855_n19505.t2 7.59513
R25311 a_15855_n19505.t4 a_15855_n19505.n3 7.59513
R25312 a_16143_n19505.n2 a_16143_n19505.n0 140.65
R25313 a_16143_n19505.n3 a_16143_n19505.n2 140.65
R25314 a_16143_n19505.n2 a_16143_n19505.n1 140.587
R25315 a_16143_n19505.n1 a_16143_n19505.t3 7.59513
R25316 a_16143_n19505.n1 a_16143_n19505.t1 7.59513
R25317 a_16143_n19505.n0 a_16143_n19505.t5 7.59513
R25318 a_16143_n19505.n0 a_16143_n19505.t4 7.59513
R25319 a_16143_n19505.n3 a_16143_n19505.t0 7.59513
R25320 a_16143_n19505.t2 a_16143_n19505.n3 7.59513
R25321 a_n19954_1406.n0 a_n19954_1406.t5 539.788
R25322 a_n19954_1406.n1 a_n19954_1406.t7 531.496
R25323 a_n19954_1406.n0 a_n19954_1406.t2 490.034
R25324 a_n19954_1406.n5 a_n19954_1406.t0 283.788
R25325 a_n19954_1406.t1 a_n19954_1406.n5 205.489
R25326 a_n19954_1406.n2 a_n19954_1406.t3 182.625
R25327 a_n19954_1406.n3 a_n19954_1406.t4 179.054
R25328 a_n19954_1406.n2 a_n19954_1406.t6 139.78
R25329 a_n19954_1406.n4 a_n19954_1406.n3 101.368
R25330 a_n19954_1406.n5 a_n19954_1406.n4 77.9135
R25331 a_n19954_1406.n4 a_n19954_1406.n1 76.1557
R25332 a_n19954_1406.n1 a_n19954_1406.n0 8.29297
R25333 a_n19954_1406.n3 a_n19954_1406.n2 3.57087
R25334 mux8_8.A0.n0 mux8_8.A0.t13 1032.02
R25335 mux8_8.A0.n0 mux8_8.A0.t14 336.962
R25336 mux8_8.A0.n0 mux8_8.A0.t12 326.154
R25337 mux8_8.A0 mux8_8.A0.n0 162.952
R25338 mux8_8.A0.n3 mux8_8.A0.n2 120.999
R25339 mux8_8.A0.n3 mux8_8.A0.n1 120.999
R25340 mux8_8.A0.n15 mux8_8.A0.n14 104.489
R25341 mux8_8.A0.n5 mux8_8.A0.n4 92.5005
R25342 mux8_8.A0.n12 mux8_8.A0.n10 86.2638
R25343 mux8_8.A0.n10 mux8_8.A0.n9 85.8873
R25344 mux8_8.A0.n10 mux8_8.A0.n7 85.724
R25345 mux8_8.A0 mux8_8.A0.n15 83.8907
R25346 mux8_8.A0.n13 mux8_8.A0.n9 75.0672
R25347 mux8_8.A0.n13 mux8_8.A0.n12 75.0672
R25348 mux8_8.A0.n7 mux8_8.A0.n6 73.1255
R25349 mux8_8.A0.n9 mux8_8.A0.n8 73.1255
R25350 mux8_8.A0.n12 mux8_8.A0.n11 73.1255
R25351 mux8_8.A0.n14 mux8_8.A0.n7 68.8946
R25352 mux8_8.A0.n15 mux8_8.A0.n5 41.9827
R25353 mux8_8.A0.n4 mux8_8.A0.t4 30.462
R25354 mux8_8.A0.n4 mux8_8.A0.t6 30.462
R25355 mux8_8.A0.n2 mux8_8.A0.t10 30.462
R25356 mux8_8.A0.n2 mux8_8.A0.t11 30.462
R25357 mux8_8.A0.n1 mux8_8.A0.t0 30.462
R25358 mux8_8.A0.n1 mux8_8.A0.t5 30.462
R25359 mux8_8.A0.n5 mux8_8.A0.n3 28.124
R25360 mux8_8.A0.n8 mux8_8.A0.t2 11.8205
R25361 mux8_8.A0.n8 mux8_8.A0.t1 11.8205
R25362 mux8_8.A0.n6 mux8_8.A0.t3 11.8205
R25363 mux8_8.A0.n6 mux8_8.A0.t8 11.8205
R25364 mux8_8.A0.n11 mux8_8.A0.t9 11.8205
R25365 mux8_8.A0.n11 mux8_8.A0.t7 11.8205
R25366 mux8_8.A0.n14 mux8_8.A0.n13 9.3005
R25367 a_n3500_1406.n0 a_n3500_1406.t3 539.788
R25368 a_n3500_1406.n1 a_n3500_1406.t2 531.496
R25369 a_n3500_1406.n0 a_n3500_1406.t7 490.034
R25370 a_n3500_1406.n5 a_n3500_1406.t0 283.788
R25371 a_n3500_1406.t1 a_n3500_1406.n5 205.489
R25372 a_n3500_1406.n2 a_n3500_1406.t6 182.625
R25373 a_n3500_1406.n3 a_n3500_1406.t5 179.054
R25374 a_n3500_1406.n2 a_n3500_1406.t4 139.78
R25375 a_n3500_1406.n4 a_n3500_1406.n3 101.368
R25376 a_n3500_1406.n5 a_n3500_1406.n4 77.9135
R25377 a_n3500_1406.n4 a_n3500_1406.n1 76.1557
R25378 a_n3500_1406.n1 a_n3500_1406.n0 8.29297
R25379 a_n3500_1406.n3 a_n3500_1406.n2 3.57087
R25380 a_n3320_2026.n7 a_n3320_2026.n1 81.2978
R25381 a_n3320_2026.n1 a_n3320_2026.n6 81.1637
R25382 a_n3320_2026.n1 a_n3320_2026.n5 81.1637
R25383 a_n3320_2026.n0 a_n3320_2026.n4 81.1637
R25384 a_n3320_2026.n0 a_n3320_2026.n3 81.1637
R25385 a_n3320_2026.n0 a_n3320_2026.n2 80.9213
R25386 a_n3320_2026.n6 a_n3320_2026.t11 11.8205
R25387 a_n3320_2026.n6 a_n3320_2026.t1 11.8205
R25388 a_n3320_2026.n5 a_n3320_2026.t10 11.8205
R25389 a_n3320_2026.n5 a_n3320_2026.t9 11.8205
R25390 a_n3320_2026.n4 a_n3320_2026.t3 11.8205
R25391 a_n3320_2026.n4 a_n3320_2026.t4 11.8205
R25392 a_n3320_2026.n3 a_n3320_2026.t7 11.8205
R25393 a_n3320_2026.n3 a_n3320_2026.t5 11.8205
R25394 a_n3320_2026.n2 a_n3320_2026.t8 11.8205
R25395 a_n3320_2026.n2 a_n3320_2026.t6 11.8205
R25396 a_n3320_2026.t2 a_n3320_2026.n7 11.8205
R25397 a_n3320_2026.n7 a_n3320_2026.t0 11.8205
R25398 a_n3320_2026.n1 a_n3320_2026.n0 0.402735
R25399 8bit_ADDER_0.S1.n0 8bit_ADDER_0.S1.t13 1032.02
R25400 8bit_ADDER_0.S1.n0 8bit_ADDER_0.S1.t12 336.962
R25401 8bit_ADDER_0.S1.n0 8bit_ADDER_0.S1.t14 326.154
R25402 mux8_2.NAND4F_3.A 8bit_ADDER_0.S1.n0 162.952
R25403 8bit_ADDER_0.S1.n3 8bit_ADDER_0.S1.n2 120.999
R25404 8bit_ADDER_0.S1.n3 8bit_ADDER_0.S1.n1 120.999
R25405 8bit_ADDER_0.S1.n15 8bit_ADDER_0.S1.n14 104.489
R25406 8bit_ADDER_0.S1.n5 8bit_ADDER_0.S1.n4 92.5005
R25407 8bit_ADDER_0.S1.n12 8bit_ADDER_0.S1.n10 86.2638
R25408 8bit_ADDER_0.S1.n10 8bit_ADDER_0.S1.n9 85.8873
R25409 8bit_ADDER_0.S1.n10 8bit_ADDER_0.S1.n7 85.724
R25410 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.Y 8bit_ADDER_0.S1.n15 83.8907
R25411 8bit_ADDER_0.S1.n13 8bit_ADDER_0.S1.n12 75.0672
R25412 8bit_ADDER_0.S1.n13 8bit_ADDER_0.S1.n9 75.0672
R25413 8bit_ADDER_0.S1.n12 8bit_ADDER_0.S1.n11 73.1255
R25414 8bit_ADDER_0.S1.n7 8bit_ADDER_0.S1.n6 73.1255
R25415 8bit_ADDER_0.S1.n9 8bit_ADDER_0.S1.n8 73.1255
R25416 8bit_ADDER_0.S1.n14 8bit_ADDER_0.S1.n7 68.8946
R25417 8bit_ADDER_0.FULL_ADDER_XORED_6.OUT mux8_2.A0 45.2041
R25418 8bit_ADDER_0.S1.n15 8bit_ADDER_0.S1.n5 41.9827
R25419 8bit_ADDER_0.S1.n4 8bit_ADDER_0.S1.t0 30.462
R25420 8bit_ADDER_0.S1.n4 8bit_ADDER_0.S1.t6 30.462
R25421 8bit_ADDER_0.S1.n2 8bit_ADDER_0.S1.t8 30.462
R25422 8bit_ADDER_0.S1.n2 8bit_ADDER_0.S1.t7 30.462
R25423 8bit_ADDER_0.S1.n1 8bit_ADDER_0.S1.t1 30.462
R25424 8bit_ADDER_0.S1.n1 8bit_ADDER_0.S1.t2 30.462
R25425 8bit_ADDER_0.S1.n5 8bit_ADDER_0.S1.n3 28.124
R25426 mux8_2.A0 mux8_2.NAND4F_3.A 15.2713
R25427 8bit_ADDER_0.S1.n6 8bit_ADDER_0.S1.t4 11.8205
R25428 8bit_ADDER_0.S1.n6 8bit_ADDER_0.S1.t10 11.8205
R25429 8bit_ADDER_0.S1.n11 8bit_ADDER_0.S1.t9 11.8205
R25430 8bit_ADDER_0.S1.n11 8bit_ADDER_0.S1.t11 11.8205
R25431 8bit_ADDER_0.S1.n8 8bit_ADDER_0.S1.t5 11.8205
R25432 8bit_ADDER_0.S1.n8 8bit_ADDER_0.S1.t3 11.8205
R25433 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.Y 8bit_ADDER_0.FULL_ADDER_XORED_6.OUT 10.6442
R25434 8bit_ADDER_0.S1.n14 8bit_ADDER_0.S1.n13 9.3005
R25435 mux8_8.NAND4F_0.C.n6 mux8_8.NAND4F_0.C.t15 978.795
R25436 mux8_8.NAND4F_0.C.n4 mux8_8.NAND4F_0.C.t9 978.795
R25437 mux8_8.NAND4F_0.C.n11 mux8_8.NAND4F_0.C.t11 978.795
R25438 mux8_8.NAND4F_0.C.n2 mux8_8.NAND4F_0.C.t13 978.795
R25439 mux8_8.NAND4F_0.C.n5 mux8_8.NAND4F_0.C.t14 308.481
R25440 mux8_8.NAND4F_0.C.n5 mux8_8.NAND4F_0.C.t12 308.481
R25441 mux8_8.NAND4F_0.C.n3 mux8_8.NAND4F_0.C.t5 308.481
R25442 mux8_8.NAND4F_0.C.n3 mux8_8.NAND4F_0.C.t4 308.481
R25443 mux8_8.NAND4F_0.C.n10 mux8_8.NAND4F_0.C.t6 308.481
R25444 mux8_8.NAND4F_0.C.n10 mux8_8.NAND4F_0.C.t7 308.481
R25445 mux8_8.NAND4F_0.C.n1 mux8_8.NAND4F_0.C.t8 308.481
R25446 mux8_8.NAND4F_0.C.n1 mux8_8.NAND4F_0.C.t10 308.481
R25447 mux8_8.NAND4F_0.C.n0 mux8_8.NAND4F_0.C.t2 256.514
R25448 mux8_8.NAND4F_0.C.n0 mux8_8.NAND4F_0.C.n8 226.258
R25449 mux8_8.NAND4F_0.C mux8_8.NAND4F_0.C.n6 161.856
R25450 mux8_8.NAND4F_0.C mux8_8.NAND4F_0.C.n4 161.847
R25451 mux8_8.NAND4F_0.C mux8_8.NAND4F_0.C.n11 161.84
R25452 mux8_8.NAND4F_0.C mux8_8.NAND4F_0.C.n2 161.831
R25453 mux8_8.NAND4F_0.C.n0 mux8_8.NAND4F_0.C.t0 83.7172
R25454 mux8_8.NAND4F_0.C.n8 mux8_8.NAND4F_0.C.t1 30.379
R25455 mux8_8.NAND4F_0.C.n8 mux8_8.NAND4F_0.C.t3 30.379
R25456 mux8_8.NAND4F_0.C.n9 mux8_8.NAND4F_0.C.n0 13.5186
R25457 mux8_8.NAND4F_0.C mux8_8.NAND4F_0.C.n12 13.0862
R25458 mux8_8.NAND4F_0.C.n7 mux8_8.NAND4F_0.C 13.0435
R25459 mux8_8.NAND4F_0.C.n12 mux8_8.NAND4F_0.C 12.4135
R25460 mux8_8.NAND4F_0.C.n7 mux8_8.NAND4F_0.C 12.4105
R25461 mux8_8.NAND4F_0.C.n6 mux8_8.NAND4F_0.C.n5 11.0463
R25462 mux8_8.NAND4F_0.C.n4 mux8_8.NAND4F_0.C.n3 11.0463
R25463 mux8_8.NAND4F_0.C.n11 mux8_8.NAND4F_0.C.n10 11.0463
R25464 mux8_8.NAND4F_0.C.n2 mux8_8.NAND4F_0.C.n1 11.0463
R25465 mux8_8.NAND4F_0.C.n12 mux8_8.NAND4F_0.C.n9 3.46056
R25466 mux8_8.NAND4F_0.C.n9 mux8_8.NAND4F_0.C.n7 1.8134
R25467 mux8_8.NAND4F_2.D.n4 mux8_8.NAND4F_2.D.t7 1388.16
R25468 mux8_8.NAND4F_2.D.n7 mux8_8.NAND4F_2.D.t12 1388.16
R25469 mux8_8.NAND4F_2.D.n10 mux8_8.NAND4F_2.D.t15 1388.16
R25470 mux8_8.NAND4F_2.D.n1 mux8_8.NAND4F_2.D.t11 1388.16
R25471 mux8_8.NAND4F_2.D.n4 mux8_8.NAND4F_2.D.t5 350.839
R25472 mux8_8.NAND4F_2.D.n7 mux8_8.NAND4F_2.D.t8 350.839
R25473 mux8_8.NAND4F_2.D.n10 mux8_8.NAND4F_2.D.t4 350.839
R25474 mux8_8.NAND4F_2.D.n1 mux8_8.NAND4F_2.D.t13 350.839
R25475 mux8_8.NAND4F_2.D.n5 mux8_8.NAND4F_2.D.t10 308.481
R25476 mux8_8.NAND4F_2.D.n8 mux8_8.NAND4F_2.D.t9 308.481
R25477 mux8_8.NAND4F_2.D.n11 mux8_8.NAND4F_2.D.t6 308.481
R25478 mux8_8.NAND4F_2.D.n2 mux8_8.NAND4F_2.D.t14 308.481
R25479 mux8_8.NAND4F_2.D.n0 mux8_8.NAND4F_2.D.t2 256.514
R25480 mux8_8.NAND4F_2.D.n0 mux8_8.NAND4F_2.D.n3 226.258
R25481 mux8_8.NAND4F_2.D mux8_8.NAND4F_2.D.n5 161.458
R25482 mux8_8.NAND4F_2.D mux8_8.NAND4F_2.D.n11 161.435
R25483 mux8_8.NAND4F_2.D mux8_8.NAND4F_2.D.n2 161.435
R25484 mux8_8.NAND4F_2.D mux8_8.NAND4F_2.D.n8 161.429
R25485 mux8_8.NAND4F_2.D.n0 mux8_8.NAND4F_2.D.t0 83.7172
R25486 mux8_8.NAND4F_2.D.n3 mux8_8.NAND4F_2.D.t1 30.379
R25487 mux8_8.NAND4F_2.D.n3 mux8_8.NAND4F_2.D.t3 30.379
R25488 mux8_8.NAND4F_2.D.n5 mux8_8.NAND4F_2.D.n4 27.752
R25489 mux8_8.NAND4F_2.D.n8 mux8_8.NAND4F_2.D.n7 27.752
R25490 mux8_8.NAND4F_2.D.n11 mux8_8.NAND4F_2.D.n10 27.752
R25491 mux8_8.NAND4F_2.D.n2 mux8_8.NAND4F_2.D.n1 27.752
R25492 mux8_8.NAND4F_2.D.n6 mux8_8.NAND4F_2.D.n0 12.759
R25493 mux8_8.NAND4F_2.D mux8_8.NAND4F_2.D.n12 10.6871
R25494 mux8_8.NAND4F_2.D.n6 mux8_8.NAND4F_2.D 9.0005
R25495 mux8_8.NAND4F_2.D.n12 mux8_8.NAND4F_2.D 9.0005
R25496 mux8_8.NAND4F_2.D.n9 mux8_8.NAND4F_2.D 9.0005
R25497 mux8_8.NAND4F_2.D.n9 mux8_8.NAND4F_2.D.n6 1.74507
R25498 mux8_8.NAND4F_2.D.n12 mux8_8.NAND4F_2.D.n9 1.69072
R25499 a_n14005_n5180.n2 a_n14005_n5180.t7 541.395
R25500 a_n14005_n5180.n3 a_n14005_n5180.t3 527.402
R25501 a_n14005_n5180.n2 a_n14005_n5180.t4 491.64
R25502 a_n14005_n5180.n5 a_n14005_n5180.t0 281.906
R25503 a_n14005_n5180.t1 a_n14005_n5180.n5 204.359
R25504 a_n14005_n5180.n0 a_n14005_n5180.t2 180.73
R25505 a_n14005_n5180.n1 a_n14005_n5180.t5 179.45
R25506 a_n14005_n5180.n0 a_n14005_n5180.t6 139.78
R25507 a_n14005_n5180.n4 a_n14005_n5180.n1 105.635
R25508 a_n14005_n5180.n4 a_n14005_n5180.n3 76.0005
R25509 a_n14005_n5180.n5 a_n14005_n5180.n4 67.9685
R25510 a_n14005_n5180.n3 a_n14005_n5180.n2 13.994
R25511 a_n14005_n5180.n1 a_n14005_n5180.n0 1.28015
R25512 a_547_1406.n2 a_547_1406.n1 121.353
R25513 a_547_1406.n2 a_547_1406.n0 121.353
R25514 a_547_1406.n3 a_547_1406.n2 121.001
R25515 a_547_1406.n1 a_547_1406.t3 30.462
R25516 a_547_1406.n1 a_547_1406.t5 30.462
R25517 a_547_1406.n0 a_547_1406.t1 30.462
R25518 a_547_1406.n0 a_547_1406.t0 30.462
R25519 a_547_1406.t2 a_547_1406.n3 30.462
R25520 a_547_1406.n3 a_547_1406.t4 30.462
R25521 mux8_3.NAND4F_0.C.n6 mux8_3.NAND4F_0.C.t8 978.795
R25522 mux8_3.NAND4F_0.C.n4 mux8_3.NAND4F_0.C.t4 978.795
R25523 mux8_3.NAND4F_0.C.n11 mux8_3.NAND4F_0.C.t15 978.795
R25524 mux8_3.NAND4F_0.C.n2 mux8_3.NAND4F_0.C.t6 978.795
R25525 mux8_3.NAND4F_0.C.n5 mux8_3.NAND4F_0.C.t12 308.481
R25526 mux8_3.NAND4F_0.C.n5 mux8_3.NAND4F_0.C.t11 308.481
R25527 mux8_3.NAND4F_0.C.n3 mux8_3.NAND4F_0.C.t7 308.481
R25528 mux8_3.NAND4F_0.C.n3 mux8_3.NAND4F_0.C.t5 308.481
R25529 mux8_3.NAND4F_0.C.n10 mux8_3.NAND4F_0.C.t13 308.481
R25530 mux8_3.NAND4F_0.C.n10 mux8_3.NAND4F_0.C.t14 308.481
R25531 mux8_3.NAND4F_0.C.n1 mux8_3.NAND4F_0.C.t9 308.481
R25532 mux8_3.NAND4F_0.C.n1 mux8_3.NAND4F_0.C.t10 308.481
R25533 mux8_3.NAND4F_0.C.n0 mux8_3.NAND4F_0.C.t1 256.514
R25534 mux8_3.NAND4F_0.C.n0 mux8_3.NAND4F_0.C.n8 226.258
R25535 mux8_3.NAND4F_0.C mux8_3.NAND4F_0.C.n6 161.856
R25536 mux8_3.NAND4F_0.C mux8_3.NAND4F_0.C.n4 161.847
R25537 mux8_3.NAND4F_0.C mux8_3.NAND4F_0.C.n11 161.84
R25538 mux8_3.NAND4F_0.C mux8_3.NAND4F_0.C.n2 161.831
R25539 mux8_3.NAND4F_0.C.n0 mux8_3.NAND4F_0.C.t0 83.7172
R25540 mux8_3.NAND4F_0.C.n8 mux8_3.NAND4F_0.C.t3 30.379
R25541 mux8_3.NAND4F_0.C.n8 mux8_3.NAND4F_0.C.t2 30.379
R25542 mux8_3.NAND4F_0.C.n9 mux8_3.NAND4F_0.C.n0 13.5186
R25543 mux8_3.NAND4F_0.C mux8_3.NAND4F_0.C.n12 13.0862
R25544 mux8_3.NAND4F_0.C.n7 mux8_3.NAND4F_0.C 13.0435
R25545 mux8_3.NAND4F_0.C.n12 mux8_3.NAND4F_0.C 12.4135
R25546 mux8_3.NAND4F_0.C.n7 mux8_3.NAND4F_0.C 12.4105
R25547 mux8_3.NAND4F_0.C.n6 mux8_3.NAND4F_0.C.n5 11.0463
R25548 mux8_3.NAND4F_0.C.n4 mux8_3.NAND4F_0.C.n3 11.0463
R25549 mux8_3.NAND4F_0.C.n11 mux8_3.NAND4F_0.C.n10 11.0463
R25550 mux8_3.NAND4F_0.C.n2 mux8_3.NAND4F_0.C.n1 11.0463
R25551 mux8_3.NAND4F_0.C.n12 mux8_3.NAND4F_0.C.n9 3.46056
R25552 mux8_3.NAND4F_0.C.n9 mux8_3.NAND4F_0.C.n7 1.8134
R25553 a_10267_n11894.t0 a_10267_n11894.t1 9.9005
R25554 a_10363_n11894.t0 a_10363_n11894.t1 9.9005
R25555 a_8400_n17350.t0 a_8400_n17350.t1 9.9005
R25556 mux8_2.NAND4F_3.Y.n7 mux8_2.NAND4F_3.Y.t11 978.795
R25557 mux8_2.NAND4F_3.Y.n6 mux8_2.NAND4F_3.Y.t9 308.481
R25558 mux8_2.NAND4F_3.Y.n6 mux8_2.NAND4F_3.Y.t10 308.481
R25559 mux8_2.NAND4F_3.Y.n0 mux8_2.NAND4F_3.Y.n1 187.373
R25560 mux8_2.NAND4F_3.Y.n0 mux8_2.NAND4F_3.Y.n2 187.192
R25561 mux8_2.NAND4F_3.Y.n0 mux8_2.NAND4F_3.Y.n3 187.192
R25562 mux8_2.NAND4F_3.Y.n5 mux8_2.NAND4F_3.Y.n4 187.192
R25563 mux8_2.NAND4F_3.Y mux8_2.NAND4F_3.Y.n7 161.839
R25564 mux8_2.NAND4F_3.Y mux8_2.NAND4F_3.Y.t4 23.4426
R25565 mux8_2.NAND4F_3.Y.n1 mux8_2.NAND4F_3.Y.t3 20.1899
R25566 mux8_2.NAND4F_3.Y.n1 mux8_2.NAND4F_3.Y.t2 20.1899
R25567 mux8_2.NAND4F_3.Y.n2 mux8_2.NAND4F_3.Y.t0 20.1899
R25568 mux8_2.NAND4F_3.Y.n2 mux8_2.NAND4F_3.Y.t1 20.1899
R25569 mux8_2.NAND4F_3.Y.n3 mux8_2.NAND4F_3.Y.t7 20.1899
R25570 mux8_2.NAND4F_3.Y.n3 mux8_2.NAND4F_3.Y.t8 20.1899
R25571 mux8_2.NAND4F_3.Y.n4 mux8_2.NAND4F_3.Y.t6 20.1899
R25572 mux8_2.NAND4F_3.Y.n4 mux8_2.NAND4F_3.Y.t5 20.1899
R25573 mux8_2.NAND4F_3.Y.n7 mux8_2.NAND4F_3.Y.n6 11.0463
R25574 mux8_2.NAND4F_3.Y mux8_2.NAND4F_3.Y.n5 0.518495
R25575 mux8_2.NAND4F_3.Y.n5 mux8_2.NAND4F_3.Y.n0 0.358709
R25576 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t17 491.64
R25577 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t13 491.64
R25578 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t23 491.64
R25579 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t19 491.64
R25580 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t16 485.221
R25581 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t18 367.928
R25582 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t14 255.588
R25583 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t20 224.478
R25584 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t21 213.688
R25585 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n0 209.19
R25586 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t22 139.78
R25587 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t12 139.78
R25588 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t15 139.78
R25589 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n10 120.999
R25590 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n11 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n9 120.999
R25591 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n22 104.489
R25592 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n12 92.5005
R25593 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n18 86.2638
R25594 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n17 85.8873
R25595 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n18 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n15 85.724
R25596 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n8 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n7 84.5046
R25597 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n23 83.8907
R25598 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n17 75.0672
R25599 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n21 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n20 75.0672
R25600 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n15 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n14 73.1255
R25601 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n17 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n16 73.1255
R25602 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n20 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n19 73.1255
R25603 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n7 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n6 72.3005
R25604 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n15 68.8946
R25605 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n8 60.9797
R25606 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n23 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n13 41.9827
R25607 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t1 30.462
R25608 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n12 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t4 30.462
R25609 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t7 30.462
R25610 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n10 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t8 30.462
R25611 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t2 30.462
R25612 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n9 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t3 30.462
R25613 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n13 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n11 28.124
R25614 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n5 19.963
R25615 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n1 17.8661
R25616 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n2 17.8661
R25617 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n3 17.1217
R25618 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t10 11.8205
R25619 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n16 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t9 11.8205
R25620 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t11 11.8205
R25621 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n14 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t6 11.8205
R25622 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t0 11.8205
R25623 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n19 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t5 11.8205
R25624 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n22 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n21 9.3005
R25625 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n4 1.8615
R25626 a_n19198_1406.n2 a_n19198_1406.n0 121.353
R25627 a_n19198_1406.n3 a_n19198_1406.n2 121.353
R25628 a_n19198_1406.n2 a_n19198_1406.n1 121.001
R25629 a_n19198_1406.n0 a_n19198_1406.t3 30.462
R25630 a_n19198_1406.n0 a_n19198_1406.t4 30.462
R25631 a_n19198_1406.n1 a_n19198_1406.t0 30.462
R25632 a_n19198_1406.n1 a_n19198_1406.t5 30.462
R25633 a_n19198_1406.n3 a_n19198_1406.t1 30.462
R25634 a_n19198_1406.t2 a_n19198_1406.n3 30.462
R25635 a_n12316_n34281.n0 a_n12316_n34281.n2 81.2978
R25636 a_n12316_n34281.n1 a_n12316_n34281.n6 81.1637
R25637 a_n12316_n34281.n1 a_n12316_n34281.n5 81.1637
R25638 a_n12316_n34281.n0 a_n12316_n34281.n4 81.1637
R25639 a_n12316_n34281.n0 a_n12316_n34281.n3 81.1637
R25640 a_n12316_n34281.n7 a_n12316_n34281.n1 80.9213
R25641 a_n12316_n34281.n6 a_n12316_n34281.t1 11.8205
R25642 a_n12316_n34281.n6 a_n12316_n34281.t11 11.8205
R25643 a_n12316_n34281.n5 a_n12316_n34281.t10 11.8205
R25644 a_n12316_n34281.n5 a_n12316_n34281.t9 11.8205
R25645 a_n12316_n34281.n4 a_n12316_n34281.t5 11.8205
R25646 a_n12316_n34281.n4 a_n12316_n34281.t4 11.8205
R25647 a_n12316_n34281.n3 a_n12316_n34281.t3 11.8205
R25648 a_n12316_n34281.n3 a_n12316_n34281.t7 11.8205
R25649 a_n12316_n34281.n2 a_n12316_n34281.t6 11.8205
R25650 a_n12316_n34281.n2 a_n12316_n34281.t8 11.8205
R25651 a_n12316_n34281.n7 a_n12316_n34281.t0 11.8205
R25652 a_n12316_n34281.t2 a_n12316_n34281.n7 11.8205
R25653 a_n12316_n34281.n1 a_n12316_n34281.n0 0.402735
R25654 a_n24048_1406.n2 a_n24048_1406.n0 121.353
R25655 a_n24048_1406.n3 a_n24048_1406.n2 121.353
R25656 a_n24048_1406.n2 a_n24048_1406.n1 121.001
R25657 a_n24048_1406.n0 a_n24048_1406.t3 30.462
R25658 a_n24048_1406.n0 a_n24048_1406.t4 30.462
R25659 a_n24048_1406.n1 a_n24048_1406.t1 30.462
R25660 a_n24048_1406.n1 a_n24048_1406.t5 30.462
R25661 a_n24048_1406.t2 a_n24048_1406.n3 30.462
R25662 a_n24048_1406.n3 a_n24048_1406.t0 30.462
R25663 MULT_0.4bit_ADDER_2.B0.n4 MULT_0.4bit_ADDER_2.B0.t18 491.64
R25664 MULT_0.4bit_ADDER_2.B0.n5 MULT_0.4bit_ADDER_2.B0.t13 491.64
R25665 MULT_0.4bit_ADDER_2.B0.n6 MULT_0.4bit_ADDER_2.B0.t12 491.64
R25666 MULT_0.4bit_ADDER_2.B0.n7 MULT_0.4bit_ADDER_2.B0.t19 491.64
R25667 MULT_0.4bit_ADDER_2.B0.n2 MULT_0.4bit_ADDER_2.B0.t23 485.221
R25668 MULT_0.4bit_ADDER_2.B0.n0 MULT_0.4bit_ADDER_2.B0.t14 367.928
R25669 MULT_0.4bit_ADDER_2.B0.n8 MULT_0.4bit_ADDER_2.B0.t17 255.588
R25670 MULT_0.4bit_ADDER_2.B0.n1 MULT_0.4bit_ADDER_2.B0.t21 224.478
R25671 MULT_0.4bit_ADDER_2.B0.n0 MULT_0.4bit_ADDER_2.B0.t22 213.688
R25672 MULT_0.4bit_ADDER_2.B0.n4 MULT_0.4bit_ADDER_2.B0.n3 209.19
R25673 MULT_0.4bit_ADDER_2.B0.n3 MULT_0.4bit_ADDER_2.B0.t15 139.78
R25674 MULT_0.4bit_ADDER_2.B0.n3 MULT_0.4bit_ADDER_2.B0.t16 139.78
R25675 MULT_0.4bit_ADDER_2.B0.n3 MULT_0.4bit_ADDER_2.B0.t20 139.78
R25676 MULT_0.4bit_ADDER_2.B0.n12 MULT_0.4bit_ADDER_2.B0.n11 120.999
R25677 MULT_0.4bit_ADDER_2.B0.n12 MULT_0.4bit_ADDER_2.B0.n10 120.999
R25678 MULT_0.4bit_ADDER_2.B0.n24 MULT_0.4bit_ADDER_2.B0.n23 104.489
R25679 MULT_0.4bit_ADDER_2.B0.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_0.A 103.258
R25680 MULT_0.4bit_ADDER_2.B0.n14 MULT_0.4bit_ADDER_2.B0.n13 92.5005
R25681 MULT_0.4bit_ADDER_2.B0.n21 MULT_0.4bit_ADDER_2.B0.n19 86.2638
R25682 MULT_0.4bit_ADDER_2.B0.n19 MULT_0.4bit_ADDER_2.B0.n18 85.8873
R25683 MULT_0.4bit_ADDER_2.B0.n19 MULT_0.4bit_ADDER_2.B0.n16 85.724
R25684 MULT_0.4bit_ADDER_2.B0.n2 MULT_0.4bit_ADDER_2.B0.n1 84.5046
R25685 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.Y MULT_0.4bit_ADDER_2.B0.n24 83.8907
R25686 MULT_0.4bit_ADDER_2.B0.n22 MULT_0.4bit_ADDER_2.B0.n18 75.0672
R25687 MULT_0.4bit_ADDER_2.B0.n22 MULT_0.4bit_ADDER_2.B0.n21 75.0672
R25688 MULT_0.4bit_ADDER_2.B0.n16 MULT_0.4bit_ADDER_2.B0.n15 73.1255
R25689 MULT_0.4bit_ADDER_2.B0.n18 MULT_0.4bit_ADDER_2.B0.n17 73.1255
R25690 MULT_0.4bit_ADDER_2.B0.n21 MULT_0.4bit_ADDER_2.B0.n20 73.1255
R25691 MULT_0.4bit_ADDER_2.B0.n1 MULT_0.4bit_ADDER_2.B0.n0 72.3005
R25692 MULT_0.4bit_ADDER_2.B0.n23 MULT_0.4bit_ADDER_2.B0.n16 68.8946
R25693 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_0.A MULT_0.4bit_ADDER_2.B0.n2 60.9816
R25694 MULT_0.4bit_ADDER_2.B0.n24 MULT_0.4bit_ADDER_2.B0.n14 41.9827
R25695 MULT_0.4bit_ADDER_2.B0.n13 MULT_0.4bit_ADDER_2.B0.t1 30.462
R25696 MULT_0.4bit_ADDER_2.B0.n13 MULT_0.4bit_ADDER_2.B0.t8 30.462
R25697 MULT_0.4bit_ADDER_2.B0.n11 MULT_0.4bit_ADDER_2.B0.t7 30.462
R25698 MULT_0.4bit_ADDER_2.B0.n11 MULT_0.4bit_ADDER_2.B0.t3 30.462
R25699 MULT_0.4bit_ADDER_2.B0.n10 MULT_0.4bit_ADDER_2.B0.t2 30.462
R25700 MULT_0.4bit_ADDER_2.B0.n10 MULT_0.4bit_ADDER_2.B0.t0 30.462
R25701 MULT_0.4bit_ADDER_2.B0.n14 MULT_0.4bit_ADDER_2.B0.n12 28.124
R25702 MULT_0.4bit_ADDER_2.B0.n5 MULT_0.4bit_ADDER_2.B0.n4 17.8661
R25703 MULT_0.4bit_ADDER_2.B0.n6 MULT_0.4bit_ADDER_2.B0.n5 17.8661
R25704 MULT_0.4bit_ADDER_2.B0.n7 MULT_0.4bit_ADDER_2.B0.n6 17.1217
R25705 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_0.A MULT_0.4bit_ADDER_2.B0.n8 15.6329
R25706 MULT_0.4bit_ADDER_2.B0.n17 MULT_0.4bit_ADDER_2.B0.t10 11.8205
R25707 MULT_0.4bit_ADDER_2.B0.n17 MULT_0.4bit_ADDER_2.B0.t11 11.8205
R25708 MULT_0.4bit_ADDER_2.B0.n15 MULT_0.4bit_ADDER_2.B0.t9 11.8205
R25709 MULT_0.4bit_ADDER_2.B0.n15 MULT_0.4bit_ADDER_2.B0.t5 11.8205
R25710 MULT_0.4bit_ADDER_2.B0.n20 MULT_0.4bit_ADDER_2.B0.t4 11.8205
R25711 MULT_0.4bit_ADDER_2.B0.n20 MULT_0.4bit_ADDER_2.B0.t6 11.8205
R25712 MULT_0.4bit_ADDER_2.B0.n9 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_0.A 10.8165
R25713 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.Y MULT_0.4bit_ADDER_1.FULL_ADDER_2.OUT 10.6476
R25714 MULT_0.4bit_ADDER_2.B0.n23 MULT_0.4bit_ADDER_2.B0.n22 9.3005
R25715 MULT_0.4bit_ADDER_2.B0.n8 MULT_0.4bit_ADDER_2.B0.n7 1.8615
R25716 MULT_0.4bit_ADDER_1.FULL_ADDER_2.OUT MULT_0.4bit_ADDER_2.FULL_ADDER_3.B 0.907191
R25717 MULT_0.4bit_ADDER_2.FULL_ADDER_3.B MULT_0.4bit_ADDER_2.B0.n9 0.868733
R25718 a_n14155_n11683.n0 a_n14155_n11683.t5 539.788
R25719 a_n14155_n11683.n1 a_n14155_n11683.t7 531.496
R25720 a_n14155_n11683.n0 a_n14155_n11683.t4 490.034
R25721 a_n14155_n11683.n5 a_n14155_n11683.t0 283.788
R25722 a_n14155_n11683.t1 a_n14155_n11683.n5 205.489
R25723 a_n14155_n11683.n2 a_n14155_n11683.t3 182.625
R25724 a_n14155_n11683.n3 a_n14155_n11683.t6 179.054
R25725 a_n14155_n11683.n2 a_n14155_n11683.t2 139.78
R25726 a_n14155_n11683.n4 a_n14155_n11683.n3 101.368
R25727 a_n14155_n11683.n5 a_n14155_n11683.n4 77.9135
R25728 a_n14155_n11683.n4 a_n14155_n11683.n1 76.1557
R25729 a_n14155_n11683.n1 a_n14155_n11683.n0 8.29297
R25730 a_n14155_n11683.n3 a_n14155_n11683.n2 3.57087
R25731 a_n13975_n11683.n2 a_n13975_n11683.n0 121.353
R25732 a_n13975_n11683.n2 a_n13975_n11683.n1 121.001
R25733 a_n13975_n11683.n3 a_n13975_n11683.n2 120.977
R25734 a_n13975_n11683.n0 a_n13975_n11683.t3 30.462
R25735 a_n13975_n11683.n0 a_n13975_n11683.t4 30.462
R25736 a_n13975_n11683.n1 a_n13975_n11683.t0 30.462
R25737 a_n13975_n11683.n1 a_n13975_n11683.t5 30.462
R25738 a_n13975_n11683.n3 a_n13975_n11683.t1 30.462
R25739 a_n13975_n11683.t2 a_n13975_n11683.n3 30.462
R25740 a_9528_n17350.t0 a_9528_n17350.t1 9.9005
R25741 mux8_4.NAND4F_1.Y.n2 mux8_4.NAND4F_1.Y.t11 978.795
R25742 mux8_4.NAND4F_1.Y.n1 mux8_4.NAND4F_1.Y.t9 308.481
R25743 mux8_4.NAND4F_1.Y.n1 mux8_4.NAND4F_1.Y.t10 308.481
R25744 mux8_4.NAND4F_1.Y.n0 mux8_4.NAND4F_1.Y.n3 187.373
R25745 mux8_4.NAND4F_1.Y.n0 mux8_4.NAND4F_1.Y.n4 187.192
R25746 mux8_4.NAND4F_1.Y.n0 mux8_4.NAND4F_1.Y.n5 187.192
R25747 mux8_4.NAND4F_1.Y.n7 mux8_4.NAND4F_1.Y.n6 187.192
R25748 mux8_4.NAND4F_1.Y mux8_4.NAND4F_1.Y.n2 161.84
R25749 mux8_4.NAND4F_1.Y mux8_4.NAND4F_1.Y.t4 23.4335
R25750 mux8_4.NAND4F_1.Y.n3 mux8_4.NAND4F_1.Y.t1 20.1899
R25751 mux8_4.NAND4F_1.Y.n3 mux8_4.NAND4F_1.Y.t0 20.1899
R25752 mux8_4.NAND4F_1.Y.n4 mux8_4.NAND4F_1.Y.t3 20.1899
R25753 mux8_4.NAND4F_1.Y.n4 mux8_4.NAND4F_1.Y.t2 20.1899
R25754 mux8_4.NAND4F_1.Y.n5 mux8_4.NAND4F_1.Y.t8 20.1899
R25755 mux8_4.NAND4F_1.Y.n5 mux8_4.NAND4F_1.Y.t7 20.1899
R25756 mux8_4.NAND4F_1.Y.n6 mux8_4.NAND4F_1.Y.t6 20.1899
R25757 mux8_4.NAND4F_1.Y.n6 mux8_4.NAND4F_1.Y.t5 20.1899
R25758 mux8_4.NAND4F_1.Y.n2 mux8_4.NAND4F_1.Y.n1 11.0463
R25759 mux8_4.NAND4F_1.Y mux8_4.NAND4F_1.Y.n7 0.527586
R25760 mux8_4.NAND4F_1.Y.n7 mux8_4.NAND4F_1.Y.n0 0.358709
R25761 a_2463_4914.n2 a_2463_4914.n0 121.353
R25762 a_2463_4914.n3 a_2463_4914.n2 121.353
R25763 a_2463_4914.n2 a_2463_4914.n1 121.001
R25764 a_2463_4914.n1 a_2463_4914.t4 30.462
R25765 a_2463_4914.n1 a_2463_4914.t0 30.462
R25766 a_2463_4914.n0 a_2463_4914.t3 30.462
R25767 a_2463_4914.n0 a_2463_4914.t5 30.462
R25768 a_2463_4914.t2 a_2463_4914.n3 30.462
R25769 a_2463_4914.n3 a_2463_4914.t1 30.462
R25770 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t10 485.221
R25771 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t7 367.928
R25772 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n5 227.526
R25773 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n4 227.266
R25774 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n6 227.266
R25775 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t9 224.478
R25776 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t8 213.688
R25777 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n2 84.5046
R25778 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n1 72.3005
R25779 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n3 61.0566
R25780 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t0 42.7747
R25781 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t5 30.379
R25782 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t4 30.379
R25783 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t2 30.379
R25784 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t1 30.379
R25785 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t3 30.379
R25786 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.t6 30.379
R25787 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A.n0 0.583137
R25788 a_n12345_n20526.n2 a_n12345_n20526.t6 541.395
R25789 a_n12345_n20526.n3 a_n12345_n20526.t3 527.402
R25790 a_n12345_n20526.n2 a_n12345_n20526.t4 491.64
R25791 a_n12345_n20526.n5 a_n12345_n20526.t0 281.906
R25792 a_n12345_n20526.t1 a_n12345_n20526.n5 204.359
R25793 a_n12345_n20526.n0 a_n12345_n20526.t7 180.73
R25794 a_n12345_n20526.n1 a_n12345_n20526.t5 179.45
R25795 a_n12345_n20526.n0 a_n12345_n20526.t2 139.78
R25796 a_n12345_n20526.n4 a_n12345_n20526.n1 105.635
R25797 a_n12345_n20526.n4 a_n12345_n20526.n3 76.0005
R25798 a_n12345_n20526.n5 a_n12345_n20526.n4 67.9685
R25799 a_n12345_n20526.n3 a_n12345_n20526.n2 13.994
R25800 a_n12345_n20526.n1 a_n12345_n20526.n0 1.28015
R25801 a_n11274_n21072.n3 a_n11274_n21072.n2 121.353
R25802 a_n11274_n21072.n2 a_n11274_n21072.n1 121.001
R25803 a_n11274_n21072.n2 a_n11274_n21072.n0 120.977
R25804 a_n11274_n21072.n0 a_n11274_n21072.t3 30.462
R25805 a_n11274_n21072.n0 a_n11274_n21072.t4 30.462
R25806 a_n11274_n21072.n1 a_n11274_n21072.t5 30.462
R25807 a_n11274_n21072.n1 a_n11274_n21072.t0 30.462
R25808 a_n11274_n21072.t2 a_n11274_n21072.n3 30.462
R25809 a_n11274_n21072.n3 a_n11274_n21072.t1 30.462
R25810 a_n12416_n7799.n7 a_n12416_n7799.n1 81.2978
R25811 a_n12416_n7799.n1 a_n12416_n7799.n6 81.1637
R25812 a_n12416_n7799.n1 a_n12416_n7799.n5 81.1637
R25813 a_n12416_n7799.n0 a_n12416_n7799.n4 81.1637
R25814 a_n12416_n7799.n0 a_n12416_n7799.n3 81.1637
R25815 a_n12416_n7799.n0 a_n12416_n7799.n2 80.9213
R25816 a_n12416_n7799.n6 a_n12416_n7799.t5 11.8205
R25817 a_n12416_n7799.n6 a_n12416_n7799.t0 11.8205
R25818 a_n12416_n7799.n5 a_n12416_n7799.t4 11.8205
R25819 a_n12416_n7799.n5 a_n12416_n7799.t3 11.8205
R25820 a_n12416_n7799.n4 a_n12416_n7799.t11 11.8205
R25821 a_n12416_n7799.n4 a_n12416_n7799.t9 11.8205
R25822 a_n12416_n7799.n3 a_n12416_n7799.t6 11.8205
R25823 a_n12416_n7799.n3 a_n12416_n7799.t10 11.8205
R25824 a_n12416_n7799.n2 a_n12416_n7799.t8 11.8205
R25825 a_n12416_n7799.n2 a_n12416_n7799.t7 11.8205
R25826 a_n12416_n7799.t2 a_n12416_n7799.n7 11.8205
R25827 a_n12416_n7799.n7 a_n12416_n7799.t1 11.8205
R25828 a_n12416_n7799.n1 a_n12416_n7799.n0 0.402735
R25829 mux8_4.NAND4F_2.D.n4 mux8_4.NAND4F_2.D.t7 1388.16
R25830 mux8_4.NAND4F_2.D.n7 mux8_4.NAND4F_2.D.t12 1388.16
R25831 mux8_4.NAND4F_2.D.n10 mux8_4.NAND4F_2.D.t4 1388.16
R25832 mux8_4.NAND4F_2.D.n1 mux8_4.NAND4F_2.D.t9 1388.16
R25833 mux8_4.NAND4F_2.D.n4 mux8_4.NAND4F_2.D.t10 350.839
R25834 mux8_4.NAND4F_2.D.n7 mux8_4.NAND4F_2.D.t13 350.839
R25835 mux8_4.NAND4F_2.D.n10 mux8_4.NAND4F_2.D.t8 350.839
R25836 mux8_4.NAND4F_2.D.n1 mux8_4.NAND4F_2.D.t5 350.839
R25837 mux8_4.NAND4F_2.D.n5 mux8_4.NAND4F_2.D.t15 308.481
R25838 mux8_4.NAND4F_2.D.n8 mux8_4.NAND4F_2.D.t14 308.481
R25839 mux8_4.NAND4F_2.D.n11 mux8_4.NAND4F_2.D.t11 308.481
R25840 mux8_4.NAND4F_2.D.n2 mux8_4.NAND4F_2.D.t6 308.481
R25841 mux8_4.NAND4F_2.D.n0 mux8_4.NAND4F_2.D.t1 256.514
R25842 mux8_4.NAND4F_2.D.n0 mux8_4.NAND4F_2.D.n3 226.258
R25843 mux8_4.NAND4F_2.D mux8_4.NAND4F_2.D.n5 161.458
R25844 mux8_4.NAND4F_2.D mux8_4.NAND4F_2.D.n11 161.435
R25845 mux8_4.NAND4F_2.D mux8_4.NAND4F_2.D.n2 161.435
R25846 mux8_4.NAND4F_2.D mux8_4.NAND4F_2.D.n8 161.429
R25847 mux8_4.NAND4F_2.D.n0 mux8_4.NAND4F_2.D.t0 83.7172
R25848 mux8_4.NAND4F_2.D.n3 mux8_4.NAND4F_2.D.t3 30.379
R25849 mux8_4.NAND4F_2.D.n3 mux8_4.NAND4F_2.D.t2 30.379
R25850 mux8_4.NAND4F_2.D.n5 mux8_4.NAND4F_2.D.n4 27.752
R25851 mux8_4.NAND4F_2.D.n8 mux8_4.NAND4F_2.D.n7 27.752
R25852 mux8_4.NAND4F_2.D.n11 mux8_4.NAND4F_2.D.n10 27.752
R25853 mux8_4.NAND4F_2.D.n2 mux8_4.NAND4F_2.D.n1 27.752
R25854 mux8_4.NAND4F_2.D.n6 mux8_4.NAND4F_2.D.n0 12.759
R25855 mux8_4.NAND4F_2.D mux8_4.NAND4F_2.D.n12 10.6871
R25856 mux8_4.NAND4F_2.D.n6 mux8_4.NAND4F_2.D 9.0005
R25857 mux8_4.NAND4F_2.D.n12 mux8_4.NAND4F_2.D 9.0005
R25858 mux8_4.NAND4F_2.D.n9 mux8_4.NAND4F_2.D 9.0005
R25859 mux8_4.NAND4F_2.D.n9 mux8_4.NAND4F_2.D.n6 1.74507
R25860 mux8_4.NAND4F_2.D.n12 mux8_4.NAND4F_2.D.n9 1.69072
R25861 MULT_0.4bit_ADDER_1.A1.n2 MULT_0.4bit_ADDER_1.A1.t14 540.38
R25862 MULT_0.4bit_ADDER_1.A1.n3 MULT_0.4bit_ADDER_1.A1.t13 491.64
R25863 MULT_0.4bit_ADDER_1.A1.n3 MULT_0.4bit_ADDER_1.A1.t15 491.64
R25864 MULT_0.4bit_ADDER_1.A1.n3 MULT_0.4bit_ADDER_1.A1.t12 491.64
R25865 MULT_0.4bit_ADDER_1.A1.n3 MULT_0.4bit_ADDER_1.A1.t7 491.64
R25866 MULT_0.4bit_ADDER_1.A1.n0 MULT_0.4bit_ADDER_1.A1.t4 367.928
R25867 MULT_0.inv_7.Y MULT_0.4bit_ADDER_1.A1.t2 256.514
R25868 MULT_0.4bit_ADDER_1.A1.n1 MULT_0.4bit_ADDER_1.A1.t6 227.356
R25869 MULT_0.inv_7.Y MULT_0.4bit_ADDER_1.A1.n7 226.204
R25870 MULT_0.4bit_ADDER_1.A1.n0 MULT_0.4bit_ADDER_1.A1.t5 213.688
R25871 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_0.B MULT_0.4bit_ADDER_1.A1.n5 162.867
R25872 MULT_0.4bit_ADDER_1.A1.n2 MULT_0.4bit_ADDER_1.A1.n1 160.439
R25873 MULT_0.4bit_ADDER_1.A1.n4 MULT_0.4bit_ADDER_1.A1.t8 139.78
R25874 MULT_0.4bit_ADDER_1.A1.n4 MULT_0.4bit_ADDER_1.A1.t11 139.78
R25875 MULT_0.4bit_ADDER_1.A1.n4 MULT_0.4bit_ADDER_1.A1.t9 139.78
R25876 MULT_0.4bit_ADDER_1.A1.n4 MULT_0.4bit_ADDER_1.A1.t10 139.78
R25877 MULT_0.4bit_ADDER_1.A1.n1 MULT_0.4bit_ADDER_1.A1.n0 94.4341
R25878 MULT_0.inv_7.Y MULT_0.4bit_ADDER_1.A1.t0 83.8101
R25879 MULT_0.4bit_ADDER_1.A1.n5 MULT_0.4bit_ADDER_1.A1.n4 38.6833
R25880 MULT_0.4bit_ADDER_1.A1.n7 MULT_0.4bit_ADDER_1.A1.t1 30.379
R25881 MULT_0.4bit_ADDER_1.A1.n7 MULT_0.4bit_ADDER_1.A1.t3 30.379
R25882 MULT_0.4bit_ADDER_1.A1.n5 MULT_0.4bit_ADDER_1.A1.n3 28.3986
R25883 MULT_0.inv_7.Y MULT_0.4bit_ADDER_1.FULL_ADDER_2.A 18.1754
R25884 MULT_0.4bit_ADDER_1.FULL_ADDER_2.A MULT_0.4bit_ADDER_1.A1.n6 16.8032
R25885 MULT_0.4bit_ADDER_1.A1.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_0.B 9.00496
R25886 MULT_0.4bit_ADDER_1.A1.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_0.B 3.87912
R25887 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_0.B MULT_0.4bit_ADDER_1.A1.n2 0.89693
R25888 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t7 540.38
R25889 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t8 367.928
R25890 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n4 227.526
R25891 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t10 227.356
R25892 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n5 227.266
R25893 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n6 227.266
R25894 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t9 213.688
R25895 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n2 160.439
R25896 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n1 94.4341
R25897 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t3 42.7944
R25898 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t5 30.379
R25899 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t6 30.379
R25900 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t0 30.379
R25901 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t4 30.379
R25902 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t2 30.379
R25903 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.t1 30.379
R25904 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n0 13.4358
R25905 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B.n3 0.821842
R25906 OR8_0.S3.n1 OR8_0.S3.t5 1032.02
R25907 OR8_0.S3.n1 OR8_0.S3.t4 336.962
R25908 OR8_0.S3.n1 OR8_0.S3.t6 326.154
R25909 OR8_0.S3.n0 OR8_0.S3.t3 256.514
R25910 OR8_0.S3.n0 OR8_0.S3.n2 226.258
R25911 mux8_4.NAND4F_2.A OR8_0.S3.n1 162.952
R25912 OR8_0.S3.n0 OR8_0.S3.t0 83.7172
R25913 OR8_0.NOT8_0.S3 mux8_4.A3 71.8617
R25914 OR8_0.S3.n2 OR8_0.S3.t1 30.379
R25915 OR8_0.S3.n2 OR8_0.S3.t2 30.379
R25916 mux8_4.A3 mux8_4.NAND4F_2.A 14.0617
R25917 OR8_0.NOT8_0.S3 OR8_0.S3.n0 1.9182
R25918 a_n12314_n29052.n7 a_n12314_n29052.n1 81.2978
R25919 a_n12314_n29052.n0 a_n12314_n29052.n3 81.1637
R25920 a_n12314_n29052.n0 a_n12314_n29052.n4 81.1637
R25921 a_n12314_n29052.n1 a_n12314_n29052.n5 81.1637
R25922 a_n12314_n29052.n1 a_n12314_n29052.n6 81.1637
R25923 a_n12314_n29052.n0 a_n12314_n29052.n2 80.9213
R25924 a_n12314_n29052.n2 a_n12314_n29052.t3 11.8205
R25925 a_n12314_n29052.n2 a_n12314_n29052.t5 11.8205
R25926 a_n12314_n29052.n3 a_n12314_n29052.t4 11.8205
R25927 a_n12314_n29052.n3 a_n12314_n29052.t9 11.8205
R25928 a_n12314_n29052.n4 a_n12314_n29052.t8 11.8205
R25929 a_n12314_n29052.n4 a_n12314_n29052.t7 11.8205
R25930 a_n12314_n29052.n5 a_n12314_n29052.t11 11.8205
R25931 a_n12314_n29052.n5 a_n12314_n29052.t6 11.8205
R25932 a_n12314_n29052.n6 a_n12314_n29052.t10 11.8205
R25933 a_n12314_n29052.n6 a_n12314_n29052.t0 11.8205
R25934 a_n12314_n29052.t2 a_n12314_n29052.n7 11.8205
R25935 a_n12314_n29052.n7 a_n12314_n29052.t1 11.8205
R25936 a_n12314_n29052.n1 a_n12314_n29052.n0 0.402735
R25937 a_n24213_n2915.t0 a_n24213_n2915.t1 19.8005
R25938 a_n15737_n11709.n2 a_n15737_n11709.t5 541.395
R25939 a_n15737_n11709.n3 a_n15737_n11709.t2 527.402
R25940 a_n15737_n11709.n2 a_n15737_n11709.t6 491.64
R25941 a_n15737_n11709.n5 a_n15737_n11709.t0 281.906
R25942 a_n15737_n11709.t1 a_n15737_n11709.n5 204.359
R25943 a_n15737_n11709.n0 a_n15737_n11709.t4 180.73
R25944 a_n15737_n11709.n1 a_n15737_n11709.t7 179.45
R25945 a_n15737_n11709.n0 a_n15737_n11709.t3 139.78
R25946 a_n15737_n11709.n4 a_n15737_n11709.n1 105.635
R25947 a_n15737_n11709.n4 a_n15737_n11709.n3 76.0005
R25948 a_n15737_n11709.n5 a_n15737_n11709.n4 67.9685
R25949 a_n15737_n11709.n3 a_n15737_n11709.n2 13.994
R25950 a_n15737_n11709.n1 a_n15737_n11709.n0 1.28015
R25951 MULT_0.NAND2_3.Y.n0 MULT_0.NAND2_3.Y.t7 393.889
R25952 MULT_0.NAND2_3.Y.n2 MULT_0.NAND2_3.Y.t8 291.829
R25953 MULT_0.NAND2_3.Y.n2 MULT_0.NAND2_3.Y.t10 291.829
R25954 MULT_0.NAND2_3.Y.n1 MULT_0.NAND2_3.Y.n3 227.526
R25955 MULT_0.NAND2_3.Y.n1 MULT_0.NAND2_3.Y.n5 227.266
R25956 MULT_0.NAND2_3.Y.n1 MULT_0.NAND2_3.Y.n4 227.266
R25957 MULT_0.NAND2_3.Y.n2 MULT_0.NAND2_3.Y.t9 221.72
R25958 MULT_0.NAND2_3.Y.n0 MULT_0.NAND2_3.Y.n2 53.4745
R25959 MULT_0.NAND2_3.Y.n1 MULT_0.NAND2_3.Y.t0 42.7333
R25960 MULT_0.NAND2_3.Y.n3 MULT_0.NAND2_3.Y.t5 30.379
R25961 MULT_0.NAND2_3.Y.n3 MULT_0.NAND2_3.Y.t4 30.379
R25962 MULT_0.NAND2_3.Y.n5 MULT_0.NAND2_3.Y.t2 30.379
R25963 MULT_0.NAND2_3.Y.n5 MULT_0.NAND2_3.Y.t1 30.379
R25964 MULT_0.NAND2_3.Y.n4 MULT_0.NAND2_3.Y.t3 30.379
R25965 MULT_0.NAND2_3.Y.n4 MULT_0.NAND2_3.Y.t6 30.379
R25966 MULT_0.NAND2_3.Y.n1 MULT_0.NAND2_3.Y.n0 0.656302
R25967 MULT_0.SO.n1 MULT_0.SO.t6 1032.02
R25968 MULT_0.SO.n1 MULT_0.SO.t5 336.962
R25969 MULT_0.SO.n1 MULT_0.SO.t4 326.154
R25970 MULT_0.SO.n0 MULT_0.SO.t1 256.514
R25971 MULT_0.SO.n0 MULT_0.SO.n2 226.251
R25972 MULT_0.SO MULT_0.SO.n1 162.952
R25973 MULT_0.SO.n0 MULT_0.SO.t0 83.7599
R25974 MULT_0.SO.n2 MULT_0.SO.t3 30.379
R25975 MULT_0.SO.n2 MULT_0.SO.t2 30.379
R25976 MULT_0.SO MULT_0.SO.n0 12.6374
R25977 NOT8_0.S0.n1 NOT8_0.S0.t5 1032.02
R25978 NOT8_0.S0.n1 NOT8_0.S0.t6 336.962
R25979 NOT8_0.S0.n1 NOT8_0.S0.t4 326.154
R25980 NOT8_0.S0.n0 NOT8_0.S0.t2 256.514
R25981 NOT8_0.S0.n0 NOT8_0.S0.n2 226.258
R25982 NOT8_0.S0 NOT8_0.S0.n1 162.952
R25983 NOT8_0.S0.n0 NOT8_0.S0.t0 83.7172
R25984 NOT8_0.S0.n2 NOT8_0.S0.t1 30.379
R25985 NOT8_0.S0.n2 NOT8_0.S0.t3 30.379
R25986 NOT8_0.S0 NOT8_0.S0.n0 1.87132
R25987 a_8400_n30006.t0 a_8400_n30006.t1 9.9005
R25988 mux8_8.NAND4F_0.Y.n1 mux8_8.NAND4F_0.Y.t9 1388.16
R25989 mux8_8.NAND4F_0.Y.n1 mux8_8.NAND4F_0.Y.t11 350.839
R25990 mux8_8.NAND4F_0.Y.n2 mux8_8.NAND4F_0.Y.t10 308.481
R25991 mux8_8.NAND4F_0.Y.n0 mux8_8.NAND4F_0.Y.n3 187.373
R25992 mux8_8.NAND4F_0.Y.n0 mux8_8.NAND4F_0.Y.n4 187.192
R25993 mux8_8.NAND4F_0.Y.n0 mux8_8.NAND4F_0.Y.n5 187.192
R25994 mux8_8.NAND4F_0.Y mux8_8.NAND4F_0.Y.n6 187.192
R25995 mux8_8.NAND4F_0.Y mux8_8.NAND4F_0.Y.n2 161.492
R25996 mux8_8.NAND4F_0.Y.n2 mux8_8.NAND4F_0.Y.n1 27.752
R25997 mux8_8.NAND4F_0.Y mux8_8.NAND4F_0.Y.t4 23.5085
R25998 mux8_8.NAND4F_0.Y.n3 mux8_8.NAND4F_0.Y.t3 20.1899
R25999 mux8_8.NAND4F_0.Y.n3 mux8_8.NAND4F_0.Y.t2 20.1899
R26000 mux8_8.NAND4F_0.Y.n4 mux8_8.NAND4F_0.Y.t1 20.1899
R26001 mux8_8.NAND4F_0.Y.n4 mux8_8.NAND4F_0.Y.t0 20.1899
R26002 mux8_8.NAND4F_0.Y.n5 mux8_8.NAND4F_0.Y.t8 20.1899
R26003 mux8_8.NAND4F_0.Y.n5 mux8_8.NAND4F_0.Y.t7 20.1899
R26004 mux8_8.NAND4F_0.Y.n6 mux8_8.NAND4F_0.Y.t6 20.1899
R26005 mux8_8.NAND4F_0.Y.n6 mux8_8.NAND4F_0.Y.t5 20.1899
R26006 mux8_8.NAND4F_0.Y mux8_8.NAND4F_0.Y.n0 0.358709
R26007 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n9 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t13 540.38
R26008 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t9 491.64
R26009 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t11 491.64
R26010 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t7 491.64
R26011 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n4 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t14 491.64
R26012 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n7 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t15 367.928
R26013 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n2 227.526
R26014 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n8 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t16 227.356
R26015 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n1 227.266
R26016 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n3 227.266
R26017 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n7 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t17 213.688
R26018 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n6 162.852
R26019 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n9 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n8 160.439
R26020 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t12 139.78
R26021 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t10 139.78
R26022 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t18 139.78
R26023 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n5 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t8 139.78
R26024 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n8 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n7 94.4341
R26025 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n0 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t0 42.7831
R26026 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n6 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n5 38.6833
R26027 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n2 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t5 30.379
R26028 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n2 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t6 30.379
R26029 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n1 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t1 30.379
R26030 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n1 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t2 30.379
R26031 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n3 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t3 30.379
R26032 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n3 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t4 30.379
R26033 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n6 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n4 28.3986
R26034 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n0 18.8832
R26035 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n10 10.7052
R26036 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n10 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 5.09176
R26037 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n10 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 4.19292
R26038 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n9 0.794268
R26039 a_n15707_n4534.n1 a_n15707_n4534.n6 81.2978
R26040 a_n15707_n4534.n1 a_n15707_n4534.n5 81.1637
R26041 a_n15707_n4534.n0 a_n15707_n4534.n4 81.1637
R26042 a_n15707_n4534.n0 a_n15707_n4534.n3 81.1637
R26043 a_n15707_n4534.n7 a_n15707_n4534.n1 81.1637
R26044 a_n15707_n4534.n0 a_n15707_n4534.n2 80.9213
R26045 a_n15707_n4534.n6 a_n15707_n4534.t1 11.8205
R26046 a_n15707_n4534.n6 a_n15707_n4534.t0 11.8205
R26047 a_n15707_n4534.n5 a_n15707_n4534.t4 11.8205
R26048 a_n15707_n4534.n5 a_n15707_n4534.t3 11.8205
R26049 a_n15707_n4534.n4 a_n15707_n4534.t11 11.8205
R26050 a_n15707_n4534.n4 a_n15707_n4534.t9 11.8205
R26051 a_n15707_n4534.n3 a_n15707_n4534.t6 11.8205
R26052 a_n15707_n4534.n3 a_n15707_n4534.t10 11.8205
R26053 a_n15707_n4534.n2 a_n15707_n4534.t8 11.8205
R26054 a_n15707_n4534.n2 a_n15707_n4534.t7 11.8205
R26055 a_n15707_n4534.n7 a_n15707_n4534.t5 11.8205
R26056 a_n15707_n4534.t2 a_n15707_n4534.n7 11.8205
R26057 a_n15707_n4534.n1 a_n15707_n4534.n0 0.402735
R26058 mux8_2.NAND4F_2.D.n4 mux8_2.NAND4F_2.D.t11 1388.16
R26059 mux8_2.NAND4F_2.D.n7 mux8_2.NAND4F_2.D.t5 1388.16
R26060 mux8_2.NAND4F_2.D.n10 mux8_2.NAND4F_2.D.t4 1388.16
R26061 mux8_2.NAND4F_2.D.n1 mux8_2.NAND4F_2.D.t6 1388.16
R26062 mux8_2.NAND4F_2.D.n4 mux8_2.NAND4F_2.D.t14 350.839
R26063 mux8_2.NAND4F_2.D.n7 mux8_2.NAND4F_2.D.t10 350.839
R26064 mux8_2.NAND4F_2.D.n10 mux8_2.NAND4F_2.D.t15 350.839
R26065 mux8_2.NAND4F_2.D.n1 mux8_2.NAND4F_2.D.t8 350.839
R26066 mux8_2.NAND4F_2.D.n5 mux8_2.NAND4F_2.D.t13 308.481
R26067 mux8_2.NAND4F_2.D.n8 mux8_2.NAND4F_2.D.t9 308.481
R26068 mux8_2.NAND4F_2.D.n11 mux8_2.NAND4F_2.D.t12 308.481
R26069 mux8_2.NAND4F_2.D.n2 mux8_2.NAND4F_2.D.t7 308.481
R26070 mux8_2.NAND4F_2.D.n0 mux8_2.NAND4F_2.D.t1 256.514
R26071 mux8_2.NAND4F_2.D.n0 mux8_2.NAND4F_2.D.n3 226.258
R26072 mux8_2.NAND4F_2.D mux8_2.NAND4F_2.D.n5 161.458
R26073 mux8_2.NAND4F_2.D mux8_2.NAND4F_2.D.n11 161.435
R26074 mux8_2.NAND4F_2.D mux8_2.NAND4F_2.D.n2 161.435
R26075 mux8_2.NAND4F_2.D mux8_2.NAND4F_2.D.n8 161.429
R26076 mux8_2.NAND4F_2.D.n0 mux8_2.NAND4F_2.D.t0 83.7172
R26077 mux8_2.NAND4F_2.D.n3 mux8_2.NAND4F_2.D.t3 30.379
R26078 mux8_2.NAND4F_2.D.n3 mux8_2.NAND4F_2.D.t2 30.379
R26079 mux8_2.NAND4F_2.D.n5 mux8_2.NAND4F_2.D.n4 27.752
R26080 mux8_2.NAND4F_2.D.n8 mux8_2.NAND4F_2.D.n7 27.752
R26081 mux8_2.NAND4F_2.D.n11 mux8_2.NAND4F_2.D.n10 27.752
R26082 mux8_2.NAND4F_2.D.n2 mux8_2.NAND4F_2.D.n1 27.752
R26083 mux8_2.NAND4F_2.D.n6 mux8_2.NAND4F_2.D.n0 12.759
R26084 mux8_2.NAND4F_2.D mux8_2.NAND4F_2.D.n12 10.6871
R26085 mux8_2.NAND4F_2.D.n6 mux8_2.NAND4F_2.D 9.0005
R26086 mux8_2.NAND4F_2.D.n12 mux8_2.NAND4F_2.D 9.0005
R26087 mux8_2.NAND4F_2.D.n9 mux8_2.NAND4F_2.D 9.0005
R26088 mux8_2.NAND4F_2.D.n9 mux8_2.NAND4F_2.D.n6 1.74507
R26089 mux8_2.NAND4F_2.D.n12 mux8_2.NAND4F_2.D.n9 1.69072
R26090 a_9336_n7266.t0 a_9336_n7266.t1 9.9005
R26091 a_n12345_n25873.n2 a_n12345_n25873.t7 541.395
R26092 a_n12345_n25873.n3 a_n12345_n25873.t5 527.402
R26093 a_n12345_n25873.n2 a_n12345_n25873.t6 491.64
R26094 a_n12345_n25873.n5 a_n12345_n25873.t0 281.906
R26095 a_n12345_n25873.t1 a_n12345_n25873.n5 204.359
R26096 a_n12345_n25873.n0 a_n12345_n25873.t2 180.73
R26097 a_n12345_n25873.n1 a_n12345_n25873.t4 179.45
R26098 a_n12345_n25873.n0 a_n12345_n25873.t3 139.78
R26099 a_n12345_n25873.n4 a_n12345_n25873.n1 105.635
R26100 a_n12345_n25873.n4 a_n12345_n25873.n3 76.0005
R26101 a_n12345_n25873.n5 a_n12345_n25873.n4 67.9685
R26102 a_n12345_n25873.n3 a_n12345_n25873.n2 13.994
R26103 a_n12345_n25873.n1 a_n12345_n25873.n0 1.28015
R26104 a_10267_n34534.t0 a_10267_n34534.t1 9.9005
R26105 a_10363_n34534.t0 a_10363_n34534.t1 9.9005
R26106 left_shifter_0.buffer_7.inv_1.A.n0 left_shifter_0.buffer_7.inv_1.A.t7 393.921
R26107 left_shifter_0.buffer_7.inv_1.A.n2 left_shifter_0.buffer_7.inv_1.A.t4 291.829
R26108 left_shifter_0.buffer_7.inv_1.A.n2 left_shifter_0.buffer_7.inv_1.A.t6 291.829
R26109 left_shifter_0.buffer_7.inv_1.A.n0 left_shifter_0.buffer_7.inv_1.A.t1 256.89
R26110 left_shifter_0.buffer_7.inv_1.A.n0 left_shifter_0.buffer_7.inv_1.A.n1 226.538
R26111 left_shifter_0.buffer_7.inv_1.A.n2 left_shifter_0.buffer_7.inv_1.A.t5 221.72
R26112 left_shifter_0.buffer_7.inv_1.A.n0 left_shifter_0.buffer_7.inv_1.A.t0 83.795
R26113 left_shifter_0.buffer_7.inv_1.A.n0 left_shifter_0.buffer_7.inv_1.A.n2 53.7938
R26114 left_shifter_0.buffer_7.inv_1.A.n1 left_shifter_0.buffer_7.inv_1.A.t2 30.379
R26115 left_shifter_0.buffer_7.inv_1.A.n1 left_shifter_0.buffer_7.inv_1.A.t3 30.379
R26116 a_3493_4914.n3 a_3493_4914.n2 121.353
R26117 a_3493_4914.n2 a_3493_4914.n1 121.001
R26118 a_3493_4914.n2 a_3493_4914.n0 120.977
R26119 a_3493_4914.n1 a_3493_4914.t4 30.462
R26120 a_3493_4914.n1 a_3493_4914.t0 30.462
R26121 a_3493_4914.n0 a_3493_4914.t3 30.462
R26122 a_3493_4914.n0 a_3493_4914.t5 30.462
R26123 a_3493_4914.t2 a_3493_4914.n3 30.462
R26124 a_3493_4914.n3 a_3493_4914.t1 30.462
R26125 a_n23404_3164.n0 a_n23404_3164.t3 539.788
R26126 a_n23404_3164.n1 a_n23404_3164.t7 531.496
R26127 a_n23404_3164.n0 a_n23404_3164.t5 490.034
R26128 a_n23404_3164.n5 a_n23404_3164.t0 283.788
R26129 a_n23404_3164.t1 a_n23404_3164.n5 205.489
R26130 a_n23404_3164.n2 a_n23404_3164.t2 182.625
R26131 a_n23404_3164.n3 a_n23404_3164.t6 179.054
R26132 a_n23404_3164.n2 a_n23404_3164.t4 139.78
R26133 a_n23404_3164.n4 a_n23404_3164.n3 101.368
R26134 a_n23404_3164.n5 a_n23404_3164.n4 77.9135
R26135 a_n23404_3164.n4 a_n23404_3164.n1 76.1557
R26136 a_n23404_3164.n1 a_n23404_3164.n0 8.29297
R26137 a_n23404_3164.n3 a_n23404_3164.n2 3.57087
R26138 a_n23992_n18833.t0 a_n23992_n18833.t1 19.8005
R26139 a_n23065_2026.n7 a_n23065_2026.n1 81.2978
R26140 a_n23065_2026.n1 a_n23065_2026.n6 81.1637
R26141 a_n23065_2026.n1 a_n23065_2026.n5 81.1637
R26142 a_n23065_2026.n0 a_n23065_2026.n4 81.1637
R26143 a_n23065_2026.n0 a_n23065_2026.n3 81.1637
R26144 a_n23065_2026.n0 a_n23065_2026.n2 80.9213
R26145 a_n23065_2026.n6 a_n23065_2026.t9 11.8205
R26146 a_n23065_2026.n6 a_n23065_2026.t0 11.8205
R26147 a_n23065_2026.n5 a_n23065_2026.t10 11.8205
R26148 a_n23065_2026.n5 a_n23065_2026.t11 11.8205
R26149 a_n23065_2026.n4 a_n23065_2026.t8 11.8205
R26150 a_n23065_2026.n4 a_n23065_2026.t6 11.8205
R26151 a_n23065_2026.n3 a_n23065_2026.t3 11.8205
R26152 a_n23065_2026.n3 a_n23065_2026.t7 11.8205
R26153 a_n23065_2026.n2 a_n23065_2026.t4 11.8205
R26154 a_n23065_2026.n2 a_n23065_2026.t5 11.8205
R26155 a_n23065_2026.t2 a_n23065_2026.n7 11.8205
R26156 a_n23065_2026.n7 a_n23065_2026.t1 11.8205
R26157 a_n23065_2026.n1 a_n23065_2026.n0 0.402735
R26158 mux8_4.NAND4F_0.Y.n1 mux8_4.NAND4F_0.Y.t9 1388.16
R26159 mux8_4.NAND4F_0.Y.n1 mux8_4.NAND4F_0.Y.t11 350.839
R26160 mux8_4.NAND4F_0.Y.n2 mux8_4.NAND4F_0.Y.t10 308.481
R26161 mux8_4.NAND4F_0.Y.n0 mux8_4.NAND4F_0.Y.n3 187.373
R26162 mux8_4.NAND4F_0.Y.n0 mux8_4.NAND4F_0.Y.n4 187.192
R26163 mux8_4.NAND4F_0.Y.n0 mux8_4.NAND4F_0.Y.n5 187.192
R26164 mux8_4.NAND4F_0.Y mux8_4.NAND4F_0.Y.n6 187.192
R26165 mux8_4.NAND4F_0.Y mux8_4.NAND4F_0.Y.n2 161.492
R26166 mux8_4.NAND4F_0.Y.n2 mux8_4.NAND4F_0.Y.n1 27.752
R26167 mux8_4.NAND4F_0.Y mux8_4.NAND4F_0.Y.t4 23.5085
R26168 mux8_4.NAND4F_0.Y.n3 mux8_4.NAND4F_0.Y.t1 20.1899
R26169 mux8_4.NAND4F_0.Y.n3 mux8_4.NAND4F_0.Y.t0 20.1899
R26170 mux8_4.NAND4F_0.Y.n4 mux8_4.NAND4F_0.Y.t3 20.1899
R26171 mux8_4.NAND4F_0.Y.n4 mux8_4.NAND4F_0.Y.t2 20.1899
R26172 mux8_4.NAND4F_0.Y.n5 mux8_4.NAND4F_0.Y.t8 20.1899
R26173 mux8_4.NAND4F_0.Y.n5 mux8_4.NAND4F_0.Y.t7 20.1899
R26174 mux8_4.NAND4F_0.Y.n6 mux8_4.NAND4F_0.Y.t5 20.1899
R26175 mux8_4.NAND4F_0.Y.n6 mux8_4.NAND4F_0.Y.t6 20.1899
R26176 mux8_4.NAND4F_0.Y mux8_4.NAND4F_0.Y.n0 0.358709
R26177 a_n14005_n11709.n2 a_n14005_n11709.t3 541.395
R26178 a_n14005_n11709.n3 a_n14005_n11709.t7 527.402
R26179 a_n14005_n11709.n2 a_n14005_n11709.t6 491.64
R26180 a_n14005_n11709.n5 a_n14005_n11709.t0 281.906
R26181 a_n14005_n11709.t1 a_n14005_n11709.n5 204.359
R26182 a_n14005_n11709.n0 a_n14005_n11709.t5 180.73
R26183 a_n14005_n11709.n1 a_n14005_n11709.t4 179.45
R26184 a_n14005_n11709.n0 a_n14005_n11709.t2 139.78
R26185 a_n14005_n11709.n4 a_n14005_n11709.n1 105.635
R26186 a_n14005_n11709.n4 a_n14005_n11709.n3 76.0005
R26187 a_n14005_n11709.n5 a_n14005_n11709.n4 67.9685
R26188 a_n14005_n11709.n3 a_n14005_n11709.n2 13.994
R26189 a_n14005_n11709.n1 a_n14005_n11709.n0 1.28015
R26190 a_8400_n30934.t0 a_8400_n30934.t1 9.9005
R26191 a_n29_2026.n0 a_n29_2026.n2 81.2978
R26192 a_n29_2026.n0 a_n29_2026.n3 81.1637
R26193 a_n29_2026.n0 a_n29_2026.n4 81.1637
R26194 a_n29_2026.n1 a_n29_2026.n5 81.1637
R26195 a_n29_2026.n1 a_n29_2026.n6 81.1637
R26196 a_n29_2026.n7 a_n29_2026.n1 80.9213
R26197 a_n29_2026.n2 a_n29_2026.t10 11.8205
R26198 a_n29_2026.n2 a_n29_2026.t8 11.8205
R26199 a_n29_2026.n3 a_n29_2026.t4 11.8205
R26200 a_n29_2026.n3 a_n29_2026.t9 11.8205
R26201 a_n29_2026.n4 a_n29_2026.t3 11.8205
R26202 a_n29_2026.n4 a_n29_2026.t5 11.8205
R26203 a_n29_2026.n5 a_n29_2026.t6 11.8205
R26204 a_n29_2026.n5 a_n29_2026.t11 11.8205
R26205 a_n29_2026.n6 a_n29_2026.t0 11.8205
R26206 a_n29_2026.n6 a_n29_2026.t7 11.8205
R26207 a_n29_2026.t2 a_n29_2026.n7 11.8205
R26208 a_n29_2026.n7 a_n29_2026.t1 11.8205
R26209 a_n29_2026.n1 a_n29_2026.n0 0.402735
R26210 left_shifter_0.S5.n1 left_shifter_0.S5.t4 1032.02
R26211 left_shifter_0.S5.n1 left_shifter_0.S5.t5 336.962
R26212 left_shifter_0.S5.n1 left_shifter_0.S5.t6 326.154
R26213 left_shifter_0.S5.n0 left_shifter_0.S5.t0 256.89
R26214 left_shifter_0.S5.n0 left_shifter_0.S5.n2 226.635
R26215 mux8_7.NAND4F_5.A left_shifter_0.S5.n1 162.952
R26216 left_shifter_0.S5.n0 left_shifter_0.S5.t1 83.7172
R26217 mux8_7.A6 left_shifter_0.S5.n0 37.144
R26218 left_shifter_0.S5.n2 left_shifter_0.S5.t3 30.379
R26219 left_shifter_0.S5.n2 left_shifter_0.S5.t2 30.379
R26220 mux8_7.A6 mux8_7.NAND4F_5.A 11.8717
R26221 a_7644_n26406.t0 a_7644_n26406.t1 9.9005
R26222 a_n10966_3190.n2 a_n10966_3190.t4 541.395
R26223 a_n10966_3190.n3 a_n10966_3190.t6 527.402
R26224 a_n10966_3190.n2 a_n10966_3190.t2 491.64
R26225 a_n10966_3190.n5 a_n10966_3190.t0 281.906
R26226 a_n10966_3190.t1 a_n10966_3190.n5 204.359
R26227 a_n10966_3190.n0 a_n10966_3190.t3 180.73
R26228 a_n10966_3190.n1 a_n10966_3190.t7 179.45
R26229 a_n10966_3190.n0 a_n10966_3190.t5 139.78
R26230 a_n10966_3190.n4 a_n10966_3190.n1 105.635
R26231 a_n10966_3190.n4 a_n10966_3190.n3 76.0005
R26232 a_n10966_3190.n5 a_n10966_3190.n4 67.9685
R26233 a_n10966_3190.n3 a_n10966_3190.n2 13.994
R26234 a_n10966_3190.n1 a_n10966_3190.n0 1.28015
R26235 a_9528_n30934.t0 a_9528_n30934.t1 9.9005
R26236 mux8_8.NAND4F_1.Y.n2 mux8_8.NAND4F_1.Y.t11 978.795
R26237 mux8_8.NAND4F_1.Y.n1 mux8_8.NAND4F_1.Y.t9 308.481
R26238 mux8_8.NAND4F_1.Y.n1 mux8_8.NAND4F_1.Y.t10 308.481
R26239 mux8_8.NAND4F_1.Y.n0 mux8_8.NAND4F_1.Y.n3 187.373
R26240 mux8_8.NAND4F_1.Y.n0 mux8_8.NAND4F_1.Y.n4 187.192
R26241 mux8_8.NAND4F_1.Y.n0 mux8_8.NAND4F_1.Y.n5 187.192
R26242 mux8_8.NAND4F_1.Y.n7 mux8_8.NAND4F_1.Y.n6 187.192
R26243 mux8_8.NAND4F_1.Y mux8_8.NAND4F_1.Y.n2 161.84
R26244 mux8_8.NAND4F_1.Y mux8_8.NAND4F_1.Y.t2 23.4335
R26245 mux8_8.NAND4F_1.Y.n3 mux8_8.NAND4F_1.Y.t1 20.1899
R26246 mux8_8.NAND4F_1.Y.n3 mux8_8.NAND4F_1.Y.t0 20.1899
R26247 mux8_8.NAND4F_1.Y.n4 mux8_8.NAND4F_1.Y.t8 20.1899
R26248 mux8_8.NAND4F_1.Y.n4 mux8_8.NAND4F_1.Y.t7 20.1899
R26249 mux8_8.NAND4F_1.Y.n5 mux8_8.NAND4F_1.Y.t6 20.1899
R26250 mux8_8.NAND4F_1.Y.n5 mux8_8.NAND4F_1.Y.t5 20.1899
R26251 mux8_8.NAND4F_1.Y.n6 mux8_8.NAND4F_1.Y.t4 20.1899
R26252 mux8_8.NAND4F_1.Y.n6 mux8_8.NAND4F_1.Y.t3 20.1899
R26253 mux8_8.NAND4F_1.Y.n2 mux8_8.NAND4F_1.Y.n1 11.0463
R26254 mux8_8.NAND4F_1.Y mux8_8.NAND4F_1.Y.n7 0.527586
R26255 mux8_8.NAND4F_1.Y.n7 mux8_8.NAND4F_1.Y.n0 0.358709
R26256 a_10267_1690.t0 a_10267_1690.t1 9.9005
R26257 a_10363_1690.t0 a_10363_1690.t1 9.9005
R26258 a_n4909_1380.n2 a_n4909_1380.t7 541.395
R26259 a_n4909_1380.n3 a_n4909_1380.t5 527.402
R26260 a_n4909_1380.n2 a_n4909_1380.t3 491.64
R26261 a_n4909_1380.n5 a_n4909_1380.t0 281.906
R26262 a_n4909_1380.t1 a_n4909_1380.n5 204.359
R26263 a_n4909_1380.n0 a_n4909_1380.t2 180.73
R26264 a_n4909_1380.n1 a_n4909_1380.t4 179.45
R26265 a_n4909_1380.n0 a_n4909_1380.t6 139.78
R26266 a_n4909_1380.n4 a_n4909_1380.n1 105.635
R26267 a_n4909_1380.n4 a_n4909_1380.n3 76.0005
R26268 a_n4909_1380.n5 a_n4909_1380.n4 67.9685
R26269 a_n4909_1380.n3 a_n4909_1380.n2 13.994
R26270 a_n4909_1380.n1 a_n4909_1380.n0 1.28015
R26271 a_n12314_n23651.n1 a_n12314_n23651.n5 81.2978
R26272 a_n12314_n23651.n0 a_n12314_n23651.n3 81.1637
R26273 a_n12314_n23651.n0 a_n12314_n23651.n4 81.1637
R26274 a_n12314_n23651.n1 a_n12314_n23651.n6 81.1637
R26275 a_n12314_n23651.n7 a_n12314_n23651.n1 81.1637
R26276 a_n12314_n23651.n0 a_n12314_n23651.n2 80.9213
R26277 a_n12314_n23651.n2 a_n12314_n23651.t3 11.8205
R26278 a_n12314_n23651.n2 a_n12314_n23651.t5 11.8205
R26279 a_n12314_n23651.n3 a_n12314_n23651.t4 11.8205
R26280 a_n12314_n23651.n3 a_n12314_n23651.t11 11.8205
R26281 a_n12314_n23651.n4 a_n12314_n23651.t10 11.8205
R26282 a_n12314_n23651.n4 a_n12314_n23651.t9 11.8205
R26283 a_n12314_n23651.n6 a_n12314_n23651.t0 11.8205
R26284 a_n12314_n23651.n6 a_n12314_n23651.t6 11.8205
R26285 a_n12314_n23651.n5 a_n12314_n23651.t8 11.8205
R26286 a_n12314_n23651.n5 a_n12314_n23651.t7 11.8205
R26287 a_n12314_n23651.t2 a_n12314_n23651.n7 11.8205
R26288 a_n12314_n23651.n7 a_n12314_n23651.t1 11.8205
R26289 a_n12314_n23651.n1 a_n12314_n23651.n0 0.402735
R26290 left_shifter_0.buffer_5.inv_1.A.n0 left_shifter_0.buffer_5.inv_1.A.t6 393.921
R26291 left_shifter_0.buffer_5.inv_1.A.n2 left_shifter_0.buffer_5.inv_1.A.t4 291.829
R26292 left_shifter_0.buffer_5.inv_1.A.n2 left_shifter_0.buffer_5.inv_1.A.t7 291.829
R26293 left_shifter_0.buffer_5.inv_1.A.n0 left_shifter_0.buffer_5.inv_1.A.t1 256.89
R26294 left_shifter_0.buffer_5.inv_1.A.n0 left_shifter_0.buffer_5.inv_1.A.n1 226.538
R26295 left_shifter_0.buffer_5.inv_1.A.n2 left_shifter_0.buffer_5.inv_1.A.t5 221.72
R26296 left_shifter_0.buffer_5.inv_1.A.n0 left_shifter_0.buffer_5.inv_1.A.t0 83.795
R26297 left_shifter_0.buffer_5.inv_1.A.n0 left_shifter_0.buffer_5.inv_1.A.n2 53.7938
R26298 left_shifter_0.buffer_5.inv_1.A.n1 left_shifter_0.buffer_5.inv_1.A.t2 30.379
R26299 left_shifter_0.buffer_5.inv_1.A.n1 left_shifter_0.buffer_5.inv_1.A.t3 30.379
R26300 a_n914_3190.n2 a_n914_3190.n0 121.353
R26301 a_n914_3190.n3 a_n914_3190.n2 121.353
R26302 a_n914_3190.n2 a_n914_3190.n1 121.001
R26303 a_n914_3190.n1 a_n914_3190.t5 30.462
R26304 a_n914_3190.n1 a_n914_3190.t0 30.462
R26305 a_n914_3190.n0 a_n914_3190.t3 30.462
R26306 a_n914_3190.n0 a_n914_3190.t4 30.462
R26307 a_n914_3190.n3 a_n914_3190.t1 30.462
R26308 a_n914_3190.t2 a_n914_3190.n3 30.462
R26309 a_n17446_n5154.n0 a_n17446_n5154.t4 539.788
R26310 a_n17446_n5154.n1 a_n17446_n5154.t7 531.496
R26311 a_n17446_n5154.n0 a_n17446_n5154.t5 490.034
R26312 a_n17446_n5154.n5 a_n17446_n5154.t0 283.788
R26313 a_n17446_n5154.t1 a_n17446_n5154.n5 205.489
R26314 a_n17446_n5154.n2 a_n17446_n5154.t2 182.625
R26315 a_n17446_n5154.n3 a_n17446_n5154.t6 179.054
R26316 a_n17446_n5154.n2 a_n17446_n5154.t3 139.78
R26317 a_n17446_n5154.n4 a_n17446_n5154.n3 101.368
R26318 a_n17446_n5154.n5 a_n17446_n5154.n4 77.9135
R26319 a_n17446_n5154.n4 a_n17446_n5154.n1 76.1557
R26320 a_n17446_n5154.n1 a_n17446_n5154.n0 8.29297
R26321 a_n17446_n5154.n3 a_n17446_n5154.n2 3.57087
R26322 a_n17266_n5154.n2 a_n17266_n5154.n0 121.353
R26323 a_n17266_n5154.n2 a_n17266_n5154.n1 121.001
R26324 a_n17266_n5154.n3 a_n17266_n5154.n2 120.977
R26325 a_n17266_n5154.n0 a_n17266_n5154.t4 30.462
R26326 a_n17266_n5154.n0 a_n17266_n5154.t5 30.462
R26327 a_n17266_n5154.n1 a_n17266_n5154.t0 30.462
R26328 a_n17266_n5154.n1 a_n17266_n5154.t3 30.462
R26329 a_n17266_n5154.t2 a_n17266_n5154.n3 30.462
R26330 a_n17266_n5154.n3 a_n17266_n5154.t1 30.462
R26331 NOT8_0.S2.n1 NOT8_0.S2.t5 1032.02
R26332 NOT8_0.S2.n1 NOT8_0.S2.t6 336.962
R26333 NOT8_0.S2.n1 NOT8_0.S2.t4 326.154
R26334 NOT8_0.S2.n0 NOT8_0.S2.t2 256.514
R26335 NOT8_0.S2.n0 NOT8_0.S2.n2 226.258
R26336 NOT8_0.S2 NOT8_0.S2.n1 162.952
R26337 NOT8_0.S2.n0 NOT8_0.S2.t0 83.7172
R26338 NOT8_0.S2.n2 NOT8_0.S2.t1 30.379
R26339 NOT8_0.S2.n2 NOT8_0.S2.t3 30.379
R26340 NOT8_0.S2 NOT8_0.S2.n0 1.91559
R26341 a_n24162_n9284.t0 a_n24162_n9284.t1 19.8005
R26342 a_7452_n7266.t0 a_7452_n7266.t1 9.9005
R26343 a_7548_n7266.t0 a_7548_n7266.t1 9.9005
R26344 mux8_2.NAND4F_6.Y.n1 mux8_2.NAND4F_6.Y.t11 933.563
R26345 mux8_2.NAND4F_6.Y.n1 mux8_2.NAND4F_6.Y.t10 367.635
R26346 mux8_2.NAND4F_6.Y.n2 mux8_2.NAND4F_6.Y.t9 308.481
R26347 mux8_2.NAND4F_6.Y.n0 mux8_2.NAND4F_6.Y.n4 187.373
R26348 mux8_2.NAND4F_6.Y.n0 mux8_2.NAND4F_6.Y.n5 187.192
R26349 mux8_2.NAND4F_6.Y.n0 mux8_2.NAND4F_6.Y.n6 187.192
R26350 mux8_2.NAND4F_6.Y.n8 mux8_2.NAND4F_6.Y.n7 187.192
R26351 mux8_2.NAND4F_6.Y mux8_2.NAND4F_6.Y.n2 162.047
R26352 mux8_2.NAND4F_6.Y.n3 mux8_2.NAND4F_6.Y.t3 22.7831
R26353 mux8_2.NAND4F_6.Y.n3 mux8_2.NAND4F_6.Y 22.171
R26354 mux8_2.NAND4F_6.Y.n4 mux8_2.NAND4F_6.Y.t0 20.1899
R26355 mux8_2.NAND4F_6.Y.n4 mux8_2.NAND4F_6.Y.t1 20.1899
R26356 mux8_2.NAND4F_6.Y.n5 mux8_2.NAND4F_6.Y.t6 20.1899
R26357 mux8_2.NAND4F_6.Y.n5 mux8_2.NAND4F_6.Y.t5 20.1899
R26358 mux8_2.NAND4F_6.Y.n6 mux8_2.NAND4F_6.Y.t7 20.1899
R26359 mux8_2.NAND4F_6.Y.n6 mux8_2.NAND4F_6.Y.t8 20.1899
R26360 mux8_2.NAND4F_6.Y.n7 mux8_2.NAND4F_6.Y.t4 20.1899
R26361 mux8_2.NAND4F_6.Y.n7 mux8_2.NAND4F_6.Y.t2 20.1899
R26362 mux8_2.NAND4F_6.Y.n2 mux8_2.NAND4F_6.Y.n1 10.955
R26363 mux8_2.NAND4F_6.Y mux8_2.NAND4F_6.Y.n3 0.781576
R26364 mux8_2.NAND4F_6.Y mux8_2.NAND4F_6.Y.n8 0.396904
R26365 mux8_2.NAND4F_6.Y.n8 mux8_2.NAND4F_6.Y.n0 0.358709
R26366 a_10459_n20950.t0 a_10459_n20950.t1 9.9005
R26367 a_n19804_1380.n2 a_n19804_1380.t7 541.395
R26368 a_n19804_1380.n3 a_n19804_1380.t4 527.402
R26369 a_n19804_1380.n2 a_n19804_1380.t3 491.64
R26370 a_n19804_1380.n5 a_n19804_1380.t0 281.906
R26371 a_n19804_1380.t1 a_n19804_1380.n5 204.359
R26372 a_n19804_1380.n0 a_n19804_1380.t2 180.73
R26373 a_n19804_1380.n1 a_n19804_1380.t5 179.45
R26374 a_n19804_1380.n0 a_n19804_1380.t6 139.78
R26375 a_n19804_1380.n4 a_n19804_1380.n1 105.635
R26376 a_n19804_1380.n4 a_n19804_1380.n3 76.0005
R26377 a_n19804_1380.n5 a_n19804_1380.n4 67.9685
R26378 a_n19804_1380.n3 a_n19804_1380.n2 13.994
R26379 a_n19804_1380.n1 a_n19804_1380.n0 1.28015
R26380 a_n21513_1406.n0 a_n21513_1406.t5 539.788
R26381 a_n21513_1406.n1 a_n21513_1406.t4 531.496
R26382 a_n21513_1406.n0 a_n21513_1406.t2 490.034
R26383 a_n21513_1406.n5 a_n21513_1406.t0 283.788
R26384 a_n21513_1406.t1 a_n21513_1406.n5 205.489
R26385 a_n21513_1406.n2 a_n21513_1406.t3 182.625
R26386 a_n21513_1406.n3 a_n21513_1406.t7 179.054
R26387 a_n21513_1406.n2 a_n21513_1406.t6 139.78
R26388 a_n21513_1406.n4 a_n21513_1406.n3 101.368
R26389 a_n21513_1406.n5 a_n21513_1406.n4 77.9135
R26390 a_n21513_1406.n4 a_n21513_1406.n1 76.1557
R26391 a_n21513_1406.n1 a_n21513_1406.n0 8.29297
R26392 a_n21513_1406.n3 a_n21513_1406.n2 3.57087
R26393 a_n6791_1406.n0 a_n6791_1406.t6 539.788
R26394 a_n6791_1406.n1 a_n6791_1406.t2 531.496
R26395 a_n6791_1406.n0 a_n6791_1406.t3 490.034
R26396 a_n6791_1406.n5 a_n6791_1406.t0 283.788
R26397 a_n6791_1406.t1 a_n6791_1406.n5 205.489
R26398 a_n6791_1406.n2 a_n6791_1406.t4 182.625
R26399 a_n6791_1406.n3 a_n6791_1406.t5 179.054
R26400 a_n6791_1406.n2 a_n6791_1406.t7 139.78
R26401 a_n6791_1406.n4 a_n6791_1406.n3 101.368
R26402 a_n6791_1406.n5 a_n6791_1406.n4 77.9135
R26403 a_n6791_1406.n4 a_n6791_1406.n1 76.1557
R26404 a_n6791_1406.n1 a_n6791_1406.n0 8.29297
R26405 a_n6791_1406.n3 a_n6791_1406.n2 3.57087
R26406 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t10 540.38
R26407 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t9 367.928
R26408 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n4 227.526
R26409 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t7 227.356
R26410 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n5 227.266
R26411 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n6 227.266
R26412 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n1 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t8 213.688
R26413 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n3 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n2 160.439
R26414 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n2 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n1 94.4341
R26415 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n0 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t0 42.7944
R26416 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t4 30.379
R26417 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n4 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t6 30.379
R26418 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t2 30.379
R26419 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n5 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t5 30.379
R26420 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t1 30.379
R26421 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n6 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.t3 30.379
R26422 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n0 13.4358
R26423 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B.n3 0.821842
R26424 AND8_0.S6.n1 AND8_0.S6.t6 1032.02
R26425 AND8_0.S6.n1 AND8_0.S6.t4 336.962
R26426 AND8_0.S6.n1 AND8_0.S6.t5 326.154
R26427 AND8_0.S6.n0 AND8_0.S6.t1 256.514
R26428 AND8_0.S6.n0 AND8_0.S6.n2 226.258
R26429 AND8_0.S6 AND8_0.S6.n1 162.945
R26430 AND8_0.S6.n0 AND8_0.S6.t3 83.7172
R26431 AND8_0.S6.n2 AND8_0.S6.t0 30.379
R26432 AND8_0.S6.n2 AND8_0.S6.t2 30.379
R26433 AND8_0.S6 AND8_0.S6.n0 1.96507
R26434 a_n18422_n11683.n2 a_n18422_n11683.n0 121.353
R26435 a_n18422_n11683.n3 a_n18422_n11683.n2 121.353
R26436 a_n18422_n11683.n2 a_n18422_n11683.n1 121.001
R26437 a_n18422_n11683.n1 a_n18422_n11683.t5 30.462
R26438 a_n18422_n11683.n1 a_n18422_n11683.t0 30.462
R26439 a_n18422_n11683.n0 a_n18422_n11683.t4 30.462
R26440 a_n18422_n11683.n0 a_n18422_n11683.t3 30.462
R26441 a_n18422_n11683.n3 a_n18422_n11683.t1 30.462
R26442 a_n18422_n11683.t2 a_n18422_n11683.n3 30.462
R26443 mux8_3.NAND4F_2.D.n4 mux8_3.NAND4F_2.D.t15 1388.16
R26444 mux8_3.NAND4F_2.D.n7 mux8_3.NAND4F_2.D.t8 1388.16
R26445 mux8_3.NAND4F_2.D.n10 mux8_3.NAND4F_2.D.t12 1388.16
R26446 mux8_3.NAND4F_2.D.n1 mux8_3.NAND4F_2.D.t5 1388.16
R26447 mux8_3.NAND4F_2.D.n4 mux8_3.NAND4F_2.D.t6 350.839
R26448 mux8_3.NAND4F_2.D.n7 mux8_3.NAND4F_2.D.t9 350.839
R26449 mux8_3.NAND4F_2.D.n10 mux8_3.NAND4F_2.D.t4 350.839
R26450 mux8_3.NAND4F_2.D.n1 mux8_3.NAND4F_2.D.t13 350.839
R26451 mux8_3.NAND4F_2.D.n5 mux8_3.NAND4F_2.D.t11 308.481
R26452 mux8_3.NAND4F_2.D.n8 mux8_3.NAND4F_2.D.t10 308.481
R26453 mux8_3.NAND4F_2.D.n11 mux8_3.NAND4F_2.D.t7 308.481
R26454 mux8_3.NAND4F_2.D.n2 mux8_3.NAND4F_2.D.t14 308.481
R26455 mux8_3.NAND4F_2.D.n0 mux8_3.NAND4F_2.D.t1 256.514
R26456 mux8_3.NAND4F_2.D.n0 mux8_3.NAND4F_2.D.n3 226.258
R26457 mux8_3.NAND4F_2.D mux8_3.NAND4F_2.D.n5 161.458
R26458 mux8_3.NAND4F_2.D mux8_3.NAND4F_2.D.n11 161.435
R26459 mux8_3.NAND4F_2.D mux8_3.NAND4F_2.D.n2 161.435
R26460 mux8_3.NAND4F_2.D mux8_3.NAND4F_2.D.n8 161.429
R26461 mux8_3.NAND4F_2.D.n0 mux8_3.NAND4F_2.D.t0 83.7172
R26462 mux8_3.NAND4F_2.D.n3 mux8_3.NAND4F_2.D.t3 30.379
R26463 mux8_3.NAND4F_2.D.n3 mux8_3.NAND4F_2.D.t2 30.379
R26464 mux8_3.NAND4F_2.D.n5 mux8_3.NAND4F_2.D.n4 27.752
R26465 mux8_3.NAND4F_2.D.n8 mux8_3.NAND4F_2.D.n7 27.752
R26466 mux8_3.NAND4F_2.D.n11 mux8_3.NAND4F_2.D.n10 27.752
R26467 mux8_3.NAND4F_2.D.n2 mux8_3.NAND4F_2.D.n1 27.752
R26468 mux8_3.NAND4F_2.D.n6 mux8_3.NAND4F_2.D.n0 12.759
R26469 mux8_3.NAND4F_2.D mux8_3.NAND4F_2.D.n12 10.6871
R26470 mux8_3.NAND4F_2.D.n6 mux8_3.NAND4F_2.D 9.0005
R26471 mux8_3.NAND4F_2.D.n12 mux8_3.NAND4F_2.D 9.0005
R26472 mux8_3.NAND4F_2.D.n9 mux8_3.NAND4F_2.D 9.0005
R26473 mux8_3.NAND4F_2.D.n9 mux8_3.NAND4F_2.D.n6 1.74507
R26474 mux8_3.NAND4F_2.D.n12 mux8_3.NAND4F_2.D.n9 1.69072
R26475 mux8_3.NAND4F_3.Y.n7 mux8_3.NAND4F_3.Y.t9 978.795
R26476 mux8_3.NAND4F_3.Y.n6 mux8_3.NAND4F_3.Y.t11 308.481
R26477 mux8_3.NAND4F_3.Y.n6 mux8_3.NAND4F_3.Y.t10 308.481
R26478 mux8_3.NAND4F_3.Y.n0 mux8_3.NAND4F_3.Y.n1 187.373
R26479 mux8_3.NAND4F_3.Y.n0 mux8_3.NAND4F_3.Y.n2 187.192
R26480 mux8_3.NAND4F_3.Y.n0 mux8_3.NAND4F_3.Y.n3 187.192
R26481 mux8_3.NAND4F_3.Y.n5 mux8_3.NAND4F_3.Y.n4 187.192
R26482 mux8_3.NAND4F_3.Y mux8_3.NAND4F_3.Y.n7 161.839
R26483 mux8_3.NAND4F_3.Y mux8_3.NAND4F_3.Y.t0 23.4426
R26484 mux8_3.NAND4F_3.Y.n1 mux8_3.NAND4F_3.Y.t4 20.1899
R26485 mux8_3.NAND4F_3.Y.n1 mux8_3.NAND4F_3.Y.t3 20.1899
R26486 mux8_3.NAND4F_3.Y.n2 mux8_3.NAND4F_3.Y.t8 20.1899
R26487 mux8_3.NAND4F_3.Y.n2 mux8_3.NAND4F_3.Y.t7 20.1899
R26488 mux8_3.NAND4F_3.Y.n3 mux8_3.NAND4F_3.Y.t6 20.1899
R26489 mux8_3.NAND4F_3.Y.n3 mux8_3.NAND4F_3.Y.t5 20.1899
R26490 mux8_3.NAND4F_3.Y.n4 mux8_3.NAND4F_3.Y.t1 20.1899
R26491 mux8_3.NAND4F_3.Y.n4 mux8_3.NAND4F_3.Y.t2 20.1899
R26492 mux8_3.NAND4F_3.Y.n7 mux8_3.NAND4F_3.Y.n6 11.0463
R26493 mux8_3.NAND4F_3.Y mux8_3.NAND4F_3.Y.n5 0.518495
R26494 mux8_3.NAND4F_3.Y.n5 mux8_3.NAND4F_3.Y.n0 0.358709
R26495 a_7644_n35462.t0 a_7644_n35462.t1 9.9005
R26496 a_n12446_n8445.n2 a_n12446_n8445.t2 541.395
R26497 a_n12446_n8445.n3 a_n12446_n8445.t5 527.402
R26498 a_n12446_n8445.n2 a_n12446_n8445.t7 491.64
R26499 a_n12446_n8445.n5 a_n12446_n8445.t0 281.906
R26500 a_n12446_n8445.t1 a_n12446_n8445.n5 204.359
R26501 a_n12446_n8445.n0 a_n12446_n8445.t3 180.73
R26502 a_n12446_n8445.n1 a_n12446_n8445.t6 179.45
R26503 a_n12446_n8445.n0 a_n12446_n8445.t4 139.78
R26504 a_n12446_n8445.n4 a_n12446_n8445.n1 105.635
R26505 a_n12446_n8445.n4 a_n12446_n8445.n3 76.0005
R26506 a_n12446_n8445.n5 a_n12446_n8445.n4 67.9685
R26507 a_n12446_n8445.n3 a_n12446_n8445.n2 13.994
R26508 a_n12446_n8445.n1 a_n12446_n8445.n0 1.28015
R26509 a_n20587_n11709.n2 a_n20587_n11709.t5 541.395
R26510 a_n20587_n11709.n3 a_n20587_n11709.t7 527.402
R26511 a_n20587_n11709.n2 a_n20587_n11709.t6 491.64
R26512 a_n20587_n11709.n5 a_n20587_n11709.t0 281.906
R26513 a_n20587_n11709.t1 a_n20587_n11709.n5 204.359
R26514 a_n20587_n11709.n0 a_n20587_n11709.t4 180.73
R26515 a_n20587_n11709.n1 a_n20587_n11709.t2 179.45
R26516 a_n20587_n11709.n0 a_n20587_n11709.t3 139.78
R26517 a_n20587_n11709.n4 a_n20587_n11709.n1 105.635
R26518 a_n20587_n11709.n4 a_n20587_n11709.n3 76.0005
R26519 a_n20587_n11709.n5 a_n20587_n11709.n4 67.9685
R26520 a_n20587_n11709.n3 a_n20587_n11709.n2 13.994
R26521 a_n20587_n11709.n1 a_n20587_n11709.n0 1.28015
R26522 a_n20557_n11683.n3 a_n20557_n11683.n2 121.353
R26523 a_n20557_n11683.n2 a_n20557_n11683.n1 121.001
R26524 a_n20557_n11683.n2 a_n20557_n11683.n0 120.977
R26525 a_n20557_n11683.n1 a_n20557_n11683.t5 30.462
R26526 a_n20557_n11683.n1 a_n20557_n11683.t0 30.462
R26527 a_n20557_n11683.n0 a_n20557_n11683.t3 30.462
R26528 a_n20557_n11683.n0 a_n20557_n11683.t4 30.462
R26529 a_n20557_n11683.n3 a_n20557_n11683.t1 30.462
R26530 a_n20557_n11683.t2 a_n20557_n11683.n3 30.462
R26531 a_n16483_1406.n2 a_n16483_1406.n0 121.353
R26532 a_n16483_1406.n2 a_n16483_1406.n1 121.001
R26533 a_n16483_1406.n3 a_n16483_1406.n2 120.977
R26534 a_n16483_1406.n0 a_n16483_1406.t3 30.462
R26535 a_n16483_1406.n0 a_n16483_1406.t4 30.462
R26536 a_n16483_1406.n1 a_n16483_1406.t1 30.462
R26537 a_n16483_1406.n1 a_n16483_1406.t5 30.462
R26538 a_n16483_1406.t2 a_n16483_1406.n3 30.462
R26539 a_n16483_1406.n3 a_n16483_1406.t0 30.462
R26540 a_664_373.t0 a_664_373.t1 19.8005
R26541 a_n20757_1406.n2 a_n20757_1406.n1 121.353
R26542 a_n20757_1406.n2 a_n20757_1406.n0 121.353
R26543 a_n20757_1406.n3 a_n20757_1406.n2 121.001
R26544 a_n20757_1406.n1 a_n20757_1406.t0 30.462
R26545 a_n20757_1406.n1 a_n20757_1406.t1 30.462
R26546 a_n20757_1406.n0 a_n20757_1406.t3 30.462
R26547 a_n20757_1406.n0 a_n20757_1406.t4 30.462
R26548 a_n20757_1406.n3 a_n20757_1406.t5 30.462
R26549 a_n20757_1406.t2 a_n20757_1406.n3 30.462
R26550 mux8_4.NAND4F_4.Y.n6 mux8_4.NAND4F_4.Y.t11 1032.02
R26551 mux8_4.NAND4F_4.Y.n6 mux8_4.NAND4F_4.Y.t9 336.962
R26552 mux8_4.NAND4F_4.Y.n6 mux8_4.NAND4F_4.Y.t10 326.154
R26553 mux8_4.NAND4F_4.Y.n0 mux8_4.NAND4F_4.Y.n1 187.373
R26554 mux8_4.NAND4F_4.Y.n0 mux8_4.NAND4F_4.Y.n2 187.192
R26555 mux8_4.NAND4F_4.Y.n0 mux8_4.NAND4F_4.Y.n3 187.192
R26556 mux8_4.NAND4F_4.Y.n5 mux8_4.NAND4F_4.Y.n4 187.192
R26557 mux8_4.NAND4F_4.Y mux8_4.NAND4F_4.Y.n6 162.942
R26558 mux8_4.NAND4F_4.Y.n7 mux8_4.NAND4F_4.Y 24.5377
R26559 mux8_4.NAND4F_4.Y.n7 mux8_4.NAND4F_4.Y.t8 22.6141
R26560 mux8_4.NAND4F_4.Y.n1 mux8_4.NAND4F_4.Y.t1 20.1899
R26561 mux8_4.NAND4F_4.Y.n1 mux8_4.NAND4F_4.Y.t0 20.1899
R26562 mux8_4.NAND4F_4.Y.n2 mux8_4.NAND4F_4.Y.t5 20.1899
R26563 mux8_4.NAND4F_4.Y.n2 mux8_4.NAND4F_4.Y.t4 20.1899
R26564 mux8_4.NAND4F_4.Y.n3 mux8_4.NAND4F_4.Y.t3 20.1899
R26565 mux8_4.NAND4F_4.Y.n3 mux8_4.NAND4F_4.Y.t2 20.1899
R26566 mux8_4.NAND4F_4.Y.n4 mux8_4.NAND4F_4.Y.t7 20.1899
R26567 mux8_4.NAND4F_4.Y.n4 mux8_4.NAND4F_4.Y.t6 20.1899
R26568 mux8_4.NAND4F_4.Y mux8_4.NAND4F_4.Y.n7 0.894894
R26569 mux8_4.NAND4F_4.Y mux8_4.NAND4F_4.Y.n5 0.452586
R26570 mux8_4.NAND4F_4.Y.n5 mux8_4.NAND4F_4.Y.n0 0.358709
R26571 a_9432_n2838.t0 a_9432_n2838.t1 9.9005
R26572 a_10363_n8193.t0 a_10363_n8193.t1 9.9005
R26573 a_10459_n8193.t0 a_10459_n8193.t1 9.9005
R26574 a_n10864_n5154.n0 a_n10864_n5154.t2 539.788
R26575 a_n10864_n5154.n1 a_n10864_n5154.t6 531.496
R26576 a_n10864_n5154.n0 a_n10864_n5154.t5 490.034
R26577 a_n10864_n5154.n5 a_n10864_n5154.t0 283.788
R26578 a_n10864_n5154.t1 a_n10864_n5154.n5 205.489
R26579 a_n10864_n5154.n2 a_n10864_n5154.t7 182.625
R26580 a_n10864_n5154.n3 a_n10864_n5154.t4 179.054
R26581 a_n10864_n5154.n2 a_n10864_n5154.t3 139.78
R26582 a_n10864_n5154.n4 a_n10864_n5154.n3 101.368
R26583 a_n10864_n5154.n5 a_n10864_n5154.n4 77.9135
R26584 a_n10864_n5154.n4 a_n10864_n5154.n1 76.1557
R26585 a_n10864_n5154.n1 a_n10864_n5154.n0 8.29297
R26586 a_n10864_n5154.n3 a_n10864_n5154.n2 3.57087
R26587 XOR8_0.S5.n0 XOR8_0.S5.t14 1032.02
R26588 XOR8_0.S5.n0 XOR8_0.S5.t12 336.962
R26589 XOR8_0.S5.n0 XOR8_0.S5.t13 326.154
R26590 XOR8_0.S5 XOR8_0.S5.n0 162.946
R26591 XOR8_0.S5.n3 XOR8_0.S5.n1 120.999
R26592 XOR8_0.S5.n3 XOR8_0.S5.n2 120.999
R26593 XOR8_0.S5.n15 XOR8_0.S5.n14 104.865
R26594 XOR8_0.S5.n5 XOR8_0.S5.n4 92.5005
R26595 XOR8_0.S5.n12 XOR8_0.S5.n10 86.2638
R26596 XOR8_0.S5.n10 XOR8_0.S5.n9 85.8873
R26597 XOR8_0.S5.n10 XOR8_0.S5.n7 85.724
R26598 XOR8_0.S5 XOR8_0.S5.n15 83.8907
R26599 XOR8_0.S5.n13 XOR8_0.S5.n12 75.0672
R26600 XOR8_0.S5.n13 XOR8_0.S5.n9 75.0672
R26601 XOR8_0.S5.n7 XOR8_0.S5.n6 73.1255
R26602 XOR8_0.S5.n12 XOR8_0.S5.n11 73.1255
R26603 XOR8_0.S5.n9 XOR8_0.S5.n8 73.1255
R26604 XOR8_0.S5.n14 XOR8_0.S5.n7 68.5181
R26605 XOR8_0.S5.n15 XOR8_0.S5.n5 41.9827
R26606 XOR8_0.S5.n4 XOR8_0.S5.t3 30.462
R26607 XOR8_0.S5.n4 XOR8_0.S5.t10 30.462
R26608 XOR8_0.S5.n1 XOR8_0.S5.t2 30.462
R26609 XOR8_0.S5.n1 XOR8_0.S5.t1 30.462
R26610 XOR8_0.S5.n2 XOR8_0.S5.t0 30.462
R26611 XOR8_0.S5.n2 XOR8_0.S5.t4 30.462
R26612 XOR8_0.S5.n5 XOR8_0.S5.n3 28.124
R26613 XOR8_0.S5.n11 XOR8_0.S5.t5 11.8205
R26614 XOR8_0.S5.n11 XOR8_0.S5.t9 11.8205
R26615 XOR8_0.S5.n6 XOR8_0.S5.t6 11.8205
R26616 XOR8_0.S5.n6 XOR8_0.S5.t11 11.8205
R26617 XOR8_0.S5.n8 XOR8_0.S5.t8 11.8205
R26618 XOR8_0.S5.n8 XOR8_0.S5.t7 11.8205
R26619 XOR8_0.S5.n14 XOR8_0.S5.n13 9.3005
R26620 XOR8_0.S2.n0 XOR8_0.S2.t13 1032.02
R26621 XOR8_0.S2.n0 XOR8_0.S2.t14 336.962
R26622 XOR8_0.S2.n0 XOR8_0.S2.t12 326.154
R26623 XOR8_0.S2 XOR8_0.S2.n0 162.946
R26624 XOR8_0.S2.n3 XOR8_0.S2.n1 120.999
R26625 XOR8_0.S2.n3 XOR8_0.S2.n2 120.999
R26626 XOR8_0.S2.n15 XOR8_0.S2.n14 104.865
R26627 XOR8_0.S2.n5 XOR8_0.S2.n4 92.5005
R26628 XOR8_0.S2.n12 XOR8_0.S2.n10 86.2638
R26629 XOR8_0.S2.n10 XOR8_0.S2.n9 85.8873
R26630 XOR8_0.S2.n10 XOR8_0.S2.n7 85.724
R26631 XOR8_0.S2 XOR8_0.S2.n15 83.8907
R26632 XOR8_0.S2.n13 XOR8_0.S2.n9 75.0672
R26633 XOR8_0.S2.n13 XOR8_0.S2.n12 75.0672
R26634 XOR8_0.S2.n9 XOR8_0.S2.n8 73.1255
R26635 XOR8_0.S2.n12 XOR8_0.S2.n11 73.1255
R26636 XOR8_0.S2.n7 XOR8_0.S2.n6 73.1255
R26637 XOR8_0.S2.n14 XOR8_0.S2.n7 68.5181
R26638 XOR8_0.S2.n15 XOR8_0.S2.n5 41.9827
R26639 XOR8_0.S2.n4 XOR8_0.S2.t2 30.462
R26640 XOR8_0.S2.n4 XOR8_0.S2.t9 30.462
R26641 XOR8_0.S2.n1 XOR8_0.S2.t0 30.462
R26642 XOR8_0.S2.n1 XOR8_0.S2.t1 30.462
R26643 XOR8_0.S2.n2 XOR8_0.S2.t10 30.462
R26644 XOR8_0.S2.n2 XOR8_0.S2.t11 30.462
R26645 XOR8_0.S2.n5 XOR8_0.S2.n3 28.124
R26646 XOR8_0.S2.n11 XOR8_0.S2.t7 11.8205
R26647 XOR8_0.S2.n11 XOR8_0.S2.t8 11.8205
R26648 XOR8_0.S2.n8 XOR8_0.S2.t5 11.8205
R26649 XOR8_0.S2.n8 XOR8_0.S2.t4 11.8205
R26650 XOR8_0.S2.n6 XOR8_0.S2.t3 11.8205
R26651 XOR8_0.S2.n6 XOR8_0.S2.t6 11.8205
R26652 XOR8_0.S2.n14 XOR8_0.S2.n13 9.3005
R26653 a_n12314_n21072.n0 a_n12314_n21072.n2 81.2978
R26654 a_n12314_n21072.n1 a_n12314_n21072.n6 81.1637
R26655 a_n12314_n21072.n1 a_n12314_n21072.n5 81.1637
R26656 a_n12314_n21072.n0 a_n12314_n21072.n4 81.1637
R26657 a_n12314_n21072.n0 a_n12314_n21072.n3 81.1637
R26658 a_n12314_n21072.n7 a_n12314_n21072.n1 80.9213
R26659 a_n12314_n21072.n6 a_n12314_n21072.t0 11.8205
R26660 a_n12314_n21072.n6 a_n12314_n21072.t8 11.8205
R26661 a_n12314_n21072.n5 a_n12314_n21072.t7 11.8205
R26662 a_n12314_n21072.n5 a_n12314_n21072.t6 11.8205
R26663 a_n12314_n21072.n4 a_n12314_n21072.t9 11.8205
R26664 a_n12314_n21072.n4 a_n12314_n21072.t10 11.8205
R26665 a_n12314_n21072.n3 a_n12314_n21072.t11 11.8205
R26666 a_n12314_n21072.n3 a_n12314_n21072.t5 11.8205
R26667 a_n12314_n21072.n2 a_n12314_n21072.t4 11.8205
R26668 a_n12314_n21072.n2 a_n12314_n21072.t3 11.8205
R26669 a_n12314_n21072.t2 a_n12314_n21072.n7 11.8205
R26670 a_n12314_n21072.n7 a_n12314_n21072.t1 11.8205
R26671 a_n12314_n21072.n1 a_n12314_n21072.n0 0.402735
R26672 a_11194_1690.t0 a_11194_1690.t1 9.9005
R26673 a_11290_1690.t0 a_11290_1690.t1 9.9005
R26674 a_n10423_n6187.t0 a_n10423_n6187.t1 19.8005
R26675 a_n12596_n5154.n0 a_n12596_n5154.t3 539.788
R26676 a_n12596_n5154.n1 a_n12596_n5154.t5 531.496
R26677 a_n12596_n5154.n0 a_n12596_n5154.t2 490.034
R26678 a_n12596_n5154.n5 a_n12596_n5154.t0 283.788
R26679 a_n12596_n5154.t1 a_n12596_n5154.n5 205.489
R26680 a_n12596_n5154.n2 a_n12596_n5154.t7 182.625
R26681 a_n12596_n5154.n3 a_n12596_n5154.t4 179.054
R26682 a_n12596_n5154.n2 a_n12596_n5154.t6 139.78
R26683 a_n12596_n5154.n4 a_n12596_n5154.n3 101.368
R26684 a_n12596_n5154.n5 a_n12596_n5154.n4 77.9135
R26685 a_n12596_n5154.n4 a_n12596_n5154.n1 76.1557
R26686 a_n12596_n5154.n1 a_n12596_n5154.n0 8.29297
R26687 a_n12596_n5154.n3 a_n12596_n5154.n2 3.57087
R26688 a_n12347_n14753.n2 a_n12347_n14753.t2 541.395
R26689 a_n12347_n14753.n3 a_n12347_n14753.t6 527.402
R26690 a_n12347_n14753.n2 a_n12347_n14753.t7 491.64
R26691 a_n12347_n14753.n5 a_n12347_n14753.t0 281.906
R26692 a_n12347_n14753.t1 a_n12347_n14753.n5 204.359
R26693 a_n12347_n14753.n0 a_n12347_n14753.t3 180.73
R26694 a_n12347_n14753.n1 a_n12347_n14753.t5 179.45
R26695 a_n12347_n14753.n0 a_n12347_n14753.t4 139.78
R26696 a_n12347_n14753.n4 a_n12347_n14753.n1 105.635
R26697 a_n12347_n14753.n4 a_n12347_n14753.n3 76.0005
R26698 a_n12347_n14753.n5 a_n12347_n14753.n4 67.9685
R26699 a_n12347_n14753.n3 a_n12347_n14753.n2 13.994
R26700 a_n12347_n14753.n1 a_n12347_n14753.n0 1.28015
R26701 a_9432_n17350.t0 a_9432_n17350.t1 9.9005
R26702 a_n17296_n11709.n2 a_n17296_n11709.t7 541.395
R26703 a_n17296_n11709.n3 a_n17296_n11709.t5 527.402
R26704 a_n17296_n11709.n2 a_n17296_n11709.t4 491.64
R26705 a_n17296_n11709.n5 a_n17296_n11709.t0 281.906
R26706 a_n17296_n11709.t1 a_n17296_n11709.n5 204.359
R26707 a_n17296_n11709.n0 a_n17296_n11709.t6 180.73
R26708 a_n17296_n11709.n1 a_n17296_n11709.t2 179.45
R26709 a_n17296_n11709.n0 a_n17296_n11709.t3 139.78
R26710 a_n17296_n11709.n4 a_n17296_n11709.n1 105.635
R26711 a_n17296_n11709.n4 a_n17296_n11709.n3 76.0005
R26712 a_n17296_n11709.n5 a_n17296_n11709.n4 67.9685
R26713 a_n17296_n11709.n3 a_n17296_n11709.n2 13.994
R26714 a_n17296_n11709.n1 a_n17296_n11709.n0 1.28015
R26715 a_n17266_n11683.n2 a_n17266_n11683.n0 121.353
R26716 a_n17266_n11683.n2 a_n17266_n11683.n1 121.001
R26717 a_n17266_n11683.n3 a_n17266_n11683.n2 120.977
R26718 a_n17266_n11683.n0 a_n17266_n11683.t4 30.462
R26719 a_n17266_n11683.n0 a_n17266_n11683.t5 30.462
R26720 a_n17266_n11683.n1 a_n17266_n11683.t1 30.462
R26721 a_n17266_n11683.n1 a_n17266_n11683.t3 30.462
R26722 a_n17266_n11683.n3 a_n17266_n11683.t0 30.462
R26723 a_n17266_n11683.t2 a_n17266_n11683.n3 30.462
R26724 a_n8432_n12716.t0 a_n8432_n12716.t1 19.8005
R26725 MULT_0.NAND2_10.Y.n5 MULT_0.NAND2_10.Y.t8 291.829
R26726 MULT_0.NAND2_10.Y.n5 MULT_0.NAND2_10.Y.t10 291.829
R26727 MULT_0.NAND2_10.Y.n0 MULT_0.NAND2_10.Y.n3 227.526
R26728 MULT_0.NAND2_10.Y.n0 MULT_0.NAND2_10.Y.n2 227.266
R26729 MULT_0.NAND2_10.Y.n0 MULT_0.NAND2_10.Y.n4 227.266
R26730 MULT_0.NAND2_10.Y.n5 MULT_0.NAND2_10.Y.t9 221.72
R26731 MULT_0.NAND2_10.Y.t7 MULT_0.NAND2_10.Y.n1 393.897
R26732 MULT_0.NAND2_10.Y.n0 MULT_0.NAND2_10.Y.t3 42.7333
R26733 MULT_0.NAND2_10.Y.n3 MULT_0.NAND2_10.Y.t1 30.379
R26734 MULT_0.NAND2_10.Y.n3 MULT_0.NAND2_10.Y.t0 30.379
R26735 MULT_0.NAND2_10.Y.n2 MULT_0.NAND2_10.Y.t5 30.379
R26736 MULT_0.NAND2_10.Y.n2 MULT_0.NAND2_10.Y.t4 30.379
R26737 MULT_0.NAND2_10.Y.n4 MULT_0.NAND2_10.Y.t6 30.379
R26738 MULT_0.NAND2_10.Y.n4 MULT_0.NAND2_10.Y.t2 30.379
R26739 MULT_0.NAND2_10.Y.n5 MULT_0.NAND2_10.Y.n1 53.491
R26740 MULT_0.NAND2_10.Y.n0 MULT_0.NAND2_10.Y.n1 0.620141
R26741 AND8_0.S2.n1 AND8_0.S2.t6 1032.02
R26742 AND8_0.S2.n1 AND8_0.S2.t4 336.962
R26743 AND8_0.S2.n1 AND8_0.S2.t5 326.154
R26744 AND8_0.S2.n0 AND8_0.S2.t1 256.514
R26745 AND8_0.S2.n0 AND8_0.S2.n2 226.258
R26746 AND8_0.S2 AND8_0.S2.n1 162.945
R26747 AND8_0.S2.n0 AND8_0.S2.t0 83.7172
R26748 AND8_0.S2.n2 AND8_0.S2.t2 30.379
R26749 AND8_0.S2.n2 AND8_0.S2.t3 30.379
R26750 AND8_0.S2 AND8_0.S2.n0 1.92145
R26751 mux8_3.NAND4F_0.Y.n1 mux8_3.NAND4F_0.Y.t9 1388.16
R26752 mux8_3.NAND4F_0.Y.n1 mux8_3.NAND4F_0.Y.t11 350.839
R26753 mux8_3.NAND4F_0.Y.n2 mux8_3.NAND4F_0.Y.t10 308.481
R26754 mux8_3.NAND4F_0.Y.n0 mux8_3.NAND4F_0.Y.n3 187.373
R26755 mux8_3.NAND4F_0.Y.n0 mux8_3.NAND4F_0.Y.n4 187.192
R26756 mux8_3.NAND4F_0.Y.n0 mux8_3.NAND4F_0.Y.n5 187.192
R26757 mux8_3.NAND4F_0.Y mux8_3.NAND4F_0.Y.n6 187.192
R26758 mux8_3.NAND4F_0.Y mux8_3.NAND4F_0.Y.n2 161.492
R26759 mux8_3.NAND4F_0.Y.n2 mux8_3.NAND4F_0.Y.n1 27.752
R26760 mux8_3.NAND4F_0.Y mux8_3.NAND4F_0.Y.t1 23.5085
R26761 mux8_3.NAND4F_0.Y.n3 mux8_3.NAND4F_0.Y.t4 20.1899
R26762 mux8_3.NAND4F_0.Y.n3 mux8_3.NAND4F_0.Y.t3 20.1899
R26763 mux8_3.NAND4F_0.Y.n4 mux8_3.NAND4F_0.Y.t6 20.1899
R26764 mux8_3.NAND4F_0.Y.n4 mux8_3.NAND4F_0.Y.t5 20.1899
R26765 mux8_3.NAND4F_0.Y.n5 mux8_3.NAND4F_0.Y.t8 20.1899
R26766 mux8_3.NAND4F_0.Y.n5 mux8_3.NAND4F_0.Y.t7 20.1899
R26767 mux8_3.NAND4F_0.Y.n6 mux8_3.NAND4F_0.Y.t0 20.1899
R26768 mux8_3.NAND4F_0.Y.n6 mux8_3.NAND4F_0.Y.t2 20.1899
R26769 mux8_3.NAND4F_0.Y mux8_3.NAND4F_0.Y.n0 0.358709
R26770 mux8_6.NAND4F_3.Y.n7 mux8_6.NAND4F_3.Y.t9 978.795
R26771 mux8_6.NAND4F_3.Y.n6 mux8_6.NAND4F_3.Y.t11 308.481
R26772 mux8_6.NAND4F_3.Y.n6 mux8_6.NAND4F_3.Y.t10 308.481
R26773 mux8_6.NAND4F_3.Y.n0 mux8_6.NAND4F_3.Y.n1 187.373
R26774 mux8_6.NAND4F_3.Y.n0 mux8_6.NAND4F_3.Y.n2 187.192
R26775 mux8_6.NAND4F_3.Y.n0 mux8_6.NAND4F_3.Y.n3 187.192
R26776 mux8_6.NAND4F_3.Y.n5 mux8_6.NAND4F_3.Y.n4 187.192
R26777 mux8_6.NAND4F_3.Y mux8_6.NAND4F_3.Y.n7 161.839
R26778 mux8_6.NAND4F_3.Y mux8_6.NAND4F_3.Y.t6 23.4426
R26779 mux8_6.NAND4F_3.Y.n1 mux8_6.NAND4F_3.Y.t1 20.1899
R26780 mux8_6.NAND4F_3.Y.n1 mux8_6.NAND4F_3.Y.t0 20.1899
R26781 mux8_6.NAND4F_3.Y.n2 mux8_6.NAND4F_3.Y.t3 20.1899
R26782 mux8_6.NAND4F_3.Y.n2 mux8_6.NAND4F_3.Y.t2 20.1899
R26783 mux8_6.NAND4F_3.Y.n3 mux8_6.NAND4F_3.Y.t5 20.1899
R26784 mux8_6.NAND4F_3.Y.n3 mux8_6.NAND4F_3.Y.t4 20.1899
R26785 mux8_6.NAND4F_3.Y.n4 mux8_6.NAND4F_3.Y.t7 20.1899
R26786 mux8_6.NAND4F_3.Y.n4 mux8_6.NAND4F_3.Y.t8 20.1899
R26787 mux8_6.NAND4F_3.Y.n7 mux8_6.NAND4F_3.Y.n6 11.0463
R26788 mux8_6.NAND4F_3.Y mux8_6.NAND4F_3.Y.n5 0.518495
R26789 mux8_6.NAND4F_3.Y.n5 mux8_6.NAND4F_3.Y.n0 0.358709
R26790 a_8400_n2838.t0 a_8400_n2838.t1 9.9005
R26791 MULT_0.NAND2_0.Y.n5 MULT_0.NAND2_0.Y.t9 291.829
R26792 MULT_0.NAND2_0.Y.n5 MULT_0.NAND2_0.Y.t7 291.829
R26793 MULT_0.NAND2_0.Y.n0 MULT_0.NAND2_0.Y.n3 227.526
R26794 MULT_0.NAND2_0.Y.n0 MULT_0.NAND2_0.Y.n2 227.266
R26795 MULT_0.NAND2_0.Y.n0 MULT_0.NAND2_0.Y.n4 227.266
R26796 MULT_0.NAND2_0.Y.n5 MULT_0.NAND2_0.Y.t10 221.72
R26797 MULT_0.NAND2_0.Y.t8 MULT_0.NAND2_0.Y.n1 393.897
R26798 MULT_0.NAND2_0.Y.n0 MULT_0.NAND2_0.Y.t3 42.7333
R26799 MULT_0.NAND2_0.Y.n3 MULT_0.NAND2_0.Y.t1 30.379
R26800 MULT_0.NAND2_0.Y.n3 MULT_0.NAND2_0.Y.t0 30.379
R26801 MULT_0.NAND2_0.Y.n2 MULT_0.NAND2_0.Y.t5 30.379
R26802 MULT_0.NAND2_0.Y.n2 MULT_0.NAND2_0.Y.t6 30.379
R26803 MULT_0.NAND2_0.Y.n4 MULT_0.NAND2_0.Y.t4 30.379
R26804 MULT_0.NAND2_0.Y.n4 MULT_0.NAND2_0.Y.t2 30.379
R26805 MULT_0.NAND2_0.Y.n5 MULT_0.NAND2_0.Y.n1 53.4907
R26806 MULT_0.NAND2_0.Y.n0 MULT_0.NAND2_0.Y.n1 0.61864
R26807 ZFLAG_0.NAND2_0.Y.n2 ZFLAG_0.NAND2_0.Y.t7 291.829
R26808 ZFLAG_0.NAND2_0.Y.n2 ZFLAG_0.NAND2_0.Y.t10 291.829
R26809 ZFLAG_0.NAND2_0.Y.n0 ZFLAG_0.NAND2_0.Y.n4 227.526
R26810 ZFLAG_0.NAND2_0.Y.n0 ZFLAG_0.NAND2_0.Y.n5 227.266
R26811 ZFLAG_0.NAND2_0.Y.n0 ZFLAG_0.NAND2_0.Y.n3 227.266
R26812 ZFLAG_0.NAND2_0.Y.n2 ZFLAG_0.NAND2_0.Y.t9 221.72
R26813 ZFLAG_0.NAND2_0.Y.t8 ZFLAG_0.NAND2_0.Y.n1 394.019
R26814 ZFLAG_0.NAND2_0.Y.n1 ZFLAG_0.NAND2_0.Y.n2 53.3945
R26815 ZFLAG_0.NAND2_0.Y.n0 ZFLAG_0.NAND2_0.Y.t4 42.7333
R26816 ZFLAG_0.NAND2_0.Y.n5 ZFLAG_0.NAND2_0.Y.t6 30.379
R26817 ZFLAG_0.NAND2_0.Y.n5 ZFLAG_0.NAND2_0.Y.t0 30.379
R26818 ZFLAG_0.NAND2_0.Y.n3 ZFLAG_0.NAND2_0.Y.t3 30.379
R26819 ZFLAG_0.NAND2_0.Y.n3 ZFLAG_0.NAND2_0.Y.t5 30.379
R26820 ZFLAG_0.NAND2_0.Y.n4 ZFLAG_0.NAND2_0.Y.t2 30.379
R26821 ZFLAG_0.NAND2_0.Y.n4 ZFLAG_0.NAND2_0.Y.t1 30.379
R26822 ZFLAG_0.NAND2_0.Y.n0 ZFLAG_0.NAND2_0.Y.n1 0.618114
R26823 Z.n2 Z.t1 256.514
R26824 Z.n1 Z.n0 226.251
R26825 Z Z.t0 83.7464
R26826 Z.n0 Z.t3 30.379
R26827 Z.n0 Z.t2 30.379
R26828 Z.n1 Z 0.0176958
R26829 Z.n2 Z.n1 0.0073109
R26830 Z Z.n2 0.00410577
R26831 a_n20659_3190.n2 a_n20659_3190.n0 121.353
R26832 a_n20659_3190.n3 a_n20659_3190.n2 121.353
R26833 a_n20659_3190.n2 a_n20659_3190.n1 121.001
R26834 a_n20659_3190.n1 a_n20659_3190.t5 30.462
R26835 a_n20659_3190.n1 a_n20659_3190.t0 30.462
R26836 a_n20659_3190.n0 a_n20659_3190.t3 30.462
R26837 a_n20659_3190.n0 a_n20659_3190.t4 30.462
R26838 a_n20659_3190.n3 a_n20659_3190.t1 30.462
R26839 a_n20659_3190.t2 a_n20659_3190.n3 30.462
R26840 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t9 540.38
R26841 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t10 367.928
R26842 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n5 227.526
R26843 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t7 227.356
R26844 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n4 227.266
R26845 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n6 227.266
R26846 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t8 213.688
R26847 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n2 160.439
R26848 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n1 94.4341
R26849 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t3 42.7944
R26850 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t0 30.379
R26851 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t1 30.379
R26852 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t4 30.379
R26853 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t5 30.379
R26854 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t6 30.379
R26855 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.t2 30.379
R26856 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n0 13.4358
R26857 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B.n3 0.821842
R26858 mux8_7.NAND4F_4.Y.n6 mux8_7.NAND4F_4.Y.t11 1032.02
R26859 mux8_7.NAND4F_4.Y.n6 mux8_7.NAND4F_4.Y.t9 336.962
R26860 mux8_7.NAND4F_4.Y.n6 mux8_7.NAND4F_4.Y.t10 326.154
R26861 mux8_7.NAND4F_4.Y.n0 mux8_7.NAND4F_4.Y.n1 187.373
R26862 mux8_7.NAND4F_4.Y.n0 mux8_7.NAND4F_4.Y.n2 187.192
R26863 mux8_7.NAND4F_4.Y.n0 mux8_7.NAND4F_4.Y.n3 187.192
R26864 mux8_7.NAND4F_4.Y.n5 mux8_7.NAND4F_4.Y.n4 187.192
R26865 mux8_7.NAND4F_4.Y mux8_7.NAND4F_4.Y.n6 162.942
R26866 mux8_7.NAND4F_4.Y.n7 mux8_7.NAND4F_4.Y 24.5377
R26867 mux8_7.NAND4F_4.Y.n7 mux8_7.NAND4F_4.Y.t0 22.6141
R26868 mux8_7.NAND4F_4.Y.n1 mux8_7.NAND4F_4.Y.t4 20.1899
R26869 mux8_7.NAND4F_4.Y.n1 mux8_7.NAND4F_4.Y.t3 20.1899
R26870 mux8_7.NAND4F_4.Y.n2 mux8_7.NAND4F_4.Y.t6 20.1899
R26871 mux8_7.NAND4F_4.Y.n2 mux8_7.NAND4F_4.Y.t5 20.1899
R26872 mux8_7.NAND4F_4.Y.n3 mux8_7.NAND4F_4.Y.t8 20.1899
R26873 mux8_7.NAND4F_4.Y.n3 mux8_7.NAND4F_4.Y.t7 20.1899
R26874 mux8_7.NAND4F_4.Y.n4 mux8_7.NAND4F_4.Y.t1 20.1899
R26875 mux8_7.NAND4F_4.Y.n4 mux8_7.NAND4F_4.Y.t2 20.1899
R26876 mux8_7.NAND4F_4.Y mux8_7.NAND4F_4.Y.n7 0.894894
R26877 mux8_7.NAND4F_4.Y mux8_7.NAND4F_4.Y.n5 0.452586
R26878 mux8_7.NAND4F_4.Y.n5 mux8_7.NAND4F_4.Y.n0 0.358709
R26879 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t10 485.221
R26880 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t8 367.928
R26881 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n5 227.526
R26882 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n6 227.266
R26883 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n4 227.266
R26884 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t7 224.478
R26885 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t9 213.688
R26886 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n3 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n2 84.5046
R26887 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n1 72.3005
R26888 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n3 61.0566
R26889 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t6 42.7747
R26890 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t3 30.379
R26891 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n6 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t0 30.379
R26892 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t4 30.379
R26893 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n4 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t5 30.379
R26894 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t2 30.379
R26895 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n5 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.t1 30.379
R26896 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A.n0 0.583137
R26897 a_n17005_n12716.t0 a_n17005_n12716.t1 19.8005
R26898 a_9528_n2838.t0 a_9528_n2838.t1 9.9005
R26899 a_n10210_3190.n2 a_n10210_3190.n0 121.353
R26900 a_n10210_3190.n3 a_n10210_3190.n2 121.001
R26901 a_n10210_3190.n2 a_n10210_3190.n1 120.977
R26902 a_n10210_3190.n1 a_n10210_3190.t0 30.462
R26903 a_n10210_3190.n1 a_n10210_3190.t1 30.462
R26904 a_n10210_3190.n0 a_n10210_3190.t3 30.462
R26905 a_n10210_3190.n0 a_n10210_3190.t4 30.462
R26906 a_n10210_3190.n3 a_n10210_3190.t5 30.462
R26907 a_n10210_3190.t2 a_n10210_3190.n3 30.462
R26908 a_n21363_1380.n2 a_n21363_1380.t6 541.395
R26909 a_n21363_1380.n3 a_n21363_1380.t4 527.402
R26910 a_n21363_1380.n2 a_n21363_1380.t3 491.64
R26911 a_n21363_1380.n5 a_n21363_1380.t0 281.906
R26912 a_n21363_1380.t1 a_n21363_1380.n5 204.359
R26913 a_n21363_1380.n0 a_n21363_1380.t5 180.73
R26914 a_n21363_1380.n1 a_n21363_1380.t7 179.45
R26915 a_n21363_1380.n0 a_n21363_1380.t2 139.78
R26916 a_n21363_1380.n4 a_n21363_1380.n1 105.635
R26917 a_n21363_1380.n4 a_n21363_1380.n3 76.0005
R26918 a_n21363_1380.n5 a_n21363_1380.n4 67.9685
R26919 a_n21363_1380.n3 a_n21363_1380.n2 13.994
R26920 a_n21363_1380.n1 a_n21363_1380.n0 1.28015
R26921 a_n21333_1406.n3 a_n21333_1406.n2 121.353
R26922 a_n21333_1406.n2 a_n21333_1406.n1 121.001
R26923 a_n21333_1406.n2 a_n21333_1406.n0 120.977
R26924 a_n21333_1406.n1 a_n21333_1406.t3 30.462
R26925 a_n21333_1406.n1 a_n21333_1406.t1 30.462
R26926 a_n21333_1406.n0 a_n21333_1406.t5 30.462
R26927 a_n21333_1406.n0 a_n21333_1406.t4 30.462
R26928 a_n21333_1406.t2 a_n21333_1406.n3 30.462
R26929 a_n21333_1406.n3 a_n21333_1406.t0 30.462
R26930 S.n1 S.t2 256.89
R26931 S.n1 S.n0 226.635
R26932 S S.t0 83.7348
R26933 S.n0 S.t1 30.379
R26934 S.n0 S.t3 30.379
R26935 S S.n1 0.0477756
R26936 a_7644_n2838.t0 a_7644_n2838.t1 9.9005
R26937 a_n24162_n4727.t0 a_n24162_n4727.t1 19.8005
R26938 MULT_0.NAND2_8.Y.n5 MULT_0.NAND2_8.Y.t7 291.829
R26939 MULT_0.NAND2_8.Y.n5 MULT_0.NAND2_8.Y.t10 291.829
R26940 MULT_0.NAND2_8.Y.n0 MULT_0.NAND2_8.Y.n3 227.526
R26941 MULT_0.NAND2_8.Y.n0 MULT_0.NAND2_8.Y.n4 227.266
R26942 MULT_0.NAND2_8.Y.n0 MULT_0.NAND2_8.Y.n2 227.266
R26943 MULT_0.NAND2_8.Y.n5 MULT_0.NAND2_8.Y.t9 221.72
R26944 MULT_0.NAND2_8.Y.t8 MULT_0.NAND2_8.Y.n1 393.897
R26945 MULT_0.NAND2_8.Y.n0 MULT_0.NAND2_8.Y.t3 42.7333
R26946 MULT_0.NAND2_8.Y.n4 MULT_0.NAND2_8.Y.t5 30.379
R26947 MULT_0.NAND2_8.Y.n4 MULT_0.NAND2_8.Y.t0 30.379
R26948 MULT_0.NAND2_8.Y.n2 MULT_0.NAND2_8.Y.t4 30.379
R26949 MULT_0.NAND2_8.Y.n2 MULT_0.NAND2_8.Y.t6 30.379
R26950 MULT_0.NAND2_8.Y.n3 MULT_0.NAND2_8.Y.t1 30.379
R26951 MULT_0.NAND2_8.Y.n3 MULT_0.NAND2_8.Y.t2 30.379
R26952 MULT_0.NAND2_8.Y.n5 MULT_0.NAND2_8.Y.n1 53.4911
R26953 MULT_0.NAND2_8.Y.n0 MULT_0.NAND2_8.Y.n1 0.620447
R26954 a_n19981_n5154.n2 a_n19981_n5154.n0 121.353
R26955 a_n19981_n5154.n3 a_n19981_n5154.n2 121.353
R26956 a_n19981_n5154.n2 a_n19981_n5154.n1 121.001
R26957 a_n19981_n5154.n0 a_n19981_n5154.t4 30.462
R26958 a_n19981_n5154.n0 a_n19981_n5154.t3 30.462
R26959 a_n19981_n5154.n1 a_n19981_n5154.t0 30.462
R26960 a_n19981_n5154.n1 a_n19981_n5154.t5 30.462
R26961 a_n19981_n5154.t2 a_n19981_n5154.n3 30.462
R26962 a_n19981_n5154.n3 a_n19981_n5154.t1 30.462
R26963 a_n14257_3190.n2 a_n14257_3190.t4 541.395
R26964 a_n14257_3190.n3 a_n14257_3190.t6 527.402
R26965 a_n14257_3190.n2 a_n14257_3190.t2 491.64
R26966 a_n14257_3190.n5 a_n14257_3190.t0 281.906
R26967 a_n14257_3190.t1 a_n14257_3190.n5 204.359
R26968 a_n14257_3190.n0 a_n14257_3190.t5 180.73
R26969 a_n14257_3190.n1 a_n14257_3190.t3 179.45
R26970 a_n14257_3190.n0 a_n14257_3190.t7 139.78
R26971 a_n14257_3190.n4 a_n14257_3190.n1 105.635
R26972 a_n14257_3190.n4 a_n14257_3190.n3 76.0005
R26973 a_n14257_3190.n5 a_n14257_3190.n4 67.9685
R26974 a_n14257_3190.n3 a_n14257_3190.n2 13.994
R26975 a_n14257_3190.n1 a_n14257_3190.n0 1.28015
R26976 Y2.n0 Y2.t6 883.668
R26977 Y2.n1 Y2.t4 740.381
R26978 Y2.n0 Y2.t5 729.428
R26979 Y2.n2 Y2.t7 700.508
R26980 Y2.n5 Y2.t1 256.514
R26981 Y2 Y2.n3 226.251
R26982 Y2 Y2.n2 162.625
R26983 Y2.n4 Y2.t0 83.7914
R26984 Y2.n1 Y2.n0 72.3005
R26985 Y2.n3 Y2.t3 30.379
R26986 Y2.n3 Y2.t2 30.379
R26987 Y2.n2 Y2.n1 16.7975
R26988 Y2.n5 Y2.n4 0.056104
R26989 Y2.n4 Y2 0.0169921
R26990 Y2 Y2.n5 0.0117434
R26991 mux8_6.NAND4F_0.Y.n1 mux8_6.NAND4F_0.Y.t9 1388.16
R26992 mux8_6.NAND4F_0.Y.n1 mux8_6.NAND4F_0.Y.t11 350.839
R26993 mux8_6.NAND4F_0.Y.n2 mux8_6.NAND4F_0.Y.t10 308.481
R26994 mux8_6.NAND4F_0.Y.n0 mux8_6.NAND4F_0.Y.n3 187.373
R26995 mux8_6.NAND4F_0.Y.n0 mux8_6.NAND4F_0.Y.n4 187.192
R26996 mux8_6.NAND4F_0.Y.n0 mux8_6.NAND4F_0.Y.n5 187.192
R26997 mux8_6.NAND4F_0.Y mux8_6.NAND4F_0.Y.n6 187.192
R26998 mux8_6.NAND4F_0.Y mux8_6.NAND4F_0.Y.n2 161.492
R26999 mux8_6.NAND4F_0.Y.n2 mux8_6.NAND4F_0.Y.n1 27.752
R27000 mux8_6.NAND4F_0.Y mux8_6.NAND4F_0.Y.t4 23.5085
R27001 mux8_6.NAND4F_0.Y.n3 mux8_6.NAND4F_0.Y.t1 20.1899
R27002 mux8_6.NAND4F_0.Y.n3 mux8_6.NAND4F_0.Y.t0 20.1899
R27003 mux8_6.NAND4F_0.Y.n4 mux8_6.NAND4F_0.Y.t3 20.1899
R27004 mux8_6.NAND4F_0.Y.n4 mux8_6.NAND4F_0.Y.t2 20.1899
R27005 mux8_6.NAND4F_0.Y.n5 mux8_6.NAND4F_0.Y.t8 20.1899
R27006 mux8_6.NAND4F_0.Y.n5 mux8_6.NAND4F_0.Y.t7 20.1899
R27007 mux8_6.NAND4F_0.Y.n6 mux8_6.NAND4F_0.Y.t6 20.1899
R27008 mux8_6.NAND4F_0.Y.n6 mux8_6.NAND4F_0.Y.t5 20.1899
R27009 mux8_6.NAND4F_0.Y mux8_6.NAND4F_0.Y.n0 0.358709
R27010 a_n18998_n4534.n7 a_n18998_n4534.n1 81.2978
R27011 a_n18998_n4534.n1 a_n18998_n4534.n6 81.1637
R27012 a_n18998_n4534.n1 a_n18998_n4534.n5 81.1637
R27013 a_n18998_n4534.n0 a_n18998_n4534.n4 81.1637
R27014 a_n18998_n4534.n0 a_n18998_n4534.n3 81.1637
R27015 a_n18998_n4534.n0 a_n18998_n4534.n2 80.9213
R27016 a_n18998_n4534.n6 a_n18998_n4534.t3 11.8205
R27017 a_n18998_n4534.n6 a_n18998_n4534.t1 11.8205
R27018 a_n18998_n4534.n5 a_n18998_n4534.t5 11.8205
R27019 a_n18998_n4534.n5 a_n18998_n4534.t4 11.8205
R27020 a_n18998_n4534.n4 a_n18998_n4534.t10 11.8205
R27021 a_n18998_n4534.n4 a_n18998_n4534.t11 11.8205
R27022 a_n18998_n4534.n3 a_n18998_n4534.t7 11.8205
R27023 a_n18998_n4534.n3 a_n18998_n4534.t9 11.8205
R27024 a_n18998_n4534.n2 a_n18998_n4534.t6 11.8205
R27025 a_n18998_n4534.n2 a_n18998_n4534.t8 11.8205
R27026 a_n18998_n4534.n7 a_n18998_n4534.t0 11.8205
R27027 a_n18998_n4534.t2 a_n18998_n4534.n7 11.8205
R27028 a_n18998_n4534.n1 a_n18998_n4534.n0 0.402735
R27029 a_n10714_n8445.n2 a_n10714_n8445.t2 541.395
R27030 a_n10714_n8445.n3 a_n10714_n8445.t4 527.402
R27031 a_n10714_n8445.n2 a_n10714_n8445.t6 491.64
R27032 a_n10714_n8445.n5 a_n10714_n8445.t0 281.906
R27033 a_n10714_n8445.t1 a_n10714_n8445.n5 204.359
R27034 a_n10714_n8445.n0 a_n10714_n8445.t3 180.73
R27035 a_n10714_n8445.n1 a_n10714_n8445.t7 179.45
R27036 a_n10714_n8445.n0 a_n10714_n8445.t5 139.78
R27037 a_n10714_n8445.n4 a_n10714_n8445.n1 105.635
R27038 a_n10714_n8445.n4 a_n10714_n8445.n3 76.0005
R27039 a_n10714_n8445.n5 a_n10714_n8445.n4 67.9685
R27040 a_n10714_n8445.n3 a_n10714_n8445.n2 13.994
R27041 a_n10714_n8445.n1 a_n10714_n8445.n0 1.28015
R27042 a_n10684_n7799.n0 a_n10684_n7799.n4 81.2978
R27043 a_n10684_n7799.n0 a_n10684_n7799.n5 81.1637
R27044 a_n10684_n7799.n0 a_n10684_n7799.n6 81.1637
R27045 a_n10684_n7799.n1 a_n10684_n7799.n3 81.1637
R27046 a_n10684_n7799.n7 a_n10684_n7799.n1 81.1637
R27047 a_n10684_n7799.n1 a_n10684_n7799.n2 80.9213
R27048 a_n10684_n7799.n4 a_n10684_n7799.t6 11.8205
R27049 a_n10684_n7799.n4 a_n10684_n7799.t5 11.8205
R27050 a_n10684_n7799.n5 a_n10684_n7799.t8 11.8205
R27051 a_n10684_n7799.n5 a_n10684_n7799.t4 11.8205
R27052 a_n10684_n7799.n6 a_n10684_n7799.t0 11.8205
R27053 a_n10684_n7799.n6 a_n10684_n7799.t7 11.8205
R27054 a_n10684_n7799.n3 a_n10684_n7799.t11 11.8205
R27055 a_n10684_n7799.n3 a_n10684_n7799.t2 11.8205
R27056 a_n10684_n7799.n2 a_n10684_n7799.t10 11.8205
R27057 a_n10684_n7799.n2 a_n10684_n7799.t9 11.8205
R27058 a_n10684_n7799.n7 a_n10684_n7799.t1 11.8205
R27059 a_n10684_n7799.t3 a_n10684_n7799.n7 11.8205
R27060 a_n10684_n7799.n1 a_n10684_n7799.n0 0.402735
R27061 a_n9155_n8445.n2 a_n9155_n8445.t2 541.395
R27062 a_n9155_n8445.n3 a_n9155_n8445.t5 527.402
R27063 a_n9155_n8445.n2 a_n9155_n8445.t7 491.64
R27064 a_n9155_n8445.n5 a_n9155_n8445.t0 281.906
R27065 a_n9155_n8445.t1 a_n9155_n8445.n5 204.359
R27066 a_n9155_n8445.n0 a_n9155_n8445.t3 180.73
R27067 a_n9155_n8445.n1 a_n9155_n8445.t6 179.45
R27068 a_n9155_n8445.n0 a_n9155_n8445.t4 139.78
R27069 a_n9155_n8445.n4 a_n9155_n8445.n1 105.635
R27070 a_n9155_n8445.n4 a_n9155_n8445.n3 76.0005
R27071 a_n9155_n8445.n5 a_n9155_n8445.n4 67.9685
R27072 a_n9155_n8445.n3 a_n9155_n8445.n2 13.994
R27073 a_n9155_n8445.n1 a_n9155_n8445.n0 1.28015
R27074 MULT_0.S2.n0 MULT_0.S2.t13 1032.02
R27075 MULT_0.S2.n0 MULT_0.S2.t12 336.962
R27076 MULT_0.S2.n0 MULT_0.S2.t14 326.154
R27077 MULT_0.S2 MULT_0.S2.n0 162.952
R27078 MULT_0.S2.n3 MULT_0.S2.n2 120.999
R27079 MULT_0.S2.n3 MULT_0.S2.n1 120.999
R27080 MULT_0.S2.n15 MULT_0.S2.n14 104.489
R27081 MULT_0.S2.n5 MULT_0.S2.n4 92.5005
R27082 MULT_0.S2.n12 MULT_0.S2.n10 86.2638
R27083 MULT_0.S2.n10 MULT_0.S2.n9 85.8873
R27084 MULT_0.S2.n10 MULT_0.S2.n7 85.724
R27085 MULT_0.S2 MULT_0.S2.n15 83.8907
R27086 MULT_0.S2.n13 MULT_0.S2.n12 75.0672
R27087 MULT_0.S2.n13 MULT_0.S2.n9 75.0672
R27088 MULT_0.S2.n12 MULT_0.S2.n11 73.1255
R27089 MULT_0.S2.n9 MULT_0.S2.n8 73.1255
R27090 MULT_0.S2.n7 MULT_0.S2.n6 73.1255
R27091 MULT_0.S2.n14 MULT_0.S2.n7 68.8946
R27092 MULT_0.S2.n15 MULT_0.S2.n5 41.9827
R27093 MULT_0.S2.n4 MULT_0.S2.t9 30.462
R27094 MULT_0.S2.n4 MULT_0.S2.t7 30.462
R27095 MULT_0.S2.n2 MULT_0.S2.t8 30.462
R27096 MULT_0.S2.n2 MULT_0.S2.t4 30.462
R27097 MULT_0.S2.n1 MULT_0.S2.t11 30.462
R27098 MULT_0.S2.n1 MULT_0.S2.t10 30.462
R27099 MULT_0.S2.n5 MULT_0.S2.n3 28.124
R27100 MULT_0.S2.n8 MULT_0.S2.t1 11.8205
R27101 MULT_0.S2.n8 MULT_0.S2.t0 11.8205
R27102 MULT_0.S2.n11 MULT_0.S2.t5 11.8205
R27103 MULT_0.S2.n11 MULT_0.S2.t6 11.8205
R27104 MULT_0.S2.n6 MULT_0.S2.t2 11.8205
R27105 MULT_0.S2.n6 MULT_0.S2.t3 11.8205
R27106 MULT_0.S2.n14 MULT_0.S2.n13 9.3005
R27107 a_n17677_n16825.n0 a_n17677_n16825.n2 231.24
R27108 a_n17677_n16825.n1 a_n17677_n16825.n5 231.24
R27109 a_n17677_n16825.n0 a_n17677_n16825.n3 231.03
R27110 a_n17677_n16825.n1 a_n17677_n16825.n4 231.03
R27111 a_n17677_n16825.n6 a_n17677_n16825.n1 231.03
R27112 a_n17677_n16825.n2 a_n17677_n16825.t6 25.395
R27113 a_n17677_n16825.n2 a_n17677_n16825.t5 25.395
R27114 a_n17677_n16825.n3 a_n17677_n16825.t9 25.395
R27115 a_n17677_n16825.n3 a_n17677_n16825.t8 25.395
R27116 a_n17677_n16825.n4 a_n17677_n16825.t7 25.395
R27117 a_n17677_n16825.n4 a_n17677_n16825.t1 25.395
R27118 a_n17677_n16825.n5 a_n17677_n16825.t3 25.395
R27119 a_n17677_n16825.n5 a_n17677_n16825.t2 25.395
R27120 a_n17677_n16825.n6 a_n17677_n16825.t0 25.395
R27121 a_n17677_n16825.t4 a_n17677_n16825.n6 25.395
R27122 a_n17677_n16825.n1 a_n17677_n16825.n0 0.421553
R27123 a_n24012_n16501.t0 a_n24012_n16501.t1 19.8005
R27124 a_n10864_n8419.n0 a_n10864_n8419.t3 539.788
R27125 a_n10864_n8419.n1 a_n10864_n8419.t6 531.496
R27126 a_n10864_n8419.n0 a_n10864_n8419.t5 490.034
R27127 a_n10864_n8419.n5 a_n10864_n8419.t0 283.788
R27128 a_n10864_n8419.t1 a_n10864_n8419.n5 205.489
R27129 a_n10864_n8419.n2 a_n10864_n8419.t7 182.625
R27130 a_n10864_n8419.n3 a_n10864_n8419.t4 179.054
R27131 a_n10864_n8419.n2 a_n10864_n8419.t2 139.78
R27132 a_n10864_n8419.n4 a_n10864_n8419.n3 101.368
R27133 a_n10864_n8419.n5 a_n10864_n8419.n4 77.9135
R27134 a_n10864_n8419.n4 a_n10864_n8419.n1 76.1557
R27135 a_n10864_n8419.n1 a_n10864_n8419.n0 8.29297
R27136 a_n10864_n8419.n3 a_n10864_n8419.n2 3.57087
R27137 a_n10684_n8419.n2 a_n10684_n8419.n1 121.353
R27138 a_n10684_n8419.n3 a_n10684_n8419.n2 121.001
R27139 a_n10684_n8419.n2 a_n10684_n8419.n0 120.977
R27140 a_n10684_n8419.n1 a_n10684_n8419.t1 30.462
R27141 a_n10684_n8419.n1 a_n10684_n8419.t0 30.462
R27142 a_n10684_n8419.n0 a_n10684_n8419.t3 30.462
R27143 a_n10684_n8419.n0 a_n10684_n8419.t5 30.462
R27144 a_n10684_n8419.n3 a_n10684_n8419.t4 30.462
R27145 a_n10684_n8419.t2 a_n10684_n8419.n3 30.462
R27146 a_7548_n26406.t0 a_7548_n26406.t1 9.9005
R27147 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t9 485.221
R27148 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t10 367.928
R27149 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n5 227.526
R27150 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n4 227.266
R27151 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n6 227.266
R27152 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t8 224.478
R27153 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t7 213.688
R27154 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n3 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n2 84.5046
R27155 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n1 72.3005
R27156 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n3 61.0566
R27157 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t3 42.7747
R27158 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t1 30.379
R27159 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n5 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t0 30.379
R27160 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t6 30.379
R27161 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n4 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t5 30.379
R27162 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t4 30.379
R27163 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n6 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.t2 30.379
R27164 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A.n0 0.583137
R27165 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t7 540.38
R27166 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t9 367.928
R27167 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n5 227.526
R27168 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t8 227.356
R27169 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n6 227.266
R27170 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n4 227.266
R27171 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t10 213.688
R27172 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n2 160.439
R27173 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n1 94.4341
R27174 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t3 42.7944
R27175 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t6 30.379
R27176 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t0 30.379
R27177 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t4 30.379
R27178 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t5 30.379
R27179 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t1 30.379
R27180 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.t2 30.379
R27181 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n0 13.4358
R27182 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B.n3 0.821842
R27183 a_n23959_n21227.t0 a_n23959_n21227.t1 19.8005
R27184 right_shifter_0.buffer_1.inv_1.A.n0 right_shifter_0.buffer_1.inv_1.A.t4 393.921
R27185 right_shifter_0.buffer_1.inv_1.A.n2 right_shifter_0.buffer_1.inv_1.A.t7 291.829
R27186 right_shifter_0.buffer_1.inv_1.A.n2 right_shifter_0.buffer_1.inv_1.A.t6 291.829
R27187 right_shifter_0.buffer_1.inv_1.A.n0 right_shifter_0.buffer_1.inv_1.A.t1 256.514
R27188 right_shifter_0.buffer_1.inv_1.A.n0 right_shifter_0.buffer_1.inv_1.A.n1 226.162
R27189 right_shifter_0.buffer_1.inv_1.A.n2 right_shifter_0.buffer_1.inv_1.A.t5 221.72
R27190 right_shifter_0.buffer_1.inv_1.A.n0 right_shifter_0.buffer_1.inv_1.A.t0 83.795
R27191 right_shifter_0.buffer_1.inv_1.A.n0 right_shifter_0.buffer_1.inv_1.A.n2 53.7938
R27192 right_shifter_0.buffer_1.inv_1.A.n1 right_shifter_0.buffer_1.inv_1.A.t3 30.379
R27193 right_shifter_0.buffer_1.inv_1.A.n1 right_shifter_0.buffer_1.inv_1.A.t2 30.379
R27194 left_shifter_0.buffer_4.inv_1.A.n0 left_shifter_0.buffer_4.inv_1.A.t5 393.921
R27195 left_shifter_0.buffer_4.inv_1.A.n2 left_shifter_0.buffer_4.inv_1.A.t6 291.829
R27196 left_shifter_0.buffer_4.inv_1.A.n2 left_shifter_0.buffer_4.inv_1.A.t4 291.829
R27197 left_shifter_0.buffer_4.inv_1.A.n0 left_shifter_0.buffer_4.inv_1.A.t3 256.89
R27198 left_shifter_0.buffer_4.inv_1.A.n0 left_shifter_0.buffer_4.inv_1.A.n1 226.538
R27199 left_shifter_0.buffer_4.inv_1.A.n2 left_shifter_0.buffer_4.inv_1.A.t7 221.72
R27200 left_shifter_0.buffer_4.inv_1.A.n0 left_shifter_0.buffer_4.inv_1.A.t0 83.795
R27201 left_shifter_0.buffer_4.inv_1.A.n0 left_shifter_0.buffer_4.inv_1.A.n2 53.7938
R27202 left_shifter_0.buffer_4.inv_1.A.n1 left_shifter_0.buffer_4.inv_1.A.t1 30.379
R27203 left_shifter_0.buffer_4.inv_1.A.n1 left_shifter_0.buffer_4.inv_1.A.t2 30.379
R27204 a_9432_n30934.t0 a_9432_n30934.t1 9.9005
R27205 a_n12345_n28794.n2 a_n12345_n28794.t2 539.788
R27206 a_n12345_n28794.n3 a_n12345_n28794.t6 531.496
R27207 a_n12345_n28794.n2 a_n12345_n28794.t4 490.034
R27208 a_n12345_n28794.n5 a_n12345_n28794.t0 283.788
R27209 a_n12345_n28794.t1 a_n12345_n28794.n5 205.489
R27210 a_n12345_n28794.n0 a_n12345_n28794.t5 182.625
R27211 a_n12345_n28794.n1 a_n12345_n28794.t3 179.054
R27212 a_n12345_n28794.n0 a_n12345_n28794.t7 139.78
R27213 a_n12345_n28794.n4 a_n12345_n28794.n1 101.368
R27214 a_n12345_n28794.n5 a_n12345_n28794.n4 77.9135
R27215 a_n12345_n28794.n4 a_n12345_n28794.n3 76.1557
R27216 a_n12345_n28794.n3 a_n12345_n28794.n2 8.29297
R27217 a_n12345_n28794.n1 a_n12345_n28794.n0 3.57087
R27218 left_shifter_0.C.n1 left_shifter_0.C.t6 1032.02
R27219 left_shifter_0.C.n1 left_shifter_0.C.t4 336.962
R27220 left_shifter_0.C.n1 left_shifter_0.C.t5 326.154
R27221 left_shifter_0.C.n0 left_shifter_0.C.t0 256.89
R27222 left_shifter_0.C.n0 left_shifter_0.C.n2 226.635
R27223 mux8_0.NAND4F_5.A left_shifter_0.C.n1 162.952
R27224 left_shifter_0.C.n0 left_shifter_0.C.t1 83.7172
R27225 mux8_0.A6 left_shifter_0.C.n0 75.289
R27226 left_shifter_0.C.n2 left_shifter_0.C.t3 30.379
R27227 left_shifter_0.C.n2 left_shifter_0.C.t2 30.379
R27228 mux8_0.A6 mux8_0.NAND4F_5.A 11.8717
R27229 MULT_0.inv_12.A.n5 MULT_0.inv_12.A.t8 291.829
R27230 MULT_0.inv_12.A.n5 MULT_0.inv_12.A.t10 291.829
R27231 MULT_0.inv_12.A.n0 MULT_0.inv_12.A.n3 227.526
R27232 MULT_0.inv_12.A.n0 MULT_0.inv_12.A.n2 227.266
R27233 MULT_0.inv_12.A.n0 MULT_0.inv_12.A.n4 227.266
R27234 MULT_0.inv_12.A.n5 MULT_0.inv_12.A.t9 221.72
R27235 MULT_0.inv_12.A.t7 MULT_0.inv_12.A.n1 393.897
R27236 MULT_0.inv_12.A.n0 MULT_0.inv_12.A.t3 42.7333
R27237 MULT_0.inv_12.A.n3 MULT_0.inv_12.A.t1 30.379
R27238 MULT_0.inv_12.A.n3 MULT_0.inv_12.A.t0 30.379
R27239 MULT_0.inv_12.A.n2 MULT_0.inv_12.A.t6 30.379
R27240 MULT_0.inv_12.A.n2 MULT_0.inv_12.A.t5 30.379
R27241 MULT_0.inv_12.A.n4 MULT_0.inv_12.A.t4 30.379
R27242 MULT_0.inv_12.A.n4 MULT_0.inv_12.A.t2 30.379
R27243 MULT_0.inv_12.A.n5 MULT_0.inv_12.A.n1 53.4913
R27244 MULT_0.inv_12.A.n0 MULT_0.inv_12.A.n1 0.621694
R27245 a_n12596_n8419.n0 a_n12596_n8419.t4 539.788
R27246 a_n12596_n8419.n1 a_n12596_n8419.t5 531.496
R27247 a_n12596_n8419.n0 a_n12596_n8419.t3 490.034
R27248 a_n12596_n8419.n5 a_n12596_n8419.t0 283.788
R27249 a_n12596_n8419.t1 a_n12596_n8419.n5 205.489
R27250 a_n12596_n8419.n2 a_n12596_n8419.t7 182.625
R27251 a_n12596_n8419.n3 a_n12596_n8419.t2 179.054
R27252 a_n12596_n8419.n2 a_n12596_n8419.t6 139.78
R27253 a_n12596_n8419.n4 a_n12596_n8419.n3 101.368
R27254 a_n12596_n8419.n5 a_n12596_n8419.n4 77.9135
R27255 a_n12596_n8419.n4 a_n12596_n8419.n1 76.1557
R27256 a_n12596_n8419.n1 a_n12596_n8419.n0 8.29297
R27257 a_n12596_n8419.n3 a_n12596_n8419.n2 3.57087
R27258 a_n12416_n8419.n2 a_n12416_n8419.n1 121.353
R27259 a_n12416_n8419.n3 a_n12416_n8419.n2 121.001
R27260 a_n12416_n8419.n2 a_n12416_n8419.n0 120.977
R27261 a_n12416_n8419.n1 a_n12416_n8419.t4 30.462
R27262 a_n12416_n8419.n1 a_n12416_n8419.t3 30.462
R27263 a_n12416_n8419.n0 a_n12416_n8419.t0 30.462
R27264 a_n12416_n8419.n0 a_n12416_n8419.t1 30.462
R27265 a_n12416_n8419.t2 a_n12416_n8419.n3 30.462
R27266 a_n12416_n8419.n3 a_n12416_n8419.t5 30.462
R27267 a_n15896_n12716.t0 a_n15896_n12716.t1 19.8005
R27268 a_n13975_n4534.n0 a_n13975_n4534.n2 81.2978
R27269 a_n13975_n4534.n0 a_n13975_n4534.n3 81.1637
R27270 a_n13975_n4534.n0 a_n13975_n4534.n4 81.1637
R27271 a_n13975_n4534.n1 a_n13975_n4534.n5 81.1637
R27272 a_n13975_n4534.n1 a_n13975_n4534.n6 81.1637
R27273 a_n13975_n4534.n7 a_n13975_n4534.n1 80.9213
R27274 a_n13975_n4534.n2 a_n13975_n4534.t9 11.8205
R27275 a_n13975_n4534.n2 a_n13975_n4534.t10 11.8205
R27276 a_n13975_n4534.n3 a_n13975_n4534.t8 11.8205
R27277 a_n13975_n4534.n3 a_n13975_n4534.t11 11.8205
R27278 a_n13975_n4534.n4 a_n13975_n4534.t7 11.8205
R27279 a_n13975_n4534.n4 a_n13975_n4534.t6 11.8205
R27280 a_n13975_n4534.n5 a_n13975_n4534.t4 11.8205
R27281 a_n13975_n4534.n5 a_n13975_n4534.t3 11.8205
R27282 a_n13975_n4534.n6 a_n13975_n4534.t0 11.8205
R27283 a_n13975_n4534.n6 a_n13975_n4534.t5 11.8205
R27284 a_n13975_n4534.n7 a_n13975_n4534.t1 11.8205
R27285 a_n13975_n4534.t2 a_n13975_n4534.n7 11.8205
R27286 a_n13975_n4534.n1 a_n13975_n4534.n0 0.402735
R27287 mux8_5.NAND4F_4.B.n10 mux8_5.NAND4F_4.B.t6 933.563
R27288 mux8_5.NAND4F_4.B.n5 mux8_5.NAND4F_4.B.t10 933.563
R27289 mux8_5.NAND4F_4.B.n3 mux8_5.NAND4F_4.B.t15 933.563
R27290 mux8_5.NAND4F_4.B.n1 mux8_5.NAND4F_4.B.t9 933.563
R27291 mux8_5.NAND4F_4.B.n10 mux8_5.NAND4F_4.B.t11 367.635
R27292 mux8_5.NAND4F_4.B.n5 mux8_5.NAND4F_4.B.t7 367.635
R27293 mux8_5.NAND4F_4.B.n3 mux8_5.NAND4F_4.B.t12 367.635
R27294 mux8_5.NAND4F_4.B.n1 mux8_5.NAND4F_4.B.t4 367.635
R27295 mux8_5.NAND4F_4.B.n11 mux8_5.NAND4F_4.B.t13 308.481
R27296 mux8_5.NAND4F_4.B.n6 mux8_5.NAND4F_4.B.t8 308.481
R27297 mux8_5.NAND4F_4.B.n4 mux8_5.NAND4F_4.B.t14 308.481
R27298 mux8_5.NAND4F_4.B.n2 mux8_5.NAND4F_4.B.t5 308.481
R27299 mux8_5.NAND4F_4.B.n0 mux8_5.NAND4F_4.B.t1 256.514
R27300 mux8_5.NAND4F_4.B.n0 mux8_5.NAND4F_4.B.n8 226.258
R27301 mux8_5.NAND4F_4.B mux8_5.NAND4F_4.B.n2 162.173
R27302 mux8_5.NAND4F_4.B mux8_5.NAND4F_4.B.n6 162.137
R27303 mux8_5.NAND4F_4.B mux8_5.NAND4F_4.B.n11 162.117
R27304 mux8_5.NAND4F_4.B.n7 mux8_5.NAND4F_4.B.n4 161.703
R27305 mux8_5.NAND4F_4.B.n0 mux8_5.NAND4F_4.B.t0 83.7172
R27306 mux8_5.NAND4F_4.B.n8 mux8_5.NAND4F_4.B.t3 30.379
R27307 mux8_5.NAND4F_4.B.n8 mux8_5.NAND4F_4.B.t2 30.379
R27308 mux8_5.NAND4F_4.B.n12 mux8_5.NAND4F_4.B 24.8912
R27309 mux8_5.NAND4F_4.B.n7 mux8_5.NAND4F_4.B 21.6618
R27310 mux8_5.NAND4F_4.B.n11 mux8_5.NAND4F_4.B.n10 10.955
R27311 mux8_5.NAND4F_4.B.n6 mux8_5.NAND4F_4.B.n5 10.955
R27312 mux8_5.NAND4F_4.B.n4 mux8_5.NAND4F_4.B.n3 10.955
R27313 mux8_5.NAND4F_4.B.n2 mux8_5.NAND4F_4.B.n1 10.955
R27314 mux8_5.NAND4F_4.B.n12 mux8_5.NAND4F_4.B.n9 3.67985
R27315 mux8_5.NAND4F_4.B.n9 mux8_5.NAND4F_4.B.n0 1.46835
R27316 mux8_5.NAND4F_4.B mux8_5.NAND4F_4.B.n12 0.502677
R27317 mux8_5.NAND4F_4.B.n9 mux8_5.NAND4F_4.B 0.498606
R27318 mux8_5.NAND4F_4.B mux8_5.NAND4F_4.B.n7 0.470197
R27319 a_n19774_1406.n2 a_n19774_1406.n1 121.353
R27320 a_n19774_1406.n3 a_n19774_1406.n2 121.001
R27321 a_n19774_1406.n2 a_n19774_1406.n0 120.977
R27322 a_n19774_1406.n1 a_n19774_1406.t0 30.462
R27323 a_n19774_1406.n1 a_n19774_1406.t1 30.462
R27324 a_n19774_1406.n0 a_n19774_1406.t5 30.462
R27325 a_n19774_1406.n0 a_n19774_1406.t3 30.462
R27326 a_n19774_1406.n3 a_n19774_1406.t4 30.462
R27327 a_n19774_1406.t2 a_n19774_1406.n3 30.462
R27328 a_n17466_1406.n2 a_n17466_1406.n0 121.353
R27329 a_n17466_1406.n3 a_n17466_1406.n2 121.353
R27330 a_n17466_1406.n2 a_n17466_1406.n1 121.001
R27331 a_n17466_1406.n1 a_n17466_1406.t5 30.462
R27332 a_n17466_1406.n1 a_n17466_1406.t0 30.462
R27333 a_n17466_1406.n0 a_n17466_1406.t3 30.462
R27334 a_n17466_1406.n0 a_n17466_1406.t4 30.462
R27335 a_n17466_1406.n3 a_n17466_1406.t1 30.462
R27336 a_n17466_1406.t2 a_n17466_1406.n3 30.462
R27337 a_7452_n25478.t0 a_7452_n25478.t1 9.9005
R27338 a_10459_n16422.t0 a_10459_n16422.t1 9.9005
R27339 left_shifter_0.buffer_0.inv_1.A.n0 left_shifter_0.buffer_0.inv_1.A.t4 393.921
R27340 left_shifter_0.buffer_0.inv_1.A.n2 left_shifter_0.buffer_0.inv_1.A.t6 291.829
R27341 left_shifter_0.buffer_0.inv_1.A.n2 left_shifter_0.buffer_0.inv_1.A.t5 291.829
R27342 left_shifter_0.buffer_0.inv_1.A.n0 left_shifter_0.buffer_0.inv_1.A.t3 256.89
R27343 left_shifter_0.buffer_0.inv_1.A.n0 left_shifter_0.buffer_0.inv_1.A.n1 226.538
R27344 left_shifter_0.buffer_0.inv_1.A.n2 left_shifter_0.buffer_0.inv_1.A.t7 221.72
R27345 left_shifter_0.buffer_0.inv_1.A.n0 left_shifter_0.buffer_0.inv_1.A.t0 83.795
R27346 left_shifter_0.buffer_0.inv_1.A.n0 left_shifter_0.buffer_0.inv_1.A.n2 53.7938
R27347 left_shifter_0.buffer_0.inv_1.A.n1 left_shifter_0.buffer_0.inv_1.A.t1 30.379
R27348 left_shifter_0.buffer_0.inv_1.A.n1 left_shifter_0.buffer_0.inv_1.A.t2 30.379
R27349 a_n7594_1406.n2 a_n7594_1406.n1 121.353
R27350 a_n7594_1406.n2 a_n7594_1406.n0 121.353
R27351 a_n7594_1406.n3 a_n7594_1406.n2 121.001
R27352 a_n7594_1406.n1 a_n7594_1406.t0 30.462
R27353 a_n7594_1406.n1 a_n7594_1406.t1 30.462
R27354 a_n7594_1406.n0 a_n7594_1406.t5 30.462
R27355 a_n7594_1406.n0 a_n7594_1406.t3 30.462
R27356 a_n7594_1406.n3 a_n7594_1406.t4 30.462
R27357 a_n7594_1406.t2 a_n7594_1406.n3 30.462
R27358 a_10363_n20950.t0 a_10363_n20950.t1 9.9005
R27359 a_8400_n3766.t0 a_8400_n3766.t1 9.9005
R27360 a_8496_n3766.t0 a_8496_n3766.t1 9.9005
R27361 a_11194_n3766.t0 a_11194_n3766.t1 9.9005
R27362 a_n10090_373.t0 a_n10090_373.t1 19.8005
R27363 a_n17677_n25225.n0 a_n17677_n25225.n2 231.24
R27364 a_n17677_n25225.n6 a_n17677_n25225.n1 231.24
R27365 a_n17677_n25225.n0 a_n17677_n25225.n3 231.03
R27366 a_n17677_n25225.n1 a_n17677_n25225.n4 231.03
R27367 a_n17677_n25225.n1 a_n17677_n25225.n5 231.03
R27368 a_n17677_n25225.n2 a_n17677_n25225.t1 25.395
R27369 a_n17677_n25225.n2 a_n17677_n25225.t0 25.395
R27370 a_n17677_n25225.n3 a_n17677_n25225.t4 25.395
R27371 a_n17677_n25225.n3 a_n17677_n25225.t3 25.395
R27372 a_n17677_n25225.n4 a_n17677_n25225.t2 25.395
R27373 a_n17677_n25225.n4 a_n17677_n25225.t6 25.395
R27374 a_n17677_n25225.n5 a_n17677_n25225.t5 25.395
R27375 a_n17677_n25225.n5 a_n17677_n25225.t9 25.395
R27376 a_n17677_n25225.t8 a_n17677_n25225.n6 25.395
R27377 a_n17677_n25225.n6 a_n17677_n25225.t7 25.395
R27378 a_n17677_n25225.n1 a_n17677_n25225.n0 0.421553
R27379 OR8_0.NOT8_0.A7.n3 OR8_0.NOT8_0.A7.t8 394.37
R27380 OR8_0.NOT8_0.A7.n2 OR8_0.NOT8_0.A7.t10 291.829
R27381 OR8_0.NOT8_0.A7.n2 OR8_0.NOT8_0.A7.t7 291.829
R27382 OR8_0.NOT8_0.A7.n0 OR8_0.NOT8_0.A7.t1 256.425
R27383 OR8_0.NOT8_0.A7.n0 OR8_0.NOT8_0.A7.n5 231.24
R27384 OR8_0.NOT8_0.A7.n0 OR8_0.NOT8_0.A7.n6 231.03
R27385 OR8_0.NOT8_0.A7.n2 OR8_0.NOT8_0.A7.t9 221.72
R27386 OR8_0.NOT8_0.A7.n4 OR8_0.NOT8_0.A7.n1 66.4763
R27387 OR8_0.NOT8_0.A7.n3 OR8_0.NOT8_0.A7.n2 53.374
R27388 OR8_0.NOT8_0.A7.n4 OR8_0.NOT8_0.A7 37.21
R27389 OR8_0.NOT8_0.A7.n5 OR8_0.NOT8_0.A7.t3 25.395
R27390 OR8_0.NOT8_0.A7.n5 OR8_0.NOT8_0.A7.t2 25.395
R27391 OR8_0.NOT8_0.A7.n6 OR8_0.NOT8_0.A7.t0 25.395
R27392 OR8_0.NOT8_0.A7.n6 OR8_0.NOT8_0.A7.t4 25.395
R27393 OR8_0.NOT8_0.A7.n1 OR8_0.NOT8_0.A7.t5 19.8005
R27394 OR8_0.NOT8_0.A7.n1 OR8_0.NOT8_0.A7.t6 19.8005
R27395 OR8_0.NOT8_0.A7 OR8_0.NOT8_0.A7.n3 1.19417
R27396 OR8_0.NOT8_0.A7 OR8_0.NOT8_0.A7.n0 0.355237
R27397 OR8_0.NOT8_0.A7 OR8_0.NOT8_0.A7.n4 0.285715
R27398 a_7548_n35462.t0 a_7548_n35462.t1 9.9005
R27399 a_8496_n12822.t0 a_8496_n12822.t1 9.9005
R27400 a_8592_n12822.t0 a_8592_n12822.t1 9.9005
R27401 a_n24162_n6019.t0 a_n24162_n6019.t1 19.8005
R27402 AND8_0.S5.n1 AND8_0.S5.t4 1032.02
R27403 AND8_0.S5.n1 AND8_0.S5.t5 336.962
R27404 AND8_0.S5.n1 AND8_0.S5.t6 326.154
R27405 AND8_0.S5.n0 AND8_0.S5.t1 256.514
R27406 AND8_0.S5.n0 AND8_0.S5.n2 226.258
R27407 AND8_0.S5 AND8_0.S5.n1 162.945
R27408 AND8_0.S5.n0 AND8_0.S5.t0 83.7172
R27409 AND8_0.S5.n2 AND8_0.S5.t2 30.379
R27410 AND8_0.S5.n2 AND8_0.S5.t3 30.379
R27411 AND8_0.S5 AND8_0.S5.n0 1.92901
R27412 a_10267_n12821.t0 a_10267_n12821.t1 9.9005
R27413 a_10363_n12821.t0 a_10363_n12821.t1 9.9005
R27414 a_1707_4914.n0 a_1707_4914.t2 539.788
R27415 a_1707_4914.n1 a_1707_4914.t7 531.496
R27416 a_1707_4914.n0 a_1707_4914.t5 490.034
R27417 a_1707_4914.n5 a_1707_4914.t0 283.788
R27418 a_1707_4914.t1 a_1707_4914.n5 205.489
R27419 a_1707_4914.n2 a_1707_4914.t6 182.625
R27420 a_1707_4914.n3 a_1707_4914.t4 179.054
R27421 a_1707_4914.n2 a_1707_4914.t3 139.78
R27422 a_1707_4914.n4 a_1707_4914.n3 101.368
R27423 a_1707_4914.n5 a_1707_4914.n4 77.9135
R27424 a_1707_4914.n4 a_1707_4914.n1 76.1557
R27425 a_1707_4914.n1 a_1707_4914.n0 8.29297
R27426 a_1707_4914.n3 a_1707_4914.n2 3.57087
R27427 AND8_0.S7.n1 AND8_0.S7.t6 1032.02
R27428 AND8_0.S7.n1 AND8_0.S7.t4 336.962
R27429 AND8_0.S7.n1 AND8_0.S7.t5 326.154
R27430 AND8_0.S7.n0 AND8_0.S7.t1 256.514
R27431 AND8_0.S7.n0 AND8_0.S7.n3 226.258
R27432 AND8_0.S7 AND8_0.S7.n1 162.945
R27433 AND8_0.S7 AND8_0.S7.n2 107.835
R27434 AND8_0.S7.n0 AND8_0.S7.t0 83.7172
R27435 AND8_0.S7.n3 AND8_0.S7.t2 30.379
R27436 AND8_0.S7.n3 AND8_0.S7.t3 30.379
R27437 AND8_0.S7.n2 AND8_0.S7 3.3505
R27438 AND8_0.S7 AND8_0.S7.n0 1.96507
R27439 AND8_0.S7.n2 AND8_0.S7 0.985794
R27440 mux8_5.NAND4F_4.Y.n6 mux8_5.NAND4F_4.Y.t11 1032.02
R27441 mux8_5.NAND4F_4.Y.n6 mux8_5.NAND4F_4.Y.t9 336.962
R27442 mux8_5.NAND4F_4.Y.n6 mux8_5.NAND4F_4.Y.t10 326.154
R27443 mux8_5.NAND4F_4.Y.n0 mux8_5.NAND4F_4.Y.n1 187.373
R27444 mux8_5.NAND4F_4.Y.n0 mux8_5.NAND4F_4.Y.n2 187.192
R27445 mux8_5.NAND4F_4.Y.n0 mux8_5.NAND4F_4.Y.n3 187.192
R27446 mux8_5.NAND4F_4.Y.n5 mux8_5.NAND4F_4.Y.n4 187.192
R27447 mux8_5.NAND4F_4.Y mux8_5.NAND4F_4.Y.n6 162.942
R27448 mux8_5.NAND4F_4.Y.n7 mux8_5.NAND4F_4.Y 24.5377
R27449 mux8_5.NAND4F_4.Y.n7 mux8_5.NAND4F_4.Y.t0 22.6141
R27450 mux8_5.NAND4F_4.Y.n1 mux8_5.NAND4F_4.Y.t6 20.1899
R27451 mux8_5.NAND4F_4.Y.n1 mux8_5.NAND4F_4.Y.t5 20.1899
R27452 mux8_5.NAND4F_4.Y.n2 mux8_5.NAND4F_4.Y.t7 20.1899
R27453 mux8_5.NAND4F_4.Y.n2 mux8_5.NAND4F_4.Y.t8 20.1899
R27454 mux8_5.NAND4F_4.Y.n3 mux8_5.NAND4F_4.Y.t4 20.1899
R27455 mux8_5.NAND4F_4.Y.n3 mux8_5.NAND4F_4.Y.t3 20.1899
R27456 mux8_5.NAND4F_4.Y.n4 mux8_5.NAND4F_4.Y.t2 20.1899
R27457 mux8_5.NAND4F_4.Y.n4 mux8_5.NAND4F_4.Y.t1 20.1899
R27458 mux8_5.NAND4F_4.Y mux8_5.NAND4F_4.Y.n7 0.894894
R27459 mux8_5.NAND4F_4.Y mux8_5.NAND4F_4.Y.n5 0.452586
R27460 mux8_5.NAND4F_4.Y.n5 mux8_5.NAND4F_4.Y.n0 0.358709
R27461 a_8400_n11894.t0 a_8400_n11894.t1 9.9005
R27462 a_n12616_1406.n2 a_n12616_1406.n0 121.353
R27463 a_n12616_1406.n3 a_n12616_1406.n2 121.353
R27464 a_n12616_1406.n2 a_n12616_1406.n1 121.001
R27465 a_n12616_1406.n1 a_n12616_1406.t3 30.462
R27466 a_n12616_1406.n1 a_n12616_1406.t1 30.462
R27467 a_n12616_1406.n0 a_n12616_1406.t4 30.462
R27468 a_n12616_1406.n0 a_n12616_1406.t5 30.462
R27469 a_n12616_1406.t2 a_n12616_1406.n3 30.462
R27470 a_n12616_1406.n3 a_n12616_1406.t0 30.462
R27471 a_n12416_n11063.n1 a_n12416_n11063.n6 81.2978
R27472 a_n12416_n11063.n1 a_n12416_n11063.n5 81.1637
R27473 a_n12416_n11063.n0 a_n12416_n11063.n4 81.1637
R27474 a_n12416_n11063.n0 a_n12416_n11063.n3 81.1637
R27475 a_n12416_n11063.n7 a_n12416_n11063.n1 81.1637
R27476 a_n12416_n11063.n0 a_n12416_n11063.n2 80.9213
R27477 a_n12416_n11063.n6 a_n12416_n11063.t6 11.8205
R27478 a_n12416_n11063.n6 a_n12416_n11063.t7 11.8205
R27479 a_n12416_n11063.n5 a_n12416_n11063.t1 11.8205
R27480 a_n12416_n11063.n5 a_n12416_n11063.t0 11.8205
R27481 a_n12416_n11063.n4 a_n12416_n11063.t4 11.8205
R27482 a_n12416_n11063.n4 a_n12416_n11063.t5 11.8205
R27483 a_n12416_n11063.n3 a_n12416_n11063.t11 11.8205
R27484 a_n12416_n11063.n3 a_n12416_n11063.t3 11.8205
R27485 a_n12416_n11063.n2 a_n12416_n11063.t9 11.8205
R27486 a_n12416_n11063.n2 a_n12416_n11063.t10 11.8205
R27487 a_n12416_n11063.t2 a_n12416_n11063.n7 11.8205
R27488 a_n12416_n11063.n7 a_n12416_n11063.t8 11.8205
R27489 a_n12416_n11063.n1 a_n12416_n11063.n0 0.402735
R27490 a_n23990_n20027.t0 a_n23990_n20027.t1 19.8005
R27491 left_shifter_0.S3.n1 left_shifter_0.S3.t4 1032.02
R27492 left_shifter_0.S3.n1 left_shifter_0.S3.t5 336.962
R27493 left_shifter_0.S3.n1 left_shifter_0.S3.t6 326.154
R27494 left_shifter_0.S3.n0 left_shifter_0.S3.t3 256.89
R27495 left_shifter_0.S3.n0 left_shifter_0.S3.n2 226.635
R27496 mux8_4.NAND4F_5.A left_shifter_0.S3.n1 162.952
R27497 left_shifter_0.S3.n0 left_shifter_0.S3.t0 83.7172
R27498 left_shifter_0.S3.n2 left_shifter_0.S3.t1 30.379
R27499 left_shifter_0.S3.n2 left_shifter_0.S3.t2 30.379
R27500 mux8_4.A6 left_shifter_0.S3.n0 27.7494
R27501 mux8_4.A6 mux8_4.NAND4F_5.A 11.8717
R27502 a_n10108_n11683.n2 a_n10108_n11683.n0 121.353
R27503 a_n10108_n11683.n3 a_n10108_n11683.n2 121.353
R27504 a_n10108_n11683.n2 a_n10108_n11683.n1 121.001
R27505 a_n10108_n11683.n1 a_n10108_n11683.t5 30.462
R27506 a_n10108_n11683.n1 a_n10108_n11683.t1 30.462
R27507 a_n10108_n11683.n0 a_n10108_n11683.t3 30.462
R27508 a_n10108_n11683.n0 a_n10108_n11683.t4 30.462
R27509 a_n10108_n11683.t2 a_n10108_n11683.n3 30.462
R27510 a_n10108_n11683.n3 a_n10108_n11683.t0 30.462
R27511 a_n2744_1406.n2 a_n2744_1406.n0 121.353
R27512 a_n2744_1406.n3 a_n2744_1406.n2 121.353
R27513 a_n2744_1406.n2 a_n2744_1406.n1 121.001
R27514 a_n2744_1406.n1 a_n2744_1406.t5 30.462
R27515 a_n2744_1406.n1 a_n2744_1406.t0 30.462
R27516 a_n2744_1406.n0 a_n2744_1406.t3 30.462
R27517 a_n2744_1406.n0 a_n2744_1406.t4 30.462
R27518 a_n2744_1406.n3 a_n2744_1406.t1 30.462
R27519 a_n2744_1406.t2 a_n2744_1406.n3 30.462
R27520 MULT_0.4bit_ADDER_2.B1.n4 MULT_0.4bit_ADDER_2.B1.t23 491.64
R27521 MULT_0.4bit_ADDER_2.B1.n5 MULT_0.4bit_ADDER_2.B1.t17 491.64
R27522 MULT_0.4bit_ADDER_2.B1.n6 MULT_0.4bit_ADDER_2.B1.t22 491.64
R27523 MULT_0.4bit_ADDER_2.B1.n7 MULT_0.4bit_ADDER_2.B1.t19 491.64
R27524 MULT_0.4bit_ADDER_2.B1.n2 MULT_0.4bit_ADDER_2.B1.t15 485.221
R27525 MULT_0.4bit_ADDER_2.B1.n0 MULT_0.4bit_ADDER_2.B1.t21 367.928
R27526 MULT_0.4bit_ADDER_2.B1.n8 MULT_0.4bit_ADDER_2.B1.t16 255.588
R27527 MULT_0.4bit_ADDER_2.B1.n1 MULT_0.4bit_ADDER_2.B1.t13 224.478
R27528 MULT_0.4bit_ADDER_2.B1.n0 MULT_0.4bit_ADDER_2.B1.t14 213.688
R27529 MULT_0.4bit_ADDER_2.B1.n4 MULT_0.4bit_ADDER_2.B1.n3 209.19
R27530 MULT_0.4bit_ADDER_2.B1.n3 MULT_0.4bit_ADDER_2.B1.t18 139.78
R27531 MULT_0.4bit_ADDER_2.B1.n3 MULT_0.4bit_ADDER_2.B1.t20 139.78
R27532 MULT_0.4bit_ADDER_2.B1.n3 MULT_0.4bit_ADDER_2.B1.t12 139.78
R27533 MULT_0.4bit_ADDER_2.B1.n12 MULT_0.4bit_ADDER_2.B1.n11 120.999
R27534 MULT_0.4bit_ADDER_2.B1.n12 MULT_0.4bit_ADDER_2.B1.n10 120.999
R27535 MULT_0.4bit_ADDER_2.B1.n24 MULT_0.4bit_ADDER_2.B1.n23 104.489
R27536 MULT_0.4bit_ADDER_2.B1.n9 MULT_0.4bit_ADDER_2.B1 103.258
R27537 MULT_0.4bit_ADDER_2.B1.n14 MULT_0.4bit_ADDER_2.B1.n13 92.5005
R27538 MULT_0.4bit_ADDER_2.B1.n21 MULT_0.4bit_ADDER_2.B1.n19 86.2638
R27539 MULT_0.4bit_ADDER_2.B1.n19 MULT_0.4bit_ADDER_2.B1.n18 85.8873
R27540 MULT_0.4bit_ADDER_2.B1.n19 MULT_0.4bit_ADDER_2.B1.n16 85.724
R27541 MULT_0.4bit_ADDER_2.B1.n2 MULT_0.4bit_ADDER_2.B1.n1 84.5046
R27542 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_2.B1.n24 83.8907
R27543 MULT_0.4bit_ADDER_2.B1.n22 MULT_0.4bit_ADDER_2.B1.n21 75.0672
R27544 MULT_0.4bit_ADDER_2.B1.n22 MULT_0.4bit_ADDER_2.B1.n18 75.0672
R27545 MULT_0.4bit_ADDER_2.B1.n21 MULT_0.4bit_ADDER_2.B1.n20 73.1255
R27546 MULT_0.4bit_ADDER_2.B1.n18 MULT_0.4bit_ADDER_2.B1.n17 73.1255
R27547 MULT_0.4bit_ADDER_2.B1.n16 MULT_0.4bit_ADDER_2.B1.n15 73.1255
R27548 MULT_0.4bit_ADDER_2.B1.n1 MULT_0.4bit_ADDER_2.B1.n0 72.3005
R27549 MULT_0.4bit_ADDER_2.B1.n23 MULT_0.4bit_ADDER_2.B1.n16 68.8946
R27550 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_2.B1.n2 60.9816
R27551 MULT_0.4bit_ADDER_2.B1.n24 MULT_0.4bit_ADDER_2.B1.n14 41.9827
R27552 MULT_0.4bit_ADDER_2.B1.n13 MULT_0.4bit_ADDER_2.B1.t0 30.462
R27553 MULT_0.4bit_ADDER_2.B1.n13 MULT_0.4bit_ADDER_2.B1.t3 30.462
R27554 MULT_0.4bit_ADDER_2.B1.n11 MULT_0.4bit_ADDER_2.B1.t4 30.462
R27555 MULT_0.4bit_ADDER_2.B1.n11 MULT_0.4bit_ADDER_2.B1.t6 30.462
R27556 MULT_0.4bit_ADDER_2.B1.n10 MULT_0.4bit_ADDER_2.B1.t1 30.462
R27557 MULT_0.4bit_ADDER_2.B1.n10 MULT_0.4bit_ADDER_2.B1.t2 30.462
R27558 MULT_0.4bit_ADDER_2.B1.n14 MULT_0.4bit_ADDER_2.B1.n12 28.124
R27559 MULT_0.4bit_ADDER_2.B1.n5 MULT_0.4bit_ADDER_2.B1.n4 17.8661
R27560 MULT_0.4bit_ADDER_2.B1.n6 MULT_0.4bit_ADDER_2.B1.n5 17.8661
R27561 MULT_0.4bit_ADDER_2.B1.n7 MULT_0.4bit_ADDER_2.B1.n6 17.1217
R27562 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_2.B1.n8 15.6329
R27563 MULT_0.4bit_ADDER_2.B1.n17 MULT_0.4bit_ADDER_2.B1.t10 11.8205
R27564 MULT_0.4bit_ADDER_2.B1.n17 MULT_0.4bit_ADDER_2.B1.t11 11.8205
R27565 MULT_0.4bit_ADDER_2.B1.n20 MULT_0.4bit_ADDER_2.B1.t7 11.8205
R27566 MULT_0.4bit_ADDER_2.B1.n20 MULT_0.4bit_ADDER_2.B1.t8 11.8205
R27567 MULT_0.4bit_ADDER_2.B1.n15 MULT_0.4bit_ADDER_2.B1.t9 11.8205
R27568 MULT_0.4bit_ADDER_2.B1.n15 MULT_0.4bit_ADDER_2.B1.t5 11.8205
R27569 MULT_0.4bit_ADDER_2.B1.n9 MULT_0.4bit_ADDER_2.B1 10.8165
R27570 MULT_0.4bit_ADDER_2.B1.n23 MULT_0.4bit_ADDER_2.B1.n22 9.3005
R27571 MULT_0.4bit_ADDER_2.B1.n8 MULT_0.4bit_ADDER_2.B1.n7 1.8615
R27572 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_2.B1.n9 0.831812
R27573 a_9528_n11894.t0 a_9528_n11894.t1 9.9005
R27574 a_n3509_373.t0 a_n3509_373.t1 19.8005
R27575 a_7548_1690.t0 a_7548_1690.t1 9.9005
R27576 a_7644_1690.t0 a_7644_1690.t1 9.9005
R27577 a_9336_n26406.t0 a_9336_n26406.t1 9.9005
R27578 a_9432_n26406.t0 a_9432_n26406.t1 9.9005
R27579 AND8_0.NOT8_0.A6.n2 AND8_0.NOT8_0.A6.t10 394.37
R27580 AND8_0.NOT8_0.A6.n1 AND8_0.NOT8_0.A6.t8 291.829
R27581 AND8_0.NOT8_0.A6.n1 AND8_0.NOT8_0.A6.t9 291.829
R27582 AND8_0.NOT8_0.A6.n0 AND8_0.NOT8_0.A6.n4 227.526
R27583 AND8_0.NOT8_0.A6.n0 AND8_0.NOT8_0.A6.n3 227.266
R27584 AND8_0.NOT8_0.A6.n0 AND8_0.NOT8_0.A6.n5 227.266
R27585 AND8_0.NOT8_0.A6.n1 AND8_0.NOT8_0.A6.t7 221.72
R27586 AND8_0.NOT8_0.A6.n2 AND8_0.NOT8_0.A6.n1 53.374
R27587 AND8_0.NOT8_0.A6.n0 AND8_0.NOT8_0.A6.t0 42.7747
R27588 AND8_0.NOT8_0.A6.n4 AND8_0.NOT8_0.A6.t5 30.379
R27589 AND8_0.NOT8_0.A6.n4 AND8_0.NOT8_0.A6.t4 30.379
R27590 AND8_0.NOT8_0.A6.n3 AND8_0.NOT8_0.A6.t2 30.379
R27591 AND8_0.NOT8_0.A6.n3 AND8_0.NOT8_0.A6.t1 30.379
R27592 AND8_0.NOT8_0.A6.n5 AND8_0.NOT8_0.A6.t3 30.379
R27593 AND8_0.NOT8_0.A6.n5 AND8_0.NOT8_0.A6.t6 30.379
R27594 AND8_0.NOT8_0.A6 AND8_0.NOT8_0.A6.n0 2.03296
R27595 AND8_0.NOT8_0.A6 AND8_0.NOT8_0.A6.n2 1.25939
R27596 left_shifter_0.S2.n1 left_shifter_0.S2.t6 1032.02
R27597 left_shifter_0.S2.n1 left_shifter_0.S2.t4 336.962
R27598 left_shifter_0.S2.n1 left_shifter_0.S2.t5 326.154
R27599 left_shifter_0.S2.n0 left_shifter_0.S2.t1 256.89
R27600 left_shifter_0.S2.n0 left_shifter_0.S2.n2 226.635
R27601 mux8_3.NAND4F_5.A left_shifter_0.S2.n1 162.952
R27602 left_shifter_0.S2.n0 left_shifter_0.S2.t0 83.7172
R27603 mux8_3.A6 left_shifter_0.S2.n0 36.2335
R27604 left_shifter_0.S2.n2 left_shifter_0.S2.t2 30.379
R27605 left_shifter_0.S2.n2 left_shifter_0.S2.t3 30.379
R27606 mux8_3.A6 mux8_3.NAND4F_5.A 11.8717
R27607 a_n18998_n11683.n3 a_n18998_n11683.n2 121.353
R27608 a_n18998_n11683.n2 a_n18998_n11683.n1 121.001
R27609 a_n18998_n11683.n2 a_n18998_n11683.n0 120.977
R27610 a_n18998_n11683.n1 a_n18998_n11683.t3 30.462
R27611 a_n18998_n11683.n1 a_n18998_n11683.t0 30.462
R27612 a_n18998_n11683.n0 a_n18998_n11683.t4 30.462
R27613 a_n18998_n11683.n0 a_n18998_n11683.t5 30.462
R27614 a_n18998_n11683.t2 a_n18998_n11683.n3 30.462
R27615 a_n18998_n11683.n3 a_n18998_n11683.t1 30.462
R27616 OR8_0.NOT8_0.A2.n3 OR8_0.NOT8_0.A2.t10 394.37
R27617 OR8_0.NOT8_0.A2.n2 OR8_0.NOT8_0.A2.t9 291.829
R27618 OR8_0.NOT8_0.A2.n2 OR8_0.NOT8_0.A2.t7 291.829
R27619 OR8_0.NOT8_0.A2.n0 OR8_0.NOT8_0.A2.t3 256.425
R27620 OR8_0.NOT8_0.A2.n0 OR8_0.NOT8_0.A2.n5 231.24
R27621 OR8_0.NOT8_0.A2.n0 OR8_0.NOT8_0.A2.n6 231.03
R27622 OR8_0.NOT8_0.A2.n2 OR8_0.NOT8_0.A2.t8 221.72
R27623 OR8_0.NOT8_0.A2.n4 OR8_0.NOT8_0.A2.n1 66.4681
R27624 OR8_0.NOT8_0.A2.n3 OR8_0.NOT8_0.A2.n2 53.374
R27625 OR8_0.NOT8_0.A2.n4 OR8_0.NOT8_0.A2 32.5766
R27626 OR8_0.NOT8_0.A2.n6 OR8_0.NOT8_0.A2.t2 25.395
R27627 OR8_0.NOT8_0.A2.n6 OR8_0.NOT8_0.A2.t1 25.395
R27628 OR8_0.NOT8_0.A2.n5 OR8_0.NOT8_0.A2.t0 25.395
R27629 OR8_0.NOT8_0.A2.n5 OR8_0.NOT8_0.A2.t4 25.395
R27630 OR8_0.NOT8_0.A2.n1 OR8_0.NOT8_0.A2.t5 19.8005
R27631 OR8_0.NOT8_0.A2.n1 OR8_0.NOT8_0.A2.t6 19.8005
R27632 OR8_0.NOT8_0.A2 OR8_0.NOT8_0.A2.n3 1.27919
R27633 OR8_0.NOT8_0.A2 OR8_0.NOT8_0.A2.n0 0.355237
R27634 OR8_0.NOT8_0.A2 OR8_0.NOT8_0.A2.n4 0.293873
R27635 OR8_0.S2.n1 OR8_0.S2.t5 1032.02
R27636 OR8_0.S2.n1 OR8_0.S2.t4 336.962
R27637 OR8_0.S2.n1 OR8_0.S2.t6 326.154
R27638 OR8_0.S2.n0 OR8_0.S2.t1 256.514
R27639 OR8_0.S2.n0 OR8_0.S2.n2 226.258
R27640 OR8_0.S2 OR8_0.S2.n1 162.952
R27641 OR8_0.S2.n0 OR8_0.S2.t0 83.7172
R27642 OR8_0.S2.n2 OR8_0.S2.t2 30.379
R27643 OR8_0.S2.n2 OR8_0.S2.t3 30.379
R27644 OR8_0.S2 OR8_0.S2.n0 1.9182
R27645 a_n15896_n9452.t0 a_n15896_n9452.t1 19.8005
R27646 a_n11199_373.t0 a_n11199_373.t1 19.8005
R27647 mux8_8.NAND4F_2.Y.n6 mux8_8.NAND4F_2.Y.t11 933.563
R27648 mux8_8.NAND4F_2.Y.n6 mux8_8.NAND4F_2.Y.t9 367.635
R27649 mux8_8.NAND4F_2.Y.n7 mux8_8.NAND4F_2.Y.t10 308.481
R27650 mux8_8.NAND4F_2.Y.n0 mux8_8.NAND4F_2.Y.n1 187.373
R27651 mux8_8.NAND4F_2.Y.n0 mux8_8.NAND4F_2.Y.n2 187.192
R27652 mux8_8.NAND4F_2.Y.n0 mux8_8.NAND4F_2.Y.n3 187.192
R27653 mux8_8.NAND4F_2.Y.n5 mux8_8.NAND4F_2.Y.n4 187.192
R27654 mux8_8.NAND4F_2.Y mux8_8.NAND4F_2.Y.n7 162.102
R27655 mux8_8.NAND4F_2.Y.n8 mux8_8.NAND4F_2.Y.t8 22.7096
R27656 mux8_8.NAND4F_2.Y.n8 mux8_8.NAND4F_2.Y 22.4285
R27657 mux8_8.NAND4F_2.Y.n1 mux8_8.NAND4F_2.Y.t1 20.1899
R27658 mux8_8.NAND4F_2.Y.n1 mux8_8.NAND4F_2.Y.t0 20.1899
R27659 mux8_8.NAND4F_2.Y.n2 mux8_8.NAND4F_2.Y.t2 20.1899
R27660 mux8_8.NAND4F_2.Y.n2 mux8_8.NAND4F_2.Y.t3 20.1899
R27661 mux8_8.NAND4F_2.Y.n3 mux8_8.NAND4F_2.Y.t5 20.1899
R27662 mux8_8.NAND4F_2.Y.n3 mux8_8.NAND4F_2.Y.t4 20.1899
R27663 mux8_8.NAND4F_2.Y.n4 mux8_8.NAND4F_2.Y.t6 20.1899
R27664 mux8_8.NAND4F_2.Y.n4 mux8_8.NAND4F_2.Y.t7 20.1899
R27665 mux8_8.NAND4F_2.Y.n7 mux8_8.NAND4F_2.Y.n6 10.955
R27666 mux8_8.NAND4F_2.Y mux8_8.NAND4F_2.Y.n8 0.799394
R27667 mux8_8.NAND4F_2.Y mux8_8.NAND4F_2.Y.n5 0.452586
R27668 mux8_8.NAND4F_2.Y.n5 mux8_8.NAND4F_2.Y.n0 0.358709
R27669 a_5017_4912.n0 a_5017_4912.t2 539.788
R27670 a_5017_4912.n1 a_5017_4912.t7 531.496
R27671 a_5017_4912.n0 a_5017_4912.t5 490.034
R27672 a_5017_4912.n5 a_5017_4912.t0 283.788
R27673 a_5017_4912.t1 a_5017_4912.n5 205.489
R27674 a_5017_4912.n2 a_5017_4912.t6 182.625
R27675 a_5017_4912.n3 a_5017_4912.t4 179.054
R27676 a_5017_4912.n2 a_5017_4912.t3 139.78
R27677 a_5017_4912.n4 a_5017_4912.n3 101.368
R27678 a_5017_4912.n5 a_5017_4912.n4 77.9135
R27679 a_5017_4912.n4 a_5017_4912.n1 76.1557
R27680 a_5017_4912.n1 a_5017_4912.n0 8.29297
R27681 a_5017_4912.n3 a_5017_4912.n2 3.57087
R27682 mux8_3.NAND4F_1.Y.n2 mux8_3.NAND4F_1.Y.t9 978.795
R27683 mux8_3.NAND4F_1.Y.n1 mux8_3.NAND4F_1.Y.t10 308.481
R27684 mux8_3.NAND4F_1.Y.n1 mux8_3.NAND4F_1.Y.t11 308.481
R27685 mux8_3.NAND4F_1.Y.n0 mux8_3.NAND4F_1.Y.n3 187.373
R27686 mux8_3.NAND4F_1.Y.n0 mux8_3.NAND4F_1.Y.n4 187.192
R27687 mux8_3.NAND4F_1.Y.n0 mux8_3.NAND4F_1.Y.n5 187.192
R27688 mux8_3.NAND4F_1.Y.n7 mux8_3.NAND4F_1.Y.n6 187.192
R27689 mux8_3.NAND4F_1.Y mux8_3.NAND4F_1.Y.n2 161.84
R27690 mux8_3.NAND4F_1.Y mux8_3.NAND4F_1.Y.t2 23.4335
R27691 mux8_3.NAND4F_1.Y.n3 mux8_3.NAND4F_1.Y.t1 20.1899
R27692 mux8_3.NAND4F_1.Y.n3 mux8_3.NAND4F_1.Y.t0 20.1899
R27693 mux8_3.NAND4F_1.Y.n4 mux8_3.NAND4F_1.Y.t8 20.1899
R27694 mux8_3.NAND4F_1.Y.n4 mux8_3.NAND4F_1.Y.t7 20.1899
R27695 mux8_3.NAND4F_1.Y.n5 mux8_3.NAND4F_1.Y.t6 20.1899
R27696 mux8_3.NAND4F_1.Y.n5 mux8_3.NAND4F_1.Y.t5 20.1899
R27697 mux8_3.NAND4F_1.Y.n6 mux8_3.NAND4F_1.Y.t3 20.1899
R27698 mux8_3.NAND4F_1.Y.n6 mux8_3.NAND4F_1.Y.t4 20.1899
R27699 mux8_3.NAND4F_1.Y.n2 mux8_3.NAND4F_1.Y.n1 11.0463
R27700 mux8_3.NAND4F_1.Y mux8_3.NAND4F_1.Y.n7 0.527586
R27701 mux8_3.NAND4F_1.Y.n7 mux8_3.NAND4F_1.Y.n0 0.358709
R27702 a_11194_n12822.t0 a_11194_n12822.t1 9.9005
R27703 a_11290_n12822.t0 a_11290_n12822.t1 9.9005
R27704 a_8400_n34534.t0 a_8400_n34534.t1 9.9005
R27705 a_n17266_n4534.n0 a_n17266_n4534.n2 81.2978
R27706 a_n17266_n4534.n0 a_n17266_n4534.n3 81.1637
R27707 a_n17266_n4534.n0 a_n17266_n4534.n4 81.1637
R27708 a_n17266_n4534.n1 a_n17266_n4534.n5 81.1637
R27709 a_n17266_n4534.n1 a_n17266_n4534.n6 81.1637
R27710 a_n17266_n4534.n7 a_n17266_n4534.n1 80.9213
R27711 a_n17266_n4534.n2 a_n17266_n4534.t4 11.8205
R27712 a_n17266_n4534.n2 a_n17266_n4534.t3 11.8205
R27713 a_n17266_n4534.n3 a_n17266_n4534.t6 11.8205
R27714 a_n17266_n4534.n3 a_n17266_n4534.t5 11.8205
R27715 a_n17266_n4534.n4 a_n17266_n4534.t8 11.8205
R27716 a_n17266_n4534.n4 a_n17266_n4534.t7 11.8205
R27717 a_n17266_n4534.n5 a_n17266_n4534.t11 11.8205
R27718 a_n17266_n4534.n5 a_n17266_n4534.t9 11.8205
R27719 a_n17266_n4534.n6 a_n17266_n4534.t0 11.8205
R27720 a_n17266_n4534.n6 a_n17266_n4534.t10 11.8205
R27721 a_n17266_n4534.t2 a_n17266_n4534.n7 11.8205
R27722 a_n17266_n4534.n7 a_n17266_n4534.t1 11.8205
R27723 a_n17266_n4534.n1 a_n17266_n4534.n0 0.402735
R27724 a_n218_373.t0 a_n218_373.t1 19.8005
R27725 a_n12345_n20814.n2 a_n12345_n20814.t6 539.788
R27726 a_n12345_n20814.n3 a_n12345_n20814.t2 531.496
R27727 a_n12345_n20814.n2 a_n12345_n20814.t7 490.034
R27728 a_n12345_n20814.n5 a_n12345_n20814.t0 283.788
R27729 a_n12345_n20814.t1 a_n12345_n20814.n5 205.489
R27730 a_n12345_n20814.n0 a_n12345_n20814.t3 182.625
R27731 a_n12345_n20814.n1 a_n12345_n20814.t5 179.054
R27732 a_n12345_n20814.n0 a_n12345_n20814.t4 139.78
R27733 a_n12345_n20814.n4 a_n12345_n20814.n1 101.368
R27734 a_n12345_n20814.n5 a_n12345_n20814.n4 77.9135
R27735 a_n12345_n20814.n4 a_n12345_n20814.n3 76.1557
R27736 a_n12345_n20814.n3 a_n12345_n20814.n2 8.29297
R27737 a_n12345_n20814.n1 a_n12345_n20814.n0 3.57087
R27738 a_5197_4912.n2 a_5197_4912.n0 121.353
R27739 a_5197_4912.n2 a_5197_4912.n1 121.001
R27740 a_5197_4912.n3 a_5197_4912.n2 120.977
R27741 a_5197_4912.n0 a_5197_4912.t5 30.462
R27742 a_5197_4912.n0 a_5197_4912.t4 30.462
R27743 a_5197_4912.n1 a_5197_4912.t1 30.462
R27744 a_5197_4912.n1 a_5197_4912.t3 30.462
R27745 a_5197_4912.n3 a_5197_4912.t0 30.462
R27746 a_5197_4912.t2 a_5197_4912.n3 30.462
R27747 a_9432_n7266.t0 a_9432_n7266.t1 9.9005
R27748 a_9528_n34534.t0 a_9528_n34534.t1 9.9005
R27749 a_10459_n17349.t0 a_10459_n17349.t1 9.9005
R27750 a_9336_n35462.t0 a_9336_n35462.t1 9.9005
R27751 a_9432_n35462.t0 a_9432_n35462.t1 9.9005
R27752 a_4069_4914.n2 a_4069_4914.n1 121.353
R27753 a_4069_4914.n2 a_4069_4914.n0 121.353
R27754 a_4069_4914.n3 a_4069_4914.n2 121.001
R27755 a_4069_4914.n1 a_4069_4914.t1 30.462
R27756 a_4069_4914.n1 a_4069_4914.t0 30.462
R27757 a_4069_4914.n0 a_4069_4914.t5 30.462
R27758 a_4069_4914.n0 a_4069_4914.t4 30.462
R27759 a_4069_4914.n3 a_4069_4914.t3 30.462
R27760 a_4069_4914.t2 a_4069_4914.n3 30.462
R27761 a_n13714_n9452.t0 a_n13714_n9452.t1 19.8005
R27762 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t10 485.221
R27763 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t8 367.928
R27764 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n4 227.526
R27765 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n5 227.266
R27766 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n6 227.266
R27767 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t9 224.478
R27768 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t7 213.688
R27769 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n2 84.5046
R27770 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n1 72.3005
R27771 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n3 61.0566
R27772 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t0 42.7747
R27773 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t5 30.379
R27774 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t6 30.379
R27775 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t2 30.379
R27776 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t4 30.379
R27777 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t3 30.379
R27778 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.t1 30.379
R27779 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A.n0 0.583137
R27780 a_n14175_1406.n2 a_n14175_1406.n0 121.353
R27781 a_n14175_1406.n3 a_n14175_1406.n2 121.353
R27782 a_n14175_1406.n2 a_n14175_1406.n1 121.001
R27783 a_n14175_1406.n0 a_n14175_1406.t4 30.462
R27784 a_n14175_1406.n0 a_n14175_1406.t5 30.462
R27785 a_n14175_1406.n1 a_n14175_1406.t0 30.462
R27786 a_n14175_1406.n1 a_n14175_1406.t3 30.462
R27787 a_n14175_1406.n3 a_n14175_1406.t1 30.462
R27788 a_n14175_1406.t2 a_n14175_1406.n3 30.462
R27789 mux8_4.NAND4F_3.Y.n7 mux8_4.NAND4F_3.Y.t9 978.795
R27790 mux8_4.NAND4F_3.Y.n6 mux8_4.NAND4F_3.Y.t11 308.481
R27791 mux8_4.NAND4F_3.Y.n6 mux8_4.NAND4F_3.Y.t10 308.481
R27792 mux8_4.NAND4F_3.Y.n0 mux8_4.NAND4F_3.Y.n1 187.373
R27793 mux8_4.NAND4F_3.Y.n0 mux8_4.NAND4F_3.Y.n2 187.192
R27794 mux8_4.NAND4F_3.Y.n0 mux8_4.NAND4F_3.Y.n3 187.192
R27795 mux8_4.NAND4F_3.Y.n5 mux8_4.NAND4F_3.Y.n4 187.192
R27796 mux8_4.NAND4F_3.Y mux8_4.NAND4F_3.Y.n7 161.839
R27797 mux8_4.NAND4F_3.Y mux8_4.NAND4F_3.Y.t6 23.4426
R27798 mux8_4.NAND4F_3.Y.n1 mux8_4.NAND4F_3.Y.t1 20.1899
R27799 mux8_4.NAND4F_3.Y.n1 mux8_4.NAND4F_3.Y.t0 20.1899
R27800 mux8_4.NAND4F_3.Y.n2 mux8_4.NAND4F_3.Y.t3 20.1899
R27801 mux8_4.NAND4F_3.Y.n2 mux8_4.NAND4F_3.Y.t2 20.1899
R27802 mux8_4.NAND4F_3.Y.n3 mux8_4.NAND4F_3.Y.t5 20.1899
R27803 mux8_4.NAND4F_3.Y.n3 mux8_4.NAND4F_3.Y.t4 20.1899
R27804 mux8_4.NAND4F_3.Y.n4 mux8_4.NAND4F_3.Y.t8 20.1899
R27805 mux8_4.NAND4F_3.Y.n4 mux8_4.NAND4F_3.Y.t7 20.1899
R27806 mux8_4.NAND4F_3.Y.n7 mux8_4.NAND4F_3.Y.n6 11.0463
R27807 mux8_4.NAND4F_3.Y mux8_4.NAND4F_3.Y.n5 0.518495
R27808 mux8_4.NAND4F_3.Y.n5 mux8_4.NAND4F_3.Y.n0 0.358709
R27809 a_n4303_1406.n2 a_n4303_1406.n1 121.353
R27810 a_n4303_1406.n2 a_n4303_1406.n0 121.353
R27811 a_n4303_1406.n3 a_n4303_1406.n2 121.001
R27812 a_n4303_1406.n1 a_n4303_1406.t0 30.462
R27813 a_n4303_1406.n1 a_n4303_1406.t1 30.462
R27814 a_n4303_1406.n0 a_n4303_1406.t3 30.462
R27815 a_n4303_1406.n0 a_n4303_1406.t5 30.462
R27816 a_n4303_1406.n3 a_n4303_1406.t4 30.462
R27817 a_n4303_1406.t2 a_n4303_1406.n3 30.462
R27818 a_n4618_373.t0 a_n4618_373.t1 19.8005
R27819 mux8_8.NAND4F_8.Y.n1 mux8_8.NAND4F_8.Y.t13 379.173
R27820 mux8_8.NAND4F_8.Y.n2 mux8_8.NAND4F_8.Y.t12 312.599
R27821 mux8_8.NAND4F_8.Y.n1 mux8_8.NAND4F_8.Y.t14 247.428
R27822 mux8_8.NAND4F_8.Y.n4 mux8_8.NAND4F_8.Y.t9 247.428
R27823 mux8_8.NAND4F_8.Y.n3 mux8_8.NAND4F_8.Y.t11 247.428
R27824 mux8_8.NAND4F_8.Y.n2 mux8_8.NAND4F_8.Y.t10 247.428
R27825 mux8_8.NAND4F_8.Y.n0 mux8_8.NAND4F_8.Y.n6 187.373
R27826 mux8_8.NAND4F_8.Y.n0 mux8_8.NAND4F_8.Y.n7 187.192
R27827 mux8_8.NAND4F_8.Y.n0 mux8_8.NAND4F_8.Y.n8 187.192
R27828 mux8_8.NAND4F_8.Y.n10 mux8_8.NAND4F_8.Y.n9 187.192
R27829 mux8_8.NAND4F_8.Y mux8_8.NAND4F_8.Y.n5 162.139
R27830 mux8_8.NAND4F_8.Y.n4 mux8_8.NAND4F_8.Y.n3 65.1723
R27831 mux8_8.NAND4F_8.Y.n3 mux8_8.NAND4F_8.Y.n2 65.1723
R27832 mux8_8.NAND4F_8.Y.n5 mux8_8.NAND4F_8.Y.n4 33.2653
R27833 mux8_8.NAND4F_8.Y.n5 mux8_8.NAND4F_8.Y.n1 31.9075
R27834 mux8_8.NAND4F_8.Y mux8_8.NAND4F_8.Y.t6 22.6141
R27835 mux8_8.NAND4F_8.Y.n6 mux8_8.NAND4F_8.Y.t2 20.1899
R27836 mux8_8.NAND4F_8.Y.n6 mux8_8.NAND4F_8.Y.t3 20.1899
R27837 mux8_8.NAND4F_8.Y.n7 mux8_8.NAND4F_8.Y.t1 20.1899
R27838 mux8_8.NAND4F_8.Y.n7 mux8_8.NAND4F_8.Y.t0 20.1899
R27839 mux8_8.NAND4F_8.Y.n8 mux8_8.NAND4F_8.Y.t5 20.1899
R27840 mux8_8.NAND4F_8.Y.n8 mux8_8.NAND4F_8.Y.t4 20.1899
R27841 mux8_8.NAND4F_8.Y.n9 mux8_8.NAND4F_8.Y.t8 20.1899
R27842 mux8_8.NAND4F_8.Y.n9 mux8_8.NAND4F_8.Y.t7 20.1899
R27843 mux8_8.NAND4F_8.Y mux8_8.NAND4F_8.Y.n10 0.452586
R27844 mux8_8.NAND4F_8.Y.n10 mux8_8.NAND4F_8.Y.n0 0.358709
R27845 a_7452_n26406.t0 a_7452_n26406.t1 9.9005
R27846 a_8400_n7266.t0 a_8400_n7266.t1 9.9005
R27847 a_n1094_3190.n2 a_n1094_3190.t7 541.395
R27848 a_n1094_3190.n3 a_n1094_3190.t2 527.402
R27849 a_n1094_3190.n2 a_n1094_3190.t5 491.64
R27850 a_n1094_3190.n5 a_n1094_3190.t0 281.906
R27851 a_n1094_3190.t1 a_n1094_3190.n5 204.359
R27852 a_n1094_3190.n0 a_n1094_3190.t6 180.73
R27853 a_n1094_3190.n1 a_n1094_3190.t4 179.45
R27854 a_n1094_3190.n0 a_n1094_3190.t3 139.78
R27855 a_n1094_3190.n4 a_n1094_3190.n1 105.635
R27856 a_n1094_3190.n4 a_n1094_3190.n3 76.0005
R27857 a_n1094_3190.n5 a_n1094_3190.n4 67.9685
R27858 a_n1094_3190.n3 a_n1094_3190.n2 13.994
R27859 a_n1094_3190.n1 a_n1094_3190.n0 1.28015
R27860 a_10363_n16422.t0 a_10363_n16422.t1 9.9005
R27861 a_n11276_n33705.n2 a_n11276_n33705.n0 121.353
R27862 a_n11276_n33705.n3 a_n11276_n33705.n2 121.353
R27863 a_n11276_n33705.n2 a_n11276_n33705.n1 121.001
R27864 a_n11276_n33705.n1 a_n11276_n33705.t0 30.462
R27865 a_n11276_n33705.n1 a_n11276_n33705.t4 30.462
R27866 a_n11276_n33705.n0 a_n11276_n33705.t3 30.462
R27867 a_n11276_n33705.n0 a_n11276_n33705.t5 30.462
R27868 a_n11276_n33705.t2 a_n11276_n33705.n3 30.462
R27869 a_n11276_n33705.n3 a_n11276_n33705.t1 30.462
R27870 a_8496_n20950.t0 a_8496_n20950.t1 9.9005
R27871 a_8592_n20950.t0 a_8592_n20950.t1 9.9005
R27872 a_9528_n7266.t0 a_9528_n7266.t1 9.9005
R27873 ZFLAG_0.nor4_1.Y.n5 ZFLAG_0.nor4_1.Y.t8 540.38
R27874 ZFLAG_0.nor4_1.Y.n3 ZFLAG_0.nor4_1.Y.t7 367.928
R27875 ZFLAG_0.nor4_1.Y.n4 ZFLAG_0.nor4_1.Y.t10 227.356
R27876 ZFLAG_0.nor4_1.Y.n3 ZFLAG_0.nor4_1.Y.t9 213.688
R27877 ZFLAG_0.nor4_1.Y.n5 ZFLAG_0.nor4_1.Y.n4 160.439
R27878 ZFLAG_0.nor4_1.Y.n2 ZFLAG_0.nor4_1.Y.t0 148.181
R27879 ZFLAG_0.nor4_1.Y.n4 ZFLAG_0.nor4_1.Y.n3 94.4341
R27880 ZFLAG_0.nor4_1.Y.n8 ZFLAG_0.nor4_1.Y.n6 66.4372
R27881 ZFLAG_0.nor4_1.Y.n8 ZFLAG_0.nor4_1.Y.n7 66.3172
R27882 ZFLAG_0.nor4_1.Y.n6 ZFLAG_0.nor4_1.Y.t4 19.8005
R27883 ZFLAG_0.nor4_1.Y.n6 ZFLAG_0.nor4_1.Y.t5 19.8005
R27884 ZFLAG_0.nor4_1.Y.n7 ZFLAG_0.nor4_1.Y.t3 19.8005
R27885 ZFLAG_0.nor4_1.Y.n7 ZFLAG_0.nor4_1.Y.t6 19.8005
R27886 ZFLAG_0.nor4_1.Y.n0 ZFLAG_0.nor4_1.Y.t2 7.59513
R27887 ZFLAG_0.nor4_1.Y.n0 ZFLAG_0.nor4_1.Y.t1 7.59513
R27888 ZFLAG_0.nor4_1.Y ZFLAG_0.nor4_1.Y.n5 0.900886
R27889 ZFLAG_0.nor4_1.Y.n1 ZFLAG_0.nor4_1.Y 0.673006
R27890 ZFLAG_0.nor4_1.Y ZFLAG_0.nor4_1.Y.n8 0.570877
R27891 ZFLAG_0.nor4_1.Y ZFLAG_0.nor4_1.Y.n2 0.0743902
R27892 ZFLAG_0.nor4_1.Y.n2 ZFLAG_0.nor4_1.Y.n1 0.00100956
R27893 ZFLAG_0.nor4_1.Y.n1 ZFLAG_0.nor4_1.Y.n0 140.589
R27894 a_7644_n7266.t0 a_7644_n7266.t1 9.9005
R27895 a_11386_n17350.t0 a_11386_n17350.t1 9.9005
R27896 a_7452_n35462.t0 a_7452_n35462.t1 9.9005
R27897 a_n11274_n28476.n2 a_n11274_n28476.n0 121.353
R27898 a_n11274_n28476.n3 a_n11274_n28476.n2 121.353
R27899 a_n11274_n28476.n2 a_n11274_n28476.n1 121.001
R27900 a_n11274_n28476.n0 a_n11274_n28476.t5 30.462
R27901 a_n11274_n28476.n0 a_n11274_n28476.t4 30.462
R27902 a_n11274_n28476.n1 a_n11274_n28476.t3 30.462
R27903 a_n11274_n28476.n1 a_n11274_n28476.t1 30.462
R27904 a_n11274_n28476.n3 a_n11274_n28476.t0 30.462
R27905 a_n11274_n28476.t2 a_n11274_n28476.n3 30.462
R27906 a_8400_n12822.t0 a_8400_n12822.t1 9.9005
R27907 a_7452_n30006.t0 a_7452_n30006.t1 9.9005
R27908 a_10459_n30933.t0 a_10459_n30933.t1 9.9005
R27909 a_n11274_n20496.n2 a_n11274_n20496.n0 121.353
R27910 a_n11274_n20496.n3 a_n11274_n20496.n2 121.353
R27911 a_n11274_n20496.n2 a_n11274_n20496.n1 121.001
R27912 a_n11274_n20496.n1 a_n11274_n20496.t1 30.462
R27913 a_n11274_n20496.n1 a_n11274_n20496.t5 30.462
R27914 a_n11274_n20496.n0 a_n11274_n20496.t4 30.462
R27915 a_n11274_n20496.n0 a_n11274_n20496.t3 30.462
R27916 a_n11274_n20496.n3 a_n11274_n20496.t0 30.462
R27917 a_n11274_n20496.t2 a_n11274_n20496.n3 30.462
R27918 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t8 540.38
R27919 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t10 367.928
R27920 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n5 227.526
R27921 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t7 227.356
R27922 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n4 227.266
R27923 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n6 227.266
R27924 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t9 213.688
R27925 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n2 160.439
R27926 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n1 94.4341
R27927 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t0 42.7944
R27928 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t5 30.379
R27929 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t6 30.379
R27930 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t2 30.379
R27931 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t1 30.379
R27932 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t3 30.379
R27933 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.t4 30.379
R27934 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n0 13.4358
R27935 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B.n3 0.821842
R27936 a_n15887_n8419.n0 a_n15887_n8419.t5 539.788
R27937 a_n15887_n8419.n1 a_n15887_n8419.t2 531.496
R27938 a_n15887_n8419.n0 a_n15887_n8419.t7 490.034
R27939 a_n15887_n8419.n5 a_n15887_n8419.t0 283.788
R27940 a_n15887_n8419.t1 a_n15887_n8419.n5 205.489
R27941 a_n15887_n8419.n2 a_n15887_n8419.t3 182.625
R27942 a_n15887_n8419.n3 a_n15887_n8419.t6 179.054
R27943 a_n15887_n8419.n2 a_n15887_n8419.t4 139.78
R27944 a_n15887_n8419.n4 a_n15887_n8419.n3 101.368
R27945 a_n15887_n8419.n5 a_n15887_n8419.n4 77.9135
R27946 a_n15887_n8419.n4 a_n15887_n8419.n1 76.1557
R27947 a_n15887_n8419.n1 a_n15887_n8419.n0 8.29297
R27948 a_n15887_n8419.n3 a_n15887_n8419.n2 3.57087
R27949 a_n15707_n7799.n1 a_n15707_n7799.n6 81.2978
R27950 a_n15707_n7799.n1 a_n15707_n7799.n5 81.1637
R27951 a_n15707_n7799.n0 a_n15707_n7799.n4 81.1637
R27952 a_n15707_n7799.n0 a_n15707_n7799.n3 81.1637
R27953 a_n15707_n7799.n7 a_n15707_n7799.n1 81.1637
R27954 a_n15707_n7799.n0 a_n15707_n7799.n2 80.9213
R27955 a_n15707_n7799.n6 a_n15707_n7799.t1 11.8205
R27956 a_n15707_n7799.n6 a_n15707_n7799.t0 11.8205
R27957 a_n15707_n7799.n5 a_n15707_n7799.t4 11.8205
R27958 a_n15707_n7799.n5 a_n15707_n7799.t3 11.8205
R27959 a_n15707_n7799.n4 a_n15707_n7799.t11 11.8205
R27960 a_n15707_n7799.n4 a_n15707_n7799.t9 11.8205
R27961 a_n15707_n7799.n3 a_n15707_n7799.t6 11.8205
R27962 a_n15707_n7799.n3 a_n15707_n7799.t10 11.8205
R27963 a_n15707_n7799.n2 a_n15707_n7799.t8 11.8205
R27964 a_n15707_n7799.n2 a_n15707_n7799.t7 11.8205
R27965 a_n15707_n7799.n7 a_n15707_n7799.t5 11.8205
R27966 a_n15707_n7799.t2 a_n15707_n7799.n7 11.8205
R27967 a_n15707_n7799.n1 a_n15707_n7799.n0 0.402735
R27968 mux8_4.inv_0.A.n1 mux8_4.inv_0.A.t9 291.829
R27969 mux8_4.inv_0.A.n1 mux8_4.inv_0.A.t7 291.829
R27970 mux8_4.inv_0.A.n0 mux8_4.inv_0.A.t3 256.425
R27971 mux8_4.inv_0.A.n0 mux8_4.inv_0.A.n2 231.24
R27972 mux8_4.inv_0.A.n0 mux8_4.inv_0.A.n3 231.03
R27973 mux8_4.inv_0.A.n1 mux8_4.inv_0.A.t10 221.72
R27974 mux8_4.inv_0.A.t8 mux8_4.inv_0.A.n0 393.959
R27975 mux8_4.inv_0.A.n4 mux8_4.inv_0.A.n0 66.6316
R27976 mux8_4.inv_0.A.n0 mux8_4.inv_0.A.n1 54.1444
R27977 mux8_4.inv_0.A.n2 mux8_4.inv_0.A.t5 25.395
R27978 mux8_4.inv_0.A.n2 mux8_4.inv_0.A.t4 25.395
R27979 mux8_4.inv_0.A.n3 mux8_4.inv_0.A.t2 25.395
R27980 mux8_4.inv_0.A.n3 mux8_4.inv_0.A.t1 25.395
R27981 mux8_4.inv_0.A.n4 mux8_4.inv_0.A.t6 19.8005
R27982 mux8_4.inv_0.A.n4 mux8_4.inv_0.A.t0 19.8005
R27983 a_11865_n16359.n1 a_11865_n16359.n4 231.24
R27984 a_11865_n16359.n0 a_11865_n16359.n2 231.24
R27985 a_11865_n16359.n1 a_11865_n16359.n5 231.03
R27986 a_11865_n16359.n0 a_11865_n16359.n3 231.03
R27987 a_11865_n16359.n6 a_11865_n16359.n1 231.03
R27988 a_11865_n16359.n4 a_11865_n16359.t4 25.395
R27989 a_11865_n16359.n4 a_11865_n16359.t1 25.395
R27990 a_11865_n16359.n5 a_11865_n16359.t3 25.395
R27991 a_11865_n16359.n5 a_11865_n16359.t0 25.395
R27992 a_11865_n16359.n3 a_11865_n16359.t5 25.395
R27993 a_11865_n16359.n3 a_11865_n16359.t9 25.395
R27994 a_11865_n16359.n2 a_11865_n16359.t7 25.395
R27995 a_11865_n16359.n2 a_11865_n16359.t6 25.395
R27996 a_11865_n16359.t8 a_11865_n16359.n6 25.395
R27997 a_11865_n16359.n6 a_11865_n16359.t2 25.395
R27998 a_11865_n16359.n1 a_11865_n16359.n0 0.421553
R27999 a_n17005_n6187.t0 a_n17005_n6187.t1 19.8005
R28000 a_n17296_n5180.n2 a_n17296_n5180.t2 541.395
R28001 a_n17296_n5180.n3 a_n17296_n5180.t6 527.402
R28002 a_n17296_n5180.n2 a_n17296_n5180.t7 491.64
R28003 a_n17296_n5180.n5 a_n17296_n5180.t0 281.906
R28004 a_n17296_n5180.t1 a_n17296_n5180.n5 204.359
R28005 a_n17296_n5180.n0 a_n17296_n5180.t3 180.73
R28006 a_n17296_n5180.n1 a_n17296_n5180.t5 179.45
R28007 a_n17296_n5180.n0 a_n17296_n5180.t4 139.78
R28008 a_n17296_n5180.n4 a_n17296_n5180.n1 105.635
R28009 a_n17296_n5180.n4 a_n17296_n5180.n3 76.0005
R28010 a_n17296_n5180.n5 a_n17296_n5180.n4 67.9685
R28011 a_n17296_n5180.n3 a_n17296_n5180.n2 13.994
R28012 a_n17296_n5180.n1 a_n17296_n5180.n0 1.28015
R28013 a_n8549_n8419.n2 a_n8549_n8419.n1 121.353
R28014 a_n8549_n8419.n2 a_n8549_n8419.n0 121.353
R28015 a_n8549_n8419.n3 a_n8549_n8419.n2 121.001
R28016 a_n8549_n8419.n1 a_n8549_n8419.t1 30.462
R28017 a_n8549_n8419.n1 a_n8549_n8419.t0 30.462
R28018 a_n8549_n8419.n0 a_n8549_n8419.t5 30.462
R28019 a_n8549_n8419.n0 a_n8549_n8419.t4 30.462
R28020 a_n8549_n8419.n3 a_n8549_n8419.t3 30.462
R28021 a_n8549_n8419.t2 a_n8549_n8419.n3 30.462
R28022 a_n59_1380.n2 a_n59_1380.t4 541.395
R28023 a_n59_1380.n3 a_n59_1380.t7 527.402
R28024 a_n59_1380.n2 a_n59_1380.t2 491.64
R28025 a_n59_1380.n5 a_n59_1380.t0 281.906
R28026 a_n59_1380.t1 a_n59_1380.n5 204.359
R28027 a_n59_1380.n0 a_n59_1380.t5 180.73
R28028 a_n59_1380.n1 a_n59_1380.t6 179.45
R28029 a_n59_1380.n0 a_n59_1380.t3 139.78
R28030 a_n59_1380.n4 a_n59_1380.n1 105.635
R28031 a_n59_1380.n4 a_n59_1380.n3 76.0005
R28032 a_n59_1380.n5 a_n59_1380.n4 67.9685
R28033 a_n59_1380.n3 a_n59_1380.n2 13.994
R28034 a_n59_1380.n1 a_n59_1380.n0 1.28015
R28035 NOT8_0.S1.n1 NOT8_0.S1.t5 1032.02
R28036 NOT8_0.S1.n1 NOT8_0.S1.t4 336.962
R28037 NOT8_0.S1.n1 NOT8_0.S1.t6 326.154
R28038 NOT8_0.S1.n0 NOT8_0.S1.t2 256.514
R28039 NOT8_0.S1.n0 NOT8_0.S1.n2 226.258
R28040 NOT8_0.S1 NOT8_0.S1.n1 162.952
R28041 NOT8_0.S1.n0 NOT8_0.S1.t0 83.7172
R28042 NOT8_0.S1.n2 NOT8_0.S1.t1 30.379
R28043 NOT8_0.S1.n2 NOT8_0.S1.t3 30.379
R28044 NOT8_0.S1 NOT8_0.S1.n0 1.89195
R28045 a_n11276_n14723.n2 a_n11276_n14723.n0 121.353
R28046 a_n11276_n14723.n3 a_n11276_n14723.n2 121.353
R28047 a_n11276_n14723.n2 a_n11276_n14723.n1 121.001
R28048 a_n11276_n14723.n1 a_n11276_n14723.t0 30.462
R28049 a_n11276_n14723.n1 a_n11276_n14723.t5 30.462
R28050 a_n11276_n14723.n0 a_n11276_n14723.t4 30.462
R28051 a_n11276_n14723.n0 a_n11276_n14723.t3 30.462
R28052 a_n11276_n14723.t2 a_n11276_n14723.n3 30.462
R28053 a_n11276_n14723.n3 a_n11276_n14723.t1 30.462
R28054 a_9432_n11894.t0 a_9432_n11894.t1 9.9005
R28055 a_n17266_n11063.n7 a_n17266_n11063.n1 81.2978
R28056 a_n17266_n11063.n1 a_n17266_n11063.n6 81.1637
R28057 a_n17266_n11063.n1 a_n17266_n11063.n5 81.1637
R28058 a_n17266_n11063.n0 a_n17266_n11063.n4 81.1637
R28059 a_n17266_n11063.n0 a_n17266_n11063.n3 81.1637
R28060 a_n17266_n11063.n0 a_n17266_n11063.n2 80.9213
R28061 a_n17266_n11063.n6 a_n17266_n11063.t4 11.8205
R28062 a_n17266_n11063.n6 a_n17266_n11063.t0 11.8205
R28063 a_n17266_n11063.n5 a_n17266_n11063.t3 11.8205
R28064 a_n17266_n11063.n5 a_n17266_n11063.t5 11.8205
R28065 a_n17266_n11063.n4 a_n17266_n11063.t8 11.8205
R28066 a_n17266_n11063.n4 a_n17266_n11063.t6 11.8205
R28067 a_n17266_n11063.n3 a_n17266_n11063.t11 11.8205
R28068 a_n17266_n11063.n3 a_n17266_n11063.t7 11.8205
R28069 a_n17266_n11063.n2 a_n17266_n11063.t9 11.8205
R28070 a_n17266_n11063.n2 a_n17266_n11063.t10 11.8205
R28071 a_n17266_n11063.n7 a_n17266_n11063.t1 11.8205
R28072 a_n17266_n11063.t2 a_n17266_n11063.n7 11.8205
R28073 a_n17266_n11063.n1 a_n17266_n11063.n0 0.402735
R28074 a_n19981_n11683.n2 a_n19981_n11683.n0 121.353
R28075 a_n19981_n11683.n3 a_n19981_n11683.n2 121.353
R28076 a_n19981_n11683.n2 a_n19981_n11683.n1 121.001
R28077 a_n19981_n11683.n1 a_n19981_n11683.t4 30.462
R28078 a_n19981_n11683.n1 a_n19981_n11683.t0 30.462
R28079 a_n19981_n11683.n0 a_n19981_n11683.t5 30.462
R28080 a_n19981_n11683.n0 a_n19981_n11683.t3 30.462
R28081 a_n19981_n11683.n3 a_n19981_n11683.t1 30.462
R28082 a_n19981_n11683.t2 a_n19981_n11683.n3 30.462
R28083 mux8_3.NAND4F_2.Y.n6 mux8_3.NAND4F_2.Y.t9 933.563
R28084 mux8_3.NAND4F_2.Y.n6 mux8_3.NAND4F_2.Y.t10 367.635
R28085 mux8_3.NAND4F_2.Y.n7 mux8_3.NAND4F_2.Y.t11 308.481
R28086 mux8_3.NAND4F_2.Y.n0 mux8_3.NAND4F_2.Y.n1 187.373
R28087 mux8_3.NAND4F_2.Y.n0 mux8_3.NAND4F_2.Y.n2 187.192
R28088 mux8_3.NAND4F_2.Y.n0 mux8_3.NAND4F_2.Y.n3 187.192
R28089 mux8_3.NAND4F_2.Y.n5 mux8_3.NAND4F_2.Y.n4 187.192
R28090 mux8_3.NAND4F_2.Y mux8_3.NAND4F_2.Y.n7 162.102
R28091 mux8_3.NAND4F_2.Y.n8 mux8_3.NAND4F_2.Y.t0 22.7096
R28092 mux8_3.NAND4F_2.Y.n8 mux8_3.NAND4F_2.Y 22.4285
R28093 mux8_3.NAND4F_2.Y.n1 mux8_3.NAND4F_2.Y.t4 20.1899
R28094 mux8_3.NAND4F_2.Y.n1 mux8_3.NAND4F_2.Y.t3 20.1899
R28095 mux8_3.NAND4F_2.Y.n2 mux8_3.NAND4F_2.Y.t5 20.1899
R28096 mux8_3.NAND4F_2.Y.n2 mux8_3.NAND4F_2.Y.t6 20.1899
R28097 mux8_3.NAND4F_2.Y.n3 mux8_3.NAND4F_2.Y.t8 20.1899
R28098 mux8_3.NAND4F_2.Y.n3 mux8_3.NAND4F_2.Y.t7 20.1899
R28099 mux8_3.NAND4F_2.Y.n4 mux8_3.NAND4F_2.Y.t2 20.1899
R28100 mux8_3.NAND4F_2.Y.n4 mux8_3.NAND4F_2.Y.t1 20.1899
R28101 mux8_3.NAND4F_2.Y.n7 mux8_3.NAND4F_2.Y.n6 10.955
R28102 mux8_3.NAND4F_2.Y mux8_3.NAND4F_2.Y.n8 0.799394
R28103 mux8_3.NAND4F_2.Y mux8_3.NAND4F_2.Y.n5 0.452586
R28104 mux8_3.NAND4F_2.Y.n5 mux8_3.NAND4F_2.Y.n0 0.358709
R28105 a_11194_n20950.t0 a_11194_n20950.t1 9.9005
R28106 a_11290_n20950.t0 a_11290_n20950.t1 9.9005
R28107 OR8_0.S6.n1 OR8_0.S6.t6 1032.02
R28108 OR8_0.S6.n1 OR8_0.S6.t4 336.962
R28109 OR8_0.S6.n1 OR8_0.S6.t5 326.154
R28110 OR8_0.S6.n0 OR8_0.S6.t2 256.514
R28111 OR8_0.S6.n0 OR8_0.S6.n2 226.258
R28112 mux8_8.NAND4F_2.A OR8_0.S6.n1 162.952
R28113 OR8_0.NOT8_0.S6 mux8_8.A3 85.08
R28114 OR8_0.S6.n0 OR8_0.S6.t0 83.7172
R28115 OR8_0.S6.n2 OR8_0.S6.t3 30.379
R28116 OR8_0.S6.n2 OR8_0.S6.t1 30.379
R28117 mux8_8.A3 mux8_8.NAND4F_2.A 14.0763
R28118 OR8_0.NOT8_0.S6 OR8_0.S6.n0 1.95466
R28119 a_n15131_n11683.n2 a_n15131_n11683.n0 121.353
R28120 a_n15131_n11683.n3 a_n15131_n11683.n2 121.353
R28121 a_n15131_n11683.n2 a_n15131_n11683.n1 121.001
R28122 a_n15131_n11683.n1 a_n15131_n11683.t5 30.462
R28123 a_n15131_n11683.n1 a_n15131_n11683.t0 30.462
R28124 a_n15131_n11683.n0 a_n15131_n11683.t3 30.462
R28125 a_n15131_n11683.n0 a_n15131_n11683.t4 30.462
R28126 a_n15131_n11683.n3 a_n15131_n11683.t1 30.462
R28127 a_n15131_n11683.t2 a_n15131_n11683.n3 30.462
R28128 a_8400_n8194.t0 a_8400_n8194.t1 9.9005
R28129 a_8496_n8194.t0 a_8496_n8194.t1 9.9005
R28130 a_11194_n8194.t0 a_11194_n8194.t1 9.9005
R28131 mux8_5.NAND4F_1.Y.n2 mux8_5.NAND4F_1.Y.t11 978.795
R28132 mux8_5.NAND4F_1.Y.n1 mux8_5.NAND4F_1.Y.t9 308.481
R28133 mux8_5.NAND4F_1.Y.n1 mux8_5.NAND4F_1.Y.t10 308.481
R28134 mux8_5.NAND4F_1.Y.n0 mux8_5.NAND4F_1.Y.n3 187.373
R28135 mux8_5.NAND4F_1.Y.n0 mux8_5.NAND4F_1.Y.n4 187.192
R28136 mux8_5.NAND4F_1.Y.n0 mux8_5.NAND4F_1.Y.n5 187.192
R28137 mux8_5.NAND4F_1.Y.n7 mux8_5.NAND4F_1.Y.n6 187.192
R28138 mux8_5.NAND4F_1.Y mux8_5.NAND4F_1.Y.n2 161.84
R28139 mux8_5.NAND4F_1.Y mux8_5.NAND4F_1.Y.t6 23.4335
R28140 mux8_5.NAND4F_1.Y.n3 mux8_5.NAND4F_1.Y.t1 20.1899
R28141 mux8_5.NAND4F_1.Y.n3 mux8_5.NAND4F_1.Y.t0 20.1899
R28142 mux8_5.NAND4F_1.Y.n4 mux8_5.NAND4F_1.Y.t3 20.1899
R28143 mux8_5.NAND4F_1.Y.n4 mux8_5.NAND4F_1.Y.t2 20.1899
R28144 mux8_5.NAND4F_1.Y.n5 mux8_5.NAND4F_1.Y.t5 20.1899
R28145 mux8_5.NAND4F_1.Y.n5 mux8_5.NAND4F_1.Y.t4 20.1899
R28146 mux8_5.NAND4F_1.Y.n6 mux8_5.NAND4F_1.Y.t8 20.1899
R28147 mux8_5.NAND4F_1.Y.n6 mux8_5.NAND4F_1.Y.t7 20.1899
R28148 mux8_5.NAND4F_1.Y.n2 mux8_5.NAND4F_1.Y.n1 11.0463
R28149 mux8_5.NAND4F_1.Y mux8_5.NAND4F_1.Y.n7 0.527586
R28150 mux8_5.NAND4F_1.Y.n7 mux8_5.NAND4F_1.Y.n0 0.358709
R28151 a_n20296_n12716.t0 a_n20296_n12716.t1 19.8005
R28152 a_n11840_n8419.n2 a_n11840_n8419.n1 121.353
R28153 a_n11840_n8419.n2 a_n11840_n8419.n0 121.353
R28154 a_n11840_n8419.n3 a_n11840_n8419.n2 121.001
R28155 a_n11840_n8419.n1 a_n11840_n8419.t1 30.462
R28156 a_n11840_n8419.n1 a_n11840_n8419.t0 30.462
R28157 a_n11840_n8419.n0 a_n11840_n8419.t5 30.462
R28158 a_n11840_n8419.n0 a_n11840_n8419.t4 30.462
R28159 a_n11840_n8419.n3 a_n11840_n8419.t3 30.462
R28160 a_n11840_n8419.t2 a_n11840_n8419.n3 30.462
R28161 a_n9125_n11063.n7 a_n9125_n11063.n1 81.2978
R28162 a_n9125_n11063.n1 a_n9125_n11063.n6 81.1637
R28163 a_n9125_n11063.n1 a_n9125_n11063.n5 81.1637
R28164 a_n9125_n11063.n0 a_n9125_n11063.n4 81.1637
R28165 a_n9125_n11063.n0 a_n9125_n11063.n3 81.1637
R28166 a_n9125_n11063.n0 a_n9125_n11063.n2 80.9213
R28167 a_n9125_n11063.n6 a_n9125_n11063.t6 11.8205
R28168 a_n9125_n11063.n6 a_n9125_n11063.t4 11.8205
R28169 a_n9125_n11063.n5 a_n9125_n11063.t7 11.8205
R28170 a_n9125_n11063.n5 a_n9125_n11063.t8 11.8205
R28171 a_n9125_n11063.n4 a_n9125_n11063.t1 11.8205
R28172 a_n9125_n11063.n4 a_n9125_n11063.t0 11.8205
R28173 a_n9125_n11063.n3 a_n9125_n11063.t11 11.8205
R28174 a_n9125_n11063.n3 a_n9125_n11063.t2 11.8205
R28175 a_n9125_n11063.n2 a_n9125_n11063.t9 11.8205
R28176 a_n9125_n11063.n2 a_n9125_n11063.t10 11.8205
R28177 a_n9125_n11063.n7 a_n9125_n11063.t3 11.8205
R28178 a_n9125_n11063.t5 a_n9125_n11063.n7 11.8205
R28179 a_n9125_n11063.n1 a_n9125_n11063.n0 0.402735
R28180 a_11386_n30934.t0 a_11386_n30934.t1 9.9005
R28181 a_n9314_n9452.t0 a_n9314_n9452.t1 19.8005
R28182 right_shifter_0.S6.n1 right_shifter_0.S6.t4 1032.02
R28183 right_shifter_0.S6.n1 right_shifter_0.S6.t5 336.962
R28184 right_shifter_0.S6.n1 right_shifter_0.S6.t6 326.154
R28185 right_shifter_0.S6.n0 right_shifter_0.S6.t1 256.514
R28186 right_shifter_0.S6.n0 right_shifter_0.S6.n2 226.258
R28187 mux8_8.NAND4F_6.A right_shifter_0.S6.n1 162.952
R28188 right_shifter_0.S6.n0 right_shifter_0.S6.t0 83.7172
R28189 mux8_8.A7 right_shifter_0.S6.n0 37.5537
R28190 right_shifter_0.S6.n2 right_shifter_0.S6.t3 30.379
R28191 right_shifter_0.S6.n2 right_shifter_0.S6.t2 30.379
R28192 mux8_8.A7 mux8_8.NAND4F_6.A 13.4456
R28193 right_shifter_0.S3.n1 right_shifter_0.S3.t4 1032.02
R28194 right_shifter_0.S3.n1 right_shifter_0.S3.t5 336.962
R28195 right_shifter_0.S3.n1 right_shifter_0.S3.t6 326.154
R28196 right_shifter_0.S3.n0 right_shifter_0.S3.t1 256.514
R28197 right_shifter_0.S3.n0 right_shifter_0.S3.n2 226.258
R28198 mux8_4.NAND4F_6.A right_shifter_0.S3.n1 162.952
R28199 right_shifter_0.S3.n0 right_shifter_0.S3.t0 83.7172
R28200 right_shifter_0.S3.n2 right_shifter_0.S3.t3 30.379
R28201 right_shifter_0.S3.n2 right_shifter_0.S3.t2 30.379
R28202 mux8_4.A7 right_shifter_0.S3.n0 23.1169
R28203 mux8_4.A7 mux8_4.NAND4F_6.A 13.4456
R28204 a_8592_n17350.t0 a_8592_n17350.t1 9.9005
R28205 a_9432_n34534.t0 a_9432_n34534.t1 9.9005
R28206 a_10363_n17349.t0 a_10363_n17349.t1 9.9005
R28207 a_n10684_n11683.n2 a_n10684_n11683.n1 121.353
R28208 a_n10684_n11683.n3 a_n10684_n11683.n2 121.001
R28209 a_n10684_n11683.n2 a_n10684_n11683.n0 120.977
R28210 a_n10684_n11683.n1 a_n10684_n11683.t3 30.462
R28211 a_n10684_n11683.n1 a_n10684_n11683.t4 30.462
R28212 a_n10684_n11683.n0 a_n10684_n11683.t0 30.462
R28213 a_n10684_n11683.n0 a_n10684_n11683.t1 30.462
R28214 a_n10684_n11683.t2 a_n10684_n11683.n3 30.462
R28215 a_n10684_n11683.n3 a_n10684_n11683.t5 30.462
R28216 left_shifter_0.buffer_1.inv_1.A.n0 left_shifter_0.buffer_1.inv_1.A.t5 393.921
R28217 left_shifter_0.buffer_1.inv_1.A.n2 left_shifter_0.buffer_1.inv_1.A.t6 291.829
R28218 left_shifter_0.buffer_1.inv_1.A.n2 left_shifter_0.buffer_1.inv_1.A.t4 291.829
R28219 left_shifter_0.buffer_1.inv_1.A.n0 left_shifter_0.buffer_1.inv_1.A.t3 256.89
R28220 left_shifter_0.buffer_1.inv_1.A.n0 left_shifter_0.buffer_1.inv_1.A.n1 226.538
R28221 left_shifter_0.buffer_1.inv_1.A.n2 left_shifter_0.buffer_1.inv_1.A.t7 221.72
R28222 left_shifter_0.buffer_1.inv_1.A.n0 left_shifter_0.buffer_1.inv_1.A.t0 83.795
R28223 left_shifter_0.buffer_1.inv_1.A.n0 left_shifter_0.buffer_1.inv_1.A.n2 53.7938
R28224 left_shifter_0.buffer_1.inv_1.A.n1 left_shifter_0.buffer_1.inv_1.A.t1 30.379
R28225 left_shifter_0.buffer_1.inv_1.A.n1 left_shifter_0.buffer_1.inv_1.A.t2 30.379
R28226 mux8_6.NAND4F_2.Y.n6 mux8_6.NAND4F_2.Y.t9 933.563
R28227 mux8_6.NAND4F_2.Y.n6 mux8_6.NAND4F_2.Y.t10 367.635
R28228 mux8_6.NAND4F_2.Y.n7 mux8_6.NAND4F_2.Y.t11 308.481
R28229 mux8_6.NAND4F_2.Y.n0 mux8_6.NAND4F_2.Y.n1 187.373
R28230 mux8_6.NAND4F_2.Y.n0 mux8_6.NAND4F_2.Y.n2 187.192
R28231 mux8_6.NAND4F_2.Y.n0 mux8_6.NAND4F_2.Y.n3 187.192
R28232 mux8_6.NAND4F_2.Y.n5 mux8_6.NAND4F_2.Y.n4 187.192
R28233 mux8_6.NAND4F_2.Y mux8_6.NAND4F_2.Y.n7 162.102
R28234 mux8_6.NAND4F_2.Y.n8 mux8_6.NAND4F_2.Y.t3 22.7096
R28235 mux8_6.NAND4F_2.Y.n8 mux8_6.NAND4F_2.Y 22.4285
R28236 mux8_6.NAND4F_2.Y.n1 mux8_6.NAND4F_2.Y.t1 20.1899
R28237 mux8_6.NAND4F_2.Y.n1 mux8_6.NAND4F_2.Y.t0 20.1899
R28238 mux8_6.NAND4F_2.Y.n2 mux8_6.NAND4F_2.Y.t5 20.1899
R28239 mux8_6.NAND4F_2.Y.n2 mux8_6.NAND4F_2.Y.t6 20.1899
R28240 mux8_6.NAND4F_2.Y.n3 mux8_6.NAND4F_2.Y.t8 20.1899
R28241 mux8_6.NAND4F_2.Y.n3 mux8_6.NAND4F_2.Y.t7 20.1899
R28242 mux8_6.NAND4F_2.Y.n4 mux8_6.NAND4F_2.Y.t2 20.1899
R28243 mux8_6.NAND4F_2.Y.n4 mux8_6.NAND4F_2.Y.t4 20.1899
R28244 mux8_6.NAND4F_2.Y.n7 mux8_6.NAND4F_2.Y.n6 10.955
R28245 mux8_6.NAND4F_2.Y mux8_6.NAND4F_2.Y.n8 0.799394
R28246 mux8_6.NAND4F_2.Y mux8_6.NAND4F_2.Y.n5 0.452586
R28247 mux8_6.NAND4F_2.Y.n5 mux8_6.NAND4F_2.Y.n0 0.358709
R28248 a_n23950_3190.n2 a_n23950_3190.n0 121.353
R28249 a_n23950_3190.n3 a_n23950_3190.n2 121.353
R28250 a_n23950_3190.n2 a_n23950_3190.n1 121.001
R28251 a_n23950_3190.n1 a_n23950_3190.t5 30.462
R28252 a_n23950_3190.n1 a_n23950_3190.t0 30.462
R28253 a_n23950_3190.n0 a_n23950_3190.t3 30.462
R28254 a_n23950_3190.n0 a_n23950_3190.t4 30.462
R28255 a_n23950_3190.n3 a_n23950_3190.t1 30.462
R28256 a_n23950_3190.t2 a_n23950_3190.n3 30.462
R28257 a_8400_762.t0 a_8400_762.t1 9.9005
R28258 a_10267_n2838.t0 a_10267_n2838.t1 9.9005
R28259 a_n11274_n17539.n2 a_n11274_n17539.n0 121.353
R28260 a_n11274_n17539.n3 a_n11274_n17539.n2 121.353
R28261 a_n11274_n17539.n2 a_n11274_n17539.n1 121.001
R28262 a_n11274_n17539.n0 a_n11274_n17539.t5 30.462
R28263 a_n11274_n17539.n0 a_n11274_n17539.t4 30.462
R28264 a_n11274_n17539.n1 a_n11274_n17539.t3 30.462
R28265 a_n11274_n17539.n1 a_n11274_n17539.t0 30.462
R28266 a_n11274_n17539.t2 a_n11274_n17539.n3 30.462
R28267 a_n11274_n17539.n3 a_n11274_n17539.t1 30.462
R28268 a_16431_n19505.n2 a_16431_n19505.n0 140.274
R28269 a_16431_n19505.n3 a_16431_n19505.n2 140.274
R28270 a_16431_n19505.n2 a_16431_n19505.n1 140.21
R28271 a_16431_n19505.n0 a_16431_n19505.t4 7.59513
R28272 a_16431_n19505.n0 a_16431_n19505.t3 7.59513
R28273 a_16431_n19505.n1 a_16431_n19505.t0 7.59513
R28274 a_16431_n19505.n1 a_16431_n19505.t5 7.59513
R28275 a_16431_n19505.t2 a_16431_n19505.n3 7.59513
R28276 a_16431_n19505.n3 a_16431_n19505.t1 7.59513
R28277 a_n2627_373.t0 a_n2627_373.t1 19.8005
R28278 a_n12605_n9452.t0 a_n12605_n9452.t1 19.8005
R28279 a_n9305_n8419.n0 a_n9305_n8419.t2 539.788
R28280 a_n9305_n8419.n1 a_n9305_n8419.t5 531.496
R28281 a_n9305_n8419.n0 a_n9305_n8419.t4 490.034
R28282 a_n9305_n8419.n5 a_n9305_n8419.t0 283.788
R28283 a_n9305_n8419.t1 a_n9305_n8419.n5 205.489
R28284 a_n9305_n8419.n2 a_n9305_n8419.t6 182.625
R28285 a_n9305_n8419.n3 a_n9305_n8419.t3 179.054
R28286 a_n9305_n8419.n2 a_n9305_n8419.t7 139.78
R28287 a_n9305_n8419.n4 a_n9305_n8419.n3 101.368
R28288 a_n9305_n8419.n5 a_n9305_n8419.n4 77.9135
R28289 a_n9305_n8419.n4 a_n9305_n8419.n1 76.1557
R28290 a_n9305_n8419.n1 a_n9305_n8419.n0 8.29297
R28291 a_n9305_n8419.n3 a_n9305_n8419.n2 3.57087
R28292 a_n9125_n8419.n2 a_n9125_n8419.n1 121.353
R28293 a_n9125_n8419.n3 a_n9125_n8419.n2 121.001
R28294 a_n9125_n8419.n2 a_n9125_n8419.n0 120.977
R28295 a_n9125_n8419.n1 a_n9125_n8419.t1 30.462
R28296 a_n9125_n8419.n1 a_n9125_n8419.t0 30.462
R28297 a_n9125_n8419.n0 a_n9125_n8419.t4 30.462
R28298 a_n9125_n8419.n0 a_n9125_n8419.t3 30.462
R28299 a_n9125_n8419.n3 a_n9125_n8419.t5 30.462
R28300 a_n9125_n8419.t2 a_n9125_n8419.n3 30.462
R28301 a_n10684_n5154.n2 a_n10684_n5154.n1 121.353
R28302 a_n10684_n5154.n3 a_n10684_n5154.n2 121.001
R28303 a_n10684_n5154.n2 a_n10684_n5154.n0 120.977
R28304 a_n10684_n5154.n1 a_n10684_n5154.t1 30.462
R28305 a_n10684_n5154.n1 a_n10684_n5154.t0 30.462
R28306 a_n10684_n5154.n0 a_n10684_n5154.t3 30.462
R28307 a_n10684_n5154.n0 a_n10684_n5154.t5 30.462
R28308 a_n10684_n5154.n3 a_n10684_n5154.t4 30.462
R28309 a_n10684_n5154.t2 a_n10684_n5154.n3 30.462
R28310 a_8496_n16422.t0 a_8496_n16422.t1 9.9005
R28311 a_8592_n16422.t0 a_8592_n16422.t1 9.9005
R28312 a_n10423_n9452.t0 a_n10423_n9452.t1 19.8005
R28313 a_8400_n20950.t0 a_8400_n20950.t1 9.9005
R28314 a_8496_762.t0 a_8496_762.t1 9.9005
R28315 a_8592_762.t0 a_8592_762.t1 9.9005
R28316 a_n12416_n5154.n2 a_n12416_n5154.n1 121.353
R28317 a_n12416_n5154.n3 a_n12416_n5154.n2 121.001
R28318 a_n12416_n5154.n2 a_n12416_n5154.n0 120.977
R28319 a_n12416_n5154.n1 a_n12416_n5154.t4 30.462
R28320 a_n12416_n5154.n1 a_n12416_n5154.t3 30.462
R28321 a_n12416_n5154.n0 a_n12416_n5154.t0 30.462
R28322 a_n12416_n5154.n0 a_n12416_n5154.t1 30.462
R28323 a_n12416_n5154.t2 a_n12416_n5154.n3 30.462
R28324 a_n12416_n5154.n3 a_n12416_n5154.t5 30.462
R28325 a_n3659_3164.n0 a_n3659_3164.t7 539.788
R28326 a_n3659_3164.n1 a_n3659_3164.t5 531.496
R28327 a_n3659_3164.n0 a_n3659_3164.t3 490.034
R28328 a_n3659_3164.n5 a_n3659_3164.t0 283.788
R28329 a_n3659_3164.t1 a_n3659_3164.n5 205.489
R28330 a_n3659_3164.n2 a_n3659_3164.t6 182.625
R28331 a_n3659_3164.n3 a_n3659_3164.t4 179.054
R28332 a_n3659_3164.n2 a_n3659_3164.t2 139.78
R28333 a_n3659_3164.n4 a_n3659_3164.n3 101.368
R28334 a_n3659_3164.n5 a_n3659_3164.n4 77.9135
R28335 a_n3659_3164.n4 a_n3659_3164.n1 76.1557
R28336 a_n3659_3164.n1 a_n3659_3164.n0 8.29297
R28337 a_n3659_3164.n3 a_n3659_3164.n2 3.57087
R28338 a_n22425_n7992.t0 a_n22425_n7992.t1 19.8005
R28339 a_11290_n17350.t0 a_11290_n17350.t1 9.9005
R28340 a_8592_n3766.t0 a_8592_n3766.t1 9.9005
R28341 a_11290_n3766.t0 a_11290_n3766.t1 9.9005
R28342 a_8592_n30934.t0 a_8592_n30934.t1 9.9005
R28343 a_10363_n30933.t0 a_10363_n30933.t1 9.9005
R28344 a_n18305_n12716.t0 a_n18305_n12716.t1 19.8005
R28345 a_n17368_3190.n2 a_n17368_3190.n0 121.353
R28346 a_n17368_3190.n3 a_n17368_3190.n2 121.353
R28347 a_n17368_3190.n2 a_n17368_3190.n1 121.001
R28348 a_n17368_3190.n1 a_n17368_3190.t3 30.462
R28349 a_n17368_3190.n1 a_n17368_3190.t0 30.462
R28350 a_n17368_3190.n0 a_n17368_3190.t5 30.462
R28351 a_n17368_3190.n0 a_n17368_3190.t4 30.462
R28352 a_n17368_3190.n3 a_n17368_3190.t1 30.462
R28353 a_n17368_3190.t2 a_n17368_3190.n3 30.462
R28354 a_n13975_n11063.n1 a_n13975_n11063.n5 81.2978
R28355 a_n13975_n11063.n1 a_n13975_n11063.n6 81.1637
R28356 a_n13975_n11063.n0 a_n13975_n11063.n4 81.1637
R28357 a_n13975_n11063.n0 a_n13975_n11063.n3 81.1637
R28358 a_n13975_n11063.n7 a_n13975_n11063.n1 81.1637
R28359 a_n13975_n11063.n0 a_n13975_n11063.n2 80.9213
R28360 a_n13975_n11063.n5 a_n13975_n11063.t8 11.8205
R28361 a_n13975_n11063.n5 a_n13975_n11063.t7 11.8205
R28362 a_n13975_n11063.n6 a_n13975_n11063.t0 11.8205
R28363 a_n13975_n11063.n6 a_n13975_n11063.t6 11.8205
R28364 a_n13975_n11063.n4 a_n13975_n11063.t10 11.8205
R28365 a_n13975_n11063.n4 a_n13975_n11063.t11 11.8205
R28366 a_n13975_n11063.n3 a_n13975_n11063.t5 11.8205
R28367 a_n13975_n11063.n3 a_n13975_n11063.t9 11.8205
R28368 a_n13975_n11063.n2 a_n13975_n11063.t3 11.8205
R28369 a_n13975_n11063.n2 a_n13975_n11063.t4 11.8205
R28370 a_n13975_n11063.n7 a_n13975_n11063.t1 11.8205
R28371 a_n13975_n11063.t2 a_n13975_n11063.n7 11.8205
R28372 a_n13975_n11063.n1 a_n13975_n11063.n0 0.402735
R28373 a_11194_n16422.t0 a_11194_n16422.t1 9.9005
R28374 a_11290_n16422.t0 a_11290_n16422.t1 9.9005
R28375 a_n8432_n9452.t0 a_n8432_n9452.t1 19.8005
R28376 a_11290_n30934.t0 a_11290_n30934.t1 9.9005
R28377 a_n13399_n8419.n2 a_n13399_n8419.n0 121.353
R28378 a_n13399_n8419.n3 a_n13399_n8419.n2 121.353
R28379 a_n13399_n8419.n2 a_n13399_n8419.n1 121.001
R28380 a_n13399_n8419.n0 a_n13399_n8419.t3 30.462
R28381 a_n13399_n8419.n0 a_n13399_n8419.t5 30.462
R28382 a_n13399_n8419.n1 a_n13399_n8419.t0 30.462
R28383 a_n13399_n8419.n1 a_n13399_n8419.t4 30.462
R28384 a_n13399_n8419.n3 a_n13399_n8419.t1 30.462
R28385 a_n13399_n8419.t2 a_n13399_n8419.n3 30.462
R28386 a_9336_1690.t0 a_9336_1690.t1 9.9005
R28387 a_n15707_n11683.n2 a_n15707_n11683.n1 121.353
R28388 a_n15707_n11683.n3 a_n15707_n11683.n2 121.001
R28389 a_n15707_n11683.n2 a_n15707_n11683.n0 120.977
R28390 a_n15707_n11683.n1 a_n15707_n11683.t5 30.462
R28391 a_n15707_n11683.n1 a_n15707_n11683.t3 30.462
R28392 a_n15707_n11683.n0 a_n15707_n11683.t0 30.462
R28393 a_n15707_n11683.n0 a_n15707_n11683.t1 30.462
R28394 a_n15707_n11683.t2 a_n15707_n11683.n3 30.462
R28395 a_n15707_n11683.n3 a_n15707_n11683.t4 30.462
R28396 a_8400_n16422.t0 a_8400_n16422.t1 9.9005
R28397 left_shifter_0.buffer_3.inv_1.A.n0 left_shifter_0.buffer_3.inv_1.A.t6 393.921
R28398 left_shifter_0.buffer_3.inv_1.A.n2 left_shifter_0.buffer_3.inv_1.A.t4 291.829
R28399 left_shifter_0.buffer_3.inv_1.A.n2 left_shifter_0.buffer_3.inv_1.A.t7 291.829
R28400 left_shifter_0.buffer_3.inv_1.A.n0 left_shifter_0.buffer_3.inv_1.A.t1 256.89
R28401 left_shifter_0.buffer_3.inv_1.A.n0 left_shifter_0.buffer_3.inv_1.A.n1 226.538
R28402 left_shifter_0.buffer_3.inv_1.A.n2 left_shifter_0.buffer_3.inv_1.A.t5 221.72
R28403 left_shifter_0.buffer_3.inv_1.A.n0 left_shifter_0.buffer_3.inv_1.A.t0 83.795
R28404 left_shifter_0.buffer_3.inv_1.A.n0 left_shifter_0.buffer_3.inv_1.A.n2 53.7938
R28405 left_shifter_0.buffer_3.inv_1.A.n1 left_shifter_0.buffer_3.inv_1.A.t2 30.379
R28406 left_shifter_0.buffer_3.inv_1.A.n1 left_shifter_0.buffer_3.inv_1.A.t3 30.379
R28407 a_11386_n11894.t0 a_11386_n11894.t1 9.9005
R28408 a_10267_n25478.t0 a_10267_n25478.t1 9.9005
R28409 a_10363_n25478.t0 a_10363_n25478.t1 9.9005
R28410 mux8_4.NAND4F_2.Y.n6 mux8_4.NAND4F_2.Y.t9 933.563
R28411 mux8_4.NAND4F_2.Y.n6 mux8_4.NAND4F_2.Y.t10 367.635
R28412 mux8_4.NAND4F_2.Y.n7 mux8_4.NAND4F_2.Y.t11 308.481
R28413 mux8_4.NAND4F_2.Y.n0 mux8_4.NAND4F_2.Y.n1 187.373
R28414 mux8_4.NAND4F_2.Y.n0 mux8_4.NAND4F_2.Y.n2 187.192
R28415 mux8_4.NAND4F_2.Y.n0 mux8_4.NAND4F_2.Y.n3 187.192
R28416 mux8_4.NAND4F_2.Y.n5 mux8_4.NAND4F_2.Y.n4 187.192
R28417 mux8_4.NAND4F_2.Y mux8_4.NAND4F_2.Y.n7 162.102
R28418 mux8_4.NAND4F_2.Y.n8 mux8_4.NAND4F_2.Y.t2 22.7096
R28419 mux8_4.NAND4F_2.Y.n8 mux8_4.NAND4F_2.Y 22.4285
R28420 mux8_4.NAND4F_2.Y.n1 mux8_4.NAND4F_2.Y.t1 20.1899
R28421 mux8_4.NAND4F_2.Y.n1 mux8_4.NAND4F_2.Y.t0 20.1899
R28422 mux8_4.NAND4F_2.Y.n2 mux8_4.NAND4F_2.Y.t6 20.1899
R28423 mux8_4.NAND4F_2.Y.n2 mux8_4.NAND4F_2.Y.t5 20.1899
R28424 mux8_4.NAND4F_2.Y.n3 mux8_4.NAND4F_2.Y.t7 20.1899
R28425 mux8_4.NAND4F_2.Y.n3 mux8_4.NAND4F_2.Y.t8 20.1899
R28426 mux8_4.NAND4F_2.Y.n4 mux8_4.NAND4F_2.Y.t4 20.1899
R28427 mux8_4.NAND4F_2.Y.n4 mux8_4.NAND4F_2.Y.t3 20.1899
R28428 mux8_4.NAND4F_2.Y.n7 mux8_4.NAND4F_2.Y.n6 10.955
R28429 mux8_4.NAND4F_2.Y mux8_4.NAND4F_2.Y.n8 0.799394
R28430 mux8_4.NAND4F_2.Y mux8_4.NAND4F_2.Y.n5 0.452586
R28431 mux8_4.NAND4F_2.Y.n5 mux8_4.NAND4F_2.Y.n0 0.358709
R28432 mux8_3.NAND4F_6.Y.n1 mux8_3.NAND4F_6.Y.t11 933.563
R28433 mux8_3.NAND4F_6.Y.n1 mux8_3.NAND4F_6.Y.t9 367.635
R28434 mux8_3.NAND4F_6.Y.n2 mux8_3.NAND4F_6.Y.t10 308.481
R28435 mux8_3.NAND4F_6.Y.n0 mux8_3.NAND4F_6.Y.n4 187.373
R28436 mux8_3.NAND4F_6.Y.n0 mux8_3.NAND4F_6.Y.n5 187.192
R28437 mux8_3.NAND4F_6.Y.n0 mux8_3.NAND4F_6.Y.n6 187.192
R28438 mux8_3.NAND4F_6.Y.n8 mux8_3.NAND4F_6.Y.n7 187.192
R28439 mux8_3.NAND4F_6.Y mux8_3.NAND4F_6.Y.n2 162.047
R28440 mux8_3.NAND4F_6.Y.n3 mux8_3.NAND4F_6.Y.t2 22.7831
R28441 mux8_3.NAND4F_6.Y.n3 mux8_3.NAND4F_6.Y 22.171
R28442 mux8_3.NAND4F_6.Y.n4 mux8_3.NAND4F_6.Y.t1 20.1899
R28443 mux8_3.NAND4F_6.Y.n4 mux8_3.NAND4F_6.Y.t0 20.1899
R28444 mux8_3.NAND4F_6.Y.n5 mux8_3.NAND4F_6.Y.t5 20.1899
R28445 mux8_3.NAND4F_6.Y.n5 mux8_3.NAND4F_6.Y.t6 20.1899
R28446 mux8_3.NAND4F_6.Y.n6 mux8_3.NAND4F_6.Y.t8 20.1899
R28447 mux8_3.NAND4F_6.Y.n6 mux8_3.NAND4F_6.Y.t7 20.1899
R28448 mux8_3.NAND4F_6.Y.n7 mux8_3.NAND4F_6.Y.t4 20.1899
R28449 mux8_3.NAND4F_6.Y.n7 mux8_3.NAND4F_6.Y.t3 20.1899
R28450 mux8_3.NAND4F_6.Y.n2 mux8_3.NAND4F_6.Y.n1 10.955
R28451 mux8_3.NAND4F_6.Y mux8_3.NAND4F_6.Y.n3 0.781576
R28452 mux8_3.NAND4F_6.Y mux8_3.NAND4F_6.Y.n8 0.396904
R28453 mux8_3.NAND4F_6.Y.n8 mux8_3.NAND4F_6.Y.n0 0.358709
R28454 OR8_0.S7.n1 OR8_0.S7.t5 1032.02
R28455 OR8_0.S7.n1 OR8_0.S7.t4 336.962
R28456 OR8_0.S7.n1 OR8_0.S7.t6 326.154
R28457 OR8_0.S7.n0 OR8_0.S7.t1 256.514
R28458 OR8_0.S7.n0 OR8_0.S7.n2 226.258
R28459 OR8_0.S7 OR8_0.S7.n1 162.952
R28460 OR8_0.S7.n0 OR8_0.S7.t0 83.7172
R28461 OR8_0.S7.n2 OR8_0.S7.t2 30.379
R28462 OR8_0.S7.n2 OR8_0.S7.t3 30.379
R28463 OR8_0.S7 OR8_0.S7.n0 1.94945
R28464 mux8_4.NAND4F_8.Y.n1 mux8_4.NAND4F_8.Y.t10 379.173
R28465 mux8_4.NAND4F_8.Y.n2 mux8_4.NAND4F_8.Y.t14 312.599
R28466 mux8_4.NAND4F_8.Y.n1 mux8_4.NAND4F_8.Y.t9 247.428
R28467 mux8_4.NAND4F_8.Y.n4 mux8_4.NAND4F_8.Y.t11 247.428
R28468 mux8_4.NAND4F_8.Y.n3 mux8_4.NAND4F_8.Y.t13 247.428
R28469 mux8_4.NAND4F_8.Y.n2 mux8_4.NAND4F_8.Y.t12 247.428
R28470 mux8_4.NAND4F_8.Y.n0 mux8_4.NAND4F_8.Y.n6 187.373
R28471 mux8_4.NAND4F_8.Y.n0 mux8_4.NAND4F_8.Y.n7 187.192
R28472 mux8_4.NAND4F_8.Y.n0 mux8_4.NAND4F_8.Y.n8 187.192
R28473 mux8_4.NAND4F_8.Y.n10 mux8_4.NAND4F_8.Y.n9 187.192
R28474 mux8_4.NAND4F_8.Y mux8_4.NAND4F_8.Y.n5 162.139
R28475 mux8_4.NAND4F_8.Y.n4 mux8_4.NAND4F_8.Y.n3 65.1723
R28476 mux8_4.NAND4F_8.Y.n3 mux8_4.NAND4F_8.Y.n2 65.1723
R28477 mux8_4.NAND4F_8.Y.n5 mux8_4.NAND4F_8.Y.n4 33.2653
R28478 mux8_4.NAND4F_8.Y.n5 mux8_4.NAND4F_8.Y.n1 31.9075
R28479 mux8_4.NAND4F_8.Y mux8_4.NAND4F_8.Y.t6 22.6141
R28480 mux8_4.NAND4F_8.Y.n6 mux8_4.NAND4F_8.Y.t4 20.1899
R28481 mux8_4.NAND4F_8.Y.n6 mux8_4.NAND4F_8.Y.t5 20.1899
R28482 mux8_4.NAND4F_8.Y.n7 mux8_4.NAND4F_8.Y.t1 20.1899
R28483 mux8_4.NAND4F_8.Y.n7 mux8_4.NAND4F_8.Y.t0 20.1899
R28484 mux8_4.NAND4F_8.Y.n8 mux8_4.NAND4F_8.Y.t3 20.1899
R28485 mux8_4.NAND4F_8.Y.n8 mux8_4.NAND4F_8.Y.t2 20.1899
R28486 mux8_4.NAND4F_8.Y.n9 mux8_4.NAND4F_8.Y.t8 20.1899
R28487 mux8_4.NAND4F_8.Y.n9 mux8_4.NAND4F_8.Y.t7 20.1899
R28488 mux8_4.NAND4F_8.Y mux8_4.NAND4F_8.Y.n10 0.452586
R28489 mux8_4.NAND4F_8.Y.n10 mux8_4.NAND4F_8.Y.n0 0.358709
R28490 a_n15014_n6187.t0 a_n15014_n6187.t1 19.8005
R28491 a_8400_n21878.t0 a_8400_n21878.t1 9.9005
R28492 a_10267_n7266.t0 a_10267_n7266.t1 9.9005
R28493 a_7644_n17350.t0 a_7644_n17350.t1 9.9005
R28494 a_9528_n21878.t0 a_9528_n21878.t1 9.9005
R28495 a_n24013_n15316.t0 a_n24013_n15316.t1 19.8005
R28496 a_n10108_n8419.n2 a_n10108_n8419.n0 121.353
R28497 a_n10108_n8419.n3 a_n10108_n8419.n2 121.353
R28498 a_n10108_n8419.n2 a_n10108_n8419.n1 121.001
R28499 a_n10108_n8419.n1 a_n10108_n8419.t3 30.462
R28500 a_n10108_n8419.n1 a_n10108_n8419.t0 30.462
R28501 a_n10108_n8419.n0 a_n10108_n8419.t5 30.462
R28502 a_n10108_n8419.n0 a_n10108_n8419.t4 30.462
R28503 a_n10108_n8419.t2 a_n10108_n8419.n3 30.462
R28504 a_n10108_n8419.n3 a_n10108_n8419.t1 30.462
R28505 a_11386_n34534.t0 a_11386_n34534.t1 9.9005
R28506 a_n24162_n11256.t0 a_n24162_n11256.t1 19.8005
R28507 a_11290_n8194.t0 a_11290_n8194.t1 9.9005
R28508 a_8592_n8194.t0 a_8592_n8194.t1 9.9005
R28509 a_8592_n11894.t0 a_8592_n11894.t1 9.9005
R28510 a_8496_1690.t0 a_8496_1690.t1 9.9005
R28511 a_8592_1690.t0 a_8592_1690.t1 9.9005
R28512 a_7452_n12822.t0 a_7452_n12822.t1 9.9005
R28513 left_shifter_0.S6.n1 left_shifter_0.S6.t4 1032.02
R28514 left_shifter_0.S6.n1 left_shifter_0.S6.t5 336.962
R28515 left_shifter_0.S6.n1 left_shifter_0.S6.t6 326.154
R28516 left_shifter_0.S6.n0 left_shifter_0.S6.t1 256.89
R28517 left_shifter_0.S6.n0 left_shifter_0.S6.n2 226.635
R28518 mux8_8.NAND4F_5.A left_shifter_0.S6.n1 162.952
R28519 left_shifter_0.S6.n0 left_shifter_0.S6.t0 83.7172
R28520 mux8_8.A6 left_shifter_0.S6.n0 41.5179
R28521 left_shifter_0.S6.n2 left_shifter_0.S6.t2 30.379
R28522 left_shifter_0.S6.n2 left_shifter_0.S6.t3 30.379
R28523 mux8_8.A6 mux8_8.NAND4F_5.A 11.8717
R28524 a_7644_n30934.t0 a_7644_n30934.t1 9.9005
R28525 a_7452_n3766.t0 a_7452_n3766.t1 9.9005
R28526 a_n17005_n9452.t0 a_n17005_n9452.t1 19.8005
R28527 a_10363_n2838.t0 a_10363_n2838.t1 9.9005
R28528 a_8592_n34534.t0 a_8592_n34534.t1 9.9005
R28529 a_11290_n11894.t0 a_11290_n11894.t1 9.9005
R28530 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t7 485.221
R28531 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t8 367.928
R28532 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n4 227.526
R28533 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n5 227.266
R28534 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n6 227.266
R28535 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t9 224.478
R28536 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t10 213.688
R28537 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n2 84.5046
R28538 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n1 72.3005
R28539 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n3 61.0566
R28540 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t0 42.7747
R28541 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t4 30.379
R28542 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t5 30.379
R28543 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t1 30.379
R28544 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t6 30.379
R28545 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t2 30.379
R28546 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.t3 30.379
R28547 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A.n0 0.583137
R28548 a_n19081_373.t0 a_n19081_373.t1 19.8005
R28549 a_15855_n18523.n2 a_15855_n18523.n0 140.274
R28550 a_15855_n18523.n3 a_15855_n18523.n2 140.274
R28551 a_15855_n18523.n2 a_15855_n18523.n1 140.21
R28552 a_15855_n18523.n1 a_15855_n18523.t3 7.59513
R28553 a_15855_n18523.n1 a_15855_n18523.t1 7.59513
R28554 a_15855_n18523.n0 a_15855_n18523.t5 7.59513
R28555 a_15855_n18523.n0 a_15855_n18523.t4 7.59513
R28556 a_15855_n18523.t2 a_15855_n18523.n3 7.59513
R28557 a_15855_n18523.n3 a_15855_n18523.t0 7.59513
R28558 a_n9155_n11709.n2 a_n9155_n11709.t2 541.395
R28559 a_n9155_n11709.n3 a_n9155_n11709.t7 527.402
R28560 a_n9155_n11709.n2 a_n9155_n11709.t6 491.64
R28561 a_n9155_n11709.n5 a_n9155_n11709.t0 281.906
R28562 a_n9155_n11709.t1 a_n9155_n11709.n5 204.359
R28563 a_n9155_n11709.n0 a_n9155_n11709.t4 180.73
R28564 a_n9155_n11709.n1 a_n9155_n11709.t3 179.45
R28565 a_n9155_n11709.n0 a_n9155_n11709.t5 139.78
R28566 a_n9155_n11709.n4 a_n9155_n11709.n1 105.635
R28567 a_n9155_n11709.n4 a_n9155_n11709.n3 76.0005
R28568 a_n9155_n11709.n5 a_n9155_n11709.n4 67.9685
R28569 a_n9155_n11709.n3 a_n9155_n11709.n2 13.994
R28570 a_n9155_n11709.n1 a_n9155_n11709.n0 1.28015
R28571 a_10267_n30006.t0 a_10267_n30006.t1 9.9005
R28572 a_7548_n17350.t0 a_7548_n17350.t1 9.9005
R28573 a_9432_n21878.t0 a_9432_n21878.t1 9.9005
R28574 a_11290_n34534.t0 a_11290_n34534.t1 9.9005
R28575 left_shifter_0.S4.n1 left_shifter_0.S4.t4 1032.02
R28576 left_shifter_0.S4.n1 left_shifter_0.S4.t5 336.962
R28577 left_shifter_0.S4.n1 left_shifter_0.S4.t6 326.154
R28578 left_shifter_0.S4.n0 left_shifter_0.S4.t1 256.89
R28579 left_shifter_0.S4.n0 left_shifter_0.S4.n2 226.635
R28580 mux8_5.NAND4F_5.A left_shifter_0.S4.n1 162.952
R28581 left_shifter_0.S4.n0 left_shifter_0.S4.t0 83.7172
R28582 mux8_5.A6 left_shifter_0.S4.n0 33.2528
R28583 left_shifter_0.S4.n2 left_shifter_0.S4.t2 30.379
R28584 left_shifter_0.S4.n2 left_shifter_0.S4.t3 30.379
R28585 mux8_5.A6 mux8_5.NAND4F_5.A 11.7469
R28586 right_shifter_0.buffer_0.inv_1.A.n0 right_shifter_0.buffer_0.inv_1.A.t4 393.921
R28587 right_shifter_0.buffer_0.inv_1.A.n2 right_shifter_0.buffer_0.inv_1.A.t7 291.829
R28588 right_shifter_0.buffer_0.inv_1.A.n2 right_shifter_0.buffer_0.inv_1.A.t6 291.829
R28589 right_shifter_0.buffer_0.inv_1.A.n0 right_shifter_0.buffer_0.inv_1.A.t1 256.514
R28590 right_shifter_0.buffer_0.inv_1.A.n0 right_shifter_0.buffer_0.inv_1.A.n1 226.162
R28591 right_shifter_0.buffer_0.inv_1.A.n2 right_shifter_0.buffer_0.inv_1.A.t5 221.72
R28592 right_shifter_0.buffer_0.inv_1.A.n0 right_shifter_0.buffer_0.inv_1.A.t0 83.795
R28593 right_shifter_0.buffer_0.inv_1.A.n0 right_shifter_0.buffer_0.inv_1.A.n2 53.7938
R28594 right_shifter_0.buffer_0.inv_1.A.n1 right_shifter_0.buffer_0.inv_1.A.t3 30.379
R28595 right_shifter_0.buffer_0.inv_1.A.n1 right_shifter_0.buffer_0.inv_1.A.t2 30.379
R28596 right_shifter_0.S1.n1 right_shifter_0.S1.t5 1032.02
R28597 right_shifter_0.S1.n1 right_shifter_0.S1.t6 336.962
R28598 right_shifter_0.S1.n1 right_shifter_0.S1.t4 326.154
R28599 right_shifter_0.S1.n0 right_shifter_0.S1.t1 256.514
R28600 right_shifter_0.S1.n0 right_shifter_0.S1.n2 226.258
R28601 mux8_2.NAND4F_6.A right_shifter_0.S1.n1 162.952
R28602 right_shifter_0.S1.n0 right_shifter_0.S1.t0 83.7172
R28603 mux8_2.A7 right_shifter_0.S1.n0 56.6316
R28604 right_shifter_0.S1.n2 right_shifter_0.S1.t3 30.379
R28605 right_shifter_0.S1.n2 right_shifter_0.S1.t2 30.379
R28606 mux8_2.A7 mux8_2.NAND4F_6.A 13.4456
R28607 a_n1327_373.t0 a_n1327_373.t1 19.8005
R28608 a_7452_1690.t0 a_7452_1690.t1 9.9005
R28609 a_7548_n30934.t0 a_7548_n30934.t1 9.9005
R28610 a_10459_1690.t0 a_10459_1690.t1 9.9005
R28611 a_9336_n17350.t0 a_9336_n17350.t1 9.9005
R28612 a_8496_n26406.t0 a_8496_n26406.t1 9.9005
R28613 a_10267_n26405.t0 a_10267_n26405.t1 9.9005
R28614 a_9528_n25478.t0 a_9528_n25478.t1 9.9005
R28615 a_8496_n35462.t0 a_8496_n35462.t1 9.9005
R28616 a_10267_n35461.t0 a_10267_n35461.t1 9.9005
R28617 a_n24007_n17714.t0 a_n24007_n17714.t1 19.8005
R28618 a_7644_n11894.t0 a_7644_n11894.t1 9.9005
R28619 a_7452_n8194.t0 a_7452_n8194.t1 9.9005
R28620 a_7452_n17350.t0 a_7452_n17350.t1 9.9005
R28621 a_11386_1690.t0 a_11386_1690.t1 9.9005
R28622 a_9336_n30934.t0 a_9336_n30934.t1 9.9005
R28623 a_11194_n26406.t0 a_11194_n26406.t1 9.9005
R28624 a_n19028_n5180.n2 a_n19028_n5180.t6 541.395
R28625 a_n19028_n5180.n3 a_n19028_n5180.t3 527.402
R28626 a_n19028_n5180.n2 a_n19028_n5180.t5 491.64
R28627 a_n19028_n5180.n5 a_n19028_n5180.t0 281.906
R28628 a_n19028_n5180.t1 a_n19028_n5180.n5 204.359
R28629 a_n19028_n5180.n0 a_n19028_n5180.t2 180.73
R28630 a_n19028_n5180.n1 a_n19028_n5180.t7 179.45
R28631 a_n19028_n5180.n0 a_n19028_n5180.t4 139.78
R28632 a_n19028_n5180.n4 a_n19028_n5180.n1 105.635
R28633 a_n19028_n5180.n4 a_n19028_n5180.n3 76.0005
R28634 a_n19028_n5180.n5 a_n19028_n5180.n4 67.9685
R28635 a_n19028_n5180.n3 a_n19028_n5180.n2 13.994
R28636 a_n19028_n5180.n1 a_n19028_n5180.n0 1.28015
R28637 a_10363_n7266.t0 a_10363_n7266.t1 9.9005
R28638 a_n9208_373.t0 a_n9208_373.t1 19.8005
R28639 a_n23254_373.t0 a_n23254_373.t1 19.8005
R28640 a_7644_n34534.t0 a_7644_n34534.t1 9.9005
R28641 a_10459_n21877.t0 a_10459_n21877.t1 9.9005
R28642 a_11194_n35462.t0 a_11194_n35462.t1 9.9005
R28643 a_7452_n30934.t0 a_7452_n30934.t1 9.9005
R28644 a_n15014_n9452.t0 a_n15014_n9452.t1 19.8005
R28645 a_8400_n26406.t0 a_8400_n26406.t1 9.9005
R28646 a_n24363_373.t0 a_n24363_373.t1 19.8005
R28647 a_11386_n21878.t0 a_11386_n21878.t1 9.9005
R28648 a_9432_n25478.t0 a_9432_n25478.t1 9.9005
R28649 a_8400_n35462.t0 a_8400_n35462.t1 9.9005
R28650 a_7548_n11894.t0 a_7548_n11894.t1 9.9005
R28651 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t7 485.221
R28652 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t8 367.928
R28653 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n5 227.526
R28654 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n4 227.266
R28655 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n6 227.266
R28656 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t9 224.478
R28657 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t10 213.688
R28658 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n2 84.5046
R28659 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n1 72.3005
R28660 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n3 61.0566
R28661 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t3 42.7747
R28662 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t0 30.379
R28663 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t1 30.379
R28664 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t4 30.379
R28665 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t6 30.379
R28666 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t5 30.379
R28667 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.t2 30.379
R28668 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A.n0 0.583137
R28669 a_9528_n30006.t0 a_9528_n30006.t1 9.9005
R28670 right_shifter_0.buffer_6.inv_1.A.n0 right_shifter_0.buffer_6.inv_1.A.t4 393.921
R28671 right_shifter_0.buffer_6.inv_1.A.n2 right_shifter_0.buffer_6.inv_1.A.t7 291.829
R28672 right_shifter_0.buffer_6.inv_1.A.n2 right_shifter_0.buffer_6.inv_1.A.t6 291.829
R28673 right_shifter_0.buffer_6.inv_1.A.n0 right_shifter_0.buffer_6.inv_1.A.t1 256.514
R28674 right_shifter_0.buffer_6.inv_1.A.n0 right_shifter_0.buffer_6.inv_1.A.n1 226.162
R28675 right_shifter_0.buffer_6.inv_1.A.n2 right_shifter_0.buffer_6.inv_1.A.t5 221.72
R28676 right_shifter_0.buffer_6.inv_1.A.n0 right_shifter_0.buffer_6.inv_1.A.t0 83.795
R28677 right_shifter_0.buffer_6.inv_1.A.n0 right_shifter_0.buffer_6.inv_1.A.n2 53.7938
R28678 right_shifter_0.buffer_6.inv_1.A.n1 right_shifter_0.buffer_6.inv_1.A.t3 30.379
R28679 right_shifter_0.buffer_6.inv_1.A.n1 right_shifter_0.buffer_6.inv_1.A.t2 30.379
R28680 a_11194_n2838.t0 a_11194_n2838.t1 9.9005
R28681 a_8496_n2838.t0 a_8496_n2838.t1 9.9005
R28682 a_7548_n34534.t0 a_7548_n34534.t1 9.9005
R28683 a_8592_n21878.t0 a_8592_n21878.t1 9.9005
R28684 a_10363_n21877.t0 a_10363_n21877.t1 9.9005
R28685 a_n18686_n2915.t0 a_n18686_n2915.t1 19.8005
R28686 a_n22425_n11256.t0 a_n22425_n11256.t1 19.8005
R28687 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t7 540.38
R28688 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t8 367.928
R28689 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n4 227.526
R28690 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t9 227.356
R28691 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n5 227.266
R28692 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n6 227.266
R28693 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t10 213.688
R28694 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n2 160.439
R28695 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n1 94.4341
R28696 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t0 42.7944
R28697 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t4 30.379
R28698 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t5 30.379
R28699 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t1 30.379
R28700 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t6 30.379
R28701 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t2 30.379
R28702 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.t3 30.379
R28703 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n0 13.4358
R28704 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B.n3 0.821842
R28705 a_9336_n11894.t0 a_9336_n11894.t1 9.9005
R28706 a_n22372_373.t0 a_n22372_373.t1 19.8005
R28707 a_11290_n21878.t0 a_11290_n21878.t1 9.9005
R28708 a_9336_n34534.t0 a_9336_n34534.t1 9.9005
R28709 a_7452_n11894.t0 a_7452_n11894.t1 9.9005
R28710 a_9432_n30006.t0 a_9432_n30006.t1 9.9005
R28711 a_n22176_n2915.t0 a_n22176_n2915.t1 19.8005
R28712 a_7452_n34534.t0 a_7452_n34534.t1 9.9005
R28713 a_n19187_n6187.t0 a_n19187_n6187.t1 19.8005
R28714 a_n19963_373.t0 a_n19963_373.t1 19.8005
R28715 a_n15014_n12716.t0 a_n15014_n12716.t1 19.8005
R28716 a_10267_n20950.t0 a_10267_n20950.t1 9.9005
R28717 a_11386_n25478.t0 a_11386_n25478.t1 9.9005
R28718 a_8496_n7266.t0 a_8496_n7266.t1 9.9005
R28719 a_11194_n7266.t0 a_11194_n7266.t1 9.9005
R28720 a_7644_n21878.t0 a_7644_n21878.t1 9.9005
R28721 a_10267_n3765.t0 a_10267_n3765.t1 9.9005
R28722 a_8592_n2838.t0 a_8592_n2838.t1 9.9005
R28723 a_11290_n2838.t0 a_11290_n2838.t1 9.9005
R28724 a_n10423_n12716.t0 a_n10423_n12716.t1 19.8005
R28725 a_10267_n16422.t0 a_10267_n16422.t1 9.9005
R28726 a_9528_762.t0 a_9528_762.t1 9.9005
R28727 a_9528_n12822.t0 a_9528_n12822.t1 9.9005
R28728 a_11386_n30006.t0 a_11386_n30006.t1 9.9005
R28729 a_9432_762.t0 a_9432_762.t1 9.9005
R28730 a_11386_n3766.t0 a_11386_n3766.t1 9.9005
R28731 a_7548_n21878.t0 a_7548_n21878.t1 9.9005
R28732 a_10459_n11894.t0 a_10459_n11894.t1 9.9005
R28733 a_8496_n17350.t0 a_8496_n17350.t1 9.9005
R28734 a_10267_763.t0 a_10267_763.t1 9.9005
R28735 a_10363_763.t0 a_10363_763.t1 9.9005
R28736 a_10267_n17349.t0 a_10267_n17349.t1 9.9005
R28737 a_10459_763.t0 a_10459_763.t1 9.9005
R28738 a_10459_n34534.t0 a_10459_n34534.t1 9.9005
R28739 a_9528_n20950.t0 a_9528_n20950.t1 9.9005
R28740 a_9336_n21878.t0 a_9336_n21878.t1 9.9005
R28741 a_11194_n17350.t0 a_11194_n17350.t1 9.9005
R28742 a_n21072_373.t0 a_n21072_373.t1 19.8005
R28743 a_8496_n30934.t0 a_8496_n30934.t1 9.9005
R28744 a_n24162_n12548.t0 a_n24162_n12548.t1 19.8005
R28745 a_10267_n30933.t0 a_10267_n30933.t1 9.9005
R28746 a_10267_n8193.t0 a_10267_n8193.t1 9.9005
R28747 a_9432_n12822.t0 a_9432_n12822.t1 9.9005
R28748 a_7644_n25478.t0 a_7644_n25478.t1 9.9005
R28749 a_11194_n30934.t0 a_11194_n30934.t1 9.9005
R28750 a_9336_n3766.t0 a_9336_n3766.t1 9.9005
R28751 a_n22426_n4727.t0 a_n22426_n4727.t1 19.8005
R28752 a_11386_n8194.t0 a_11386_n8194.t1 9.9005
R28753 a_9528_n16422.t0 a_9528_n16422.t1 9.9005
R28754 a_7548_n3766.t0 a_7548_n3766.t1 9.9005
R28755 a_10459_n2838.t0 a_10459_n2838.t1 9.9005
R28756 a_n22426_n6019.t0 a_n22426_n6019.t1 19.8005
R28757 a_7548_n25478.t0 a_7548_n25478.t1 9.9005
R28758 a_n6800_373.t0 a_n6800_373.t1 19.8005
R28759 a_7644_n30006.t0 a_7644_n30006.t1 9.9005
R28760 a_10459_n12821.t0 a_10459_n12821.t1 9.9005
R28761 a_n13714_n6187.t0 a_n13714_n6187.t1 19.8005
R28762 a_8496_n11894.t0 a_8496_n11894.t1 9.9005
R28763 a_n16672_373.t0 a_n16672_373.t1 19.8005
R28764 a_9336_n25478.t0 a_9336_n25478.t1 9.9005
R28765 a_11386_n12822.t0 a_11386_n12822.t1 9.9005
R28766 a_8496_n34534.t0 a_8496_n34534.t1 9.9005
R28767 a_11194_n11894.t0 a_11194_n11894.t1 9.9005
R28768 a_n17781_373.t0 a_n17781_373.t1 19.8005
R28769 a_9336_n8194.t0 a_9336_n8194.t1 9.9005
R28770 a_11194_n34534.t0 a_11194_n34534.t1 9.9005
R28771 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t7 485.221
R28772 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t10 367.928
R28773 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n4 227.526
R28774 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n5 227.266
R28775 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n6 227.266
R28776 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t8 224.478
R28777 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n1 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t9 213.688
R28778 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n3 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n2 84.5046
R28779 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n2 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n1 72.3005
R28780 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n3 61.0566
R28781 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t0 42.7747
R28782 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t4 30.379
R28783 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n4 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t5 30.379
R28784 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t2 30.379
R28785 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n5 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t6 30.379
R28786 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t3 30.379
R28787 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n6 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.t1 30.379
R28788 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A.n0 0.583137
R28789 a_n9314_n6187.t0 a_n9314_n6187.t1 19.8005
R28790 a_7548_n30006.t0 a_7548_n30006.t1 9.9005
R28791 a_7548_n8194.t0 a_7548_n8194.t1 9.9005
R28792 a_10459_n7266.t0 a_10459_n7266.t1 9.9005
R28793 a_n12605_n6187.t0 a_n12605_n6187.t1 19.8005
R28794 a_11386_n20950.t0 a_11386_n20950.t1 9.9005
R28795 a_9432_n3766.t0 a_9432_n3766.t1 9.9005
R28796 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t7 540.38
R28797 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t8 367.928
R28798 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n5 227.526
R28799 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t9 227.356
R28800 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n4 227.266
R28801 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n6 227.266
R28802 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n1 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t10 213.688
R28803 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n3 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n2 160.439
R28804 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n2 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n1 94.4341
R28805 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n0 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t3 42.7944
R28806 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t0 30.379
R28807 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n5 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t1 30.379
R28808 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t6 30.379
R28809 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n4 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t4 30.379
R28810 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t5 30.379
R28811 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n6 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.t2 30.379
R28812 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n0 13.4358
R28813 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B.n3 0.821842
R28814 a_9336_n30006.t0 a_9336_n30006.t1 9.9005
R28815 a_9528_n3766.t0 a_9528_n3766.t1 9.9005
R28816 a_7644_n3766.t0 a_7644_n3766.t1 9.9005
R28817 a_n8432_n6187.t0 a_n8432_n6187.t1 19.8005
R28818 a_n22425_n12548.t0 a_n22425_n12548.t1 19.8005
R28819 a_17528_n18777.t0 a_17528_n18777.t1 19.8005
R28820 a_7452_762.t0 a_7452_762.t1 9.9005
R28821 a_7644_762.t0 a_7644_762.t1 9.9005
R28822 a_n11723_n6187.t0 a_n11723_n6187.t1 19.8005
R28823 a_11386_n16422.t0 a_11386_n16422.t1 9.9005
R28824 a_7548_762.t0 a_7548_762.t1 9.9005
R28825 a_n15790_373.t0 a_n15790_373.t1 19.8005
R28826 a_9528_n26406.t0 a_9528_n26406.t1 9.9005
R28827 a_9336_762.t0 a_9336_762.t1 9.9005
R28828 a_7644_n12822.t0 a_7644_n12822.t1 9.9005
R28829 a_9432_n8194.t0 a_9432_n8194.t1 9.9005
R28830 a_9528_n35462.t0 a_9528_n35462.t1 9.9005
R28831 a_10459_n25478.t0 a_10459_n25478.t1 9.9005
R28832 a_8496_n21878.t0 a_8496_n21878.t1 9.9005
R28833 a_10267_n21877.t0 a_10267_n21877.t1 9.9005
R28834 a_7644_n20950.t0 a_7644_n20950.t1 9.9005
R28835 a_11194_n21878.t0 a_11194_n21878.t1 9.9005
R28836 a_7548_n12822.t0 a_7548_n12822.t1 9.9005
R28837 a_n20296_n6187.t0 a_n20296_n6187.t1 19.8005
C0 mux8_6.NAND4F_4.B mux8_6.NAND4F_3.Y 0.223331f
C1 mux8_5.A1 mux8_5.NAND4F_6.Y 8.98e-23
C2 mux8_3.NAND4F_9.Y Y2 7.08e-19
C3 mux8_4.NAND4F_4.Y mux8_4.NAND4F_5.Y 0.087643f
C4 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 0.012283f
C5 OR8_0.S1 mux8_2.NAND4F_3.Y 2.56e-19
C6 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 0.00162f
C7 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 0.644048f
C8 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 0.792412f
C9 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT 1.58859f
C10 V_FLAG_0.XOR2_2.B mux8_6.A0 0.060245f
C11 mux8_4.NAND4F_4.Y XOR8_0.S3 2.3e-19
C12 mux8_3.NAND4F_5.Y mux8_4.NAND4F_4.Y 0.002218f
C13 B7 B0 0.096009f
C14 MULT_0.SO mux8_1.NAND4F_8.Y 1.16e-22
C15 AND8_0.S7 B6 0.039068f
C16 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 1.58859f
C17 mux8_8.A1 SEL0 1.1712f
C18 OR8_0.S1 NOT8_0.S2 1.41e-19
C19 mux8_4.A1 AND8_0.S3 6.65362f
C20 mux8_6.NAND4F_0.C SEL1 1.13389f
C21 mux8_0.NAND4F_4.B 8bit_ADDER_0.C 1.52147f
C22 MULT_0.4bit_ADDER_0.A2 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A 0.00194f
C23 mux8_7.NAND4F_4.Y mux8_7.NAND4F_5.Y 0.087643f
C24 AND8_0.S6 OR8_0.NOT8_0.A7 0.05959f
C25 mux8_6.A1 mux8_6.NAND4F_1.Y 8.98e-23
C26 XOR8_0.S5 B7 0.082103f
C27 mux8_1.NAND4F_2.Y mux8_1.NAND4F_5.Y 4.33e-19
C28 NOT8_0.S4 mux8_5.NAND4F_4.B 0.105153f
C29 AND8_0.S1 mux8_2.NAND4F_5.Y 5.23e-19
C30 8bit_ADDER_0.S2 XOR8_0.S1 0.030205f
C31 MULT_0.4bit_ADDER_0.B2 A1 0.214949f
C32 mux8_4.NAND4F_3.Y mux8_4.NAND4F_4.Y 0.102178f
C33 mux8_4.NAND4F_0.Y mux8_4.NAND4F_8.Y 0.249057f
C34 MULT_0.4bit_ADDER_2.B2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT 0.119906f
C35 mux8_4.NAND4F_6.Y SEL0 0.353714f
C36 mux8_8.A1 mux8_8.NAND4F_4.B 0.039141f
C37 MULT_0.4bit_ADDER_1.B3 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A 0.257603f
C38 VDD Y2 0.974072f
C39 mux8_4.A0 8bit_ADDER_0.S0 0.055875f
C40 mux8_8.NAND4F_0.Y mux8_8.NAND4F_5.Y 4.32e-19
C41 NOT8_0.S6 mux8_8.NAND4F_0.Y 5.24e-19
C42 MULT_0.S2 mux8_3.NAND4F_2.D 0.107639f
C43 mux8_1.NAND4F_5.Y VDD 2.20007f
C44 mux8_7.NAND4F_4.B mux8_7.NAND4F_4.Y 0.275773f
C45 mux8_7.A0 mux8_3.NAND4F_0.C 1.67e-19
C46 mux8_1.NAND4F_9.Y SEL0 2.8e-19
C47 MULT_0.4bit_ADDER_1.A2 MULT_0.inv_9.Y 0.001794f
C48 NOT8_0.S7 mux8_6.NAND4F_0.Y 5.24e-19
C49 mux8_3.NAND4F_6.Y SEL0 0.353735f
C50 mux8_2.NAND4F_5.Y mux8_2.NAND4F_1.Y 0.110562f
C51 XOR8_0.S7 mux8_6.NAND4F_6.Y 0.520706f
C52 mux8_6.NAND4F_4.Y mux8_6.NAND4F_1.Y 4.33e-19
C53 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT A1 0.003441f
C54 XOR8_0.S5 SEL0 0.16904f
C55 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A 0.118063f
C56 NOT8_0.S7 B6 0.465474f
C57 mux8_5.NAND4F_0.C mux8_7.NAND4F_0.C 0.001594f
C58 mux8_7.A0 mux8_7.NAND4F_3.Y 0.406267f
C59 NOT8_0.S5 NOT8_0.S6 1.65673f
C60 Y4 Y7 0.023368f
C61 Y5 Y6 3.20366f
C62 mux8_1.NAND4F_4.B mux8_1.NAND4F_6.Y 0.187883f
C63 8bit_ADDER_0.S2 mux8_3.NAND4F_2.D 0.105158f
C64 OR8_0.S7 mux8_6.NAND4F_2.Y 0.402593f
C65 OR8_0.NOT8_0.A3 A2 0.205927f
C66 AND8_0.S1 B1 0.037104f
C67 mux8_2.NAND4F_0.Y mux8_2.NAND4F_4.Y 0.28646f
C68 mux8_2.NAND4F_3.Y mux8_2.NAND4F_2.Y 1.63543f
C69 mux8_2.NAND4F_0.C mux8_2.NAND4F_5.Y 0.051024f
C70 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A 8.33e-19
C71 left_shifter_0.S0 XOR8_0.S2 0.025839f
C72 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A SEL3 6.99e-19
C73 mux8_2.NAND4F_4.B XOR8_0.S1 0.96335f
C74 NOT8_0.S3 B5 0.004141f
C75 mux8_7.A1 XOR8_0.S4 2.06613f
C76 A7 B7 51.2456f
C77 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A 0.248556f
C78 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B 0.209959f
C79 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A 8bit_ADDER_0.S2 0.200037f
C80 mux8_2.NAND4F_4.Y mux8_2.NAND4F_7.Y 4.32e-19
C81 XOR8_0.S1 A1 0.558628f
C82 NOT8_0.S4 mux8_5.NAND4F_0.Y 5.24e-19
C83 mux8_7.NAND4F_2.Y XOR8_0.S5 1.49e-19
C84 mux8_7.NAND4F_4.B mux8_7.NAND4F_5.Y 0.248856f
C85 mux8_8.NAND4F_5.Y VDD 2.19984f
C86 NOT8_0.S6 VDD 0.946576f
C87 mux8_4.A0 left_shifter_0.S0 0.016512f
C88 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A mux8_6.A1 0.186718f
C89 mux8_1.NAND4F_3.Y NOT8_0.S0 3.24e-22
C90 OR8_0.S7 A2 0.01362f
C91 mux8_8.A0 XOR8_0.S1 0.025513f
C92 MULT_0.S2 mux8_3.NAND4F_6.Y 8.98e-23
C93 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A 2.56e-19
C94 mux8_4.NAND4F_4.B AND8_0.S3 1.04047f
C95 mux8_4.A0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 0.007337f
C96 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A 0.001379f
C97 VDD A0 13.4333f
C98 mux8_7.NAND4F_0.C mux8_7.NAND4F_0.Y 0.223896f
C99 mux8_0.NAND4F_4.B mux8_0.NAND4F_1.Y 0.222551f
C100 MULT_0.inv_9.Y A1 0.009951f
C101 MULT_0.S2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B 0.005184f
C102 mux8_2.NAND4F_0.C mux8_3.NAND4F_0.C 0.001477f
C103 mux8_7.A1 mux8_6.A1 1.83e-20
C104 AND8_0.S3 AND8_0.NOT8_0.A2 0.266381f
C105 mux8_6.NAND4F_4.B mux8_6.NAND4F_1.Y 0.222551f
C106 mux8_6.A0 NOT8_0.S6 0.026415f
C107 mux8_8.NAND4F_0.Y SEL2 2.97e-20
C108 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B VDD 1.8288f
C109 mux8_0.NAND4F_1.Y mux8_0.NAND4F_7.Y 0.617483f
C110 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A VDD 1.35225f
C111 AND8_0.NOT8_0.A0 AND8_0.NOT8_0.A2 1.5e-19
C112 mux8_3.NAND4F_4.Y mux8_3.NAND4F_1.Y 4.33e-19
C113 mux8_6.NAND4F_7.Y SEL0 0.234594f
C114 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT A3 0.003441f
C115 mux8_0.NAND4F_0.C SEL0 12.4679f
C116 mux8_6.A0 A0 0.004911f
C117 mux8_0.NAND4F_2.Y mux8_0.NAND4F_9.Y 2.96e-20
C118 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B 0.008371f
C119 mux8_5.NAND4F_4.B mux8_5.NAND4F_3.Y 0.223331f
C120 8bit_ADDER_0.S2 mux8_3.NAND4F_6.Y 2.97e-22
C121 mux8_0.NAND4F_4.Y mux8_0.NAND4F_5.Y 0.087643f
C122 mux8_4.NAND4F_0.C mux8_4.NAND4F_4.Y 0.049743f
C123 mux8_5.NAND4F_4.B XOR8_0.S4 0.963496f
C124 mux8_3.NAND4F_3.Y NOT8_0.S2 3.24e-22
C125 mux8_8.A0 mux8_3.NAND4F_2.D 1.11e-19
C126 8bit_ADDER_0.S0 AND8_0.S0 0.059486f
C127 NOT8_0.S5 SEL2 0.122807f
C128 NOT8_0.S1 VDD 0.984917f
C129 mux8_3.NAND4F_9.Y SEL2 1.49e-20
C130 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 0.001075f
C131 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A A1 0.008956f
C132 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y B0 0.005392f
C133 mux8_5.NAND4F_1.Y SEL1 2.35e-20
C134 mux8_6.NAND4F_2.D SEL0 0.147146f
C135 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y B0 0.005392f
C136 NOT8_0.S5 mux8_7.NAND4F_1.Y 0.55011f
C137 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y B0 0.005392f
C138 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y B0 0.122687f
C139 mux8_5.NAND4F_2.Y SEL2 3.61e-20
C140 mux8_7.A0 AND8_0.S3 0.020481f
C141 mux8_5.NAND4F_8.Y mux8_5.NAND4F_6.Y 2.96e-20
C142 mux8_7.A1 AND8_0.S5 2.06602f
C143 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A mux8_8.A0 1.08e-19
C144 A6 A0 0.02576f
C145 B0 A4 0.033653f
C146 mux8_8.NAND4F_0.C mux8_6.NAND4F_0.C 0.001594f
C147 mux8_6.A0 NOT8_0.S1 0.017056f
C148 mux8_8.NAND4F_8.Y mux8_8.NAND4F_6.Y 2.96e-20
C149 mux8_1.NAND4F_2.Y SEL2 3.61e-20
C150 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_1.A2 7.1e-19
C151 OR8_0.S2 SEL0 1.09976f
C152 XOR8_0.S5 A4 0.033738f
C153 MULT_0.inv_15.Y VDD 1.9283f
C154 VDD SEL2 11.024f
C155 mux8_8.NAND4F_4.Y SEL1 0.30433f
C156 AND8_0.S6 mux8_8.NAND4F_4.Y 0.402481f
C157 mux8_2.NAND4F_4.Y SEL0 0.116692f
C158 NOT8_0.S3 B6 9.03e-21
C159 AND8_0.S4 left_shifter_0.S7 0.227279f
C160 mux8_7.NAND4F_1.Y VDD 2.1816f
C161 SEL3 A3 0.256157f
C162 mux8_8.A0 mux8_8.A1 4.73956f
C163 mux8_3.NAND4F_0.Y mux8_3.NAND4F_3.Y 0.616159f
C164 B0 A1 2.05905f
C165 mux8_4.NAND4F_9.Y mux8_4.NAND4F_7.Y 0.248336f
C166 AND8_0.S1 AND8_0.S3 1.49e-19
C167 mux8_2.NAND4F_9.Y mux8_2.NAND4F_5.Y 0.402985f
C168 OR8_0.NOT8_0.A2 A2 0.332742f
C169 mux8_6.NAND4F_3.Y mux8_6.NAND4F_8.Y 0.222524f
C170 mux8_5.NAND4F_0.Y mux8_5.NAND4F_3.Y 0.616159f
C171 mux8_6.A0 SEL2 0.988007f
C172 AND8_0.S1 AND8_0.NOT8_0.A0 0.266264f
C173 B2 A2 45.9863f
C174 MULT_0.4bit_ADDER_1.B3 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT 0.004585f
C175 mux8_0.NAND4F_2.D VDD 1.39778f
C176 AND8_0.S0 left_shifter_0.S0 0.009169f
C177 mux8_4.NAND4F_2.D mux8_4.NAND4F_0.Y 0.184536f
C178 XOR8_0.S2 A0 5.26e-19
C179 AND8_0.S6 B7 0.055265f
C180 AND8_0.NOT8_0.A1 AND8_0.NOT8_0.A2 1.81366f
C181 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B 1.2618f
C182 NOT8_0.S6 AND8_0.S7 0.222534f
C183 mux8_4.NAND4F_0.Y NOT8_0.S3 5.24e-19
C184 mux8_8.A0 XOR8_0.S5 0.050803f
C185 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y A7 2.72778f
C186 mux8_1.NAND4F_0.Y mux8_1.NAND4F_3.Y 0.616159f
C187 mux8_2.NAND4F_5.Y mux8_3.NAND4F_4.Y 0.002062f
C188 V_FLAG_0.XOR2_0.Y V 3.99e-19
C189 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A 1.01138f
C190 AND8_0.S3 AND8_0.NOT8_0.A4 6.32e-21
C191 A7 A4 0.079269f
C192 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A A3 0.008956f
C193 mux8_5.NAND4F_4.B AND8_0.S5 0.001198f
C194 NOT8_0.S5 mux8_7.NAND4F_9.Y 3.17e-20
C195 NOT8_0.S4 mux8_5.NAND4F_5.Y 0.288211f
C196 mux8_4.A0 A0 1.23e-19
C197 SEL1 SEL0 33.598602f
C198 AND8_0.S6 SEL0 0.12865f
C199 mux8_2.NAND4F_3.Y XOR8_0.S1 5.23e-19
C200 OR8_0.NOT8_0.A5 B4 0.037481f
C201 MULT_0.S2 OR8_0.S2 0.283233f
C202 mux8_3.NAND4F_2.Y SEL0 0.296538f
C203 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT SEL3 1.92e-19
C204 AND8_0.NOT8_0.A5 VDD 2.28564f
C205 mux8_4.A0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 0.005184f
C206 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A 8.34e-19
C207 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A A1 0.006225f
C208 XOR8_0.S1 NOT8_0.S2 2.29e-19
C209 NOT8_0.S1 XOR8_0.S2 0.020433f
C210 mux8_8.NAND4F_4.B SEL1 4.36064f
C211 MULT_0.S2 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A 0.002364f
C212 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT 0.001576f
C213 AND8_0.S6 mux8_8.NAND4F_4.B 1.04047f
C214 OR8_0.NOT8_0.A0 A0 0.310325f
C215 A7 A1 0.04706f
C216 8bit_ADDER_0.C SEL0 0.672462f
C217 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A VDD 1.66874f
C218 NOT8_0.S6 NOT8_0.S7 2.17011f
C219 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 8bit_ADDER_0.S2 0.716167f
C220 XOR8_0.S6 B3 5.28e-19
C221 mux8_0.NAND4F_2.D mux8_0.NAND4F_8.Y 4.88e-20
C222 ZFLAG_0.nor4_1.Y Y6 0.045114f
C223 mux8_3.NAND4F_0.C mux8_3.NAND4F_4.Y 0.049743f
C224 mux8_7.NAND4F_9.Y VDD 2.28759f
C225 AND8_0.S4 OR8_0.NOT8_0.A4 0.036355f
C226 mux8_5.NAND4F_0.Y mux8_5.NAND4F_7.Y 0.08762f
C227 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A 5.18e-20
C228 AND8_0.S4 A3 0.337327f
C229 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT mux8_6.A1 0.127992f
C230 8bit_ADDER_0.S2 OR8_0.S2 0.059957f
C231 mux8_4.A0 NOT8_0.S1 0.017991f
C232 AND8_0.S0 mux8_1.NAND4F_5.Y 5.23e-19
C233 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A 0.005938f
C234 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 0.119902f
C235 mux8_7.NAND4F_2.Y SEL1 0.222331f
C236 mux8_5.NAND4F_9.Y mux8_5.NAND4F_6.Y 0.222562f
C237 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 0.511769f
C238 OR8_0.NOT8_0.A2 OR8_0.NOT8_0.A3 0.221546f
C239 XOR8_0.S2 SEL2 0.196197f
C240 B3 A5 0.021359f
C241 OR8_0.NOT8_0.A3 B2 0.004191f
C242 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 2.43e-19
C243 mux8_4.A1 SEL0 1.17111f
C244 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A 0.186684f
C245 mux8_3.NAND4F_2.D NOT8_0.S2 4.43e-19
C246 mux8_6.NAND4F_3.Y VDD 2.17571f
C247 AND8_0.S1 AND8_0.NOT8_0.A1 0.396894f
C248 XOR8_0.S3 NOT8_0.S5 0.318864f
C249 mux8_4.NAND4F_2.Y mux8_4.NAND4F_9.Y 2.96e-20
C250 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT VDD 3.5013f
C251 mux8_3.NAND4F_9.Y mux8_3.NAND4F_5.Y 0.402985f
C252 mux8_0.NAND4F_3.Y VDD 2.17543f
C253 MULT_0.S2 SEL1 0.070061f
C254 AND8_0.NOT8_0.A5 A6 5.25e-21
C255 AND8_0.S7 SEL2 0.02143f
C256 mux8_4.A0 SEL2 0.647036f
C257 MULT_0.4bit_ADDER_1.B3 MULT_0.4bit_ADDER_1.A2 0.120212f
C258 MULT_0.S2 mux8_3.NAND4F_2.Y 1.16938f
C259 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B 0.007216f
C260 XOR8_0.S0 SEL0 0.168116f
C261 OR8_0.S7 B2 8.55e-19
C262 8bit_ADDER_0.S0 mux8_1.NAND4F_4.Y 0.047022f
C263 mux8_6.A0 mux8_6.NAND4F_3.Y 0.406267f
C264 mux8_8.NAND4F_8.Y mux8_8.NAND4F_9.Y 0.696806f
C265 mux8_4.NAND4F_5.Y VDD 2.19962f
C266 mux8_6.A1 mux8_6.NAND4F_2.Y 1.16938f
C267 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT A1 0.129004f
C268 AND8_0.NOT8_0.A1 AND8_0.NOT8_0.A4 7.07e-22
C269 mux8_1.NAND4F_7.Y mux8_2.NAND4F_8.Y 1.02e-21
C270 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B 0.087175f
C271 mux8_2.NAND4F_4.B mux8_2.NAND4F_4.Y 0.275773f
C272 8bit_ADDER_0.S0 mux8_1.NAND4F_1.Y 5.23e-19
C273 XOR8_0.S3 VDD 1.60555f
C274 mux8_3.NAND4F_5.Y VDD 2.19984f
C275 mux8_8.NAND4F_0.C mux8_8.NAND4F_4.Y 0.049743f
C276 8bit_ADDER_0.S2 SEL1 0.339028f
C277 mux8_8.A1 NOT8_0.S2 0.114085f
C278 mux8_1.NAND4F_2.D mux8_1.NAND4F_3.Y 0.397922f
C279 OR8_0.S2 A1 0.01629f
C280 mux8_6.NAND4F_0.Y mux8_6.NAND4F_9.Y 2.96e-20
C281 mux8_3.NAND4F_2.D mux8_3.NAND4F_0.Y 0.184536f
C282 8bit_ADDER_0.S2 mux8_3.NAND4F_2.Y 0.200461f
C283 mux8_1.NAND4F_9.Y mux8_2.NAND4F_3.Y 1.02e-21
C284 mux8_5.NAND4F_3.Y mux8_5.NAND4F_5.Y 4.33e-19
C285 NOT8_0.S7 SEL2 0.052754f
C286 mux8_4.NAND4F_3.Y VDD 2.17571f
C287 mux8_6.NAND4F_2.Y mux8_6.NAND4F_4.Y 2.04463f
C288 mux8_4.NAND4F_4.Y mux8_4.NAND4F_7.Y 4.32e-19
C289 OR8_0.NOT8_0.A5 B5 0.0271f
C290 AND8_0.S0 A0 0.054687f
C291 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A SEL3 6.99e-19
C292 mux8_8.A0 OR8_0.S2 0.024803f
C293 OR8_0.NOT8_0.A1 A0 0.242779f
C294 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.A2 0.001881f
C295 mux8_6.A1 A2 0.854441f
C296 XOR8_0.S4 mux8_5.NAND4F_5.Y 0.602406f
C297 mux8_6.A0 XOR8_0.S3 0.031775f
C298 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A MULT_0.inv_9.Y 0.001139f
C299 mux8_0.NAND4F_1.Y SEL0 0.339784f
C300 MULT_0.S2 mux8_4.A1 0.018575f
C301 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B 0.001328f
C302 8bit_ADDER_0.C 8bit_ADDER_0.S2 0.169203f
C303 NOT8_0.S2 B0 0.229233f
C304 mux8_0.NAND4F_2.Y mux8_0.NAND4F_4.Y 2.04463f
C305 mux8_0.NAND4F_3.Y mux8_0.NAND4F_8.Y 0.222524f
C306 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A 0.127125f
C307 NOT8_0.S2 mux8_3.NAND4F_6.Y 0.79864f
C308 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A 8bit_ADDER_0.S2 7.38e-19
C309 mux8_7.NAND4F_4.Y mux8_7.NAND4F_7.Y 4.32e-19
C310 AND8_0.S6 A4 0.354428f
C311 XOR8_0.S6 B4 0.136287f
C312 mux8_2.NAND4F_0.Y mux8_2.NAND4F_1.Y 5.28e-20
C313 AND8_0.NOT8_0.A5 AND8_0.S7 1.15e-19
C314 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 8bit_ADDER_0.C 0.002397f
C315 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_1.B0 9.98e-20
C316 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 8bit_ADDER_0.C 0.002397f
C317 mux8_8.A1 mux8_8.NAND4F_8.Y 1.16e-22
C318 XOR8_0.S0 MULT_0.S2 0.024477f
C319 mux8_4.NAND4F_4.B SEL0 1.61022f
C320 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 8bit_ADDER_0.C 0.002397f
C321 mux8_8.NAND4F_0.Y mux8_8.NAND4F_7.Y 0.08762f
C322 mux8_1.NAND4F_7.Y VDD 2.14088f
C323 mux8_1.NAND4F_4.Y left_shifter_0.S0 5.23e-19
C324 mux8_2.NAND4F_4.B SEL1 4.36079f
C325 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y 8bit_ADDER_0.C 0.107163f
C326 MULT_0.4bit_ADDER_1.B3 A1 0.076319f
C327 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y VDD 1.58634f
C328 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A 0.248956f
C329 mux8_5.A0 mux8_5.NAND4F_2.Y 0.200461f
C330 mux8_7.NAND4F_4.Y mux8_7.NAND4F_8.Y 0.404949f
C331 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y VDD 1.58635f
C332 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A 0.001379f
C333 mux8_8.NAND4F_0.C SEL0 12.484799f
C334 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y VDD 1.58591f
C335 AND8_0.S0 NOT8_0.S1 7.01e-20
C336 mux8_4.A0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 0.002366f
C337 8bit_ADDER_0.C A4 0.036554f
C338 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y VDD 1.58864f
C339 mux8_2.NAND4F_1.Y mux8_2.NAND4F_7.Y 0.617483f
C340 B4 A5 0.056561f
C341 SEL3 B0 1.85665f
C342 AND8_0.S5 A2 0.03008f
C343 mux8_2.NAND4F_0.C mux8_2.NAND4F_0.Y 0.223896f
C344 mux8_3.NAND4F_8.Y mux8_3.NAND4F_9.Y 0.696806f
C345 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B VDD 1.8288f
C346 mux8_5.A0 VDD 1.46858f
C347 mux8_8.NAND4F_2.D mux8_8.NAND4F_0.Y 0.184536f
C348 mux8_8.NAND4F_0.C mux8_8.NAND4F_4.B 2.13077f
C349 V_FLAG_0.XOR2_2.Y V 0.001141f
C350 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT A3 0.129004f
C351 mux8_1.NAND4F_6.Y OR8_0.S1 1.02e-21
C352 8bit_ADDER_0.S2 XOR8_0.S0 0.022861f
C353 mux8_8.A0 SEL1 0.334092f
C354 mux8_7.NAND4F_6.Y SEL2 0.419676f
C355 mux8_5.NAND4F_6.Y mux8_5.NAND4F_1.Y 2.45057f
C356 mux8_5.NAND4F_5.Y mux8_5.NAND4F_7.Y 0.235079f
C357 mux8_8.A0 AND8_0.S6 0.135403f
C358 NOT8_0.S4 B2 2.89e-19
C359 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 0.01866f
C360 mux8_6.NAND4F_1.Y VDD 2.18132f
C361 OR8_0.NOT8_0.A2 B2 0.051675f
C362 8bit_ADDER_0.C A1 0.042413f
C363 mux8_2.NAND4F_0.C mux8_2.NAND4F_7.Y 0.224691f
C364 mux8_6.NAND4F_4.B mux8_6.NAND4F_2.Y 0.112019f
C365 AND8_0.S0 MULT_0.inv_15.Y 1.78e-19
C366 mux8_7.NAND4F_6.Y mux8_7.NAND4F_1.Y 2.45057f
C367 AND8_0.S0 SEL2 0.066981f
C368 mux8_7.NAND4F_5.Y mux8_7.NAND4F_7.Y 0.235079f
C369 mux8_4.NAND4F_8.Y mux8_4.NAND4F_5.Y 0.001122f
C370 B3 B1 0.083105f
C371 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_2.B1 0.019641f
C372 OR8_0.S1 mux8_2.NAND4F_2.Y 0.402593f
C373 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A A1 0.685441f
C374 XOR8_0.S4 OR8_0.S7 0.102447f
C375 mux8_6.A0 mux8_5.A0 0.032998f
C376 8bit_ADDER_0.C mux8_8.A0 0.229998f
C377 XOR8_0.S2 mux8_3.NAND4F_5.Y 0.602392f
C378 mux8_6.A1 OR8_0.NOT8_0.A3 0.149096f
C379 mux8_3.NAND4F_8.Y VDD 3.39068f
C380 mux8_7.A0 SEL0 0.675782f
C381 mux8_8.NAND4F_7.Y VDD 2.14052f
C382 MULT_0.SO SEL0 1.17077f
C383 mux8_6.A0 mux8_6.NAND4F_1.Y 5.23e-19
C384 mux8_7.NAND4F_8.Y mux8_7.NAND4F_5.Y 0.001122f
C385 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A mux8_8.A0 1.08e-19
C386 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y A6 2.7267f
C387 mux8_1.NAND4F_4.Y mux8_1.NAND4F_5.Y 0.087643f
C388 mux8_0.NAND4F_0.C mux8_1.NAND4F_4.B 0.002598f
C389 mux8_4.A0 mux8_4.NAND4F_5.Y 2.08e-19
C390 mux8_4.NAND4F_2.Y mux8_4.NAND4F_4.Y 2.04463f
C391 mux8_4.NAND4F_3.Y mux8_4.NAND4F_8.Y 0.222524f
C392 AND8_0.S2 mux8_5.A1 0.014518f
C393 XOR8_0.S3 AND8_0.S7 0.165168f
C394 mux8_8.NAND4F_3.Y mux8_8.NAND4F_5.Y 4.33e-19
C395 mux8_4.NAND4F_0.C VDD 1.39701f
C396 mux8_4.A0 XOR8_0.S3 0.009216f
C397 NOT8_0.S6 mux8_8.NAND4F_3.Y 3.24e-22
C398 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT mux8_7.A0 0.152872f
C399 mux8_1.NAND4F_5.Y mux8_1.NAND4F_1.Y 0.110562f
C400 mux8_8.A1 AND8_0.S4 0.02448f
C401 NOT8_0.S7 mux8_6.NAND4F_3.Y 3.24e-22
C402 A7 SEL3 0.108426f
C403 mux8_8.A0 mux8_4.A1 0.047055f
C404 mux8_8.NAND4F_2.D VDD 1.37792f
C405 MULT_0.4bit_ADDER_1.B1 VDD 1.98218f
C406 mux8_6.A1 OR8_0.S7 0.334678f
C407 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 0.132282f
C408 MULT_0.4bit_ADDER_2.B1 mux8_7.A1 0.018669f
C409 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A mux8_5.A1 0.001005f
C410 mux8_4.NAND4F_2.D SEL2 0.481923f
C411 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A 0.118063f
C412 AND8_0.S1 SEL0 0.128375f
C413 MULT_0.4bit_ADDER_2.B2 mux8_6.A1 0.012283f
C414 mux8_4.A0 mux8_4.NAND4F_3.Y 0.406267f
C415 mux8_1.NAND4F_6.Y mux8_2.NAND4F_2.Y 0.0024f
C416 mux8_7.A1 NOT8_0.S5 0.019926f
C417 NOT8_0.S3 SEL2 0.09821f
C418 XOR8_0.S6 B5 0.157786f
C419 mux8_7.A0 mux8_7.NAND4F_2.Y 0.200461f
C420 mux8_8.A0 XOR8_0.S0 0.024063f
C421 mux8_2.NAND4F_1.Y SEL0 0.339784f
C422 mux8_6.A0 mux8_8.NAND4F_2.D 0.001114f
C423 left_shifter_0.S7 mux8_6.NAND4F_5.Y 0.402437f
C424 OR8_0.S7 mux8_6.NAND4F_4.Y 0.526611f
C425 ZFLAG_0.nor4_0.Y Y0 0.595568f
C426 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT 1.58859f
C427 mux8_2.NAND4F_3.Y mux8_2.NAND4F_4.Y 0.102178f
C428 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A VDD 1.34488f
C429 XOR8_0.S3 NOT8_0.S7 0.044014f
C430 mux8_5.NAND4F_6.Y SEL0 0.353719f
C431 OR8_0.S2 NOT8_0.S2 0.001232f
C432 mux8_7.NAND4F_9.Y mux8_7.NAND4F_6.Y 0.222562f
C433 mux8_7.A0 MULT_0.S2 0.024275f
C434 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B 0.209959f
C435 B5 A5 48.7118f
C436 mux8_0.NAND4F_5.Y VDD 2.19984f
C437 mux8_1.NAND4F_4.B mux8_2.NAND4F_4.Y 1.02e-21
C438 OR8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B 7.29e-19
C439 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A A3 0.685441f
C440 mux8_5.A0 XOR8_0.S2 0.022511f
C441 mux8_7.A1 VDD 1.21165f
C442 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y mux8_4.A0 2.76e-19
C443 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y mux8_4.A0 0.018656f
C444 NOT8_0.S4 mux8_5.NAND4F_3.Y 3.24e-22
C445 mux8_7.NAND4F_4.Y XOR8_0.S5 2.3e-19
C446 AND8_0.S5 OR8_0.S7 0.026409f
C447 mux8_2.NAND4F_0.C SEL0 12.9172f
C448 mux8_1.NAND4F_2.Y NOT8_0.S0 1.43e-19
C449 NOT8_0.S4 XOR8_0.S4 10.0763f
C450 mux8_2.NAND4F_0.Y mux8_2.NAND4F_9.Y 2.96e-20
C451 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT SEL3 1.92e-19
C452 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.inv_9.Y 0.002003f
C453 MULT_0.4bit_ADDER_0.A2 A1 0.173675f
C454 NOT8_0.S0 VDD 0.973991f
C455 AND8_0.NOT8_0.A6 AND8_0.S6 0.393091f
C456 B4 B1 0.021378f
C457 mux8_7.NAND4F_0.C mux8_7.NAND4F_3.Y 0.399921f
C458 mux8_5.A0 mux8_4.A0 10.5707f
C459 mux8_7.A0 8bit_ADDER_0.S2 2.14e-19
C460 mux8_6.A0 mux8_7.A1 0.028646f
C461 8bit_ADDER_0.S2 MULT_0.SO 0.015825f
C462 AND8_0.S1 MULT_0.S2 0.022274f
C463 mux8_2.NAND4F_2.D mux8_2.NAND4F_8.Y 4.88e-20
C464 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 8bit_ADDER_0.S2 0.01942f
C465 mux8_5.NAND4F_6.Y mux8_7.NAND4F_2.Y 0.002218f
C466 mux8_8.NAND4F_3.Y SEL2 2.96e-20
C467 mux8_2.NAND4F_9.Y mux8_2.NAND4F_7.Y 0.248336f
C468 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A VDD 1.66874f
C469 AND8_0.NOT8_0.A2 A1 0.1594f
C470 AND8_0.S3 B3 0.059452f
C471 mux8_7.NAND4F_1.Y mux8_8.NAND4F_3.Y 0.002218f
C472 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y mux8_7.A0 1.53e-19
C473 mux8_3.NAND4F_0.C AND8_0.S2 0.037277f
C474 AND8_0.S2 B1 0.042801f
C475 mux8_6.A0 NOT8_0.S0 0.014029f
C476 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y mux8_7.A0 1.53e-19
C477 mux8_1.NAND4F_4.B SEL1 4.36064f
C478 mux8_0.NAND4F_4.Y mux8_0.NAND4F_9.Y 5.28e-19
C479 AND8_0.NOT8_0.A0 B3 0.001171f
C480 mux8_5.NAND4F_4.B mux8_5.NAND4F_2.Y 0.112019f
C481 NOT8_0.S2 SEL1 0.074941f
C482 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 0.00162f
C483 mux8_0.NAND4F_8.Y mux8_0.NAND4F_5.Y 0.001122f
C484 mux8_6.A1 NOT8_0.S4 0.040875f
C485 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 0.511769f
C486 mux8_8.A0 mux8_8.NAND4F_0.C 0.084171f
C487 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A mux8_7.A0 0.200037f
C488 OR8_0.S7 mux8_6.NAND4F_4.B 0.079695f
C489 Y2 Y3 1.32577f
C490 mux8_6.A1 OR8_0.NOT8_0.A2 0.06222f
C491 mux8_7.A0 A4 0.431687f
C492 8bit_ADDER_0.S2 AND8_0.S1 0.031696f
C493 mux8_3.NAND4F_2.Y NOT8_0.S2 1.43e-19
C494 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 1.58859f
C495 XOR8_0.S5 mux8_7.NAND4F_5.Y 0.602392f
C496 mux8_6.A1 B2 0.223574f
C497 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B 0.792412f
C498 mux8_1.NAND4F_0.C mux8_2.NAND4F_0.Y 9.03e-22
C499 mux8_5.NAND4F_4.B VDD 1.19888f
C500 mux8_8.NAND4F_5.Y mux8_8.NAND4F_1.Y 0.110562f
C501 V_FLAG_0.XOR2_0.Y VDD 0.933222f
C502 NOT8_0.S6 mux8_8.NAND4F_1.Y 0.55011f
C503 NOT8_0.S4 mux8_5.NAND4F_7.Y 0.431664f
C504 mux8_5.NAND4F_4.Y SEL2 8.74e-20
C505 NOT8_0.S7 mux8_6.NAND4F_1.Y 0.55011f
C506 mux8_4.A0 mux8_4.NAND4F_0.C 0.099535f
C507 mux8_7.NAND4F_4.B XOR8_0.S5 0.96335f
C508 mux8_5.NAND4F_0.C SEL2 1.4681f
C509 XOR8_0.S6 B6 0.30186f
C510 mux8_2.NAND4F_2.D VDD 1.37507f
C511 mux8_1.NAND4F_4.Y SEL2 8.74e-20
C512 mux8_7.A0 A1 6.44e-20
C513 OR8_0.S1 XOR8_0.S1 14.392499f
C514 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B 1.2618f
C515 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A MULT_0.inv_9.Y 0.019351f
C516 SEL3 SEL1 1.44e-20
C517 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT A1 0.010334f
C518 mux8_6.A0 V_FLAG_0.XOR2_0.Y 0.566275f
C519 mux8_1.NAND4F_1.Y SEL2 0.37854f
C520 mux8_4.NAND4F_2.D mux8_4.NAND4F_5.Y 9.34e-20
C521 NOT8_0.S4 AND8_0.S5 0.358937f
C522 mux8_4.A1 NOT8_0.S2 0.025378f
C523 B6 A5 29.372f
C524 8bit_ADDER_0.S2 mux8_2.NAND4F_0.C 3.31e-19
C525 mux8_8.A0 mux8_7.A0 9.321071f
C526 mux8_2.NAND4F_4.B AND8_0.S1 1.04047f
C527 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A 0.009176f
C528 mux8_8.A0 MULT_0.SO 0.02831f
C529 OR8_0.S1 MULT_0.inv_9.Y 1.69e-20
C530 mux8_3.NAND4F_0.Y mux8_3.NAND4F_2.Y 0.170507f
C531 mux8_7.A1 XOR8_0.S2 0.158511f
C532 mux8_6.A0 mux8_2.NAND4F_2.D 9.02e-20
C533 mux8_4.NAND4F_2.D XOR8_0.S3 4.4e-19
C534 NOT8_0.S3 mux8_4.NAND4F_5.Y 0.288211f
C535 OR8_0.NOT8_0.A4 A3 0.264441f
C536 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT mux8_8.A0 5.1e-19
C537 AND8_0.S5 B2 0.028098f
C538 8bit_ADDER_0.C SEL3 0.218848f
C539 XOR8_0.S0 mux8_2.NAND4F_3.Y 1.02e-21
C540 OR8_0.S2 AND8_0.S4 0.003669f
C541 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B 0.007216f
C542 mux8_5.NAND4F_0.Y mux8_5.NAND4F_2.Y 0.170507f
C543 mux8_6.NAND4F_2.Y mux8_6.NAND4F_8.Y 0.222339f
C544 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT 0.012283f
C545 XOR8_0.S3 NOT8_0.S3 5.98547f
C546 AND8_0.S1 A1 0.040754f
C547 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A SEL3 6.99e-19
C548 mux8_6.NAND4F_0.C XOR8_0.S7 0.094395f
C549 8bit_ADDER_0.S2 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 0.006051f
C550 AND8_0.NOT8_0.A4 A4 0.954517f
C551 mux8_2.NAND4F_4.B mux8_2.NAND4F_1.Y 0.222551f
C552 mux8_1.NAND4F_4.B XOR8_0.S0 0.963376f
C553 mux8_5.NAND4F_3.Y XOR8_0.S4 5.23e-19
C554 mux8_4.NAND4F_0.Y mux8_4.NAND4F_1.Y 5.28e-20
C555 mux8_4.NAND4F_2.D mux8_4.NAND4F_3.Y 0.397922f
C556 XOR8_0.S0 NOT8_0.S2 1.01e-19
C557 NOT8_0.S0 XOR8_0.S2 0.032144f
C558 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B 0.005184f
C559 mux8_6.NAND4F_6.Y SEL2 0.419676f
C560 mux8_2.NAND4F_9.Y SEL0 2.8e-19
C561 B5 B1 0.020952f
C562 AND8_0.S5 mux8_7.NAND4F_2.D 0.097092f
C563 mux8_7.NAND4F_0.Y SEL2 2.97e-20
C564 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A 1.01138f
C565 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A 8bit_ADDER_0.S2 4.24e-19
C566 mux8_5.NAND4F_0.Y VDD 2.13487f
C567 mux8_8.A0 AND8_0.S1 0.016924f
C568 mux8_6.NAND4F_9.Y SEL2 1.49e-20
C569 mux8_3.NAND4F_9.Y mux8_3.NAND4F_7.Y 0.248336f
C570 OR8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A 1.07e-19
C571 mux8_4.NAND4F_3.Y NOT8_0.S3 3.24e-22
C572 mux8_5.A0 AND8_0.S0 0.012292f
C573 mux8_1.NAND4F_0.Y mux8_1.NAND4F_2.Y 0.170507f
C574 AND8_0.NOT8_0.A1 B3 0.053928f
C575 mux8_7.NAND4F_0.Y mux8_7.NAND4F_1.Y 5.28e-20
C576 mux8_1.NAND4F_0.Y VDD 2.21066f
C577 AND8_0.S3 B4 0.007432f
C578 mux8_4.A0 NOT8_0.S0 0.013094f
C579 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A mux8_8.A1 4.9e-19
C580 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B 0.007216f
C581 mux8_2.NAND4F_0.C mux8_2.NAND4F_4.B 2.13077f
C582 mux8_2.NAND4F_2.Y XOR8_0.S1 1.49e-19
C583 mux8_8.NAND4F_1.Y SEL2 0.37854f
C584 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A 0.001379f
C585 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A 0.009047f
C586 mux8_4.NAND4F_7.Y VDD 2.14052f
C587 MULT_0.4bit_ADDER_0.B2 A3 0.381547f
C588 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B 0.001328f
C589 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT VDD 3.30054f
C590 mux8_3.NAND4F_4.Y SEL0 0.116487f
C591 OR8_0.S1 mux8_8.A1 0.03966f
C592 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A 2.56e-19
C593 mux8_3.NAND4F_7.Y VDD 2.14052f
C594 AND8_0.S2 AND8_0.S3 1.87639f
C595 mux8_6.A1 XOR8_0.S4 0.032804f
C596 AND8_0.S4 SEL1 0.111612f
C597 AND8_0.S4 AND8_0.S6 0.004135f
C598 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT A3 0.010334f
C599 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B VDD 1.8288f
C600 AND8_0.S2 AND8_0.NOT8_0.A0 1.3e-19
C601 mux8_1.NAND4F_0.C SEL0 13.0495f
C602 mux8_5.NAND4F_3.Y mux8_5.NAND4F_7.Y 5.28e-20
C603 OR8_0.S1 B0 0.070158f
C604 XOR8_0.S4 mux8_5.NAND4F_7.Y 9.74e-20
C605 MULT_0.4bit_ADDER_1.A2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B 0.950228f
C606 mux8_7.NAND4F_4.Y SEL1 0.30433f
C607 mux8_5.A0 NOT8_0.S3 0.018524f
C608 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B 0.087175f
C609 mux8_8.A0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 0.001899f
C610 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 0.005377f
C611 OR8_0.NOT8_0.A7 B4 0.015736f
C612 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B 0.001075f
C613 mux8_6.NAND4F_2.Y VDD 2.1749f
C614 mux8_4.NAND4F_4.Y mux8_4.NAND4F_9.Y 5.28e-19
C615 mux8_2.NAND4F_8.Y mux8_2.NAND4F_6.Y 2.96e-20
C616 mux8_4.A0 mux8_2.NAND4F_2.D 3.06e-19
C617 mux8_4.NAND4F_5.Y mux8_5.NAND4F_4.Y 0.002218f
C618 AND8_0.NOT8_0.A7 VDD 2.17472f
C619 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A mux8_8.A0 1.08e-19
C620 mux8_0.NAND4F_2.Y VDD 2.1746f
C621 mux8_5.NAND4F_2.D SEL1 3.38949f
C622 OR8_0.NOT8_0.A3 OR8_0.NOT8_0.A6 1.07e-20
C623 mux8_8.NAND4F_9.Y mux8_8.NAND4F_6.Y 0.222562f
C624 AND8_0.S5 XOR8_0.S4 0.024843f
C625 left_shifter_0.S0 mux8_5.A1 0.02473f
C626 mux8_7.NAND4F_0.Y mux8_7.NAND4F_9.Y 2.96e-20
C627 MULT_0.S2 mux8_3.NAND4F_4.Y 0.157118f
C628 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A 0.127125f
C629 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A 2.06e-19
C630 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT mux8_7.A0 0.697477f
C631 mux8_6.A0 mux8_6.NAND4F_2.Y 0.200461f
C632 mux8_7.A1 mux8_7.NAND4F_6.Y 8.98e-23
C633 mux8_6.A1 mux8_6.NAND4F_4.Y 0.157118f
C634 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B 0.087175f
C635 AND8_0.NOT8_0.A3 A2 0.335175f
C636 mux8_4.NAND4F_2.D mux8_4.NAND4F_0.C 1.55302f
C637 VDD A2 6.49764f
C638 B6 B1 0.020758f
C639 mux8_1.NAND4F_9.Y mux8_1.NAND4F_6.Y 0.222562f
C640 MULT_0.inv_9.Y A3 0.243265f
C641 AND8_0.S0 mux8_7.A1 0.149616f
C642 OR8_0.NOT8_0.A6 OR8_0.S7 0.34431f
C643 AND8_0.NOT8_0.A1 B4 6.46e-22
C644 mux8_4.NAND4F_0.C NOT8_0.S3 0.054353f
C645 mux8_7.A0 NOT8_0.S2 0.016346f
C646 mux8_1.NAND4F_2.D mux8_1.NAND4F_2.Y 0.339934f
C647 mux8_1.NAND4F_4.B MULT_0.SO 0.039141f
C648 left_shifter_0.S7 XOR8_0.S5 0.032772f
C649 V_FLAG_0.XOR2_2.Y VDD 1.1264f
C650 mux8_7.NAND4F_5.Y SEL1 0.306449f
C651 mux8_3.NAND4F_2.D mux8_3.NAND4F_3.Y 0.397922f
C652 8bit_ADDER_0.S2 mux8_3.NAND4F_4.Y 0.047022f
C653 mux8_1.NAND4F_2.D VDD 1.66929f
C654 mux8_5.NAND4F_2.Y mux8_5.NAND4F_5.Y 4.33e-19
C655 mux8_1.NAND4F_9.Y mux8_2.NAND4F_2.Y 1.02e-21
C656 mux8_6.A1 AND8_0.S5 0.01978f
C657 mux8_4.NAND4F_2.Y VDD 2.17488f
C658 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_1.A2 7.68e-20
C659 mux8_4.NAND4F_8.Y mux8_4.NAND4F_7.Y 9.84e-20
C660 MULT_0.4bit_ADDER_0.A2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A 1.19e-19
C661 AND8_0.S0 NOT8_0.S0 8.06e-19
C662 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT MULT_0.inv_9.Y 0.134332f
C663 8bit_ADDER_0.S2 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 4.24e-19
C664 mux8_7.NAND4F_4.B SEL1 4.36064f
C665 mux8_2.NAND4F_6.Y VDD 2.17807f
C666 mux8_8.NAND4F_1.Y mux8_6.NAND4F_3.Y 0.002218f
C667 AND8_0.NOT8_0.A7 A6 0.169207f
C668 AND8_0.S2 AND8_0.NOT8_0.A1 0.338686f
C669 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A 0.002364f
C670 mux8_0.NAND4F_2.Y mux8_0.NAND4F_8.Y 0.222339f
C671 XOR8_0.S2 mux8_3.NAND4F_7.Y 9.74e-20
C672 V_FLAG_0.XOR2_2.Y mux8_6.A0 0.28638f
C673 8bit_ADDER_0.S2 mux8_1.NAND4F_0.C 3.31e-19
C674 mux8_7.NAND4F_8.Y mux8_7.NAND4F_7.Y 9.84e-20
C675 OR8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 9.14e-19
C676 mux8_5.NAND4F_5.Y VDD 2.19984f
C677 mux8_8.A1 mux8_8.NAND4F_6.Y 8.98e-23
C678 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B 0.792412f
C679 AND8_0.S1 NOT8_0.S2 1.07e-19
C680 AND8_0.NOT8_0.A4 AND8_0.NOT8_0.A6 2.48e-20
C681 mux8_1.NAND4F_4.Y mux8_1.NAND4F_7.Y 4.32e-19
C682 mux8_2.NAND4F_3.Y mux8_2.NAND4F_1.Y 0.086984f
C683 mux8_7.A0 SEL3 6.44e-20
C684 XOR8_0.S6 mux8_8.NAND4F_5.Y 0.602392f
C685 NOT8_0.S6 XOR8_0.S6 8.6694f
C686 B7 B3 0.090874f
C687 mux8_8.NAND4F_3.Y mux8_8.NAND4F_7.Y 5.28e-20
C688 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT SEL3 0.128176f
C689 mux8_6.NAND4F_5.Y Y7 0.001312f
C690 A6 A2 0.023553f
C691 mux8_1.NAND4F_1.Y mux8_1.NAND4F_7.Y 0.617483f
C692 mux8_5.A0 mux8_5.NAND4F_4.Y 0.047022f
C693 mux8_7.A1 NOT8_0.S3 0.019628f
C694 mux8_5.A0 mux8_5.NAND4F_0.C 0.099709f
C695 mux8_6.A1 mux8_6.NAND4F_4.B 0.039141f
C696 OR8_0.NOT8_0.A7 B5 0.023973f
C697 mux8_8.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B 0.003836f
C698 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A VDD 1.34628f
C699 mux8_2.NAND4F_0.C mux8_2.NAND4F_3.Y 0.399921f
C700 XOR8_0.S7 B7 0.330439f
C701 mux8_8.NAND4F_2.D mux8_8.NAND4F_3.Y 0.397922f
C702 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A VDD 1.66874f
C703 left_shifter_0.S0 B1 0.001444f
C704 OR8_0.NOT8_0.A3 VDD 0.942836f
C705 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT mux8_8.A1 0.014376f
C706 mux8_1.NAND4F_0.C mux8_2.NAND4F_4.B 0.003147f
C707 B0 A3 1.03436f
C708 A5 A0 0.024581f
C709 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 0.51175f
C710 OR8_0.S1 OR8_0.S2 1.87533f
C711 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT 0.003009f
C712 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A mux8_7.A0 3.29e-19
C713 mux8_6.NAND4F_4.B mux8_6.NAND4F_4.Y 0.275773f
C714 AND8_0.S7 mux8_6.NAND4F_2.Y 1.24e-19
C715 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A 0.009055f
C716 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A 0.118063f
C717 XOR8_0.S5 A3 4.61e-19
C718 OR8_0.S1 mux8_2.NAND4F_4.Y 0.526611f
C719 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A 0.186684f
C720 AND8_0.NOT8_0.A7 AND8_0.S7 0.393091f
C721 XOR8_0.S7 SEL0 0.121026f
C722 mux8_8.A0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 1.08e-19
C723 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT 0.119903f
C724 XOR8_0.S2 A2 0.558891f
C725 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A 3.34e-19
C726 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B 2.43e-19
C727 left_shifter_0.S7 mux8_6.NAND4F_2.D 4.32e-19
C728 OR8_0.S7 VDD 1.38602f
C729 mux8_4.NAND4F_0.C mux8_5.NAND4F_0.C 0.001594f
C730 MULT_0.4bit_ADDER_2.B2 VDD 1.97689f
C731 mux8_5.A1 A0 2.44e-19
C732 mux8_1.NAND4F_8.Y mux8_1.NAND4F_5.Y 0.001122f
C733 mux8_4.NAND4F_2.Y mux8_4.NAND4F_8.Y 0.222339f
C734 mux8_4.A0 A2 0.43851f
C735 AND8_0.S7 A2 0.00167f
C736 MULT_0.4bit_ADDER_0.B2 B0 0.088893f
C737 mux8_6.NAND4F_6.Y mux8_6.NAND4F_1.Y 2.45057f
C738 mux8_6.NAND4F_5.Y mux8_6.NAND4F_7.Y 0.235079f
C739 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B 0.209959f
C740 mux8_8.NAND4F_2.Y mux8_8.NAND4F_5.Y 4.33e-19
C741 NOT8_0.S6 mux8_8.NAND4F_2.Y 1.43e-19
C742 mux8_6.NAND4F_9.Y mux8_6.NAND4F_1.Y 0.222572f
C743 mux8_7.A0 AND8_0.S4 0.022627f
C744 NOT8_0.S7 mux8_6.NAND4F_2.Y 1.43e-19
C745 XOR8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A 9.55e-20
C746 XOR8_0.S6 SEL2 0.236671f
C747 mux8_6.A0 OR8_0.S7 0.061252f
C748 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A 0.118063f
C749 mux8_4.NAND4F_1.Y SEL2 0.37854f
C750 mux8_2.NAND4F_9.Y Y1 6.43e-19
C751 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B SEL3 0.209959f
C752 mux8_4.A0 mux8_1.NAND4F_2.D 3.06e-19
C753 mux8_4.A0 mux8_4.NAND4F_2.Y 0.200461f
C754 A7 A3 0.055695f
C755 OR8_0.S1 SEL1 0.105609f
C756 OR8_0.NOT8_0.A0 A2 5.81e-19
C757 mux8_3.NAND4F_1.Y SEL2 0.37854f
C758 mux8_6.NAND4F_2.D mux8_6.NAND4F_5.Y 9.34e-20
C759 mux8_7.A0 mux8_7.NAND4F_4.Y 0.047022f
C760 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B 1.2618f
C761 B7 B4 0.117301f
C762 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A SEL3 1.58984f
C763 NOT8_0.S1 mux8_5.A1 0.015097f
C764 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT 0.094762f
C765 mux8_0.NAND4F_0.Y mux8_0.NAND4F_7.Y 0.08762f
C766 mux8_7.NAND4F_0.C SEL0 12.6702f
C767 8bit_ADDER_0.S2 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 0.023419f
C768 XOR8_0.S1 mux8_8.A1 0.022349f
C769 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT 1.58859f
C770 mux8_6.NAND4F_0.C mux8_6.NAND4F_0.Y 0.223896f
C771 mux8_2.NAND4F_2.Y mux8_2.NAND4F_4.Y 2.04463f
C772 XOR8_0.S5 mux8_7.NAND4F_7.Y 9.74e-20
C773 mux8_0.NAND4F_5.Y mux8_1.NAND4F_4.Y 0.002218f
C774 AND8_0.S1 AND8_0.S4 2.1e-20
C775 OR8_0.S7 A6 0.00176f
C776 mux8_0.NAND4F_9.Y VDD 2.28341f
C777 mux8_7.A1 mux8_5.NAND4F_0.C 3.1e-20
C778 NOT8_0.S4 NOT8_0.S5 1.70891f
C779 mux8_8.NAND4F_1.Y mux8_8.NAND4F_7.Y 0.617483f
C780 mux8_7.NAND4F_0.C mux8_8.NAND4F_4.B 0.002598f
C781 OR8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A 4.2e-20
C782 OR8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A 1.25e-19
C783 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A 0.013169f
C784 OR8_0.NOT8_0.A7 B6 0.037892f
C785 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 0.139263f
C786 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B 0.001075f
C787 XOR8_0.S1 B0 0.143834f
C788 NOT8_0.S4 mux8_5.NAND4F_2.Y 1.43e-19
C789 MULT_0.inv_9.Y mux8_8.A1 4.71e-19
C790 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A 2.56e-19
C791 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y B3 0.202041f
C792 mux8_5.A1 SEL2 0.075829f
C793 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 1.2618f
C794 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A 0.001379f
C795 mux8_1.NAND4F_4.Y NOT8_0.S0 2.18e-19
C796 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y B3 0.001047f
C797 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.A2 4.15e-20
C798 left_shifter_0.S7 SEL1 0.069384f
C799 AND8_0.NOT8_0.A4 AND8_0.S4 0.395881f
C800 mux8_8.NAND4F_2.D mux8_8.NAND4F_1.Y 2.96e-20
C801 AND8_0.S6 left_shifter_0.S7 0.030124f
C802 mux8_1.NAND4F_6.Y SEL1 0.222306f
C803 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B 0.005184f
C804 OR8_0.S1 mux8_4.A1 0.017872f
C805 B3 A4 0.053474f
C806 AND8_0.S2 SEL0 0.128342f
C807 NOT8_0.S5 mux8_7.NAND4F_2.D 4.43e-19
C808 mux8_7.NAND4F_0.C mux8_7.NAND4F_2.Y 0.122872f
C809 mux8_4.NAND4F_2.D mux8_4.NAND4F_7.Y 2.97e-20
C810 NOT8_0.S0 mux8_1.NAND4F_1.Y 0.55011f
C811 NOT8_0.S4 VDD 0.966965f
C812 left_shifter_0.S0 AND8_0.S3 0.006997f
C813 mux8_7.A0 mux8_7.NAND4F_5.Y 2.08e-19
C814 OR8_0.NOT8_0.A2 VDD 0.930405f
C815 AND8_0.NOT8_0.A3 B2 0.017454f
C816 mux8_8.NAND4F_2.Y SEL2 3.61e-20
C817 VDD B2 8.39797f
C818 NOT8_0.S3 mux8_4.NAND4F_7.Y 0.431664f
C819 mux8_8.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A 2.52e-19
C820 NOT8_0.S1 mux8_2.NAND4F_5.Y 0.288211f
C821 mux8_2.NAND4F_2.Y SEL1 0.222332f
C822 mux8_0.NAND4F_6.Y SEL2 0.419676f
C823 OR8_0.S2 mux8_3.NAND4F_3.Y 2.56e-19
C824 B1 A0 36.8088f
C825 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B VDD 1.96375f
C826 mux8_7.A1 mux8_7.NAND4F_0.Y 0.43187f
C827 AND8_0.NOT8_0.A5 A5 0.932489f
C828 OR8_0.S2 A3 2.37e-19
C829 mux8_7.A0 mux8_7.NAND4F_4.B 1.52147f
C830 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B A1 0.950228f
C831 XOR8_0.S0 OR8_0.S1 0.05719f
C832 mux8_0.NAND4F_8.Y mux8_0.NAND4F_9.Y 0.696806f
C833 ZFLAG_0.nor4_0.Y VDD 0.647593f
C834 B3 A1 1.88729f
C835 mux8_6.A0 NOT8_0.S4 0.015765f
C836 mux8_3.NAND4F_2.D mux8_3.NAND4F_6.Y 2.96e-20
C837 mux8_5.NAND4F_4.B mux8_5.NAND4F_4.Y 0.275773f
C838 MULT_0.4bit_ADDER_1.A2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B 0.00981f
C839 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B 0.001328f
C840 mux8_5.NAND4F_2.D mux8_5.NAND4F_6.Y 2.96e-20
C841 mux8_6.NAND4F_5.Y SEL1 0.306282f
C842 AND8_0.S7 OR8_0.S7 25.2186f
C843 mux8_7.NAND4F_2.D VDD 1.36772f
C844 mux8_5.NAND4F_0.C mux8_5.NAND4F_4.B 2.13074f
C845 AND8_0.S0 A2 0.031741f
C846 mux8_3.NAND4F_4.Y NOT8_0.S2 2.18e-19
C847 OR8_0.NOT8_0.A1 A2 0.055854f
C848 mux8_8.A0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 0.001899f
C849 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B 0.021215f
C850 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A B6 0.001945f
C851 mux8_0.NAND4F_2.D mux8_0.NAND4F_6.Y 2.96e-20
C852 mux8_1.NAND4F_0.C mux8_2.NAND4F_3.Y 1.02e-21
C853 mux8_2.NAND4F_5.Y SEL2 0.323263f
C854 mux8_1.NAND4F_2.D AND8_0.S0 0.076916f
C855 mux8_1.NAND4F_0.C mux8_1.NAND4F_4.B 2.13077f
C856 NOT8_0.S1 B1 0.429815f
C857 mux8_8.NAND4F_6.Y SEL1 0.222305f
C858 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B 0.087175f
C859 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT mux8_7.A0 0.007796f
C860 B7 B5 0.174581f
C861 mux8_1.NAND4F_1.Y mux8_2.NAND4F_2.D 1.02e-21
C862 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT 0.003012f
C863 MULT_0.S2 AND8_0.S2 11.979f
C864 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A 1.01138f
C865 mux8_8.A1 B0 0.008754f
C866 VDD Y0 0.947402f
C867 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 0.132279f
C868 mux8_6.A1 mux8_6.NAND4F_8.Y 1.16e-22
C869 MULT_0.4bit_ADDER_1.B3 A3 1.78e-19
C870 B2 A6 0.019948f
C871 NOT8_0.S7 OR8_0.S7 0.040898f
C872 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B A6 0.950228f
C873 XOR8_0.S0 mux8_1.NAND4F_6.Y 0.520706f
C874 mux8_4.NAND4F_5.Y mux8_4.NAND4F_1.Y 0.110562f
C875 mux8_3.NAND4F_4.B VDD 1.19881f
C876 mux8_8.A1 XOR8_0.S5 0.031392f
C877 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A SEL3 1.01138f
C878 AND8_0.S6 A3 0.035568f
C879 mux8_4.NAND4F_9.Y VDD 2.28291f
C880 mux8_3.NAND4F_3.Y mux8_3.NAND4F_2.Y 1.63543f
C881 mux8_3.NAND4F_0.Y mux8_3.NAND4F_4.Y 0.28646f
C882 XOR8_0.S3 mux8_4.NAND4F_1.Y 0.404949f
C883 NOT8_0.S5 XOR8_0.S4 0.032894f
C884 mux8_3.NAND4F_0.C SEL2 1.46809f
C885 MULT_0.inv_9.Y MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 0.950228f
C886 mux8_5.NAND4F_0.Y mux8_5.NAND4F_4.Y 0.28646f
C887 mux8_5.NAND4F_3.Y mux8_5.NAND4F_2.Y 1.63543f
C888 mux8_6.NAND4F_4.Y mux8_6.NAND4F_8.Y 0.404949f
C889 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A 0.127125f
C890 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y B4 0.001436f
C891 8bit_ADDER_0.S2 AND8_0.S2 0.060472f
C892 mux8_3.NAND4F_5.Y mux8_3.NAND4F_1.Y 0.110562f
C893 Y4 Y5 1.63112f
C894 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 0.087175f
C895 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y B4 3.28e-19
C896 mux8_5.NAND4F_0.C mux8_5.NAND4F_0.Y 0.223896f
C897 mux8_5.NAND4F_2.Y XOR8_0.S4 1.49e-19
C898 8bit_ADDER_0.S2 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 0.009025f
C899 mux8_4.NAND4F_3.Y mux8_4.NAND4F_1.Y 0.086984f
C900 mux8_4.NAND4F_2.D mux8_4.NAND4F_2.Y 0.339934f
C901 8bit_ADDER_0.C A3 0.037264f
C902 AND8_0.S5 OR8_0.NOT8_0.A6 0.024124f
C903 B4 A4 43.4211f
C904 MULT_0.4bit_ADDER_1.B0 VDD 1.99314f
C905 mux8_7.NAND4F_3.Y SEL2 2.96e-20
C906 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_1.B3 0.012283f
C907 mux8_5.NAND4F_3.Y VDD 2.17571f
C908 mux8_3.NAND4F_1.Y mux8_4.NAND4F_3.Y 0.002218f
C909 mux8_4.NAND4F_2.Y NOT8_0.S3 1.43e-19
C910 mux8_1.NAND4F_3.Y mux8_1.NAND4F_2.Y 1.63543f
C911 mux8_1.NAND4F_0.Y mux8_1.NAND4F_4.Y 0.28646f
C912 OR8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 2.91e-22
C913 XOR8_0.S2 B2 0.252983f
C914 mux8_7.NAND4F_3.Y mux8_7.NAND4F_1.Y 0.086984f
C915 XOR8_0.S4 VDD 0.893611f
C916 OR8_0.NOT8_0.A1 OR8_0.NOT8_0.A3 5.54e-19
C917 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B 2.43e-19
C918 XOR8_0.S1 OR8_0.S2 0.051936f
C919 mux8_1.NAND4F_3.Y VDD 2.30196f
C920 mux8_6.A1 NOT8_0.S5 0.043273f
C921 mux8_1.NAND4F_0.Y mux8_1.NAND4F_1.Y 5.28e-20
C922 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_2.B1 9.98e-20
C923 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A 0.127125f
C924 mux8_2.NAND4F_4.Y XOR8_0.S1 2.3e-19
C925 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A 0.186684f
C926 mux8_6.NAND4F_5.Y S 2.73e-20
C927 B4 A1 0.024551f
C928 mux8_5.A1 XOR8_0.S3 0.049315f
C929 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A 0.002364f
C930 AND8_0.S7 B2 0.002823f
C931 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A B0 0.001042f
C932 AND8_0.S3 A0 0.232489f
C933 mux8_6.A0 XOR8_0.S4 0.025752f
C934 mux8_4.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B 0.005184f
C935 mux8_7.A0 OR8_0.S1 0.023842f
C936 AND8_0.NOT8_0.A0 A0 0.979725f
C937 OR8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT 1.69e-20
C938 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT 0.125439f
C939 A7 B0 0.587667f
C940 mux8_8.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 0.003836f
C941 AND8_0.S0 MULT_0.4bit_ADDER_2.B2 5.07e-19
C942 AND8_0.S2 A1 0.043756f
C943 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A VDD 1.68257f
C944 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT 0.119905f
C945 mux8_6.A1 VDD 3.53964f
C946 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A 1.77e-19
C947 OR8_0.NOT8_0.A0 OR8_0.NOT8_0.A2 3.11e-19
C948 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y A5 5.82e-19
C949 mux8_3.NAND4F_2.D OR8_0.S2 0.08162f
C950 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 0.511767f
C951 OR8_0.NOT8_0.A0 B2 0.056989f
C952 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A mux8_7.A0 1.53e-19
C953 MULT_0.4bit_ADDER_1.A2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A 0.00194f
C954 NOT8_0.S4 NOT8_0.S7 0.004712f
C955 XOR8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B 0.001619f
C956 B7 B6 5.46351f
C957 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A VDD 1.35602f
C958 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 1.58859f
C959 mux8_8.A0 AND8_0.S2 0.016924f
C960 NOT8_0.S5 AND8_0.S5 0.017209f
C961 mux8_8.A0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 1.08e-19
C962 mux8_5.NAND4F_7.Y VDD 2.14052f
C963 AND8_0.S1 OR8_0.S1 32.287598f
C964 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A 0.008333f
C965 mux8_3.NAND4F_4.B XOR8_0.S2 0.96335f
C966 NOT8_0.S1 AND8_0.S3 0.041013f
C967 mux8_6.NAND4F_0.Y SEL0 0.236427f
C968 XOR8_0.S1 SEL1 0.093735f
C969 mux8_6.A0 mux8_6.A1 4.77685f
C970 mux8_6.NAND4F_4.Y VDD 2.21738f
C971 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B 0.792412f
C972 mux8_4.NAND4F_8.Y mux8_4.NAND4F_9.Y 0.696806f
C973 mux8_0.NAND4F_0.Y SEL0 0.236427f
C974 XOR8_0.S6 mux8_8.NAND4F_7.Y 9.74e-20
C975 mux8_0.NAND4F_4.Y VDD 2.21695f
C976 MULT_0.4bit_ADDER_1.B3 MULT_0.inv_9.Y 0.001146f
C977 MULT_0.SO mux8_1.NAND4F_6.Y 8.98e-23
C978 VDD V 0.832878f
C979 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A 0.118063f
C980 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y B5 0.202041f
C981 OR8_0.S2 mux8_8.A1 0.016473f
C982 mux8_8.NAND4F_0.C mux8_8.NAND4F_6.Y 0.142729f
C983 mux8_6.A0 mux8_6.NAND4F_4.Y 0.047022f
C984 AND8_0.S5 VDD 1.40455f
C985 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A B5 0.001945f
C986 MULT_0.4bit_ADDER_0.A2 A3 0.003697f
C987 mux8_5.A0 mux8_5.A1 4.79045f
C988 mux8_4.NAND4F_0.C mux8_4.NAND4F_1.Y 0.402437f
C989 mux8_8.NAND4F_2.D XOR8_0.S6 4.4e-19
C990 AND8_0.S3 SEL2 0.078529f
C991 8bit_ADDER_0.S0 SEL0 0.671967f
C992 B5 A4 35.9488f
C993 mux8_3.NAND4F_2.D SEL1 3.36943f
C994 mux8_6.NAND4F_2.Y mux8_6.NAND4F_6.Y 0.08709f
C995 mux8_2.NAND4F_0.C OR8_0.S1 0.051105f
C996 mux8_6.A0 V 1.33e-20
C997 mux8_1.NAND4F_2.D mux8_1.NAND4F_4.Y 0.349681f
C998 mux8_6.NAND4F_2.Y mux8_6.NAND4F_9.Y 2.96e-20
C999 OR8_0.S2 B0 0.309528f
C1000 SEL3 B3 1.18462f
C1001 mux8_3.NAND4F_2.D mux8_3.NAND4F_2.Y 0.339934f
C1002 OR8_0.S2 mux8_3.NAND4F_6.Y 5.23e-19
C1003 mux8_6.A0 AND8_0.S5 0.015328f
C1004 mux8_4.NAND4F_0.Y SEL0 0.236427f
C1005 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B 0.209959f
C1006 mux8_1.NAND4F_9.Y mux8_2.NAND4F_4.Y 1.02e-21
C1007 AND8_0.NOT8_0.A2 A3 0.088115f
C1008 XOR8_0.S1 mux8_4.A1 0.020135f
C1009 mux8_5.NAND4F_4.Y mux8_5.NAND4F_5.Y 0.087643f
C1010 MULT_0.inv_9.Y MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A 0.685441f
C1011 mux8_4.NAND4F_4.Y VDD 2.21738f
C1012 mux8_1.NAND4F_2.D mux8_1.NAND4F_1.Y 2.96e-20
C1013 mux8_3.NAND4F_0.C mux8_3.NAND4F_5.Y 0.051024f
C1014 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A 0.118063f
C1015 AND8_0.NOT8_0.A1 A0 0.181031f
C1016 8bit_ADDER_0.S2 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 0.005184f
C1017 mux8_5.NAND4F_0.C mux8_5.NAND4F_5.Y 0.051024f
C1018 B5 A1 0.024059f
C1019 AND8_0.S1 mux8_2.NAND4F_2.Y 1.24e-19
C1020 mux8_0.NAND4F_4.B SEL2 0.734118f
C1021 mux8_0.NAND4F_4.Y mux8_0.NAND4F_8.Y 0.404949f
C1022 XOR8_0.S4 AND8_0.S7 0.037626f
C1023 OR8_0.NOT8_0.A1 OR8_0.NOT8_0.A2 1.16238f
C1024 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B 0.792412f
C1025 AND8_0.S0 B2 0.148218f
C1026 OR8_0.NOT8_0.A1 B2 0.046436f
C1027 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_0.A2 2.90168f
C1028 OR8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A 8.58e-21
C1029 mux8_0.NAND4F_7.Y SEL2 0.176544f
C1030 mux8_6.NAND4F_4.B VDD 1.19723f
C1031 XOR8_0.S0 XOR8_0.S1 0.009902f
C1032 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 0.008371f
C1033 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_1.A2 2.3109f
C1034 mux8_1.NAND4F_8.Y mux8_1.NAND4F_7.Y 9.84e-20
C1035 mux8_2.NAND4F_2.Y mux8_2.NAND4F_1.Y 3.31e-22
C1036 mux8_8.A1 SEL1 0.06839f
C1037 mux8_7.NAND4F_2.D mux8_7.NAND4F_6.Y 2.96e-20
C1038 XOR8_0.S2 mux8_6.A1 0.1811f
C1039 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A 0.001379f
C1040 mux8_8.A1 AND8_0.S6 2.18427f
C1041 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A 2.56e-19
C1042 V_FLAG_0.XOR2_2.B B7 0.55689f
C1043 AND8_0.NOT8_0.A6 B4 2.23e-20
C1044 mux8_6.NAND4F_0.C SEL2 1.48751f
C1045 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 0.209959f
C1046 mux8_0.NAND4F_2.D mux8_0.NAND4F_4.B 1.27138f
C1047 mux8_5.NAND4F_9.Y SEL2 1.49e-20
C1048 left_shifter_0.S0 SEL0 0.130208f
C1049 mux8_7.A0 A3 6.44e-20
C1050 mux8_4.NAND4F_6.Y SEL1 0.222305f
C1051 mux8_6.A0 mux8_6.NAND4F_4.B 1.52147f
C1052 mux8_0.NAND4F_2.D mux8_0.NAND4F_7.Y 2.97e-20
C1053 mux8_4.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A 0.002364f
C1054 NOT8_0.S7 XOR8_0.S4 0.051787f
C1055 mux8_6.A1 AND8_0.S7 3.5423f
C1056 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y B1 0.001436f
C1057 mux8_6.NAND4F_2.D mux8_6.NAND4F_7.Y 2.97e-20
C1058 mux8_3.NAND4F_6.Y SEL1 0.222305f
C1059 mux8_2.NAND4F_0.C mux8_2.NAND4F_2.Y 0.122872f
C1060 mux8_8.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A 2.52e-19
C1061 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A MULT_0.inv_15.Y 7.7e-20
C1062 mux8_8.NAND4F_2.D mux8_8.NAND4F_2.Y 0.339934f
C1063 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y B1 6.57e-19
C1064 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A mux8_8.A1 2.52e-19
C1065 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y B1 6.57e-19
C1066 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B 1.2618f
C1067 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B MULT_0.inv_9.Y 0.001496f
C1068 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B VDD 1.82538f
C1069 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y B1 6.57e-19
C1070 XOR8_0.S5 SEL1 0.09541f
C1071 mux8_3.NAND4F_2.Y mux8_3.NAND4F_6.Y 0.08709f
C1072 ZFLAG_0.nor4_1.Y Y4 0.006226f
C1073 AND8_0.S6 XOR8_0.S5 2.30403f
C1074 NOT8_0.S3 NOT8_0.S4 0.137019f
C1075 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A 0.001571f
C1076 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B A1 0.00981f
C1077 ZFLAG_0.nor4_0.Y Y6 2.06e-19
C1078 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A 8.33e-19
C1079 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT 0.127988f
C1080 8bit_ADDER_0.S2 8bit_ADDER_0.S0 0.056298f
C1081 NOT8_0.S3 B2 0.389001f
C1082 XOR8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A 2.35e-19
C1083 AND8_0.S7 mux8_6.NAND4F_4.Y 0.402481f
C1084 mux8_6.A1 OR8_0.NOT8_0.A0 0.006068f
C1085 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B 0.005184f
C1086 AND8_0.S1 A3 1.3e-20
C1087 8bit_ADDER_0.C B0 0.08296f
C1088 mux8_5.A0 mux8_3.NAND4F_0.C 1.95e-19
C1089 XOR8_0.S2 AND8_0.S5 0.001841f
C1090 AND8_0.S4 B3 1.15815f
C1091 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y B6 0.001436f
C1092 mux8_7.A1 mux8_5.A1 8.87622f
C1093 mux8_8.A1 mux8_4.A1 4e-19
C1094 AND8_0.S2 NOT8_0.S2 6.31e-19
C1095 mux8_8.A0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 0.001899f
C1096 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B 0.005184f
C1097 B6 A4 0.024758f
C1098 mux8_2.NAND4F_1.Y mux8_3.NAND4F_3.Y 0.002062f
C1099 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B 8.3e-19
C1100 MULT_0.SO MULT_0.4bit_ADDER_0.B2 9.08e-19
C1101 mux8_6.A1 NOT8_0.S7 0.093275f
C1102 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_1.B3 0.186718f
C1103 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT 7.81e-20
C1104 mux8_4.A1 mux8_4.NAND4F_6.Y 8.98e-23
C1105 AND8_0.S5 AND8_0.S7 0.006182f
C1106 mux8_0.NAND4F_5.Y mux8_0.NAND4F_6.Y 1.93433f
C1107 SEL3 B4 1.17767f
C1108 NOT8_0.S0 mux8_5.A1 0.01556f
C1109 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT mux8_7.A0 6.44e-20
C1110 mux8_4.NAND4F_4.Y mux8_4.NAND4F_8.Y 0.404949f
C1111 XOR8_0.S0 mux8_8.A1 0.266966f
C1112 mux8_2.NAND4F_0.Y NOT8_0.S1 5.24e-19
C1113 left_shifter_0.S0 MULT_0.S2 0.034637f
C1114 AND8_0.NOT8_0.A4 A3 0.189069f
C1115 mux8_1.NAND4F_5.Y SEL0 0.123423f
C1116 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT VDD 3.50211f
C1117 mux8_8.NAND4F_4.Y mux8_8.NAND4F_5.Y 0.087643f
C1118 NOT8_0.S6 mux8_8.NAND4F_4.Y 2.18e-19
C1119 NOT8_0.S7 mux8_6.NAND4F_4.Y 2.18e-19
C1120 B6 A1 0.023945f
C1121 AND8_0.S3 mux8_4.NAND4F_5.Y 5.23e-19
C1122 mux8_8.NAND4F_0.C mux8_8.NAND4F_9.Y 4.79e-21
C1123 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B A6 0.00981f
C1124 NOT8_0.S1 mux8_2.NAND4F_7.Y 0.431664f
C1125 AND8_0.S3 XOR8_0.S3 1.69e-19
C1126 mux8_4.A0 mux8_4.NAND4F_4.Y 0.047022f
C1127 mux8_3.NAND4F_0.C mux8_4.NAND4F_0.C 0.001594f
C1128 OR8_0.S7 mux8_6.NAND4F_6.Y 5.23e-19
C1129 XOR8_0.S0 B0 0.227887f
C1130 mux8_0.NAND4F_4.B mux8_0.NAND4F_3.Y 0.223331f
C1131 mux8_8.A0 B6 5.02e-19
C1132 8bit_ADDER_0.S2 left_shifter_0.S0 0.016749f
C1133 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT 1.58859f
C1134 MULT_0.inv_9.Y MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 0.00981f
C1135 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A 0.001568f
C1136 NOT8_0.S7 AND8_0.S5 0.018894f
C1137 mux8_2.NAND4F_0.Y SEL2 3.06e-20
C1138 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A 1.01138f
C1139 8bit_ADDER_0.C A7 0.2109f
C1140 mux8_0.NAND4F_3.Y mux8_0.NAND4F_7.Y 5.28e-20
C1141 AND8_0.NOT8_0.A6 B5 0.050259f
C1142 NOT8_0.S6 B7 0.035606f
C1143 mux8_0.NAND4F_0.C SEL1 1.12331f
C1144 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A B4 0.001945f
C1145 mux8_7.A0 XOR8_0.S1 0.024552f
C1146 mux8_4.NAND4F_9.Y NOT8_0.S3 3.17e-20
C1147 mux8_6.NAND4F_0.C mux8_6.NAND4F_3.Y 0.399921f
C1148 8bit_ADDER_0.S2 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 0.002364f
C1149 AND8_0.S7 mux8_6.NAND4F_4.B 1.04047f
C1150 mux8_5.A1 mux8_5.NAND4F_4.B 0.039141f
C1151 mux8_8.A0 8bit_ADDER_0.S0 0.059367f
C1152 B7 A0 0.07108f
C1153 mux8_2.NAND4F_7.Y SEL2 0.176544f
C1154 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B 0.001075f
C1155 AND8_0.S0 mux8_6.A1 0.160455f
C1156 mux8_5.NAND4F_1.Y SEL2 0.37854f
C1157 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 0.005938f
C1158 mux8_6.A1 OR8_0.NOT8_0.A1 0.11437f
C1159 NOT8_0.S6 SEL0 1.10257f
C1160 mux8_8.NAND4F_5.Y SEL0 0.122083f
C1161 mux8_6.NAND4F_2.D SEL1 3.26355f
C1162 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 0.792412f
C1163 mux8_0.NAND4F_0.C 8bit_ADDER_0.C 0.083755f
C1164 NOT8_0.S4 mux8_5.NAND4F_4.Y 2.18e-19
C1165 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 0.087175f
C1166 MULT_0.inv_9.Y MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT 0.010334f
C1167 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A 1.01138f
C1168 NOT8_0.S4 mux8_5.NAND4F_0.C 0.053254f
C1169 AND8_0.S1 XOR8_0.S1 8.21e-19
C1170 mux8_2.NAND4F_2.Y mux8_2.NAND4F_9.Y 2.96e-20
C1171 mux8_8.A1 mux8_8.NAND4F_0.C 0.065359f
C1172 mux8_8.NAND4F_4.B mux8_8.NAND4F_5.Y 0.248856f
C1173 NOT8_0.S6 mux8_8.NAND4F_4.B 0.105153f
C1174 MULT_0.4bit_ADDER_0.A2 B0 0.001412f
C1175 mux8_7.A0 mux8_3.NAND4F_2.D 1.75e-19
C1176 mux8_4.NAND4F_1.Y mux8_4.NAND4F_7.Y 0.617483f
C1177 mux8_7.NAND4F_0.C mux8_7.NAND4F_4.Y 0.049743f
C1178 left_shifter_0.S0 mux8_2.NAND4F_4.B 3.2e-21
C1179 AND8_0.S4 B4 0.105122f
C1180 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A 0.248556f
C1181 NOT8_0.S7 mux8_6.NAND4F_4.B 0.105153f
C1182 mux8_4.NAND4F_4.B mux8_4.NAND4F_6.Y 0.187883f
C1183 OR8_0.S2 SEL1 0.105682f
C1184 XOR8_0.S1 mux8_2.NAND4F_1.Y 0.404949f
C1185 mux8_8.NAND4F_4.Y SEL2 8.74e-20
C1186 mux8_8.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 0.017894f
C1187 mux8_2.NAND4F_4.Y SEL1 0.304331f
C1188 OR8_0.S2 mux8_3.NAND4F_2.Y 0.402593f
C1189 AND8_0.S1 MULT_0.inv_9.Y 7.17e-20
C1190 NOT8_0.S0 B1 7.06e-20
C1191 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A 0.127125f
C1192 mux8_5.A0 AND8_0.S3 0.057074f
C1193 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A VDD 1.66874f
C1194 mux8_7.A1 mux8_7.NAND4F_3.Y 0.541275f
C1195 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 0.511769f
C1196 mux8_5.NAND4F_0.C mux8_7.NAND4F_2.D 4.54e-19
C1197 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 0.119902f
C1198 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A mux8_7.A0 1.53e-19
C1199 mux8_3.NAND4F_1.Y mux8_3.NAND4F_7.Y 0.617483f
C1200 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A 1.16e-19
C1201 AND8_0.S2 AND8_0.S4 2.82e-19
C1202 SEL3 B5 1.17298f
C1203 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A A1 0.00194f
C1204 mux8_1.NAND4F_0.C mux8_1.NAND4F_6.Y 0.142729f
C1205 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A 0.186684f
C1206 mux8_5.A1 mux8_5.NAND4F_0.Y 0.43187f
C1207 mux8_8.A0 left_shifter_0.S0 0.01811f
C1208 OR8_0.NOT8_0.A6 VDD 0.924276f
C1209 XOR8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 6.68e-20
C1210 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A 0.002364f
C1211 NOT8_0.S1 SEL0 1.10219f
C1212 mux8_2.NAND4F_2.D mux8_2.NAND4F_5.Y 9.34e-20
C1213 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B A5 0.950228f
C1214 mux8_2.NAND4F_0.C XOR8_0.S1 0.0799f
C1215 mux8_8.A0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 1.08e-19
C1216 mux8_6.NAND4F_8.Y VDD 3.38852f
C1217 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A 0.002364f
C1218 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A 1.21e-19
C1219 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.inv_15.Y 4.16e-20
C1220 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT mux8_8.A1 0.003904f
C1221 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B VDD 1.98049f
C1222 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_0.A2 0.022087f
C1223 OR8_0.NOT8_0.A5 OR8_0.S7 1.23e-19
C1224 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT 8.9e-19
C1225 mux8_7.NAND4F_0.C mux8_7.NAND4F_5.Y 0.051024f
C1226 OR8_0.S2 mux8_4.A1 0.109227f
C1227 AND8_0.NOT8_0.A6 B6 0.1517f
C1228 mux8_1.NAND4F_5.Y mux8_2.NAND4F_4.B 1.02e-21
C1229 SEL2 SEL0 1.07663f
C1230 AND8_0.S6 SEL1 0.112904f
C1231 AND8_0.NOT8_0.A7 A5 0.086332f
C1232 mux8_4.NAND4F_0.C AND8_0.S3 0.038301f
C1233 MULT_0.SO B0 0.006498f
C1234 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A mux8_4.A1 2.28e-19
C1235 mux8_8.NAND4F_0.Y VDD 2.13488f
C1236 mux8_7.NAND4F_2.D mux8_7.NAND4F_0.Y 0.184536f
C1237 mux8_7.NAND4F_0.C mux8_7.NAND4F_4.B 2.13077f
C1238 mux8_0.NAND4F_0.C mux8_0.NAND4F_1.Y 0.402437f
C1239 mux8_3.NAND4F_2.Y SEL1 0.222331f
C1240 mux8_7.NAND4F_1.Y SEL0 0.339784f
C1241 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A A6 0.00194f
C1242 mux8_2.NAND4F_8.Y VDD 3.39057f
C1243 AND8_0.S1 mux8_8.A1 0.069201f
C1244 mux8_7.A0 XOR8_0.S5 0.009372f
C1245 mux8_8.NAND4F_4.B SEL2 0.734121f
C1246 mux8_6.NAND4F_0.C mux8_6.NAND4F_1.Y 0.402437f
C1247 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.B3 0.127992f
C1248 XOR8_0.S0 OR8_0.S2 0.005012f
C1249 mux8_3.NAND4F_3.Y mux8_3.NAND4F_4.Y 0.102178f
C1250 OR8_0.NOT8_0.A6 A6 0.256456f
C1251 MULT_0.4bit_ADDER_2.B1 VDD 1.96352f
C1252 8bit_ADDER_0.C SEL1 0.332878f
C1253 8bit_ADDER_0.S2 A0 1.72e-19
C1254 mux8_5.NAND4F_3.Y mux8_5.NAND4F_4.Y 0.102178f
C1255 mux8_0.NAND4F_2.D SEL0 0.228824f
C1256 MULT_0.inv_9.Y MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A 0.00194f
C1257 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A 1.16e-19
C1258 A5 A2 0.022564f
C1259 NOT8_0.S5 VDD 1.00406f
C1260 MULT_0.S2 NOT8_0.S1 0.033848f
C1261 mux8_5.NAND4F_0.C mux8_5.NAND4F_3.Y 0.399921f
C1262 AND8_0.S1 B0 0.066184f
C1263 mux8_5.NAND4F_4.Y XOR8_0.S4 2.3e-19
C1264 mux8_3.NAND4F_9.Y VDD 2.28477f
C1265 mux8_4.NAND4F_2.D mux8_4.NAND4F_4.Y 0.349681f
C1266 mux8_4.NAND4F_2.Y mux8_4.NAND4F_1.Y 3.31e-22
C1267 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y A0 0.001406f
C1268 mux8_5.NAND4F_0.C XOR8_0.S4 0.08068f
C1269 8bit_ADDER_0.S0 mux8_1.NAND4F_4.B 1.52147f
C1270 mux8_7.NAND4F_2.Y SEL2 3.61e-20
C1271 AND8_0.S4 B5 0.050103f
C1272 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y A0 0.00101f
C1273 mux8_5.NAND4F_2.Y VDD 2.1749f
C1274 mux8_4.NAND4F_4.Y NOT8_0.S3 2.18e-19
C1275 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B 2.43e-19
C1276 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y A0 0.00101f
C1277 mux8_1.NAND4F_3.Y mux8_1.NAND4F_4.Y 0.102178f
C1278 mux8_1.NAND4F_0.Y mux8_1.NAND4F_8.Y 0.249057f
C1279 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y A0 0.007226f
C1280 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B 0.792412f
C1281 mux8_4.A1 SEL1 0.069249f
C1282 mux8_7.NAND4F_2.Y mux8_7.NAND4F_1.Y 3.31e-22
C1283 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 0.001075f
C1284 mux8_6.A0 NOT8_0.S5 0.019218f
C1285 mux8_7.A1 AND8_0.S3 0.030658f
C1286 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A 0.001379f
C1287 mux8_1.NAND4F_2.Y VDD 2.27924f
C1288 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 0.139263f
C1289 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A 0.248956f
C1290 A4 A0 0.024733f
C1291 mux8_1.NAND4F_3.Y mux8_1.NAND4F_1.Y 0.086984f
C1292 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT 8.89e-19
C1293 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A 0.118063f
C1294 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A B3 0.001945f
C1295 AND8_0.NOT8_0.A3 VDD 2.34754f
C1296 8bit_ADDER_0.S2 NOT8_0.S1 0.021247f
C1297 MULT_0.S2 SEL2 0.076698f
C1298 mux8_8.NAND4F_0.C mux8_6.NAND4F_2.D 4.54e-19
C1299 SEL3 B6 1.18486f
C1300 ZFLAG_0.nor4_0.Y Y3 0.006286f
C1301 mux8_0.NAND4F_2.Y mux8_0.NAND4F_6.Y 0.08709f
C1302 NOT8_0.S0 AND8_0.S3 0.027753f
C1303 XOR8_0.S0 SEL1 0.095831f
C1304 mux8_0.NAND4F_4.B mux8_0.NAND4F_5.Y 0.248856f
C1305 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A 0.248556f
C1306 8bit_ADDER_0.S0 SEL3 0.881449f
C1307 A1 A0 1.28004f
C1308 mux8_7.NAND4F_9.Y SEL0 2.8e-19
C1309 mux8_8.A0 mux8_8.NAND4F_5.Y 2.08e-19
C1310 mux8_8.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A 0.007358f
C1311 mux8_1.NAND4F_7.Y mux8_2.NAND4F_0.Y 0.002399f
C1312 mux8_8.A0 NOT8_0.S6 1.18e-19
C1313 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A 0.248556f
C1314 mux8_6.A0 VDD 1.96111f
C1315 OR8_0.NOT8_0.A6 AND8_0.S7 0.068695f
C1316 mux8_0.NAND4F_5.Y mux8_0.NAND4F_7.Y 0.235079f
C1317 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B MULT_0.inv_9.Y 0.013749f
C1318 mux8_5.NAND4F_4.Y mux8_5.NAND4F_7.Y 4.32e-19
C1319 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 0.209959f
C1320 mux8_3.NAND4F_0.C mux8_3.NAND4F_7.Y 0.224691f
C1321 8bit_ADDER_0.S2 SEL2 1.13198f
C1322 mux8_5.NAND4F_0.C mux8_5.NAND4F_7.Y 0.224691f
C1323 mux8_5.A1 mux8_5.NAND4F_5.Y 1.57e-19
C1324 XOR8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A 1.6e-20
C1325 mux8_1.NAND4F_4.B left_shifter_0.S0 1.01693f
C1326 Y1 Y2 5.77433f
C1327 Y0 Y3 0.023358f
C1328 left_shifter_0.S0 NOT8_0.S2 0.077778f
C1329 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A B0 0.001945f
C1330 mux8_2.NAND4F_4.B NOT8_0.S1 0.105153f
C1331 mux8_6.NAND4F_3.Y SEL0 0.360934f
C1332 mux8_8.A0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 0.001899f
C1333 mux8_0.NAND4F_1.Y SEL1 2.35e-20
C1334 left_shifter_0.S7 XOR8_0.S7 0.056737f
C1335 mux8_0.NAND4F_3.Y SEL0 0.360934f
C1336 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 0.001075f
C1337 MULT_0.4bit_ADDER_0.A2 MULT_0.4bit_ADDER_1.B3 0.003441f
C1338 OR8_0.S7 XOR8_0.S6 0.035853f
C1339 mux8_0.NAND4F_8.Y VDD 3.38852f
C1340 VDD A6 2.08508f
C1341 mux8_4.NAND4F_9.Y Y3 9.11e-19
C1342 XOR8_0.S3 B7 0.144817f
C1343 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A 0.001571f
C1344 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT mux8_7.A0 6.44e-20
C1345 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A VDD 1.69318f
C1346 XOR8_0.S0 mux8_4.A1 0.022578f
C1347 mux8_5.NAND4F_0.Y mux8_5.NAND4F_8.Y 0.249057f
C1348 mux8_5.NAND4F_0.C AND8_0.S5 6.54e-20
C1349 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT 1.69e-20
C1350 mux8_7.NAND4F_2.Y mux8_7.NAND4F_9.Y 2.96e-20
C1351 mux8_6.A1 mux8_6.NAND4F_6.Y 8.98e-23
C1352 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 0.132279f
C1353 mux8_3.NAND4F_9.Y mux8_4.NAND4F_8.Y 0.001427f
C1354 mux8_4.NAND4F_5.Y SEL0 0.122346f
C1355 8bit_ADDER_0.C mux8_0.NAND4F_1.Y 5.23e-19
C1356 mux8_5.A0 mux8_5.NAND4F_1.Y 5.23e-19
C1357 mux8_8.A0 NOT8_0.S1 0.017307f
C1358 mux8_7.A0 OR8_0.S2 0.023842f
C1359 OR8_0.S7 A5 0.007828f
C1360 mux8_4.NAND4F_4.B SEL1 4.36064f
C1361 mux8_2.NAND4F_4.B SEL2 0.734122f
C1362 mux8_6.A0 A6 0.439146f
C1363 XOR8_0.S3 SEL0 0.167762f
C1364 mux8_3.NAND4F_5.Y SEL0 0.12371f
C1365 mux8_8.NAND4F_0.C SEL1 1.12431f
C1366 AND8_0.S4 B6 0.055449f
C1367 mux8_5.NAND4F_7.Y mux8_7.NAND4F_0.Y 0.002217f
C1368 AND8_0.S6 mux8_8.NAND4F_0.C 0.039158f
C1369 mux8_2.NAND4F_5.Y mux8_2.NAND4F_6.Y 1.93433f
C1370 AND8_0.S2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A 1.54e-19
C1371 mux8_6.NAND4F_4.Y mux8_6.NAND4F_6.Y 4.33e-19
C1372 XOR8_0.S7 mux8_6.NAND4F_5.Y 0.602392f
C1373 V_FLAG_0.XOR2_0.Y mux8_0.NAND4F_4.B 3.87e-21
C1374 mux8_1.NAND4F_2.D mux8_1.NAND4F_8.Y 4.88e-20
C1375 mux8_6.NAND4F_4.Y mux8_6.NAND4F_9.Y 5.28e-19
C1376 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_0.A2 0.135871f
C1377 mux8_3.NAND4F_2.D mux8_3.NAND4F_4.Y 0.349681f
C1378 V_FLAG_0.XOR2_2.B SEL3 0.311554f
C1379 mux8_4.NAND4F_3.Y SEL0 0.360934f
C1380 B1 A2 1.31978f
C1381 mux8_4.NAND4F_8.Y VDD 3.3899f
C1382 OR8_0.NOT8_0.A4 B3 0.012105f
C1383 XOR8_0.S2 VDD 1.22139f
C1384 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A 0.186684f
C1385 mux8_1.NAND4F_4.B mux8_1.NAND4F_5.Y 0.248856f
C1386 OR8_0.S1 AND8_0.S2 2.77078f
C1387 mux8_8.A0 SEL2 0.950299f
C1388 B3 A3 43.1059f
C1389 AND8_0.S1 mux8_2.NAND4F_4.Y 0.402481f
C1390 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y B7 0.001436f
C1391 OR8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A 1.07e-19
C1392 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B 0.001075f
C1393 mux8_4.A0 VDD 1.56041f
C1394 AND8_0.S7 VDD 1.24685f
C1395 mux8_6.A0 XOR8_0.S2 0.025261f
C1396 mux8_4.A1 mux8_4.NAND4F_4.B 0.039141f
C1397 AND8_0.NOT8_0.A5 A4 0.268713f
C1398 mux8_2.NAND4F_4.Y mux8_2.NAND4F_1.Y 4.33e-19
C1399 NOT8_0.S5 NOT8_0.S7 3.53e-19
C1400 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 2.43e-19
C1401 mux8_7.A0 SEL1 0.340165f
C1402 mux8_1.NAND4F_7.Y SEL0 0.234595f
C1403 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT 1.69e-20
C1404 MULT_0.SO SEL1 0.070206f
C1405 mux8_8.NAND4F_4.Y mux8_8.NAND4F_7.Y 4.32e-19
C1406 MULT_0.S2 mux8_3.NAND4F_5.Y 1.57e-19
C1407 mux8_6.A0 mux8_4.A0 0.033668f
C1408 mux8_6.A0 AND8_0.S7 0.062091f
C1409 OR8_0.NOT8_0.A0 VDD 0.909904f
C1410 8bit_ADDER_0.C mux8_7.A0 0.091956f
C1411 mux8_5.A0 SEL0 0.680478f
C1412 mux8_2.NAND4F_0.C mux8_2.NAND4F_4.Y 0.049743f
C1413 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 0.007216f
C1414 mux8_8.NAND4F_2.D mux8_8.NAND4F_4.Y 0.349681f
C1415 mux8_6.NAND4F_4.B mux8_6.NAND4F_6.Y 0.187883f
C1416 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 0.012283f
C1417 mux8_8.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B 0.005184f
C1418 MULT_0.SO MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT 1.74e-19
C1419 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 0.007216f
C1420 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 0.428846f
C1421 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A mux8_7.A0 1.53e-19
C1422 NOT8_0.S7 VDD 0.905602f
C1423 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 0.00162f
C1424 AND8_0.S1 SEL1 0.111539f
C1425 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A 1.01138f
C1426 mux8_3.NAND4F_4.Y mux8_3.NAND4F_6.Y 4.33e-19
C1427 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A MULT_0.inv_9.Y 0.001123f
C1428 mux8_6.NAND4F_1.Y SEL0 0.339784f
C1429 NOT8_0.S0 mux8_2.NAND4F_0.Y 9.03e-22
C1430 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 0.007227f
C1431 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT 1.58859f
C1432 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 1.58859f
C1433 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 0.007216f
C1434 mux8_0.NAND4F_7.Y mux8_1.NAND4F_0.Y 0.002217f
C1435 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 0.007216f
C1436 8bit_ADDER_0.S2 mux8_3.NAND4F_5.Y 2.08e-19
C1437 B2 A5 0.019069f
C1438 mux8_5.NAND4F_0.Y mux8_5.NAND4F_9.Y 2.96e-20
C1439 mux8_2.NAND4F_1.Y SEL1 2.35e-20
C1440 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 0.007216f
C1441 AND8_0.S7 A6 0.001321f
C1442 mux8_1.NAND4F_0.C mux8_1.NAND4F_9.Y 4.79e-21
C1443 mux8_7.A0 mux8_4.A1 0.027035f
C1444 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B A5 0.00981f
C1445 mux8_3.NAND4F_8.Y SEL0 4.08e-19
C1446 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT 0.001576f
C1447 mux8_6.A0 NOT8_0.S7 1.33e-19
C1448 mux8_8.A0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 1.08e-19
C1449 mux8_0.NAND4F_9.Y C 5.24e-19
C1450 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT mux8_4.A1 0.145602f
C1451 mux8_8.NAND4F_7.Y SEL0 0.234594f
C1452 mux8_5.NAND4F_6.Y SEL1 0.222305f
C1453 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A 1.6e-19
C1454 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT 0.001576f
C1455 AND8_0.S0 MULT_0.4bit_ADDER_2.B1 5.07e-19
C1456 NOT8_0.S5 mux8_7.NAND4F_6.Y 0.79864f
C1457 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A 1.6e-19
C1458 mux8_0.NAND4F_9.Y mux8_0.NAND4F_6.Y 0.222562f
C1459 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT 0.012283f
C1460 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A 1.16e-19
C1461 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B VDD 1.97529f
C1462 mux8_5.NAND4F_8.Y mux8_5.NAND4F_5.Y 0.001122f
C1463 mux8_5.A1 NOT8_0.S4 0.009276f
C1464 mux8_7.A0 XOR8_0.S0 0.023194f
C1465 mux8_2.NAND4F_3.Y NOT8_0.S1 3.24e-22
C1466 mux8_4.NAND4F_0.C SEL0 12.684f
C1467 MULT_0.SO XOR8_0.S0 3.04e-20
C1468 OR8_0.NOT8_0.A4 B4 0.037671f
C1469 mux8_2.NAND4F_0.C SEL1 1.12028f
C1470 mux8_8.NAND4F_8.Y mux8_8.NAND4F_5.Y 0.001122f
C1471 mux8_8.NAND4F_2.D SEL0 0.229432f
C1472 B4 A3 23.923698f
C1473 AND8_0.S1 mux8_4.A1 0.018036f
C1474 NOT8_0.S1 NOT8_0.S2 0.326531f
C1475 SEL3 A0 0.349328f
C1476 mux8_5.A0 MULT_0.S2 0.022235f
C1477 OR8_0.NOT8_0.A5 AND8_0.S5 0.127774f
C1478 AND8_0.S3 A2 0.063218f
C1479 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A 8.34e-19
C1480 mux8_7.NAND4F_6.Y VDD 2.17811f
C1481 mux8_2.NAND4F_2.D mux8_2.NAND4F_0.Y 0.184536f
C1482 AND8_0.S0 mux8_1.NAND4F_2.Y 1.24e-19
C1483 mux8_4.A0 XOR8_0.S2 0.028931f
C1484 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 8bit_ADDER_0.S2 4.24e-19
C1485 AND8_0.NOT8_0.A0 A2 0.09976f
C1486 mux8_0.NAND4F_4.B mux8_0.NAND4F_2.Y 0.112019f
C1487 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT 8.9e-19
C1488 mux8_8.NAND4F_2.D mux8_8.NAND4F_4.B 1.27138f
C1489 MULT_0.inv_9.Y B3 0.457564f
C1490 mux8_4.NAND4F_9.Y mux8_4.NAND4F_1.Y 0.222572f
C1491 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A 0.001568f
C1492 AND8_0.S0 VDD 1.05196f
C1493 AND8_0.S2 A3 0.020867f
C1494 mux8_3.NAND4F_4.B mux8_3.NAND4F_1.Y 0.222551f
C1495 mux8_2.NAND4F_3.Y SEL2 3.06e-20
C1496 XOR8_0.S0 AND8_0.S1 3.53069f
C1497 OR8_0.NOT8_0.A1 VDD 0.970678f
C1498 mux8_0.NAND4F_9.Y mux8_1.NAND4F_8.Y 0.001427f
C1499 mux8_5.NAND4F_4.B mux8_5.NAND4F_1.Y 0.222551f
C1500 AND8_0.S3 mux8_4.NAND4F_2.Y 1.24e-19
C1501 mux8_2.NAND4F_2.D mux8_2.NAND4F_7.Y 2.97e-20
C1502 mux8_6.NAND4F_0.C mux8_6.NAND4F_2.Y 0.122872f
C1503 mux8_1.NAND4F_4.B SEL2 0.734121f
C1504 MULT_0.S2 mux8_3.NAND4F_8.Y 1.16e-22
C1505 NOT8_0.S2 SEL2 0.109565f
C1506 mux8_5.A0 8bit_ADDER_0.S2 3.21e-19
C1507 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 0.050843f
C1508 mux8_0.NAND4F_5.Y SEL0 0.123636f
C1509 mux8_8.A0 XOR8_0.S3 0.02968f
C1510 AND8_0.S2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT 6.95e-20
C1511 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B 0.792412f
C1512 mux8_6.A0 AND8_0.S0 0.021856f
C1513 mux8_7.A1 SEL0 1.17116f
C1514 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B 2.43e-19
C1515 mux8_4.NAND4F_1.Y mux8_5.NAND4F_3.Y 0.002218f
C1516 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A 5.19e-20
C1517 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A 2.56e-19
C1518 MULT_0.SO MULT_0.4bit_ADDER_0.A2 4.77e-19
C1519 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A 0.001379f
C1520 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B 0.087175f
C1521 XOR8_0.S4 XOR8_0.S6 0.017216f
C1522 mux8_7.NAND4F_0.C mux8_7.NAND4F_7.Y 0.224691f
C1523 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y A4 2.72669f
C1524 V_FLAG_0.XOR2_2.Y mux8_0.NAND4F_4.B 1.61e-20
C1525 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_2.B2 2.27e-19
C1526 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y mux8_5.A0 2.04e-19
C1527 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 0.008371f
C1528 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y mux8_5.A0 0.018423f
C1529 mux8_0.NAND4F_0.C mux8_1.NAND4F_0.C 0.001594f
C1530 VDD Y6 0.962594f
C1531 NOT8_0.S0 SEL0 1.10214f
C1532 mux8_2.NAND4F_4.Y mux8_2.NAND4F_9.Y 5.28e-19
C1533 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B A4 0.950228f
C1534 mux8_4.NAND4F_2.D VDD 1.36905f
C1535 NOT8_0.S7 AND8_0.S7 0.062526f
C1536 AND8_0.NOT8_0.A5 AND8_0.NOT8_0.A6 0.147743f
C1537 SEL3 SEL2 0.26782f
C1538 NOT8_0.S6 AND8_0.S4 0.0184f
C1539 mux8_8.A1 B3 8.04e-21
C1540 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y A1 0.001095f
C1541 NOT8_0.S3 VDD 1.35031f
C1542 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y A1 5.14e-19
C1543 mux8_8.NAND4F_0.Y mux8_8.NAND4F_3.Y 0.616159f
C1544 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y A1 5.14e-19
C1545 mux8_3.NAND4F_0.Y SEL2 2.97e-20
C1546 mux8_8.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A 0.002364f
C1547 OR8_0.S2 mux8_3.NAND4F_4.Y 0.526611f
C1548 mux8_6.A1 XOR8_0.S6 0.036502f
C1549 mux8_7.A1 mux8_7.NAND4F_2.Y 1.16938f
C1550 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B MULT_0.inv_9.Y 0.013749f
C1551 NOT8_0.S4 B1 2.87e-21
C1552 mux8_5.NAND4F_0.Y mux8_5.NAND4F_1.Y 5.28e-20
C1553 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y mux8_8.A0 1.08e-19
C1554 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y mux8_8.A0 1.08e-19
C1555 OR8_0.NOT8_0.A2 B1 0.005656f
C1556 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A VDD 1.35016f
C1557 mux8_5.A0 A1 9.63e-20
C1558 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y mux8_8.A0 1.08e-19
C1559 mux8_5.A1 mux8_5.NAND4F_3.Y 0.541275f
C1560 B2 B1 1.50454f
C1561 mux8_0.NAND4F_2.D SEL3 0.002782f
C1562 B3 B0 0.121184f
C1563 AND8_0.S1 AND8_0.NOT8_0.A2 9.72e-21
C1564 mux8_6.A0 NOT8_0.S3 0.015495f
C1565 AND8_0.NOT8_0.A1 A2 0.043465f
C1566 mux8_5.NAND4F_9.Y mux8_5.NAND4F_5.Y 0.402985f
C1567 mux8_5.A1 XOR8_0.S4 6.83e-20
C1568 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A A5 0.00194f
C1569 B5 A3 0.026323f
C1570 XOR8_0.S5 B3 0.168302f
C1571 mux8_5.NAND4F_4.B SEL0 1.60998f
C1572 mux8_8.A0 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 0.001899f
C1573 V_FLAG_0.XOR2_0.Y SEL0 4.29e-19
C1574 mux8_8.A0 mux8_5.A0 0.004073f
C1575 mux8_7.A0 MULT_0.SO 0.024039f
C1576 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 0.001201f
C1577 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT mux8_7.A0 8.09e-19
C1578 XOR8_0.S1 AND8_0.S2 3.64355f
C1579 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A VDD 1.6936f
C1580 mux8_2.NAND4F_2.D SEL0 0.229162f
C1581 AND8_0.S0 XOR8_0.S2 3.62e-20
C1582 NOT8_0.S0 MULT_0.S2 0.020734f
C1583 left_shifter_0.S7 B6 0.005473f
C1584 XOR8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A 9.55e-20
C1585 mux8_8.NAND4F_3.Y VDD 2.17571f
C1586 mux8_7.NAND4F_2.D mux8_7.NAND4F_3.Y 0.397922f
C1587 mux8_3.NAND4F_4.Y SEL1 0.30433f
C1588 mux8_7.A0 AND8_0.S1 0.015963f
C1589 mux8_6.NAND4F_8.Y mux8_6.NAND4F_6.Y 2.96e-20
C1590 mux8_1.NAND4F_1.Y mux8_2.NAND4F_8.Y 1.02e-21
C1591 mux8_4.A0 AND8_0.S0 0.013336f
C1592 mux8_6.NAND4F_8.Y mux8_6.NAND4F_9.Y 0.696806f
C1593 8bit_ADDER_0.S0 mux8_1.NAND4F_6.Y 2.97e-22
C1594 mux8_3.NAND4F_2.Y mux8_3.NAND4F_4.Y 2.04463f
C1595 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT 7.17e-20
C1596 mux8_6.NAND4F_0.Y mux8_6.NAND4F_5.Y 4.32e-19
C1597 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT 1.69e-20
C1598 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A 1.16e-19
C1599 AND8_0.S5 A5 0.006872f
C1600 AND8_0.S4 SEL2 0.076881f
C1601 8bit_ADDER_0.S2 NOT8_0.S0 0.013311f
C1602 mux8_5.NAND4F_2.Y mux8_5.NAND4F_4.Y 2.04463f
C1603 mux8_3.NAND4F_2.D AND8_0.S2 0.076916f
C1604 mux8_3.NAND4F_0.C mux8_3.NAND4F_4.B 2.13077f
C1605 A7 B3 0.047631f
C1606 left_shifter_0.S0 OR8_0.S1 0.019711f
C1607 mux8_5.A1 mux8_5.NAND4F_7.Y 5.24e-19
C1608 mux8_1.NAND4F_0.C SEL1 1.11929f
C1609 mux8_7.NAND4F_9.Y mux8_8.NAND4F_8.Y 0.001427f
C1610 mux8_5.NAND4F_0.C mux8_5.NAND4F_2.Y 0.122872f
C1611 mux8_4.NAND4F_4.Y mux8_4.NAND4F_1.Y 4.33e-19
C1612 mux8_4.NAND4F_2.D mux8_4.NAND4F_8.Y 4.88e-20
C1613 AND8_0.S0 OR8_0.NOT8_0.A0 0.001422f
C1614 mux8_8.A0 mux8_8.NAND4F_2.D 0.105266f
C1615 OR8_0.NOT8_0.A0 OR8_0.NOT8_0.A1 1.02549f
C1616 OR8_0.S7 mux8_6.NAND4F_0.C 0.065599f
C1617 OR8_0.NOT8_0.A7 OR8_0.S7 0.393091f
C1618 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 0.013137f
C1619 mux8_5.NAND4F_0.Y SEL0 0.236427f
C1620 mux8_7.NAND4F_4.Y SEL2 8.74e-20
C1621 mux8_5.NAND4F_4.Y VDD 2.21741f
C1622 mux8_1.NAND4F_3.Y mux8_1.NAND4F_8.Y 0.222524f
C1623 mux8_1.NAND4F_2.Y mux8_1.NAND4F_4.Y 2.04463f
C1624 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B 0.001075f
C1625 NOT8_0.S2 mux8_3.NAND4F_5.Y 0.288211f
C1626 mux8_7.NAND4F_4.Y mux8_7.NAND4F_1.Y 4.33e-19
C1627 mux8_5.NAND4F_0.C VDD 1.39921f
C1628 mux8_1.NAND4F_0.Y SEL0 0.236427f
C1629 XOR8_0.S7 A7 0.560993f
C1630 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A 0.186684f
C1631 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A 0.118063f
C1632 mux8_7.A0 mux8_2.NAND4F_0.C 1.67e-19
C1633 mux8_1.NAND4F_4.Y VDD 2.31569f
C1634 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 0.792412f
C1635 mux8_1.NAND4F_2.Y mux8_1.NAND4F_1.Y 3.31e-22
C1636 mux8_4.A0 mux8_4.NAND4F_2.D 0.132792f
C1637 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A 0.005938f
C1638 mux8_7.NAND4F_0.C XOR8_0.S5 0.081526f
C1639 mux8_4.NAND4F_7.Y SEL0 0.234594f
C1640 mux8_5.NAND4F_2.D SEL2 0.481922f
C1641 mux8_8.NAND4F_0.Y mux8_8.NAND4F_1.Y 5.28e-20
C1642 mux8_1.NAND4F_1.Y VDD 2.18282f
C1643 mux8_0.NAND4F_4.Y mux8_0.NAND4F_6.Y 4.33e-19
C1644 mux8_4.A0 NOT8_0.S3 1.11e-19
C1645 AND8_0.S2 mux8_8.A1 0.036917f
C1646 NOT8_0.S0 mux8_2.NAND4F_4.B 2.74e-21
C1647 NOT8_0.S5 mux8_7.NAND4F_0.Y 5.24e-19
C1648 B4 B0 0.045405f
C1649 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_2.B2 0.200037f
C1650 mux8_3.NAND4F_7.Y SEL0 0.234594f
C1651 mux8_7.A0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 0.002498f
C1652 mux8_2.NAND4F_6.Y mux8_2.NAND4F_7.Y 0.14618f
C1653 XOR8_0.S7 mux8_6.NAND4F_7.Y 9.74e-20
C1654 left_shifter_0.S0 mux8_1.NAND4F_6.Y 1.2e-19
C1655 B6 A3 0.024914f
C1656 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 1.2618f
C1657 mux8_8.A0 mux8_7.A1 0.253207f
C1658 XOR8_0.S5 B4 0.118792f
C1659 AND8_0.S3 OR8_0.NOT8_0.A2 0.002366f
C1660 mux8_0.NAND4F_9.Y mux8_0.NAND4F_7.Y 0.248336f
C1661 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 0.119902f
C1662 8bit_ADDER_0.S2 mux8_2.NAND4F_2.D 4.83e-19
C1663 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A mux8_8.A1 2.52e-19
C1664 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 1.2618f
C1665 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A mux8_7.A0 1.53e-19
C1666 mux8_2.NAND4F_0.C AND8_0.S1 0.037374f
C1667 AND8_0.S3 B2 0.077522f
C1668 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 1.2618f
C1669 AND8_0.S2 B0 0.51406f
C1670 AND8_0.NOT8_0.A7 B7 0.149348f
C1671 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A MULT_0.inv_9.Y 0.001123f
C1672 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A 0.186684f
C1673 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 1.2618f
C1674 AND8_0.NOT8_0.A0 B2 0.04157f
C1675 mux8_3.NAND4F_0.Y mux8_3.NAND4F_5.Y 4.32e-19
C1676 mux8_5.NAND4F_5.Y mux8_5.NAND4F_1.Y 0.110562f
C1677 mux8_7.NAND4F_5.Y SEL2 0.323263f
C1678 mux8_4.NAND4F_9.Y mux8_5.NAND4F_8.Y 0.001427f
C1679 mux8_8.A0 NOT8_0.S0 0.014216f
C1680 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 1.2618f
C1681 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT mux8_5.A0 0.156073f
C1682 mux8_6.NAND4F_6.Y VDD 2.17784f
C1683 mux8_6.NAND4F_2.D XOR8_0.S7 4.4e-19
C1684 OR8_0.S2 B3 0.008979f
C1685 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_1.B2 0.019892f
C1686 mux8_2.NAND4F_0.C mux8_2.NAND4F_1.Y 0.402437f
C1687 mux8_7.NAND4F_0.Y VDD 2.13487f
C1688 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 1.2618f
C1689 mux8_1.NAND4F_0.C XOR8_0.S0 0.07976f
C1690 mux8_6.NAND4F_9.Y VDD 2.28057f
C1691 mux8_7.NAND4F_5.Y mux8_7.NAND4F_1.Y 0.110562f
C1692 mux8_6.A1 B1 0.041208f
C1693 OR8_0.NOT8_0.A5 OR8_0.NOT8_0.A6 0.523978f
C1694 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B 1.2618f
C1695 mux8_6.NAND4F_2.Y SEL0 0.296519f
C1696 mux8_7.NAND4F_4.B SEL2 0.734121f
C1697 mux8_8.A0 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A 1.08e-19
C1698 mux8_0.NAND4F_2.Y SEL0 0.296554f
C1699 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A 0.001571f
C1700 B7 A2 0.084795f
C1701 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A 1.76e-19
C1702 mux8_5.A0 NOT8_0.S2 0.014305f
C1703 mux8_7.NAND4F_4.B mux8_7.NAND4F_1.Y 0.222551f
C1704 mux8_6.A0 mux8_6.NAND4F_6.Y 2.97e-22
C1705 mux8_8.NAND4F_1.Y VDD 2.1816f
C1706 mux8_5.NAND4F_3.Y mux8_5.NAND4F_8.Y 0.222524f
C1707 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B VDD 1.97601f
C1708 mux8_7.NAND4F_4.Y mux8_7.NAND4F_9.Y 5.28e-19
C1709 mux8_2.NAND4F_2.D mux8_2.NAND4F_4.B 1.27138f
C1710 A7 B4 0.060656f
C1711 NOT8_0.S4 mux8_5.NAND4F_9.Y 3.17e-20
C1712 MULT_0.S2 mux8_3.NAND4F_7.Y 5.24e-19
C1713 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y SEL3 0.733054f
C1714 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y SEL3 0.732311f
C1715 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y SEL3 0.73352f
C1716 mux8_1.NAND4F_5.Y mux8_1.NAND4F_6.Y 1.93433f
C1717 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y SEL3 0.737337f
C1718 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A mux8_8.A1 2.28e-19
C1719 V_FLAG_0.XOR2_2.Y SEL0 0.004151f
C1720 MULT_0.4bit_ADDER_0.A2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A 0.685441f
C1721 mux8_5.A0 SEL3 9.63e-20
C1722 mux8_8.A0 mux8_2.NAND4F_2.D 1.11e-19
C1723 mux8_1.NAND4F_2.D SEL0 0.229191f
C1724 AND8_0.S6 B3 0.09025f
C1725 mux8_4.NAND4F_2.Y SEL0 0.296548f
C1726 OR8_0.S1 A0 0.054686f
C1727 XOR8_0.S3 AND8_0.S4 0.029711f
C1728 VDD Y3 1.51167f
C1729 mux8_2.NAND4F_6.Y SEL0 0.353704f
C1730 B5 B0 0.045125f
C1731 AND8_0.S2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 4.5e-19
C1732 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 0.017305f
C1733 mux8_5.NAND4F_5.Y SEL0 0.12244f
C1734 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 0.087175f
C1735 mux8_7.NAND4F_9.Y mux8_7.NAND4F_5.Y 0.402985f
C1736 MULT_0.4bit_ADDER_1.B2 MULT_0.inv_9.Y 0.001146f
C1737 8bit_ADDER_0.C B3 0.001969f
C1738 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A 0.248956f
C1739 AND8_0.NOT8_0.A1 B2 0.020457f
C1740 XOR8_0.S7 SEL1 0.036401f
C1741 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B 2.43e-19
C1742 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 0.087175f
C1743 XOR8_0.S5 B5 0.28542f
C1744 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B 0.792412f
C1745 mux8_5.NAND4F_8.Y mux8_5.NAND4F_7.Y 9.84e-20
C1746 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 0.087175f
C1747 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 0.001075f
C1748 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 0.087175f
C1749 NOT8_0.S6 left_shifter_0.S7 0.029835f
C1750 mux8_3.NAND4F_0.Y mux8_3.NAND4F_8.Y 0.249057f
C1751 mux8_8.NAND4F_8.Y mux8_8.NAND4F_7.Y 9.84e-20
C1752 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 0.139263f
C1753 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 0.087175f
C1754 Y5 Y7 0.010732f
C1755 OR8_0.S1 NOT8_0.S1 7.92e-19
C1756 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A mux8_5.A0 0.200037f
C1757 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 0.087175f
C1758 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B A4 0.00981f
C1759 OR8_0.NOT8_0.A5 VDD 0.913999f
C1760 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B 0.087175f
C1761 mux8_7.A0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 1.53e-19
C1762 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B 0.087175f
C1763 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 0.127125f
C1764 MULT_0.4bit_ADDER_1.B3 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B 0.139263f
C1765 mux8_2.NAND4F_9.Y mux8_2.NAND4F_1.Y 0.222572f
C1766 MULT_0.4bit_ADDER_1.A2 A2 0.001538f
C1767 mux8_8.NAND4F_2.D mux8_8.NAND4F_8.Y 4.88e-20
C1768 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_2.B1 2.27e-19
C1769 MULT_0.SO MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A 8.21e-19
C1770 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 0.127125f
C1771 mux8_7.A1 NOT8_0.S2 0.077313f
C1772 mux8_7.A0 mux8_1.NAND4F_0.C 1.67e-19
C1773 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT 0.127988f
C1774 mux8_4.NAND4F_2.D NOT8_0.S3 4.43e-19
C1775 mux8_1.NAND4F_0.C MULT_0.SO 0.06328f
C1776 OR8_0.S7 B7 0.053529f
C1777 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 0.127125f
C1778 AND8_0.S2 OR8_0.S2 18.415499f
C1779 mux8_6.A1 AND8_0.S3 0.060145f
C1780 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 0.127125f
C1781 OR8_0.S1 SEL2 0.095695f
C1782 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A 0.127125f
C1783 A7 B5 0.092166f
C1784 mux8_1.NAND4F_4.B NOT8_0.S0 0.105156f
C1785 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.B2 0.697999f
C1786 AND8_0.NOT8_0.A7 A4 0.00584f
C1787 mux8_5.A0 AND8_0.S4 0.059486f
C1788 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A 0.127125f
C1789 NOT8_0.S0 NOT8_0.S2 7.42e-19
C1790 mux8_7.NAND4F_0.C SEL1 1.12184f
C1791 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A 0.127125f
C1792 mux8_2.NAND4F_0.C mux8_2.NAND4F_9.Y 4.79e-21
C1793 OR8_0.S7 SEL0 1.05469f
C1794 mux8_8.A0 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 0.02828f
C1795 8bit_ADDER_0.S2 mux8_1.NAND4F_2.D 4.83e-19
C1796 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y A2 5.91e-19
C1797 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A 2.56e-19
C1798 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A 1.16e-19
C1799 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B 0.001322f
C1800 left_shifter_0.S0 XOR8_0.S1 0.022426f
C1801 OR8_0.NOT8_0.A6 A5 0.270837f
C1802 mux8_8.NAND4F_5.Y mux8_8.NAND4F_6.Y 1.93433f
C1803 NOT8_0.S6 mux8_8.NAND4F_6.Y 0.79864f
C1804 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y A2 0.001931f
C1805 NOT8_0.S4 mux8_5.NAND4F_1.Y 0.55011f
C1806 NOT8_0.S7 mux8_6.NAND4F_6.Y 0.79864f
C1807 MULT_0.4bit_ADDER_1.B2 B0 1.58e-19
C1808 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A VDD 1.69389f
C1809 AND8_0.S6 B4 0.086459f
C1810 NOT8_0.S7 mux8_6.NAND4F_9.Y 3.17e-20
C1811 A4 A2 0.023674f
C1812 mux8_2.NAND4F_2.Y NOT8_0.S1 1.43e-19
C1813 AND8_0.S3 AND8_0.S5 0.00307f
C1814 left_shifter_0.S7 SEL2 0.097411f
C1815 mux8_5.A0 mux8_5.NAND4F_2.D 0.138011f
C1816 B6 B0 0.044886f
C1817 mux8_6.A1 mux8_6.NAND4F_0.C 0.078065f
C1818 mux8_1.NAND4F_6.Y SEL2 0.419676f
C1819 AND8_0.S2 SEL1 0.111612f
C1820 8bit_ADDER_0.C B4 0.001202f
C1821 mux8_2.NAND4F_2.D mux8_2.NAND4F_3.Y 0.397922f
C1822 AND8_0.S0 mux8_1.NAND4F_4.Y 0.402481f
C1823 mux8_0.NAND4F_4.B mux8_0.NAND4F_4.Y 0.275773f
C1824 XOR8_0.S5 B6 0.072816f
C1825 A3 A0 0.725741f
C1826 A2 A1 0.854639f
C1827 AND8_0.S2 mux8_3.NAND4F_2.Y 1.24e-19
C1828 mux8_2.NAND4F_2.Y SEL2 3.71e-20
C1829 8bit_ADDER_0.S0 B0 5.02e-19
C1830 mux8_1.NAND4F_0.C mux8_2.NAND4F_0.C 0.00173f
C1831 mux8_0.NAND4F_4.Y mux8_0.NAND4F_7.Y 4.32e-19
C1832 AND8_0.S3 mux8_4.NAND4F_4.Y 0.402481f
C1833 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 0.792412f
C1834 mux8_5.NAND4F_9.Y mux8_5.NAND4F_7.Y 0.248336f
C1835 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B A3 0.950228f
C1836 mux8_6.NAND4F_0.C mux8_6.NAND4F_4.Y 0.049743f
C1837 mux8_0.NAND4F_9.Y SEL0 2.8e-19
C1838 mux8_2.NAND4F_4.B mux8_2.NAND4F_6.Y 0.187883f
C1839 AND8_0.NOT8_0.A2 B3 0.052101f
C1840 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 0.001913f
C1841 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT A0 7.25e-19
C1842 mux8_6.NAND4F_5.Y SEL2 0.323173f
C1843 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_1.B2 0.200037f
C1844 AND8_0.S2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A 1.98e-19
C1845 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 0.118063f
C1846 NOT8_0.S4 B7 0.023656f
C1847 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 0.118063f
C1848 mux8_3.NAND4F_9.Y mux8_3.NAND4F_1.Y 0.222572f
C1849 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B 0.001075f
C1850 MULT_0.4bit_ADDER_0.A2 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT 0.010334f
C1851 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 0.118063f
C1852 B7 B2 0.077735f
C1853 mux8_8.A0 mux8_1.NAND4F_2.D 1.8e-19
C1854 mux8_4.NAND4F_0.C mux8_5.NAND4F_2.D 4.6e-19
C1855 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 2.43e-19
C1856 OR8_0.NOT8_0.A5 AND8_0.S7 0.082749f
C1857 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 0.118063f
C1858 AND8_0.S5 OR8_0.NOT8_0.A7 0.041298f
C1859 MULT_0.4bit_ADDER_0.B2 A0 0.02313f
C1860 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A 0.118063f
C1861 AND8_0.S2 mux8_4.A1 0.038541f
C1862 XOR8_0.S6 VDD 0.938484f
C1863 left_shifter_0.S0 mux8_8.A1 0.046467f
C1864 mux8_8.NAND4F_6.Y SEL2 0.419676f
C1865 MULT_0.4bit_ADDER_1.A2 MULT_0.4bit_ADDER_2.B2 0.451291f
C1866 mux8_4.NAND4F_1.Y VDD 2.1816f
C1867 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A 0.118063f
C1868 A7 B6 0.180404f
C1869 NOT8_0.S4 SEL0 1.10123f
C1870 mux8_7.A1 AND8_0.S4 0.028565f
C1871 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A A4 0.00194f
C1872 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A 0.118063f
C1873 mux8_7.A0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 0.002498f
C1874 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 0.012305f
C1875 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A 0.118063f
C1876 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 0.00162f
C1877 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A mux8_4.A1 0.200075f
C1878 mux8_3.NAND4F_1.Y VDD 2.1816f
C1879 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 0.209959f
C1880 mux8_6.NAND4F_0.Y mux8_6.NAND4F_7.Y 0.08762f
C1881 mux8_8.NAND4F_0.Y mux8_8.NAND4F_2.Y 0.170507f
C1882 VDD A5 2.18833f
C1883 mux8_3.NAND4F_3.Y SEL2 2.96e-20
C1884 mux8_6.A0 XOR8_0.S6 0.088001f
C1885 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 0.209959f
C1886 XOR8_0.S0 AND8_0.S2 0.08216f
C1887 left_shifter_0.S0 B0 0.962264f
C1888 mux8_0.NAND4F_0.C mux8_0.NAND4F_0.Y 0.223896f
C1889 MULT_0.inv_15.Y A3 0.010751f
C1890 mux8_7.A1 mux8_7.NAND4F_4.Y 0.157118f
C1891 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 0.209959f
C1892 mux8_5.NAND4F_3.Y mux8_5.NAND4F_1.Y 0.086984f
C1893 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 0.209959f
C1894 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT mux8_5.A0 0.699206f
C1895 AND8_0.S6 B5 0.067804f
C1896 ZFLAG_0.nor4_0.Y Y4 6.55e-20
C1897 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 0.209959f
C1898 mux8_5.A1 mux8_5.NAND4F_2.Y 1.16938f
C1899 mux8_7.NAND4F_2.D SEL0 0.229596f
C1900 AND8_0.NOT8_0.A1 AND8_0.S5 8.31e-22
C1901 XOR8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A 2.35e-19
C1902 XOR8_0.S4 mux8_5.NAND4F_1.Y 0.404949f
C1903 OR8_0.S7 A4 0.102316f
C1904 mux8_6.NAND4F_2.D mux8_6.NAND4F_0.Y 0.184536f
C1905 mux8_6.NAND4F_0.C mux8_6.NAND4F_4.B 2.13077f
C1906 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B 0.209959f
C1907 mux8_6.A0 A5 1.52e-19
C1908 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B 0.209959f
C1909 AND8_0.S1 B3 0.030859f
C1910 NOT8_0.S2 mux8_3.NAND4F_7.Y 0.431664f
C1911 mux8_8.A0 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A 0.01036f
C1912 mux8_7.NAND4F_0.C mux8_8.NAND4F_0.C 0.001594f
C1913 MULT_0.SO MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT 4.62e-19
C1914 XOR8_0.S1 A0 0.070954f
C1915 mux8_5.A1 VDD 1.13834f
C1916 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A 2.37e-19
C1917 XOR8_0.S6 A6 0.559495f
C1918 mux8_2.NAND4F_8.Y mux8_2.NAND4F_5.Y 0.001122f
C1919 ZFLAG_0.nor4_1.Y Y7 0.592953f
C1920 AND8_0.NOT8_0.A6 AND8_0.NOT8_0.A7 0.248603f
C1921 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B VDD 1.97106f
C1922 mux8_8.NAND4F_9.Y mux8_8.NAND4F_5.Y 0.402985f
C1923 NOT8_0.S6 mux8_8.NAND4F_9.Y 3.17e-20
C1924 mux8_5.NAND4F_4.B AND8_0.S4 1.04047f
C1925 VDD C 0.862192f
C1926 mux8_0.NAND4F_6.Y mux8_1.NAND4F_2.Y 0.002218f
C1927 A6 A5 0.062934f
C1928 MULT_0.inv_9.Y A0 2.76e-19
C1929 AND8_0.NOT8_0.A4 B3 0.013409f
C1930 mux8_3.NAND4F_4.B SEL0 1.61043f
C1931 mux8_7.NAND4F_2.D mux8_7.NAND4F_2.Y 0.339934f
C1932 mux8_8.NAND4F_2.Y VDD 2.1749f
C1933 mux8_6.A0 mux8_5.A1 0.026863f
C1934 mux8_7.A1 mux8_7.NAND4F_5.Y 1.57e-19
C1935 mux8_0.NAND4F_6.Y VDD 2.17811f
C1936 mux8_4.NAND4F_9.Y SEL0 2.8e-19
C1937 mux8_1.NAND4F_9.Y mux8_1.NAND4F_5.Y 0.402985f
C1938 XOR8_0.S3 left_shifter_0.S7 1.28e-20
C1939 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT 0.119902f
C1940 mux8_6.NAND4F_3.Y mux8_6.NAND4F_5.Y 4.33e-19
C1941 XOR8_0.S1 NOT8_0.S1 19.954601f
C1942 mux8_3.NAND4F_0.Y mux8_3.NAND4F_7.Y 0.08762f
C1943 mux8_5.NAND4F_1.Y mux8_5.NAND4F_7.Y 0.617483f
C1944 mux8_7.NAND4F_7.Y SEL2 0.176544f
C1945 mux8_7.A1 mux8_7.NAND4F_4.B 0.039141f
C1946 MULT_0.4bit_ADDER_1.A2 B2 0.001982f
C1947 XOR8_0.S4 B7 0.037005f
C1948 AND8_0.S2 AND8_0.NOT8_0.A2 0.396516f
C1949 mux8_7.A0 mux8_7.NAND4F_0.C 0.083261f
C1950 V_FLAG_0.XOR2_2.B A7 0.31537f
C1951 mux8_7.NAND4F_1.Y mux8_7.NAND4F_7.Y 0.617483f
C1952 mux8_5.NAND4F_0.C mux8_5.NAND4F_4.Y 0.049743f
C1953 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 0.001075f
C1954 8bit_ADDER_0.S2 B2 5.02e-19
C1955 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_1.B3 0.184903f
C1956 mux8_5.NAND4F_2.D mux8_5.NAND4F_4.B 1.27138f
C1957 mux8_2.NAND4F_5.Y VDD 2.19971f
C1958 mux8_5.NAND4F_3.Y SEL0 0.360934f
C1959 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A 2.57e-19
C1960 AND8_0.S2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 9.92e-19
C1961 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 0.017305f
C1962 mux8_5.A0 OR8_0.S1 0.021801f
C1963 XOR8_0.S2 mux8_3.NAND4F_1.Y 0.404949f
C1964 mux8_1.NAND4F_2.Y mux8_1.NAND4F_8.Y 0.222339f
C1965 mux8_3.NAND4F_0.C mux8_3.NAND4F_9.Y 4.79e-21
C1966 XOR8_0.S4 SEL0 0.171969f
C1967 NOT8_0.S5 B1 8.31e-22
C1968 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B 0.792412f
C1969 AND8_0.S7 XOR8_0.S6 1.8592f
C1970 mux8_8.A1 mux8_8.NAND4F_5.Y 1.57e-19
C1971 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B 2.43e-19
C1972 mux8_1.NAND4F_3.Y SEL0 0.360934f
C1973 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A VDD 1.30818f
C1974 mux8_8.A1 NOT8_0.S6 0.051334f
C1975 XOR8_0.S1 SEL2 0.195221f
C1976 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y B2 0.001436f
C1977 mux8_1.NAND4F_8.Y VDD 3.42138f
C1978 mux8_4.A0 mux8_4.NAND4F_1.Y 5.23e-19
C1979 mux8_1.NAND4F_4.Y mux8_1.NAND4F_1.Y 4.33e-19
C1980 mux8_1.NAND4F_2.D mux8_1.NAND4F_4.B 1.27138f
C1981 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A mux8_5.A0 4.03e-19
C1982 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y B2 0.001926f
C1983 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B 0.008371f
C1984 mux8_6.A1 B7 0.277106f
C1985 mux8_8.A1 A0 0.013504f
C1986 mux8_8.NAND4F_3.Y mux8_8.NAND4F_1.Y 0.086984f
C1987 mux8_0.NAND4F_8.Y mux8_0.NAND4F_6.Y 2.96e-20
C1988 AND8_0.S6 B6 0.049377f
C1989 mux8_1.NAND4F_6.Y mux8_1.NAND4F_7.Y 0.14618f
C1990 MULT_0.S2 mux8_3.NAND4F_4.B 0.039141f
C1991 B2 A4 0.019383f
C1992 mux8_7.A0 AND8_0.S2 0.015963f
C1993 NOT8_0.S5 mux8_7.NAND4F_3.Y 3.24e-22
C1994 AND8_0.S7 A5 0.042001f
C1995 MULT_0.inv_15.Y MULT_0.inv_9.Y 0.002801f
C1996 mux8_7.A0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 1.53e-19
C1997 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A 0.200037f
C1998 mux8_8.NAND4F_9.Y SEL2 1.49e-20
C1999 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.B2 0.69756f
C2000 AND8_0.NOT8_0.A3 B1 1.51e-22
C2001 SEL3 A2 0.284203f
C2002 mux8_3.NAND4F_0.C VDD 1.40145f
C2003 VDD B1 8.25688f
C2004 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 1.01138f
C2005 8bit_ADDER_0.S0 SEL1 0.334783f
C2006 NOT8_0.S6 XOR8_0.S5 0.023818f
C2007 mux8_5.A1 XOR8_0.S2 0.138392f
C2008 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 1.01138f
C2009 B0 A0 57.079395f
C2010 mux8_6.A1 SEL0 1.13725f
C2011 left_shifter_0.S0 OR8_0.S2 0.024846f
C2012 NOT8_0.S7 XOR8_0.S6 0.030191f
C2013 mux8_5.NAND4F_4.B mux8_7.NAND4F_4.B 0.001581f
C2014 mux8_3.NAND4F_2.D SEL2 0.481313f
C2015 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A 0.186684f
C2016 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 1.01138f
C2017 V_FLAG_0.XOR2_2.Y SEL3 0.240956f
C2018 OR8_0.NOT8_0.A2 A1 0.219668f
C2019 left_shifter_0.S0 mux8_2.NAND4F_4.Y 1.02e-21
C2020 mux8_3.NAND4F_3.Y mux8_3.NAND4F_5.Y 4.33e-19
C2021 B2 A1 35.928f
C2022 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A 1.01138f
C2023 XOR8_0.S3 A3 0.585343f
C2024 8bit_ADDER_0.S2 mux8_3.NAND4F_4.B 1.52147f
C2025 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A 1.01138f
C2026 NOT8_0.S1 mux8_8.A1 0.017326f
C2027 mux8_7.NAND4F_3.Y VDD 2.17571f
C2028 AND8_0.S1 AND8_0.S2 6.94501f
C2029 mux8_8.A0 NOT8_0.S4 0.015234f
C2030 mux8_5.NAND4F_2.D mux8_5.NAND4F_0.Y 0.184536f
C2031 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A 1.01138f
C2032 mux8_5.NAND4F_7.Y SEL0 0.234594f
C2033 8bit_ADDER_0.C 8bit_ADDER_0.S0 0.055679f
C2034 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A A6 0.008956f
C2035 mux8_7.NAND4F_9.Y mux8_7.NAND4F_7.Y 0.248336f
C2036 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A 1.01138f
C2037 mux8_6.NAND4F_4.Y SEL0 0.111961f
C2038 AND8_0.NOT8_0.A4 B4 0.245546f
C2039 AND8_0.S5 B7 0.050098f
C2040 mux8_8.A0 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B 0.005184f
C2041 mux8_0.NAND4F_4.Y SEL0 0.117031f
C2042 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A 1.21e-19
C2043 NOT8_0.S1 B0 0.576725f
C2044 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A mux8_7.A1 0.200037f
C2045 mux8_5.NAND4F_2.Y mux8_5.NAND4F_8.Y 0.222339f
C2046 mux8_7.NAND4F_8.Y mux8_7.NAND4F_9.Y 0.696806f
C2047 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A VDD 1.69307f
C2048 mux8_8.A1 SEL2 0.077532f
C2049 AND8_0.S5 SEL0 0.134346f
C2050 mux8_6.NAND4F_5.Y mux8_6.NAND4F_1.Y 0.110562f
C2051 B1 A6 0.022403f
C2052 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A A0 0.002461f
C2053 mux8_6.NAND4F_9.Y mux8_6.NAND4F_6.Y 0.222562f
C2054 OR8_0.S1 mux8_7.A1 0.010804f
C2055 mux8_5.NAND4F_8.Y VDD 3.38981f
C2056 left_shifter_0.S0 SEL1 0.115279f
C2057 mux8_2.NAND4F_4.B mux8_3.NAND4F_4.B 0.001468f
C2058 mux8_4.NAND4F_6.Y SEL2 0.419676f
C2059 A7 A0 0.100898f
C2060 mux8_4.A1 mux8_4.NAND4F_0.Y 0.43187f
C2061 mux8_7.A0 B5 5.02e-19
C2062 mux8_1.NAND4F_9.Y SEL2 1.49e-20
C2063 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y A3 3.97e-19
C2064 mux8_1.NAND4F_5.Y mux8_2.NAND4F_4.Y 0.0024f
C2065 8bit_ADDER_0.S0 XOR8_0.S0 0.009216f
C2066 OR8_0.NOT8_0.A6 OR8_0.NOT8_0.A7 1.2593f
C2067 mux8_3.NAND4F_6.Y SEL2 0.419676f
C2068 mux8_4.NAND4F_4.Y SEL0 0.117021f
C2069 NOT8_0.S0 OR8_0.S1 0.018734f
C2070 AND8_0.S4 A2 0.057817f
C2071 XOR8_0.S5 SEL2 0.236391f
C2072 mux8_0.NAND4F_0.Y mux8_0.NAND4F_1.Y 5.28e-20
C2073 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 2.43e-19
C2074 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B A0 0.001659f
C2075 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B A3 0.00981f
C2076 mux8_5.A0 A3 0.433667f
C2077 XOR8_0.S4 A4 0.558383f
C2078 XOR8_0.S5 mux8_7.NAND4F_1.Y 0.404949f
C2079 AND8_0.S5 mux8_7.NAND4F_2.Y 1.24e-19
C2080 MULT_0.4bit_ADDER_0.A2 MULT_0.4bit_ADDER_1.B2 0.446124f
C2081 AND8_0.S2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A 1.55e-19
C2082 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 0.001913f
C2083 mux8_6.NAND4F_4.B SEL0 1.57298f
C2084 mux8_3.NAND4F_0.C XOR8_0.S2 0.079804f
C2085 mux8_8.NAND4F_6.Y mux8_8.NAND4F_7.Y 0.14618f
C2086 XOR8_0.S2 B1 0.133881f
C2087 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B 0.001075f
C2088 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B 0.792412f
C2089 mux8_3.NAND4F_3.Y mux8_3.NAND4F_8.Y 0.222524f
C2090 left_shifter_0.S0 mux8_4.A1 0.030877f
C2091 mux8_8.NAND4F_4.B mux8_6.NAND4F_4.B 0.001581f
C2092 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A 0.005938f
C2093 AND8_0.S3 AND8_0.NOT8_0.A3 0.396187f
C2094 AND8_0.S4 mux8_5.NAND4F_5.Y 5.23e-19
C2095 AND8_0.S3 VDD 1.94628f
C2096 mux8_4.A0 mux8_3.NAND4F_0.C 2.46e-19
C2097 ZFLAG_0.nor4_0.Y Y1 0.045328f
C2098 mux8_8.NAND4F_2.D mux8_8.NAND4F_6.Y 2.96e-20
C2099 AND8_0.NOT8_0.A0 AND8_0.NOT8_0.A3 3e-19
C2100 mux8_1.NAND4F_5.Y SEL1 0.30645f
C2101 AND8_0.NOT8_0.A0 VDD 2.36084f
C2102 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 0.120014f
C2103 mux8_7.A0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 0.002498f
C2104 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT A0 0.003441f
C2105 NOT8_0.S0 mux8_1.NAND4F_6.Y 0.79864f
C2106 mux8_4.NAND4F_2.D mux8_4.NAND4F_1.Y 2.96e-20
C2107 AND8_0.S0 mux8_5.A1 0.106725f
C2108 mux8_8.A0 XOR8_0.S4 0.024828f
C2109 A7 SEL2 4.95e-19
C2110 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT VDD 3.25348f
C2111 left_shifter_0.S0 XOR8_0.S0 0.008943f
C2112 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT 1.58859f
C2113 mux8_5.NAND4F_5.Y mux8_7.NAND4F_4.Y 0.002218f
C2114 OR8_0.S2 A0 0.350579f
C2115 NOT8_0.S3 mux8_4.NAND4F_1.Y 0.55011f
C2116 mux8_2.NAND4F_2.D OR8_0.S1 0.08162f
C2117 mux8_6.A0 AND8_0.S3 0.043559f
C2118 OR8_0.NOT8_0.A0 B1 0.02617f
C2119 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT mux8_5.A0 0.008948f
C2120 ZFLAG_0.nor4_1.Y Z 0.001454f
C2121 mux8_7.NAND4F_6.Y mux8_8.NAND4F_2.Y 0.002218f
C2122 mux8_0.NAND4F_4.B VDD 1.20108f
C2123 mux8_3.NAND4F_2.D mux8_3.NAND4F_5.Y 9.34e-20
C2124 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_2.B2 9.98e-20
C2125 mux8_6.A1 A1 0.048792f
C2126 mux8_5.NAND4F_2.D mux8_5.NAND4F_5.Y 9.34e-20
C2127 mux8_5.NAND4F_2.Y mux8_5.NAND4F_9.Y 2.96e-20
C2128 mux8_6.NAND4F_7.Y SEL2 0.176544f
C2129 mux8_0.NAND4F_2.D A7 5.07e-19
C2130 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 0.703381f
C2131 OR8_0.NOT8_0.A3 AND8_0.S4 0.08086f
C2132 Y0 Y1 6.22215f
C2133 mux8_0.NAND4F_0.C SEL2 1.46809f
C2134 mux8_0.NAND4F_7.Y VDD 2.14052f
C2135 mux8_8.A0 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A 0.002364f
C2136 NOT8_0.S2 B2 0.436881f
C2137 mux8_6.NAND4F_0.C VDD 1.3868f
C2138 OR8_0.NOT8_0.A7 VDD 0.731063f
C2139 AND8_0.S5 A4 0.474703f
C2140 NOT8_0.S1 OR8_0.S2 0.014964f
C2141 mux8_5.NAND4F_9.Y VDD 2.28309f
C2142 mux8_6.NAND4F_2.D SEL2 0.445231f
C2143 mux8_8.NAND4F_5.Y SEL1 0.306449f
C2144 NOT8_0.S6 SEL1 0.072828f
C2145 mux8_2.NAND4F_4.Y NOT8_0.S1 2.18e-19
C2146 AND8_0.S6 mux8_8.NAND4F_5.Y 5.23e-19
C2147 NOT8_0.S6 AND8_0.S6 0.031344f
C2148 mux8_0.NAND4F_2.D mux8_0.NAND4F_0.C 1.55301f
C2149 mux8_5.A0 XOR8_0.S1 0.022511f
C2150 mux8_1.NAND4F_6.Y mux8_2.NAND4F_2.D 1.02e-21
C2151 mux8_5.A1 NOT8_0.S3 0.027789f
C2152 AND8_0.S4 OR8_0.S7 0.001081f
C2153 mux8_7.A0 8bit_ADDER_0.S0 0.057335f
C2154 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT A6 0.129004f
C2155 mux8_8.A1 XOR8_0.S3 0.039623f
C2156 mux8_8.NAND4F_3.Y XOR8_0.S6 5.23e-19
C2157 8bit_ADDER_0.S0 MULT_0.SO 10.241f
C2158 mux8_6.A0 mux8_6.NAND4F_0.C 0.097437f
C2159 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A 0.186684f
C2160 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A VDD 1.35444f
C2161 XOR8_0.S0 mux8_1.NAND4F_5.Y 0.602395f
C2162 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 8bit_ADDER_0.S0 0.179046f
C2163 mux8_4.NAND4F_5.Y mux8_4.NAND4F_6.Y 1.93433f
C2164 mux8_7.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B 0.005343f
C2165 mux8_2.NAND4F_2.D mux8_2.NAND4F_2.Y 0.339934f
C2166 SEL3 B2 1.20652f
C2167 OR8_0.S2 SEL2 0.096671f
C2168 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT A2 0.003452f
C2169 AND8_0.S2 mux8_3.NAND4F_4.Y 0.402481f
C2170 XOR8_0.S3 mux8_4.NAND4F_6.Y 0.520706f
C2171 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT mux8_7.A1 0.711947f
C2172 AND8_0.NOT8_0.A1 AND8_0.NOT8_0.A3 9.06e-20
C2173 AND8_0.NOT8_0.A1 VDD 2.39075f
C2174 mux8_2.NAND4F_4.Y SEL2 8.84e-20
C2175 mux8_0.NAND4F_8.Y mux8_0.NAND4F_7.Y 9.84e-20
C2176 mux8_8.A0 AND8_0.S5 0.017059f
C2177 8bit_ADDER_0.C A0 0.050713f
C2178 mux8_2.NAND4F_0.Y mux8_2.NAND4F_8.Y 0.249057f
C2179 mux8_3.NAND4F_5.Y mux8_3.NAND4F_6.Y 1.93433f
C2180 XOR8_0.S2 AND8_0.S3 0.187998f
C2181 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A A0 8.48e-19
C2182 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A A3 0.00194f
C2183 mux8_5.A0 mux8_3.NAND4F_2.D 2.18e-19
C2184 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A 0.248956f
C2185 XOR8_0.S3 XOR8_0.S5 0.121318f
C2186 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A A0 0.008956f
C2187 OR8_0.NOT8_0.A7 A6 0.260106f
C2188 AND8_0.S2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B 0.001185f
C2189 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 0.017305f
C2190 AND8_0.S0 B1 0.049026f
C2191 OR8_0.NOT8_0.A1 B1 0.053203f
C2192 mux8_3.NAND4F_4.B NOT8_0.S2 0.105153f
C2193 NOT8_0.S1 SEL1 0.074865f
C2194 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A VDD 1.33101f
C2195 mux8_2.NAND4F_8.Y mux8_2.NAND4F_7.Y 9.84e-20
C2196 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B 2.43e-19
C2197 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B 0.792412f
C2198 mux8_8.NAND4F_9.Y mux8_8.NAND4F_7.Y 0.248336f
C2199 mux8_4.A0 AND8_0.S3 0.059486f
C2200 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT MULT_0.S2 0.14546f
C2201 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A mux8_5.A0 2.04e-19
C2202 mux8_7.A0 left_shifter_0.S0 0.017149f
C2203 mux8_3.NAND4F_2.D mux8_3.NAND4F_8.Y 4.88e-20
C2204 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B 0.139263f
C2205 MULT_0.SO left_shifter_0.S0 1.34e-21
C2206 mux8_7.A1 mux8_7.NAND4F_7.Y 5.24e-19
C2207 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A 6.39e-19
C2208 mux8_7.A0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 1.53e-19
C2209 OR8_0.NOT8_0.A0 AND8_0.S3 0.035283f
C2210 SEL2 SEL1 52.0979f
C2211 mux8_1.NAND4F_9.Y mux8_1.NAND4F_7.Y 0.248336f
C2212 AND8_0.S6 SEL2 0.086808f
C2213 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y B0 0.207433f
C2214 mux8_6.NAND4F_3.Y mux8_6.NAND4F_7.Y 5.28e-20
C2215 XOR8_0.S0 A0 0.558361f
C2216 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y B0 0.005392f
C2217 mux8_8.NAND4F_0.Y mux8_8.NAND4F_4.Y 0.28646f
C2218 mux8_8.NAND4F_3.Y mux8_8.NAND4F_2.Y 1.63543f
C2219 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y B0 0.005392f
C2220 mux8_3.NAND4F_2.Y SEL2 3.61e-20
C2221 mux8_7.NAND4F_1.Y SEL1 2.35e-20
C2222 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y B0 0.005392f
C2223 mux8_1.NAND4F_4.B mux8_1.NAND4F_3.Y 0.223331f
C2224 mux8_3.NAND4F_0.C mux8_4.NAND4F_2.D 4.59e-19
C2225 mux8_2.NAND4F_0.Y VDD 2.13551f
C2226 mux8_0.NAND4F_0.C mux8_0.NAND4F_3.Y 0.399921f
C2227 mux8_7.A1 mux8_7.NAND4F_8.Y 1.16e-22
C2228 mux8_5.NAND4F_2.Y mux8_5.NAND4F_1.Y 3.31e-22
C2229 NOT8_0.S4 AND8_0.S4 0.018009f
C2230 NOT8_0.S1 mux8_4.A1 0.019183f
C2231 8bit_ADDER_0.S0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 0.005184f
C2232 left_shifter_0.S0 AND8_0.S1 0.170311f
C2233 OR8_0.NOT8_0.A2 AND8_0.S4 0.005052f
C2234 NOT8_0.S3 B1 0.002954f
C2235 8bit_ADDER_0.C SEL2 0.113055f
C2236 mux8_5.A1 mux8_5.NAND4F_4.Y 0.157118f
C2237 XOR8_0.S1 mux8_7.A1 0.012f
C2238 OR8_0.S1 A2 0.036777f
C2239 AND8_0.S4 B2 0.114462f
C2240 mux8_0.NAND4F_2.D SEL1 3.36948f
C2241 mux8_2.NAND4F_7.Y VDD 2.14031f
C2242 mux8_6.NAND4F_2.D mux8_6.NAND4F_3.Y 0.397922f
C2243 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A A6 0.685441f
C2244 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A MULT_0.inv_9.Y 0.001189f
C2245 mux8_5.A1 mux8_5.NAND4F_0.C 0.063475f
C2246 AND8_0.S7 mux8_6.NAND4F_0.C 0.051868f
C2247 mux8_6.NAND4F_8.Y SEL0 4.08e-19
C2248 OR8_0.NOT8_0.A7 AND8_0.S7 0.04483f
C2249 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A 8bit_ADDER_0.S0 0.200075f
C2250 mux8_5.NAND4F_1.Y VDD 2.1816f
C2251 mux8_8.A1 mux8_8.NAND4F_7.Y 5.24e-19
C2252 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A A2 0.008967f
C2253 XOR8_0.S0 NOT8_0.S1 2.33e-19
C2254 NOT8_0.S0 XOR8_0.S1 0.023433f
C2255 MULT_0.inv_9.Y mux8_7.A1 0.447782f
C2256 XOR8_0.S6 mux8_8.NAND4F_1.Y 0.404949f
C2257 mux8_0.NAND4F_2.D 8bit_ADDER_0.C 0.104289f
C2258 mux8_4.A1 SEL2 0.077261f
C2259 OR8_0.S1 mux8_2.NAND4F_6.Y 5.23e-19
C2260 MULT_0.SO mux8_1.NAND4F_5.Y 1.57e-19
C2261 NOT8_0.S4 mux8_5.NAND4F_2.D 4.43e-19
C2262 mux8_3.NAND4F_8.Y mux8_3.NAND4F_6.Y 2.96e-20
C2263 MULT_0.4bit_ADDER_0.A2 A0 6.05e-19
C2264 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.B1 0.178362f
C2265 mux8_8.A1 mux8_8.NAND4F_2.D 0.107639f
C2266 mux8_8.NAND4F_0.Y SEL0 0.236427f
C2267 NOT8_0.S5 B7 0.023713f
C2268 mux8_8.NAND4F_0.C mux8_8.NAND4F_5.Y 0.051024f
C2269 mux8_8.NAND4F_4.Y VDD 2.21738f
C2270 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B 0.139263f
C2271 NOT8_0.S6 mux8_8.NAND4F_0.C 0.05521f
C2272 left_shifter_0.S0 mux8_2.NAND4F_0.C 3.2e-21
C2273 mux8_2.NAND4F_8.Y SEL0 4.08e-19
C2274 mux8_7.NAND4F_2.D mux8_7.NAND4F_4.Y 0.349681f
C2275 NOT8_0.S7 mux8_6.NAND4F_0.C 0.067919f
C2276 AND8_0.S5 AND8_0.NOT8_0.A6 1e-19
C2277 AND8_0.NOT8_0.A5 AND8_0.S6 0.47388f
C2278 mux8_4.NAND4F_0.C mux8_4.NAND4F_6.Y 0.142729f
C2279 B4 B3 3.73881f
C2280 mux8_7.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A 3.63e-19
C2281 XOR8_0.S0 SEL2 0.191879f
C2282 mux8_6.NAND4F_2.Y mux8_6.NAND4F_5.Y 4.33e-19
C2283 mux8_3.NAND4F_3.Y mux8_3.NAND4F_7.Y 5.28e-20
C2284 mux8_1.NAND4F_5.Y AND8_0.S1 1.02e-21
C2285 NOT8_0.S5 SEL0 1.1026f
C2286 OR8_0.S2 mux8_3.NAND4F_5.Y 2.34e-19
C2287 AND8_0.S0 AND8_0.S3 1.26e-19
C2288 mux8_3.NAND4F_9.Y SEL0 2.8e-19
C2289 AND8_0.S3 OR8_0.NOT8_0.A1 0.159746f
C2290 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A mux8_8.A1 0.200037f
C2291 mux8_1.NAND4F_2.D mux8_1.NAND4F_6.Y 2.96e-20
C2292 AND8_0.S2 B3 0.19125f
C2293 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 0.792412f
C2294 AND8_0.S0 AND8_0.NOT8_0.A0 0.397836f
C2295 VDD B7 5.21f
C2296 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT 0.127988f
C2297 mux8_5.NAND4F_2.Y SEL0 0.296538f
C2298 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT VDD 3.56168f
C2299 mux8_8.NAND4F_6.Y mux8_6.NAND4F_2.Y 0.002218f
C2300 AND8_0.S2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A 2.07e-19
C2301 mux8_2.NAND4F_2.D XOR8_0.S1 4.4e-19
C2302 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 0.001913f
C2303 mux8_8.A1 mux8_7.A1 12.6993f
C2304 mux8_1.NAND4F_4.Y mux8_1.NAND4F_8.Y 0.404949f
C2305 mux8_1.NAND4F_2.Y SEL0 0.296533f
C2306 mux8_0.NAND4F_1.Y SEL2 0.37854f
C2307 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B 0.001075f
C2308 mux8_2.NAND4F_2.Y mux8_2.NAND4F_6.Y 0.08709f
C2309 mux8_6.A0 B7 0.006767f
C2310 mux8_7.NAND4F_2.D mux8_7.NAND4F_5.Y 9.34e-20
C2311 VDD SEL0 9.39487f
C2312 mux8_6.NAND4F_1.Y mux8_6.NAND4F_7.Y 0.617483f
C2313 NOT8_0.S0 mux8_8.A1 0.099863f
C2314 MULT_0.4bit_ADDER_2.B2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A 0.248556f
C2315 mux8_7.A0 A0 6.44e-20
C2316 mux8_8.NAND4F_2.Y mux8_8.NAND4F_1.Y 3.31e-22
C2317 VDD Y4 1.52229f
C2318 mux8_7.A1 B0 0.006586f
C2319 MULT_0.SO A0 0.008355f
C2320 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 0.012283f
C2321 NOT8_0.S5 mux8_7.NAND4F_2.Y 1.43e-19
C2322 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT 0.00162f
C2323 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT A0 0.129004f
C2324 AND8_0.S4 XOR8_0.S4 1.69e-19
C2325 mux8_4.NAND4F_2.D AND8_0.S3 0.076916f
C2326 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_1.B2 9.98e-20
C2327 mux8_8.NAND4F_4.B VDD 1.19418f
C2328 mux8_4.NAND4F_5.Y SEL1 0.306449f
C2329 mux8_7.A0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 0.002498f
C2330 mux8_7.NAND4F_2.D mux8_7.NAND4F_4.B 1.27138f
C2331 mux8_0.NAND4F_2.D mux8_0.NAND4F_1.Y 2.96e-20
C2332 mux8_4.NAND4F_4.B SEL2 0.734121f
C2333 mux8_7.A1 XOR8_0.S5 0.037095f
C2334 8bit_ADDER_0.C mux8_0.NAND4F_3.Y 0.406267f
C2335 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT VDD 3.19832f
C2336 MULT_0.SO MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A 8.21e-19
C2337 mux8_6.A0 SEL0 0.633835f
C2338 mux8_1.NAND4F_9.Y NOT8_0.S0 3.17e-20
C2339 AND8_0.S3 NOT8_0.S3 9.87e-19
C2340 OR8_0.NOT8_0.A6 A4 0.025544f
C2341 XOR8_0.S3 SEL1 0.094489f
C2342 mux8_6.NAND4F_2.D mux8_6.NAND4F_1.Y 2.96e-20
C2343 NOT8_0.S0 B0 0.461519f
C2344 mux8_8.NAND4F_0.C SEL2 1.4681f
C2345 mux8_3.NAND4F_5.Y SEL1 0.306449f
C2346 XOR8_0.S3 AND8_0.S6 0.154477f
C2347 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT mux8_5.A0 9.63e-20
C2348 OR8_0.NOT8_0.A5 A5 0.255811f
C2349 B7 A6 23.1575f
C2350 mux8_3.NAND4F_2.Y mux8_3.NAND4F_5.Y 4.33e-19
C2351 A3 A2 4.69018f
C2352 AND8_0.S1 A0 0.043694f
C2353 mux8_6.A0 mux8_8.NAND4F_4.B 7.13e-21
C2354 8bit_ADDER_0.S0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 0.002364f
C2355 mux8_7.A0 NOT8_0.S1 0.016346f
C2356 mux8_5.A0 OR8_0.S2 0.021801f
C2357 mux8_7.NAND4F_2.Y VDD 2.1749f
C2358 mux8_5.NAND4F_2.D mux8_5.NAND4F_3.Y 0.397922f
C2359 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 0.012122f
C2360 mux8_6.A1 AND8_0.S4 3.14041f
C2361 mux8_5.NAND4F_2.D XOR8_0.S4 4.4e-19
C2362 8bit_ADDER_0.S0 mux8_1.NAND4F_0.C 0.081597f
C2363 mux8_0.NAND4F_8.Y SEL0 4.08e-19
C2364 B5 B3 0.020297f
C2365 left_shifter_0.S7 OR8_0.S7 0.031747f
C2366 MULT_0.S2 VDD 0.940197f
C2367 AND8_0.S0 AND8_0.NOT8_0.A1 1.13e-20
C2368 mux8_5.NAND4F_4.Y mux8_5.NAND4F_8.Y 0.404949f
C2369 mux8_4.A1 mux8_4.NAND4F_5.Y 1.57e-19
C2370 mux8_7.A0 SEL2 1.48878f
C2371 AND8_0.S1 NOT8_0.S1 5.33e-19
C2372 mux8_4.A1 XOR8_0.S3 3.04e-20
C2373 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT A6 0.010334f
C2374 MULT_0.4bit_ADDER_0.B2 A2 0.442058f
C2375 MULT_0.SO SEL2 0.076839f
C2376 XOR8_0.S2 B7 5.3e-19
C2377 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT MULT_0.inv_9.Y 0.004135f
C2378 AND8_0.S2 B4 1.28e-21
C2379 mux8_7.NAND4F_0.Y mux8_7.NAND4F_3.Y 0.616159f
C2380 MULT_0.4bit_ADDER_1.A2 VDD 3.3429f
C2381 mux8_7.A0 mux8_7.NAND4F_1.Y 5.23e-19
C2382 mux8_6.A0 MULT_0.S2 0.024985f
C2383 mux8_0.NAND4F_0.C mux8_0.NAND4F_5.Y 0.050993f
C2384 NOT8_0.S1 mux8_2.NAND4F_1.Y 0.55011f
C2385 mux8_7.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 0.02137f
C2386 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT A2 0.129026f
C2387 8bit_ADDER_0.S2 VDD 1.28098f
C2388 mux8_4.A1 mux8_4.NAND4F_3.Y 0.541275f
C2389 AND8_0.S4 AND8_0.S5 0.160471f
C2390 OR8_0.S7 mux8_6.NAND4F_5.Y 2.34e-19
C2391 mux8_5.A0 SEL1 0.356866f
C2392 AND8_0.S7 B7 0.044989f
C2393 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B A0 0.950228f
C2394 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 8bit_ADDER_0.C 0.002397f
C2395 mux8_4.NAND4F_8.Y SEL0 4.08e-19
C2396 XOR8_0.S2 SEL0 0.167406f
C2397 mux8_3.NAND4F_2.D mux8_3.NAND4F_7.Y 2.97e-20
C2398 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 8bit_ADDER_0.C 0.002397f
C2399 AND8_0.S1 MULT_0.inv_15.Y 5.74e-20
C2400 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 8bit_ADDER_0.C 0.002397f
C2401 AND8_0.S1 SEL2 0.076988f
C2402 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 8bit_ADDER_0.C 0.014679f
C2403 mux8_5.NAND4F_2.D mux8_5.NAND4F_7.Y 2.97e-20
C2404 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A 2.56e-19
C2405 OR8_0.NOT8_0.A3 OR8_0.NOT8_0.A4 0.098402f
C2406 mux8_0.NAND4F_3.Y mux8_0.NAND4F_1.Y 0.086984f
C2407 mux8_6.NAND4F_1.Y SEL1 2.35e-20
C2408 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y VDD 1.58631f
C2409 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 0.001075f
C2410 OR8_0.S1 OR8_0.NOT8_0.A2 1.27e-20
C2411 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A A0 0.685441f
C2412 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y VDD 1.58631f
C2413 mux8_1.NAND4F_0.C left_shifter_0.S0 0.037495f
C2414 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y VDD 1.58515f
C2415 OR8_0.NOT8_0.A3 A3 0.26083f
C2416 OR8_0.S1 B2 0.092075f
C2417 mux8_6.A0 8bit_ADDER_0.S2 0.031212f
C2418 AND8_0.S5 mux8_7.NAND4F_4.Y 0.402481f
C2419 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y VDD 1.57295f
C2420 mux8_2.NAND4F_0.C NOT8_0.S1 0.053425f
C2421 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 0.017305f
C2422 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A VDD 1.30818f
C2423 AND8_0.NOT8_0.A3 A4 1.27e-19
C2424 8bit_ADDER_0.C mux8_5.A0 0.102978f
C2425 mux8_2.NAND4F_1.Y SEL2 0.37854f
C2426 AND8_0.S7 SEL0 0.093941f
C2427 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A MULT_0.S2 2.27e-19
C2428 mux8_4.A0 SEL0 0.67918f
C2429 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT 0.012283f
C2430 VDD A4 2.75842f
C2431 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B 0.792412f
C2432 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A mux8_5.A0 2.04e-19
C2433 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B 2.43e-19
C2434 mux8_5.NAND4F_6.Y SEL2 0.419676f
C2435 V_FLAG_0.XOR2_0.Y A7 0.199941f
C2436 mux8_3.NAND4F_2.Y mux8_3.NAND4F_8.Y 0.222339f
C2437 mux8_8.A0 NOT8_0.S5 0.040367f
C2438 NOT8_0.S7 B7 0.477109f
C2439 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 3.6e-19
C2440 mux8_2.NAND4F_4.B VDD 1.19433f
C2441 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT mux8_8.A1 0.706883f
C2442 OR8_0.S7 A3 0.092942f
C2443 OR8_0.S2 mux8_7.A1 0.012559f
C2444 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A 3.6e-19
C2445 mux8_1.NAND4F_0.Y mux8_1.NAND4F_9.Y 2.96e-20
C2446 mux8_4.NAND4F_0.C SEL1 1.12237f
C2447 XOR8_0.S0 mux8_1.NAND4F_7.Y 9.74e-20
C2448 mux8_4.NAND4F_6.Y mux8_4.NAND4F_7.Y 0.14618f
C2449 mux8_5.A0 mux8_4.A1 0.057604f
C2450 mux8_2.NAND4F_0.C SEL2 1.4681f
C2451 NOT8_0.S4 left_shifter_0.S7 0.026056f
C2452 VDD A1 6.65557f
C2453 mux8_7.A0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 1.53e-19
C2454 mux8_4.NAND4F_4.B mux8_4.NAND4F_5.Y 0.248856f
C2455 MULT_0.inv_9.Y A2 0.372254f
C2456 mux8_8.NAND4F_2.D SEL1 3.38942f
C2457 AND8_0.S6 mux8_8.NAND4F_2.D 0.084271f
C2458 XOR8_0.S6 A5 0.031827f
C2459 NOT8_0.S7 SEL0 1.06748f
C2460 NOT8_0.S0 OR8_0.S2 0.017476f
C2461 XOR8_0.S1 mux8_2.NAND4F_6.Y 0.520706f
C2462 B5 B4 6.40189f
C2463 V_FLAG_0.XOR2_0.Y mux8_0.NAND4F_0.C 2.74e-20
C2464 mux8_4.NAND4F_4.B XOR8_0.S3 0.96337f
C2465 B6 B3 0.019887f
C2466 MULT_0.S2 XOR8_0.S2 3.04e-20
C2467 mux8_8.A0 VDD 1.30471f
C2468 AND8_0.S5 mux8_7.NAND4F_5.Y 5.23e-19
C2469 mux8_3.NAND4F_6.Y mux8_3.NAND4F_7.Y 0.14618f
C2470 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y A6 3.98e-19
C2471 mux8_5.A0 XOR8_0.S0 0.021342f
C2472 MULT_0.4bit_ADDER_2.B2 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT 0.001576f
C2473 MULT_0.4bit_ADDER_1.B3 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A 5.19e-20
C2474 mux8_1.NAND4F_0.C mux8_1.NAND4F_5.Y 0.051024f
C2475 mux8_4.NAND4F_4.B mux8_4.NAND4F_3.Y 0.223331f
C2476 mux8_5.NAND4F_4.Y mux8_5.NAND4F_9.Y 5.28e-19
C2477 A6 A4 0.026988f
C2478 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.B1 0.167796f
C2479 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A 0.186684f
C2480 mux8_4.A0 MULT_0.S2 0.027398f
C2481 AND8_0.S5 mux8_7.NAND4F_4.B 1.04124f
C2482 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A 5.19e-20
C2483 mux8_5.NAND4F_0.C mux8_5.NAND4F_9.Y 4.79e-21
C2484 XOR8_0.S7 B6 0.016229f
C2485 MULT_0.SO MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT 4.62e-19
C2486 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A A2 0.685441f
C2487 mux8_6.A0 mux8_8.A0 21.160301f
C2488 mux8_0.NAND4F_5.Y SEL1 0.306449f
C2489 8bit_ADDER_0.S2 XOR8_0.S2 0.009242f
C2490 mux8_4.A1 mux8_4.NAND4F_0.C 0.064499f
C2491 mux8_7.A1 SEL1 0.069436f
C2492 AND8_0.NOT8_0.A4 AND8_0.NOT8_0.A5 0.165325f
C2493 A6 A1 0.026095f
C2494 mux8_4.A0 8bit_ADDER_0.S2 5.86054f
C2495 8bit_ADDER_0.C mux8_0.NAND4F_5.Y 2.08e-19
C2496 mux8_8.NAND4F_2.Y XOR8_0.S6 1.49e-19
C2497 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B 0.008371f
C2498 mux8_7.A0 XOR8_0.S3 0.03518f
C2499 NOT8_0.S0 SEL1 0.074562f
C2500 mux8_7.NAND4F_6.Y SEL0 0.353718f
C2501 mux8_7.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A 0.00837f
C2502 mux8_2.NAND4F_2.D mux8_2.NAND4F_4.Y 0.349681f
C2503 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A mux8_7.A1 6.44e-19
C2504 mux8_6.NAND4F_0.C mux8_6.NAND4F_6.Y 0.142729f
C2505 AND8_0.S0 SEL0 0.128281f
C2506 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y mux8_4.A0 2.76e-19
C2507 mux8_6.NAND4F_0.C mux8_6.NAND4F_9.Y 4.79e-21
C2508 B0 A2 1.47839f
C2509 mux8_2.NAND4F_9.Y NOT8_0.S1 3.17e-20
C2510 mux8_5.A0 mux8_4.NAND4F_4.B 6.94e-21
C2511 OR8_0.NOT8_0.A2 A3 0.002952f
C2512 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 0.007216f
C2513 mux8_2.NAND4F_3.Y mux8_2.NAND4F_8.Y 0.222524f
C2514 B2 A3 2.13584f
C2515 VDD Y1 0.957559f
C2516 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 2.43e-19
C2517 AND8_0.S7 A4 0.130309f
C2518 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B 0.139263f
C2519 mux8_4.NAND4F_2.Y mux8_4.NAND4F_6.Y 0.08709f
C2520 mux8_7.A1 mux8_4.A1 8.29e-19
C2521 XOR8_0.S2 A1 0.024666f
C2522 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A 0.001913f
C2523 OR8_0.S1 mux8_6.A1 0.02887f
C2524 mux8_3.NAND4F_6.Y mux8_4.NAND4F_2.Y 0.002218f
C2525 mux8_5.NAND4F_4.B SEL1 4.36064f
C2526 V_FLAG_0.XOR2_0.Y SEL1 4.88e-20
C2527 mux8_7.NAND4F_2.Y mux8_7.NAND4F_6.Y 0.08709f
C2528 left_shifter_0.S7 XOR8_0.S4 0.036861f
C2529 B6 B4 0.021624f
C2530 mux8_2.NAND4F_9.Y SEL2 1.49e-20
C2531 mux8_8.A0 XOR8_0.S2 0.025513f
C2532 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y mux8_7.A0 1.53e-19
C2533 MULT_0.SO mux8_1.NAND4F_7.Y 5.24e-19
C2534 NOT8_0.S0 mux8_4.A1 0.018964f
C2535 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y mux8_7.A0 1.53e-19
C2536 MULT_0.4bit_ADDER_2.B2 MULT_0.inv_9.Y 0.070904f
C2537 AND8_0.NOT8_0.A7 A7 0.932478f
C2538 mux8_4.A0 A1 1.23e-19
C2539 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y mux8_7.A0 0.018349f
C2540 XOR8_0.S0 mux8_7.A1 0.06411f
C2541 Y4 Y6 0.017762f
C2542 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 0.119902f
C2543 mux8_4.NAND4F_2.D SEL0 0.229117f
C2544 mux8_8.NAND4F_0.C mux8_8.NAND4F_7.Y 0.224691f
C2545 AND8_0.NOT8_0.A3 AND8_0.NOT8_0.A6 1.07e-20
C2546 mux8_3.NAND4F_9.Y NOT8_0.S2 3.17e-20
C2547 mux8_2.NAND4F_2.D SEL1 3.39097f
C2548 AND8_0.NOT8_0.A6 VDD 2.31897f
C2549 mux8_4.NAND4F_0.C mux8_4.NAND4F_4.B 2.13077f
C2550 NOT8_0.S3 SEL0 1.10252f
C2551 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT VDD 3.18262f
C2552 mux8_7.A0 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 0.013109f
C2553 mux8_7.A0 mux8_5.A0 19.278698f
C2554 mux8_8.A0 mux8_4.A0 0.004466f
C2555 XOR8_0.S0 NOT8_0.S0 23.7059f
C2556 mux8_5.A0 MULT_0.SO 0.0201f
C2557 mux8_8.NAND4F_3.Y mux8_8.NAND4F_4.Y 0.102178f
C2558 mux8_8.NAND4F_0.Y mux8_8.NAND4F_8.Y 0.249057f
C2559 AND8_0.S0 MULT_0.S2 0.061873f
C2560 mux8_3.NAND4F_4.Y SEL2 8.74e-20
C2561 mux8_2.NAND4F_3.Y VDD 2.17641f
C2562 mux8_1.NAND4F_4.B mux8_1.NAND4F_2.Y 0.112019f
C2563 OR8_0.NOT8_0.A0 A1 0.033992f
C2564 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT mux8_5.A0 0.001145f
C2565 A7 A2 0.049852f
C2566 mux8_0.NAND4F_0.C mux8_0.NAND4F_2.Y 0.122872f
C2567 mux8_8.NAND4F_2.D mux8_8.NAND4F_0.C 1.55303f
C2568 mux8_6.A1 left_shifter_0.S7 0.092597f
C2569 mux8_3.NAND4F_4.B mux8_3.NAND4F_3.Y 0.223331f
C2570 mux8_5.NAND4F_4.Y mux8_5.NAND4F_1.Y 4.33e-19
C2571 mux8_0.NAND4F_5.Y mux8_0.NAND4F_1.Y 0.110562f
C2572 mux8_1.NAND4F_4.B VDD 1.25748f
C2573 mux8_3.NAND4F_0.C mux8_3.NAND4F_1.Y 0.402437f
C2574 V_FLAG_0.XOR2_2.Y A7 0.083561f
C2575 NOT8_0.S2 VDD 1.39906f
C2576 mux8_5.NAND4F_0.C mux8_5.NAND4F_1.Y 0.402437f
C2577 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 1.52e-19
C2578 B1 A5 0.02148f
C2579 mux8_6.NAND4F_2.D mux8_6.NAND4F_2.Y 0.339934f
C2580 MULT_0.inv_15.Y MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B 0.955489f
C2581 mux8_1.NAND4F_0.C SEL2 1.4681f
C2582 mux8_8.A1 OR8_0.S7 0.050427f
C2583 mux8_5.A0 AND8_0.S1 0.013922f
C2584 8bit_ADDER_0.S2 AND8_0.S0 0.013528f
C2585 mux8_3.NAND4F_0.Y mux8_3.NAND4F_9.Y 2.96e-20
C2586 left_shifter_0.S7 mux8_6.NAND4F_4.Y 5.23e-19
C2587 AND8_0.S4 OR8_0.NOT8_0.A6 0.001469f
C2588 MULT_0.4bit_ADDER_2.B2 mux8_8.A1 0.018513f
C2589 mux8_6.A0 NOT8_0.S2 0.017056f
C2590 mux8_7.NAND4F_2.D mux8_7.NAND4F_7.Y 2.97e-20
C2591 V_FLAG_0.XOR2_2.Y mux8_0.NAND4F_0.C 1.61e-20
C2592 AND8_0.NOT8_0.A6 A6 0.932826f
C2593 mux8_6.A1 mux8_6.NAND4F_5.Y 1.57e-19
C2594 OR8_0.NOT8_0.A5 OR8_0.NOT8_0.A7 0.001703f
C2595 mux8_0.NAND4F_0.C mux8_1.NAND4F_2.D 4.58e-19
C2596 mux8_1.NAND4F_7.Y mux8_2.NAND4F_0.C 9.03e-22
C2597 XOR8_0.S1 B2 2.98e-21
C2598 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_2.B1 0.200037f
C2599 VDD SEL3 11.1678f
C2600 mux8_8.NAND4F_3.Y SEL0 0.360934f
C2601 AND8_0.S5 left_shifter_0.S7 0.024011f
C2602 mux8_5.A0 mux8_5.NAND4F_6.Y 2.97e-22
C2603 XOR8_0.S4 A3 0.009017f
C2604 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT 0.127988f
C2605 mux8_8.NAND4F_8.Y VDD 3.38984f
C2606 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A 0.005938f
C2607 mux8_7.NAND4F_2.D mux8_7.NAND4F_8.Y 4.88e-20
C2608 OR8_0.S7 XOR8_0.S5 0.032453f
C2609 mux8_3.NAND4F_0.Y VDD 2.13518f
C2610 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT A2 0.010334f
C2611 mux8_7.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 0.005184f
C2612 NOT8_0.S6 B3 3.98e-20
C2613 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 0.139263f
C2614 MULT_0.inv_9.Y B2 7.23e-19
C2615 mux8_8.NAND4F_4.B mux8_8.NAND4F_3.Y 0.223331f
C2616 mux8_6.NAND4F_4.Y mux8_6.NAND4F_5.Y 0.087643f
C2617 mux8_5.A0 mux8_2.NAND4F_0.C 1.95e-19
C2618 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A MULT_0.S2 0.200075f
C2619 left_shifter_0.S0 AND8_0.S2 0.0268f
C2620 mux8_6.A0 SEL3 0.523993f
C2621 OR8_0.S2 A2 0.06804f
C2622 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B A0 0.00981f
C2623 B6 B5 4.64638f
C2624 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A 0.248956f
C2625 B3 A0 1.16482f
C2626 AND8_0.S0 A1 0.056154f
C2627 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A VDD 1.35672f
C2628 mux8_5.A0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 0.003184f
C2629 OR8_0.NOT8_0.A1 A1 0.307892f
C2630 mux8_5.NAND4F_4.Y SEL0 0.116703f
C2631 mux8_6.A1 A3 0.014943f
C2632 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A VDD 1.30818f
C2633 mux8_7.A0 mux8_7.A1 5.83179f
C2634 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 0.017305f
C2635 mux8_5.NAND4F_0.C SEL0 12.981099f
C2636 NOT8_0.S5 AND8_0.S4 0.017028f
C2637 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A mux8_5.A0 2.04e-19
C2638 left_shifter_0.S7 mux8_6.NAND4F_4.B 1.01693f
C2639 mux8_6.NAND4F_2.Y SEL1 0.222331f
C2640 mux8_1.NAND4F_4.Y SEL0 0.116386f
C2641 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT mux8_7.A1 0.018349f
C2642 mux8_4.A1 mux8_4.NAND4F_7.Y 5.24e-19
C2643 mux8_8.A0 AND8_0.S0 0.014485f
C2644 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A B2 0.001945f
C2645 mux8_4.NAND4F_4.B mux8_5.NAND4F_4.B 0.001581f
C2646 SEL3 A6 0.264979f
C2647 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B 0.792412f
C2648 mux8_0.NAND4F_2.Y SEL1 0.222331f
C2649 AND8_0.S6 AND8_0.NOT8_0.A7 1.56e-20
C2650 AND8_0.NOT8_0.A6 AND8_0.S7 0.339564f
C2651 mux8_2.NAND4F_4.Y mux8_2.NAND4F_6.Y 4.33e-19
C2652 mux8_1.NAND4F_1.Y SEL0 0.339784f
C2653 AND8_0.S4 mux8_5.NAND4F_2.Y 1.24e-19
C2654 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A 1.77e-19
C2655 XOR8_0.S2 NOT8_0.S2 11.484401f
C2656 mux8_7.A0 NOT8_0.S0 0.013529f
C2657 mux8_5.A1 mux8_5.NAND4F_8.Y 1.16e-22
C2658 mux8_8.NAND4F_4.Y mux8_8.NAND4F_1.Y 4.33e-19
C2659 MULT_0.SO NOT8_0.S0 0.009258f
C2660 mux8_8.A1 NOT8_0.S4 0.017073f
C2661 NOT8_0.S5 mux8_7.NAND4F_4.Y 2.18e-19
C2662 MULT_0.4bit_ADDER_1.B3 A2 0.001271f
C2663 mux8_8.A1 B2 5.17e-20
C2664 AND8_0.S1 mux8_7.A1 0.011083f
C2665 mux8_7.A0 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A 0.005588f
C2666 AND8_0.NOT8_0.A3 AND8_0.S4 0.339801f
C2667 8bit_ADDER_0.C mux8_0.NAND4F_2.Y 0.200461f
C2668 OR8_0.NOT8_0.A4 AND8_0.S5 0.004157f
C2669 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A 0.186684f
C2670 AND8_0.S4 VDD 1.52651f
C2671 AND8_0.S6 A2 0.003632f
C2672 mux8_4.A0 NOT8_0.S2 0.020205f
C2673 AND8_0.S5 A3 0.043157f
C2674 mux8_6.NAND4F_4.B mux8_6.NAND4F_5.Y 0.248856f
C2675 V_FLAG_0.XOR2_2.Y SEL1 0.003933f
C2676 mux8_3.NAND4F_4.Y mux8_3.NAND4F_5.Y 0.087643f
C2677 NOT8_0.S0 AND8_0.S1 0.845202f
C2678 mux8_6.NAND4F_6.Y SEL0 0.353704f
C2679 mux8_3.NAND4F_2.D mux8_3.NAND4F_4.B 1.27138f
C2680 mux8_7.NAND4F_0.Y SEL0 0.236427f
C2681 B2 B0 0.121796f
C2682 MULT_0.inv_15.Y B3 0.026111f
C2683 mux8_1.NAND4F_2.D SEL1 3.38955f
C2684 mux8_6.NAND4F_9.Y SEL0 2.8e-19
C2685 mux8_5.NAND4F_2.D mux8_5.NAND4F_2.Y 0.339934f
C2686 mux8_4.NAND4F_2.Y SEL1 0.222331f
C2687 mux8_7.NAND4F_4.Y VDD 2.2174f
C2688 OR8_0.S2 OR8_0.NOT8_0.A3 1.1e-20
C2689 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT A5 0.003441f
C2690 8bit_ADDER_0.C A2 0.03881f
C2691 mux8_6.A0 AND8_0.S4 0.018672f
C2692 OR8_0.S7 mux8_6.NAND4F_2.D 0.08162f
C2693 mux8_8.A0 NOT8_0.S3 0.014315f
C2694 mux8_2.NAND4F_6.Y SEL1 0.222305f
C2695 mux8_7.A0 mux8_5.NAND4F_4.B 6.92e-21
C2696 XOR8_0.S5 B2 0.003568f
C2697 mux8_2.NAND4F_6.Y mux8_3.NAND4F_2.Y 0.002062f
C2698 mux8_8.NAND4F_1.Y SEL0 0.339784f
C2699 mux8_5.NAND4F_5.Y SEL1 0.306449f
C2700 mux8_5.NAND4F_2.D VDD 1.37379f
C2701 NOT8_0.S6 B4 1.54e-19
C2702 mux8_4.A0 SEL3 1.23e-19
C2703 mux8_5.A1 AND8_0.S3 0.035792f
C2704 NOT8_0.S5 mux8_7.NAND4F_5.Y 0.288211f
C2705 XOR8_0.S7 SEL2 0.127804f
C2706 mux8_7.A0 mux8_2.NAND4F_2.D 1.75e-19
C2707 ZFLAG_0.nor4_1.Y Y5 0.013249f
C2708 mux8_7.NAND4F_2.D XOR8_0.S5 4.4e-19
C2709 ZFLAG_0.nor4_0.Y Y7 0.002702f
C2710 B4 A0 0.027224f
C2711 mux8_8.NAND4F_4.B mux8_8.NAND4F_1.Y 0.222551f
C2712 NOT8_0.S5 mux8_7.NAND4F_4.B 0.105153f
C2713 mux8_7.NAND4F_0.Y mux8_7.NAND4F_2.Y 0.170507f
C2714 NOT8_0.S0 mux8_2.NAND4F_0.C 2.74e-21
C2715 OR8_0.NOT8_0.A7 A5 0.029621f
C2716 mux8_0.NAND4F_0.C mux8_0.NAND4F_9.Y 4.79e-21
C2717 mux8_1.NAND4F_9.Y Y0 9.11e-19
C2718 mux8_4.A1 mux8_4.NAND4F_2.Y 1.16938f
C2719 mux8_7.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A 0.002364f
C2720 mux8_2.NAND4F_2.D AND8_0.S1 0.076916f
C2721 AND8_0.S2 A0 0.180193f
C2722 mux8_7.NAND4F_5.Y VDD 2.19984f
C2723 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A A0 0.00194f
C2724 A7 B2 0.042119f
C2725 mux8_4.NAND4F_9.Y mux8_4.NAND4F_6.Y 0.222562f
C2726 mux8_1.NAND4F_0.C mux8_1.NAND4F_7.Y 0.224691f
C2727 mux8_3.NAND4F_4.B mux8_3.NAND4F_6.Y 0.187883f
C2728 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_2.B1 0.697944f
C2729 mux8_2.NAND4F_9.Y mux8_3.NAND4F_8.Y 0.001328f
C2730 mux8_0.NAND4F_2.Y mux8_0.NAND4F_1.Y 3.31e-22
C2731 mux8_5.NAND4F_4.B mux8_5.NAND4F_6.Y 0.187883f
C2732 mux8_8.A0 mux8_8.NAND4F_3.Y 0.406267f
C2733 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 1.2618f
C2734 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B MULT_0.inv_15.Y 0.001496f
C2735 Y2 Y5 0.020883f
C2736 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A MULT_0.inv_9.Y 7.7e-20
C2737 Y0 Y7 0.020761f
C2738 Y3 Y4 0.020883f
C2739 Y1 Y6 0.020883f
C2740 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B 0.008371f
C2741 mux8_7.NAND4F_4.B VDD 1.19458f
C2742 mux8_2.NAND4F_2.D mux8_2.NAND4F_1.Y 2.96e-20
C2743 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 0.792412f
C2744 mux8_1.NAND4F_2.D XOR8_0.S0 4.4e-19
C2745 mux8_5.A0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 2.04e-19
C2746 mux8_0.NAND4F_4.B mux8_0.NAND4F_6.Y 0.187883f
C2747 mux8_8.A1 XOR8_0.S4 0.032842f
C2748 mux8_7.NAND4F_0.C SEL2 1.4681f
C2749 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A 0.001913f
C2750 XOR8_0.S2 AND8_0.S4 0.075659f
C2751 MULT_0.SO mux8_1.NAND4F_0.Y 0.43187f
C2752 mux8_5.A0 mux8_1.NAND4F_0.C 1.95e-19
C2753 OR8_0.S7 SEL1 0.049574f
C2754 mux8_7.NAND4F_0.C mux8_7.NAND4F_1.Y 0.402437f
C2755 AND8_0.S6 OR8_0.S7 0.016954f
C2756 mux8_0.NAND4F_6.Y mux8_0.NAND4F_7.Y 0.14618f
C2757 mux8_1.NAND4F_4.B AND8_0.S0 1.04047f
C2758 NOT8_0.S1 AND8_0.S2 2.04025f
C2759 AND8_0.S0 NOT8_0.S2 4.06e-20
C2760 mux8_3.NAND4F_4.Y mux8_3.NAND4F_8.Y 0.404949f
C2761 mux8_2.NAND4F_2.D mux8_2.NAND4F_0.C 1.55302f
C2762 mux8_1.NAND4F_1.Y mux8_2.NAND4F_4.B 1.02e-21
C2763 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B 0.139263f
C2764 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_1.A2 0.001492f
C2765 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A A5 0.008956f
C2766 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT VDD 3.5613f
C2767 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 1.58859f
C2768 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A 0.001568f
C2769 MULT_0.4bit_ADDER_0.A2 A2 0.00325f
C2770 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT VDD 3.18261f
C2771 XOR8_0.S4 XOR8_0.S5 0.10055f
C2772 mux8_7.A0 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 0.005184f
C2773 mux8_8.A1 mux8_6.A1 0.259054f
C2774 AND8_0.S3 B1 0.486525f
C2775 AND8_0.S2 SEL2 0.077523f
C2776 NOT8_0.S6 B5 0.61009f
C2777 AND8_0.NOT8_0.A0 B1 0.025364f
C2778 8bit_ADDER_0.S0 left_shifter_0.S0 8.02e-22
C2779 OR8_0.S2 OR8_0.NOT8_0.A2 0.399606f
C2780 AND8_0.NOT8_0.A2 A2 0.976024f
C2781 AND8_0.S1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT 1.75e-19
C2782 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A 2.56e-19
C2783 OR8_0.S2 B2 0.017919f
C2784 mux8_6.NAND4F_3.Y XOR8_0.S7 5.23e-19
C2785 B5 A0 0.024607f
C2786 mux8_4.NAND4F_4.B mux8_4.NAND4F_2.Y 0.112019f
C2787 mux8_6.A1 B0 0.037358f
C2788 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_1.B1 0.200037f
C2789 NOT8_0.S7 AND8_0.S4 0.022994f
C2790 XOR8_0.S3 B3 0.637585f
C2791 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT 0.127988f
C2792 OR8_0.S1 MULT_0.4bit_ADDER_2.B1 1.31e-19
C2793 NOT8_0.S2 NOT8_0.S3 0.041063f
C2794 mux8_6.A1 XOR8_0.S5 0.029956f
C2795 mux8_7.NAND4F_0.C mux8_7.NAND4F_9.Y 4.79e-21
C2796 mux8_8.A1 AND8_0.S5 0.016959f
C2797 AND8_0.NOT8_0.A5 B4 0.02593f
C2798 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A VDD 1.34493f
C2799 mux8_7.A0 A2 6.44e-20
C2800 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B 0.087175f
C2801 mux8_8.NAND4F_4.Y XOR8_0.S6 2.3e-19
C2802 MULT_0.4bit_ADDER_1.B3 B2 6.2e-19
C2803 NOT8_0.S4 SEL1 0.07293f
C2804 mux8_6.NAND4F_8.Y mux8_6.NAND4F_5.Y 0.001122f
C2805 mux8_1.NAND4F_6.Y mux8_2.NAND4F_8.Y 1.02e-21
C2806 mux8_8.A0 mux8_8.NAND4F_1.Y 5.23e-19
C2807 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 0.008371f
C2808 8bit_ADDER_0.S0 mux8_1.NAND4F_5.Y 2.08e-19
C2809 OR8_0.S1 VDD 1.22306f
C2810 mux8_7.A0 mux8_1.NAND4F_2.D 1.75e-19
C2811 AND8_0.S6 B2 0.005132f
C2812 mux8_1.NAND4F_2.D MULT_0.SO 0.107639f
C2813 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y B3 0.00144f
C2814 mux8_3.NAND4F_4.B OR8_0.S2 0.079695f
C2815 AND8_0.S5 XOR8_0.S5 1.69e-19
C2816 mux8_2.NAND4F_2.Y mux8_2.NAND4F_8.Y 0.222339f
C2817 NOT8_0.S5 left_shifter_0.S7 0.031305f
C2818 mux8_5.A1 mux8_5.NAND4F_1.Y 8.98e-23
C2819 AND8_0.S1 A2 0.171509f
C2820 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A 0.127125f
C2821 XOR8_0.S6 B7 0.092419f
C2822 mux8_1.NAND4F_0.C NOT8_0.S0 0.053145f
C2823 mux8_4.NAND4F_4.Y mux8_4.NAND4F_6.Y 4.33e-19
C2824 MULT_0.4bit_ADDER_1.B1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A 0.005938f
C2825 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A VDD 1.30818f
C2826 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 0.001078f
C2827 mux8_5.A0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 0.003184f
C2828 mux8_7.NAND4F_2.D SEL1 3.38953f
C2829 OR8_0.NOT8_0.A4 OR8_0.NOT8_0.A6 2.48e-20
C2830 mux8_6.A0 OR8_0.S1 0.024551f
C2831 8bit_ADDER_0.C B2 0.003774f
C2832 AND8_0.NOT8_0.A1 B1 0.180048f
C2833 OR8_0.NOT8_0.A1 AND8_0.S4 3.06e-22
C2834 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B 0.02452f
C2835 OR8_0.NOT8_0.A6 A3 0.006343f
C2836 mux8_7.NAND4F_4.Y mux8_7.NAND4F_6.Y 4.33e-19
C2837 MULT_0.4bit_ADDER_1.B2 A0 1.17e-19
C2838 mux8_6.A1 mux8_6.NAND4F_7.Y 5.24e-19
C2839 B7 A5 0.137003f
C2840 OR8_0.NOT8_0.A5 A4 0.203525f
C2841 NOT8_0.S6 B6 0.475307f
C2842 XOR8_0.S6 SEL0 0.168096f
C2843 mux8_1.NAND4F_2.Y mux8_1.NAND4F_6.Y 0.08709f
C2844 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT mux8_4.A0 0.152545f
C2845 mux8_2.NAND4F_0.Y mux8_2.NAND4F_5.Y 4.32e-19
C2846 left_shifter_0.S7 VDD 0.88095f
C2847 mux8_4.NAND4F_1.Y SEL0 0.339784f
C2848 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT MULT_0.inv_9.Y 4.16e-20
C2849 mux8_5.NAND4F_8.Y mux8_5.NAND4F_9.Y 0.696806f
C2850 mux8_1.NAND4F_6.Y VDD 2.1782f
C2851 B6 A0 0.024505f
C2852 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A 1.16e-19
C2853 mux8_8.NAND4F_4.B XOR8_0.S6 0.963395f
C2854 mux8_3.NAND4F_1.Y SEL0 0.339784f
C2855 XOR8_0.S3 B4 0.115748f
C2856 AND8_0.NOT8_0.A0 AND8_0.S3 1.03e-19
C2857 MULT_0.SO MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A 0.008733f
C2858 mux8_2.NAND4F_6.Y mux8_2.NAND4F_1.Y 2.45057f
C2859 mux8_2.NAND4F_5.Y mux8_2.NAND4F_7.Y 0.235079f
C2860 mux8_6.A1 mux8_6.NAND4F_2.D 0.107639f
C2861 left_shifter_0.S0 mux8_1.NAND4F_5.Y 0.402437f
C2862 XOR8_0.S7 mux8_6.NAND4F_1.Y 0.404949f
C2863 mux8_6.NAND4F_4.Y mux8_6.NAND4F_7.Y 4.32e-19
C2864 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A mux8_7.A1 2.28e-19
C2865 mux8_7.A0 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A 0.002364f
C2866 mux8_8.NAND4F_3.Y mux8_8.NAND4F_8.Y 0.222524f
C2867 mux8_3.NAND4F_4.B SEL1 4.36049f
C2868 mux8_8.NAND4F_2.Y mux8_8.NAND4F_4.Y 2.04463f
C2869 mux8_2.NAND4F_2.Y VDD 2.175f
C2870 mux8_1.NAND4F_4.B mux8_1.NAND4F_4.Y 0.275773f
C2871 mux8_0.NAND4F_9.Y mux8_0.NAND4F_1.Y 0.222572f
C2872 mux8_6.A0 left_shifter_0.S7 1.4e-20
C2873 mux8_0.NAND4F_0.C mux8_0.NAND4F_4.Y 0.049713f
C2874 mux8_1.NAND4F_1.Y mux8_2.NAND4F_3.Y 0.0024f
C2875 mux8_3.NAND4F_4.B mux8_3.NAND4F_2.Y 0.112019f
C2876 MULT_0.4bit_ADDER_2.B2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 0.139263f
C2877 mux8_1.NAND4F_0.C mux8_2.NAND4F_2.D 5.98e-19
C2878 mux8_1.NAND4F_4.B mux8_1.NAND4F_1.Y 0.222551f
C2879 mux8_5.NAND4F_5.Y mux8_5.NAND4F_6.Y 1.93433f
C2880 AND8_0.S2 mux8_3.NAND4F_5.Y 5.23e-19
C2881 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT A5 0.129004f
C2882 ZFLAG_0.nor4_0.Y Z 4.72e-19
C2883 AND8_0.NOT8_0.A5 B5 0.152578f
C2884 mux8_6.NAND4F_5.Y VDD 2.19904f
C2885 mux8_6.NAND4F_2.D mux8_6.NAND4F_4.Y 0.349681f
C2886 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B B0 0.021678f
C2887 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT 8.89e-19
C2888 OR8_0.S2 mux8_6.A1 0.139471f
C2889 mux8_2.NAND4F_0.C mux8_2.NAND4F_6.Y 0.142729f
C2890 mux8_7.NAND4F_5.Y mux8_7.NAND4F_6.Y 1.93433f
C2891 mux8_5.A1 SEL0 1.17085f
C2892 OR8_0.S1 XOR8_0.S2 1.14e-19
C2893 mux8_7.NAND4F_4.B mux8_7.NAND4F_6.Y 0.187883f
C2894 XOR8_0.S4 SEL1 0.106019f
C2895 mux8_7.NAND4F_9.Y Y5 5.66e-19
C2896 mux8_6.A0 mux8_6.NAND4F_5.Y 2.08e-19
C2897 AND8_0.S6 XOR8_0.S4 0.086618f
C2898 mux8_8.NAND4F_6.Y VDD 2.17811f
C2899 mux8_6.NAND4F_0.Y SEL2 2.97e-20
C2900 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT 0.119909f
C2901 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y B4 0.202041f
C2902 mux8_0.NAND4F_0.Y SEL2 2.97e-20
C2903 mux8_8.NAND4F_2.Y SEL0 0.296545f
C2904 MULT_0.S2 mux8_3.NAND4F_1.Y 8.98e-23
C2905 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.B1 0.697859f
C2906 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A 0.118063f
C2907 Y1 Y3 0.017734f
C2908 mux8_0.NAND4F_6.Y SEL0 0.353737f
C2909 OR8_0.NOT8_0.A4 VDD 0.988795f
C2910 mux8_4.A0 OR8_0.S1 0.02521f
C2911 mux8_3.NAND4F_3.Y VDD 2.17569f
C2912 AND8_0.NOT8_0.A3 A3 1.00515f
C2913 VDD A3 7.76967f
C2914 mux8_5.A0 B4 5.02e-19
C2915 mux8_5.NAND4F_1.Y mux8_7.NAND4F_3.Y 0.002218f
C2916 AND8_0.S1 MULT_0.4bit_ADDER_2.B2 1.77e-19
C2917 mux8_8.NAND4F_4.B mux8_8.NAND4F_2.Y 0.112019f
C2918 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 0.005938f
C2919 mux8_1.NAND4F_0.C mux8_1.NAND4F_0.Y 0.223896f
C2920 mux8_3.NAND4F_4.Y mux8_3.NAND4F_7.Y 4.32e-19
C2921 mux8_0.NAND4F_2.D mux8_0.NAND4F_0.Y 0.184536f
C2922 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B 1.2618f
C2923 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A B7 0.001945f
C2924 mux8_7.NAND4F_7.Y mux8_8.NAND4F_0.Y 0.002217f
C2925 8bit_ADDER_0.S0 SEL2 0.099336f
C2926 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B VDD 1.8478f
C2927 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A mux8_4.A0 0.200037f
C2928 mux8_6.A1 SEL1 0.025591f
C2929 mux8_6.A1 AND8_0.S6 0.026017f
C2930 AND8_0.S3 AND8_0.NOT8_0.A1 1.11e-19
C2931 OR8_0.S1 OR8_0.NOT8_0.A0 0.269009f
C2932 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B A7 0.950228f
C2933 8bit_ADDER_0.S2 mux8_3.NAND4F_1.Y 5.23e-19
C2934 AND8_0.NOT8_0.A2 B2 0.176303f
C2935 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT VDD 3.30026f
C2936 mux8_5.A0 AND8_0.S2 0.013922f
C2937 mux8_2.NAND4F_5.Y SEL0 0.121352f
C2938 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B 0.209959f
C2939 AND8_0.NOT8_0.A0 AND8_0.NOT8_0.A1 0.854726f
C2940 mux8_6.NAND4F_2.D mux8_6.NAND4F_4.B 1.27138f
C2941 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 2.43e-19
C2942 mux8_5.A0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 2.04e-19
C2943 mux8_4.NAND4F_0.Y SEL2 2.97e-20
C2944 XOR8_0.S3 B5 0.103013f
C2945 mux8_8.NAND4F_9.Y mux8_6.NAND4F_8.Y 0.001427f
C2946 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A 0.001913f
C2947 XOR8_0.S6 A4 2.38e-19
C2948 mux8_7.NAND4F_0.C mux8_8.NAND4F_2.D 4.62e-19
C2949 NOT8_0.S5 mux8_7.NAND4F_7.Y 0.431664f
C2950 mux8_6.NAND4F_4.Y SEL1 0.30433f
C2951 mux8_1.NAND4F_8.Y SEL0 4.08e-19
C2952 left_shifter_0.S7 AND8_0.S7 0.039174f
C2953 B7 B1 0.07542f
C2954 left_shifter_0.S0 NOT8_0.S1 0.021223f
C2955 MULT_0.4bit_ADDER_0.B2 VDD 3.43894f
C2956 mux8_0.NAND4F_4.Y SEL1 0.30433f
C2957 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y A5 2.72689f
C2958 AND8_0.S4 mux8_5.NAND4F_4.Y 0.402481f
C2959 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A A5 0.685441f
C2960 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A 0.001571f
C2961 mux8_1.NAND4F_3.Y XOR8_0.S0 5.23e-19
C2962 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A 0.186684f
C2963 mux8_7.A0 NOT8_0.S4 0.015109f
C2964 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B 0.008371f
C2965 A6 A3 0.028017f
C2966 A5 A4 0.059017f
C2967 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_1.A2 0.009698f
C2968 mux8_5.NAND4F_0.C AND8_0.S4 0.037277f
C2969 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT VDD 3.18247f
C2970 AND8_0.S5 SEL1 0.12468f
C2971 mux8_8.NAND4F_0.Y mux8_8.NAND4F_9.Y 2.96e-20
C2972 mux8_3.NAND4F_0.C SEL0 12.9904f
C2973 AND8_0.S5 AND8_0.S6 6.54236f
C2974 8bit_ADDER_0.C mux8_0.NAND4F_4.Y 0.047022f
C2975 mux8_7.NAND4F_7.Y VDD 2.14052f
C2976 mux8_3.NAND4F_4.B mux8_4.NAND4F_4.B 0.001581f
C2977 left_shifter_0.S0 SEL2 0.154834f
C2978 mux8_2.NAND4F_9.Y mux8_2.NAND4F_6.Y 0.222562f
C2979 NOT8_0.S7 left_shifter_0.S7 8.37271f
C2980 AND8_0.S7 mux8_6.NAND4F_5.Y 5.23e-19
C2981 mux8_8.A0 XOR8_0.S6 0.009235f
C2982 MULT_0.4bit_ADDER_2.B1 MULT_0.inv_9.Y 2.33128f
C2983 mux8_7.A1 mux8_7.NAND4F_0.C 0.064711f
C2984 A5 A1 0.024888f
C2985 mux8_7.A0 mux8_7.NAND4F_2.D 0.104891f
C2986 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A 2.06e-19
C2987 mux8_7.NAND4F_3.Y SEL0 0.360934f
C2988 mux8_7.NAND4F_8.Y VDD 3.39014f
C2989 mux8_4.NAND4F_4.Y SEL1 0.30433f
C2990 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A 0.001568f
C2991 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y B5 0.001436f
C2992 mux8_5.NAND4F_2.D mux8_5.NAND4F_4.Y 0.349681f
C2993 mux8_6.NAND4F_0.Y mux8_6.NAND4F_3.Y 0.616159f
C2994 mux8_0.NAND4F_1.Y mux8_1.NAND4F_3.Y 0.002218f
C2995 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT 1.69e-20
C2996 AND8_0.S1 B2 0.043732f
C2997 mux8_5.NAND4F_2.D mux8_5.NAND4F_0.C 1.55303f
C2998 mux8_3.NAND4F_3.Y XOR8_0.S2 5.23e-19
C2999 XOR8_0.S1 VDD 1.00237f
C3000 mux8_8.A0 A5 0.445204f
C3001 mux8_0.NAND4F_0.Y mux8_0.NAND4F_3.Y 0.616159f
C3002 AND8_0.S0 OR8_0.S1 3.99e-19
C3003 OR8_0.S1 OR8_0.NOT8_0.A1 0.399126f
C3004 AND8_0.S2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A 1.54e-19
C3005 mux8_6.NAND4F_4.B SEL1 4.36059f
C3006 NOT8_0.S6 mux8_8.NAND4F_5.Y 0.288211f
C3007 NOT8_0.S4 mux8_5.NAND4F_6.Y 0.79864f
C3008 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B 0.087175f
C3009 NOT8_0.S7 mux8_6.NAND4F_5.Y 0.288211f
C3010 mux8_1.NAND4F_2.D mux8_1.NAND4F_0.C 1.55302f
C3011 MULT_0.inv_9.Y VDD 3.03477f
C3012 mux8_8.A1 mux8_8.NAND4F_0.Y 0.43187f
C3013 mux8_8.NAND4F_9.Y VDD 2.28324f
C3014 mux8_6.A0 XOR8_0.S1 0.025261f
C3015 AND8_0.S2 mux8_7.A1 0.011199f
C3016 AND8_0.S7 A3 0.091313f
C3017 MULT_0.S2 mux8_3.NAND4F_0.C 0.063475f
C3018 mux8_7.NAND4F_3.Y mux8_7.NAND4F_2.Y 1.63543f
C3019 mux8_7.NAND4F_0.Y mux8_7.NAND4F_4.Y 0.28646f
C3020 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B A1 0.016771f
C3021 mux8_5.NAND4F_8.Y SEL0 4.08e-19
C3022 mux8_8.A0 mux8_5.A1 0.027484f
C3023 mux8_1.NAND4F_5.Y SEL2 0.323263f
C3024 XOR8_0.S3 B6 0.092822f
C3025 mux8_3.NAND4F_2.D VDD 1.37487f
C3026 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A mux8_7.A1 3.63e-19
C3027 MULT_0.4bit_ADDER_2.B1 mux8_8.A1 2.52e-19
C3028 mux8_4.A1 mux8_4.NAND4F_4.Y 0.157118f
C3029 MULT_0.4bit_ADDER_2.B2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B 0.001328f
C3030 NOT8_0.S0 AND8_0.S2 0.01861f
C3031 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 0.139263f
C3032 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A 0.127125f
C3033 mux8_1.NAND4F_9.Y mux8_2.NAND4F_8.Y 0.001543f
C3034 mux8_5.NAND4F_0.C mux8_7.NAND4F_4.B 0.002598f
C3035 mux8_8.A1 NOT8_0.S5 0.021181f
C3036 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A VDD 1.67061f
C3037 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A 0.248956f
C3038 mux8_0.NAND4F_4.Y mux8_0.NAND4F_1.Y 4.33e-19
C3039 mux8_8.A0 mux8_8.NAND4F_2.Y 0.200461f
C3040 8bit_ADDER_0.S2 mux8_3.NAND4F_0.C 0.082259f
C3041 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A VDD 1.30818f
C3042 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A 1.01138f
C3043 mux8_5.NAND4F_9.Y mux8_5.NAND4F_1.Y 0.222572f
C3044 MULT_0.SO MULT_0.4bit_ADDER_1.B0 1.73e-22
C3045 mux8_6.A0 mux8_3.NAND4F_2.D 9.02e-20
C3046 mux8_2.NAND4F_4.B mux8_2.NAND4F_5.Y 0.248856f
C3047 mux8_5.A0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 0.003184f
C3048 mux8_4.NAND4F_0.Y mux8_4.NAND4F_5.Y 4.32e-19
C3049 mux8_7.A0 XOR8_0.S4 0.031573f
C3050 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B 1.28945f
C3051 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y B1 0.202698f
C3052 MULT_0.SO mux8_1.NAND4F_3.Y 0.541275f
C3053 mux8_3.NAND4F_9.Y mux8_3.NAND4F_6.Y 0.222562f
C3054 mux8_4.NAND4F_6.Y mux8_5.NAND4F_2.Y 0.002218f
C3055 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y B1 6.57e-19
C3056 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B mux8_6.A1 0.007216f
C3057 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y B1 6.57e-19
C3058 mux8_8.A1 VDD 1.21295f
C3059 NOT8_0.S5 XOR8_0.S5 10.3278f
C3060 mux8_7.NAND4F_0.Y mux8_7.NAND4F_5.Y 4.32e-19
C3061 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT mux8_4.A0 0.700777f
C3062 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y B1 0.004464f
C3063 AND8_0.S3 SEL0 0.128583f
C3064 B1 A4 0.021666f
C3065 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A 1.16e-19
C3066 mux8_4.NAND4F_0.Y mux8_4.NAND4F_3.Y 0.616159f
C3067 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A 0.005938f
C3068 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_1.A2 7.1e-19
C3069 mux8_1.NAND4F_2.Y mux8_1.NAND4F_9.Y 2.96e-20
C3070 mux8_8.NAND4F_5.Y SEL2 0.323263f
C3071 NOT8_0.S6 SEL2 0.099477f
C3072 mux8_4.NAND4F_6.Y VDD 2.17811f
C3073 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y B6 0.202041f
C3074 mux8_6.NAND4F_8.Y mux8_6.NAND4F_7.Y 9.84e-20
C3075 XOR8_0.S1 XOR8_0.S2 0.160302f
C3076 mux8_1.NAND4F_9.Y VDD 2.28375f
C3077 VDD B0 23.3322f
C3078 mux8_2.NAND4F_0.C mux8_3.NAND4F_4.B 0.002116f
C3079 mux8_6.A0 mux8_8.A1 0.061632f
C3080 mux8_3.NAND4F_6.Y VDD 2.17811f
C3081 mux8_6.NAND4F_0.Y mux8_6.NAND4F_1.Y 5.28e-20
C3082 XOR8_0.S5 VDD 1.07195f
C3083 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B VDD 1.98127f
C3084 AND8_0.S4 OR8_0.NOT8_0.A5 0.00377f
C3085 AND8_0.NOT8_0.A6 A5 0.163408f
C3086 MULT_0.4bit_ADDER_2.B2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B 0.008371f
C3087 OR8_0.NOT8_0.A7 B7 0.032763f
C3088 B1 A1 46.231396f
C3089 mux8_0.NAND4F_4.B SEL0 1.61041f
C3090 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT A5 0.010334f
C3091 mux8_6.NAND4F_2.Y XOR8_0.S7 1.49e-19
C3092 VDD Y7 1.30105f
C3093 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT 8.9e-19
C3094 mux8_6.NAND4F_2.D mux8_6.NAND4F_8.Y 4.88e-20
C3095 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A 8.34e-19
C3096 mux8_4.A0 XOR8_0.S1 0.026197f
C3097 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 0.132279f
C3098 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A 1.16e-19
C3099 B3 A2 30.294699f
C3100 mux8_6.A0 B0 0.006923f
C3101 mux8_4.NAND4F_4.B mux8_4.NAND4F_4.Y 0.275773f
C3102 mux8_5.A0 8bit_ADDER_0.S0 0.054131f
C3103 mux8_0.NAND4F_7.Y SEL0 0.234594f
C3104 XOR8_0.S4 mux8_5.NAND4F_6.Y 0.520706f
C3105 OR8_0.NOT8_0.A1 OR8_0.NOT8_0.A4 7.07e-22
C3106 mux8_8.NAND4F_7.Y mux8_6.NAND4F_0.Y 0.002217f
C3107 OR8_0.NOT8_0.A1 A3 3.27e-22
C3108 mux8_6.A0 XOR8_0.S5 0.028419f
C3109 NOT8_0.S2 mux8_3.NAND4F_1.Y 0.55011f
C3110 mux8_3.NAND4F_2.D XOR8_0.S2 4.4e-19
C3111 AND8_0.S1 mux8_6.A1 0.027533f
C3112 mux8_6.NAND4F_0.C SEL0 10.590401f
C3113 mux8_5.NAND4F_9.Y SEL0 2.8e-19
C3114 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 0.139263f
C3115 NOT8_0.S1 SEL2 0.108557f
C3116 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT 1.58859f
C3117 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B 0.00323f
C3118 mux8_2.NAND4F_0.Y mux8_2.NAND4F_7.Y 0.08762f
C3119 mux8_5.NAND4F_9.Y Y4 9.13e-19
C3120 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A 0.118063f
C3121 mux8_8.NAND4F_0.C mux8_6.NAND4F_4.B 0.002598f
C3122 mux8_7.A0 AND8_0.S5 0.128516f
C3123 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT 0.094647f
C3124 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A VDD 1.35001f
C3125 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT 8.89e-19
C3126 B0 A6 0.034249f
C3127 mux8_4.A0 mux8_3.NAND4F_2.D 3.06e-19
C3128 VDD A7 2.61467f
C3129 AND8_0.S2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT 1.53e-19
C3130 mux8_5.A1 NOT8_0.S2 0.108577f
C3131 SEL3 A5 0.264725f
C3132 mux8_8.A1 XOR8_0.S2 0.020459f
C3133 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A mux8_4.A0 5.13e-19
C3134 mux8_3.NAND4F_0.Y mux8_3.NAND4F_1.Y 5.28e-20
C3135 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B 0.209959f
C3136 mux8_5.NAND4F_6.Y mux8_5.NAND4F_7.Y 0.14618f
C3137 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B VDD 1.85269f
C3138 mux8_7.NAND4F_1.Y SEL2 0.37854f
C3139 mux8_6.A0 A7 1.13856f
C3140 mux8_6.NAND4F_7.Y VDD 2.13996f
C3141 mux8_5.A0 left_shifter_0.S0 0.015108f
C3142 mux8_2.NAND4F_4.Y mux8_2.NAND4F_8.Y 0.404949f
C3143 mux8_0.NAND4F_0.C VDD 1.40563f
C3144 mux8_7.NAND4F_6.Y mux8_7.NAND4F_7.Y 0.14618f
C3145 mux8_4.NAND4F_8.Y mux8_4.NAND4F_6.Y 2.96e-20
C3146 mux8_0.NAND4F_0.Y mux8_0.NAND4F_5.Y 4.32e-19
C3147 mux8_4.NAND4F_0.C mux8_4.NAND4F_0.Y 0.223896f
C3148 AND8_0.S6 OR8_0.NOT8_0.A6 0.018856f
C3149 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 0.792412f
C3150 mux8_5.A0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A 2.04e-19
C3151 mux8_0.NAND4F_2.D SEL2 0.473378f
C3152 mux8_8.A1 AND8_0.S7 0.041279f
C3153 XOR8_0.S2 B0 0.225356f
C3154 OR8_0.NOT8_0.A3 B3 0.077815f
C3155 XOR8_0.S2 mux8_3.NAND4F_6.Y 0.520706f
C3156 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A 0.129047f
C3157 AND8_0.S3 A4 4.36e-21
C3158 mux8_6.NAND4F_2.D VDD 1.37926f
C3159 mux8_7.NAND4F_8.Y mux8_7.NAND4F_6.Y 2.96e-20
C3160 mux8_6.A0 mux8_0.NAND4F_0.C 4.16e-19
C3161 AND8_0.NOT8_0.A4 AND8_0.S5 0.463698f
C3162 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 0.012283f
C3163 mux8_4.A0 mux8_4.NAND4F_6.Y 2.97e-22
C3164 A7 A6 0.424409f
C3165 mux8_1.NAND4F_4.Y mux8_1.NAND4F_6.Y 4.33e-19
C3166 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT 0.00162f
C3167 mux8_2.NAND4F_3.Y mux8_2.NAND4F_5.Y 4.33e-19
C3168 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 1.58859f
C3169 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT VDD 3.18262f
C3170 mux8_8.A1 OR8_0.NOT8_0.A0 0.054715f
C3171 mux8_1.NAND4F_6.Y mux8_1.NAND4F_1.Y 2.45057f
C3172 mux8_1.NAND4F_5.Y mux8_1.NAND4F_7.Y 0.235079f
C3173 B4 A2 0.023198f
C3174 OR8_0.S7 B3 0.122066f
C3175 mux8_6.A0 mux8_6.NAND4F_2.D 0.105154f
C3176 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT 1.58859f
C3177 AND8_0.S7 XOR8_0.S5 0.03359f
C3178 OR8_0.S2 VDD 1.40834f
C3179 AND8_0.S3 A1 0.084364f
C3180 XOR8_0.S3 NOT8_0.S6 0.220929f
C3181 mux8_8.NAND4F_2.Y mux8_8.NAND4F_8.Y 0.222339f
C3182 mux8_2.NAND4F_0.Y SEL0 0.236428f
C3183 mux8_2.NAND4F_4.Y VDD 2.21756f
C3184 AND8_0.NOT8_0.A0 A1 0.028106f
C3185 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_1.A2 0.022379f
C3186 OR8_0.NOT8_0.A0 B0 0.059885f
C3187 8bit_ADDER_0.S0 NOT8_0.S0 1.11e-19
C3188 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A VDD 1.69318f
C3189 mux8_3.NAND4F_4.B mux8_3.NAND4F_4.Y 0.275773f
C3190 AND8_0.S2 A2 0.049803f
C3191 MULT_0.4bit_ADDER_2.B2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A 0.005938f
C3192 mux8_8.A0 AND8_0.S3 0.018509f
C3193 AND8_0.S0 MULT_0.inv_9.Y 0.013822f
C3194 mux8_2.NAND4F_7.Y SEL0 0.234594f
C3195 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT 1.69e-20
C3196 OR8_0.S7 XOR8_0.S7 0.278732f
C3197 mux8_6.A0 OR8_0.S2 0.024551f
C3198 mux8_7.NAND4F_9.Y SEL2 1.49e-20
C3199 left_shifter_0.S7 mux8_6.NAND4F_6.Y 1.2e-19
C3200 NOT8_0.S5 SEL1 0.074201f
C3201 OR8_0.NOT8_0.A7 A4 0.059207f
C3202 mux8_5.NAND4F_1.Y SEL0 0.339784f
C3203 mux8_7.NAND4F_9.Y mux8_7.NAND4F_1.Y 0.222572f
C3204 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT mux8_8.A0 0.152506f
C3205 mux8_3.NAND4F_2.Y mux8_3.NAND4F_9.Y 2.96e-20
C3206 mux8_3.NAND4F_0.C NOT8_0.S2 0.053329f
C3207 NOT8_0.S7 XOR8_0.S5 0.029405f
C3208 NOT8_0.S2 B1 0.492218f
C3209 mux8_5.NAND4F_2.Y SEL1 0.222331f
C3210 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A SEL3 6.08e-19
C3211 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A 2.59e-19
C3212 MULT_0.4bit_ADDER_1.B3 VDD 3.54648f
C3213 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A 0.248556f
C3214 mux8_6.NAND4F_3.Y SEL2 2.96e-20
C3215 mux8_1.NAND4F_2.Y SEL1 0.222331f
C3216 mux8_0.NAND4F_3.Y SEL2 2.96e-20
C3217 left_shifter_0.S0 mux8_7.A1 0.019566f
C3218 mux8_8.NAND4F_9.Y Y6 6.01e-19
C3219 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT 1.69e-20
C3220 VDD SEL1 8.470441f
C3221 mux8_5.A1 AND8_0.S4 5.71322f
C3222 mux8_8.NAND4F_4.Y SEL0 0.117162f
C3223 AND8_0.S6 VDD 1.11727f
C3224 mux8_6.NAND4F_5.Y mux8_6.NAND4F_6.Y 1.93433f
C3225 mux8_6.NAND4F_9.Y mux8_6.NAND4F_5.Y 0.402985f
C3226 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y A0 2.7267f
C3227 mux8_3.NAND4F_2.Y VDD 2.17486f
C3228 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y A0 0.00101f
C3229 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y A0 0.00101f
C3230 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y A0 0.00101f
C3231 left_shifter_0.S0 NOT8_0.S0 18.388302f
C3232 AND8_0.NOT8_0.A7 B5 0.051933f
C3233 mux8_4.NAND4F_5.Y SEL2 0.323263f
C3234 mux8_8.NAND4F_4.B mux8_8.NAND4F_4.Y 0.275773f
C3235 SEL3 B1 1.23276f
C3236 AND8_0.S0 mux8_8.A1 0.519575f
C3237 mux8_1.NAND4F_0.C mux8_1.NAND4F_3.Y 0.399921f
C3238 MULT_0.4bit_ADDER_2.B2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B 0.005184f
C3239 mux8_0.NAND4F_2.D mux8_0.NAND4F_3.Y 0.397922f
C3240 mux8_6.A0 SEL1 0.290639f
C3241 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 0.008381f
C3242 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A 2.56e-19
C3243 8bit_ADDER_0.C VDD 2.59355f
C3244 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A 1.01138f
C3245 mux8_3.NAND4F_0.C mux8_3.NAND4F_0.Y 0.223896f
C3246 XOR8_0.S3 SEL2 0.211062f
C3247 mux8_6.A0 AND8_0.S6 0.31448f
C3248 mux8_3.NAND4F_5.Y SEL2 0.323263f
C3249 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A VDD 1.67098f
C3250 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT VDD 3.56186f
C3251 mux8_5.A0 A0 9.63e-20
C3252 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A VDD 1.30818f
C3253 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A VDD 1.34441f
C3254 NOT8_0.S4 B3 0.484306f
C3255 OR8_0.NOT8_0.A2 B3 0.011308f
C3256 AND8_0.NOT8_0.A1 A1 0.975547f
C3257 mux8_5.A1 mux8_5.NAND4F_2.D 0.107639f
C3258 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 0.001075f
C3259 AND8_0.S7 mux8_6.NAND4F_2.D 0.076916f
C3260 B5 A2 0.021258f
C3261 AND8_0.S0 B0 0.050348f
C3262 mux8_4.NAND4F_3.Y SEL2 2.96e-20
C3263 OR8_0.NOT8_0.A1 B0 0.006833f
C3264 mux8_5.A0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 0.015199f
C3265 B3 B2 3.08006f
C3266 XOR8_0.S5 mux8_7.NAND4F_6.Y 0.520706f
C3267 OR8_0.S7 B4 0.23402f
C3268 OR8_0.S2 XOR8_0.S2 9.08794f
C3269 mux8_6.A0 8bit_ADDER_0.C 0.416721f
C3270 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B 0.001328f
C3271 mux8_8.NAND4F_5.Y mux8_8.NAND4F_7.Y 0.235079f
C3272 mux8_8.NAND4F_6.Y mux8_8.NAND4F_1.Y 2.45057f
C3273 NOT8_0.S6 mux8_8.NAND4F_7.Y 0.431664f
C3274 mux8_4.A1 VDD 0.947472f
C3275 NOT8_0.S7 mux8_6.NAND4F_7.Y 0.431664f
C3276 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT mux8_4.A0 0.010519f
C3277 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B mux8_6.A1 1.26434f
C3278 mux8_1.NAND4F_2.Y XOR8_0.S0 1.49e-19
C3279 mux8_5.A0 NOT8_0.S1 0.014305f
C3280 mux8_4.A0 OR8_0.S2 0.026964f
C3281 VDD Z 0.892677f
C3282 mux8_8.NAND4F_4.B SEL0 1.6099f
C3283 XOR8_0.S0 VDD 0.869808f
C3284 mux8_8.NAND4F_2.D mux8_8.NAND4F_5.Y 9.34e-20
C3285 mux8_6.A0 mux8_4.A1 0.046296f
C3286 AND8_0.S3 AND8_0.NOT8_0.A6 9.03e-21
C3287 mux8_8.A1 NOT8_0.S3 0.018739f
C3288 MULT_0.4bit_ADDER_2.B2 AND8_0.S2 1.54e-19
C3289 NOT8_0.S6 mux8_8.NAND4F_2.D 4.43e-19
C3290 mux8_1.NAND4F_7.Y SEL2 0.176544f
C3291 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A mux8_8.A0 0.200037f
C3292 8bit_ADDER_0.C A6 0.038798f
C3293 NOT8_0.S7 mux8_6.NAND4F_2.D 4.43e-19
C3294 NOT8_0.S0 mux8_1.NAND4F_5.Y 0.288211f
C3295 mux8_4.NAND4F_2.D mux8_4.NAND4F_6.Y 2.96e-20
C3296 V_FLAG_0.XOR2_2.B V_FLAG_0.XOR2_0.Y 1.03e-20
C3297 mux8_8.NAND4F_0.C mux8_8.NAND4F_0.Y 0.223896f
C3298 OR8_0.S2 OR8_0.NOT8_0.A0 1.26e-19
C3299 NOT8_0.S3 mux8_4.NAND4F_6.Y 0.79864f
C3300 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B VDD 1.976f
C3301 mux8_6.A0 XOR8_0.S0 0.023832f
C3302 VDD S 0.885561f
C3303 mux8_7.NAND4F_2.Y SEL0 0.296545f
C3304 Y6 Y7 4.56471f
C3305 mux8_5.A0 SEL2 0.979616f
C3306 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B A2 0.950228f
C3307 AND8_0.S4 B1 0.002254f
C3308 NOT8_0.S2 AND8_0.S3 0.127907f
C3309 XOR8_0.S2 SEL1 0.093809f
C3310 mux8_6.NAND4F_0.Y mux8_6.NAND4F_2.Y 0.170507f
C3311 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_1.B1 9.98e-20
C3312 mux8_4.NAND4F_0.Y mux8_4.NAND4F_7.Y 0.08762f
C3313 mux8_6.NAND4F_1.Y SEL2 0.37854f
C3314 mux8_3.NAND4F_2.Y XOR8_0.S2 1.49e-19
C3315 mux8_0.NAND4F_1.Y VDD 2.1816f
C3316 mux8_3.NAND4F_7.Y mux8_4.NAND4F_0.Y 0.002217f
C3317 mux8_0.NAND4F_0.Y mux8_0.NAND4F_2.Y 0.170507f
C3318 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B 0.139263f
C3319 MULT_0.S2 SEL0 1.17083f
C3320 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.A2 0.13595f
C3321 AND8_0.NOT8_0.A7 B6 0.062492f
C3322 mux8_7.NAND4F_0.Y mux8_7.NAND4F_7.Y 0.08762f
C3323 mux8_4.A0 SEL1 0.35149f
C3324 AND8_0.S7 SEL1 0.066504f
C3325 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B 0.087175f
C3326 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 0.008371f
C3327 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 0.00323f
C3328 AND8_0.S6 AND8_0.S7 3.97946f
C3329 MULT_0.4bit_ADDER_0.A2 VDD 3.13158f
C3330 mux8_0.NAND4F_4.B mux8_1.NAND4F_4.B 0.001581f
C3331 mux8_7.A1 A0 0.00125f
C3332 mux8_8.NAND4F_7.Y SEL2 0.176544f
C3333 mux8_8.A1 mux8_8.NAND4F_3.Y 0.541275f
C3334 NOT8_0.S4 B4 0.448605f
C3335 mux8_4.NAND4F_4.B VDD 1.19644f
C3336 mux8_1.NAND4F_5.Y mux8_2.NAND4F_2.D 1.02e-21
C3337 mux8_7.NAND4F_3.Y mux8_7.NAND4F_4.Y 0.102178f
C3338 mux8_7.NAND4F_0.Y mux8_7.NAND4F_8.Y 0.249057f
C3339 AND8_0.NOT8_0.A2 AND8_0.NOT8_0.A3 1.03801f
C3340 mux8_8.NAND4F_0.C VDD 1.403f
C3341 B6 A2 0.020989f
C3342 mux8_7.NAND4F_2.D mux8_7.NAND4F_0.C 1.553f
C3343 8bit_ADDER_0.C mux8_4.A0 0.117789f
C3344 B4 B2 0.019483f
C3345 XOR8_0.S4 B3 0.010513f
C3346 8bit_ADDER_0.S2 SEL0 0.674821f
C3347 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y B7 0.202041f
C3348 mux8_4.NAND4F_0.C SEL2 1.4681f
C3349 OR8_0.S7 B5 0.054115f
C3350 AND8_0.NOT8_0.A2 VDD 2.32492f
C3351 mux8_4.A1 mux8_4.NAND4F_8.Y 1.16e-22
C3352 OR8_0.NOT8_0.A4 OR8_0.NOT8_0.A5 0.118909f
C3353 mux8_4.A1 XOR8_0.S2 0.044778f
C3354 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT SEL3 2e-19
C3355 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A mux8_4.A0 2.76e-19
C3356 mux8_8.NAND4F_2.D SEL2 0.481921f
C3357 MULT_0.4bit_ADDER_2.B2 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A 0.002364f
C3358 B7 A4 0.120508f
C3359 OR8_0.NOT8_0.A5 A3 0.018817f
C3360 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT 0.001576f
C3361 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 0.005944f
C3362 XOR8_0.S3 mux8_4.NAND4F_5.Y 0.602392f
C3363 mux8_7.A0 NOT8_0.S5 2.42e-19
C3364 NOT8_0.S7 SEL1 0.029144f
C3365 NOT8_0.S7 AND8_0.S6 0.028963f
C3366 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B VDD 1.84917f
C3367 AND8_0.S2 B2 0.045987f
C3368 mux8_6.A0 mux8_8.NAND4F_0.C 3.32e-19
C3369 mux8_8.A0 mux8_8.NAND4F_4.Y 0.047022f
C3370 NOT8_0.S1 mux8_7.A1 0.011468f
C3371 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.B0 0.181943f
C3372 mux8_4.A0 mux8_4.A1 4.87148f
C3373 mux8_4.NAND4F_3.Y mux8_4.NAND4F_5.Y 4.33e-19
C3374 XOR8_0.S0 XOR8_0.S2 9.46e-20
C3375 OR8_0.S2 OR8_0.NOT8_0.A1 0.341185f
C3376 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B 2.43e-19
C3377 mux8_5.A0 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A 0.006336f
C3378 8bit_ADDER_0.S0 mux8_1.NAND4F_2.D 0.104289f
C3379 AND8_0.S1 MULT_0.4bit_ADDER_2.B1 1.6e-19
C3380 mux8_6.A1 B3 0.231823f
C3381 B7 A1 0.087613f
C3382 MULT_0.inv_15.Y MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A 0.685441f
C3383 mux8_4.NAND4F_3.Y XOR8_0.S3 5.23e-19
C3384 MULT_0.SO mux8_1.NAND4F_2.Y 1.16938f
C3385 NOT8_0.S0 NOT8_0.S1 0.463276f
C3386 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 0.119902f
C3387 mux8_7.A0 VDD 1.35857f
C3388 mux8_0.NAND4F_5.Y SEL2 0.323263f
C3389 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A mux8_6.A1 0.127125f
C3390 mux8_7.NAND4F_3.Y mux8_7.NAND4F_5.Y 4.33e-19
C3391 mux8_8.NAND4F_9.Y mux8_8.NAND4F_1.Y 0.222572f
C3392 MULT_0.SO VDD 1.69589f
C3393 mux8_2.NAND4F_4.B SEL0 1.61012f
C3394 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A 0.186684f
C3395 mux8_4.A0 XOR8_0.S0 0.022627f
C3396 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT VDD 3.26516f
C3397 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT VDD 3.16726f
C3398 mux8_1.NAND4F_0.Y mux8_1.NAND4F_5.Y 4.32e-19
C3399 left_shifter_0.S7 XOR8_0.S6 0.039982f
C3400 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT A4 0.003441f
C3401 mux8_7.A1 SEL2 0.142863f
C3402 mux8_4.NAND4F_0.Y mux8_4.NAND4F_2.Y 0.170507f
C3403 mux8_5.NAND4F_2.D mux8_5.NAND4F_8.Y 4.88e-20
C3404 mux8_1.NAND4F_4.Y mux8_1.NAND4F_9.Y 5.28e-19
C3405 mux8_7.A1 mux8_7.NAND4F_1.Y 8.98e-23
C3406 8bit_ADDER_0.S2 MULT_0.S2 4.77555f
C3407 mux8_7.NAND4F_4.B mux8_7.NAND4F_3.Y 0.223331f
C3408 mux8_6.A1 XOR8_0.S7 0.080024f
C3409 OR8_0.S1 mux8_5.A1 0.014137f
C3410 mux8_1.NAND4F_9.Y mux8_1.NAND4F_1.Y 0.222572f
C3411 mux8_6.A0 mux8_7.A0 0.030611f
C3412 mux8_6.A0 MULT_0.SO 0.049217f
C3413 mux8_0.NAND4F_2.D mux8_0.NAND4F_5.Y 9.34e-20
C3414 mux8_6.NAND4F_3.Y mux8_6.NAND4F_1.Y 0.086984f
C3415 NOT8_0.S0 SEL2 0.098454f
C3416 AND8_0.S3 AND8_0.S4 0.090083f
C3417 AND8_0.S1 AND8_0.NOT8_0.A3 2.47e-21
C3418 mux8_8.A0 SEL0 0.672711f
C3419 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT 0.001099f
C3420 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B 0.007216f
C3421 mux8_7.NAND4F_6.Y SEL1 0.222305f
C3422 AND8_0.S1 VDD 1.03516f
C3423 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A VDD 1.6936f
C3424 mux8_3.NAND4F_4.B AND8_0.S2 1.04047f
C3425 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A 0.009047f
C3426 AND8_0.S5 B3 0.090106f
C3427 AND8_0.S0 SEL1 0.111325f
C3428 mux8_5.NAND4F_2.Y mux8_5.NAND4F_6.Y 0.08709f
C3429 mux8_6.NAND4F_4.Y XOR8_0.S7 2.3e-19
C3430 mux8_8.A0 mux8_8.NAND4F_4.B 1.52147f
C3431 mux8_2.NAND4F_1.Y VDD 2.18156f
C3432 NOT8_0.S4 B5 0.034463f
C3433 mux8_1.NAND4F_2.D left_shifter_0.S0 4.32e-19
C3434 mux8_5.A0 XOR8_0.S3 0.037309f
C3435 mux8_2.NAND4F_0.Y mux8_2.NAND4F_3.Y 0.616159f
C3436 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT mux8_8.A0 0.720724f
C3437 MULT_0.4bit_ADDER_1.B2 MULT_0.4bit_ADDER_2.B2 0.019679f
C3438 mux8_2.NAND4F_2.D NOT8_0.S1 4.43e-19
C3439 mux8_6.A0 AND8_0.S1 0.016672f
C3440 B5 B2 0.018375f
C3441 mux8_5.NAND4F_6.Y VDD 2.17811f
C3442 AND8_0.NOT8_0.A3 AND8_0.NOT8_0.A4 0.376986f
C3443 XOR8_0.S4 B4 0.240846f
C3444 mux8_8.A1 mux8_8.NAND4F_1.Y 8.98e-23
C3445 V_FLAG_0.XOR2_2.B V_FLAG_0.XOR2_2.Y 0.5618f
C3446 OR8_0.S7 B6 0.049746f
C3447 AND8_0.NOT8_0.A4 VDD 2.32032f
C3448 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A SEL3 7.03e-19
C3449 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y 8bit_ADDER_0.S2 0.018758f
C3450 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A 0.005938f
C3451 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A 0.118063f
C3452 mux8_2.NAND4F_3.Y mux8_2.NAND4F_7.Y 5.28e-20
C3453 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A 2.59e-19
C3454 XOR8_0.S6 mux8_8.NAND4F_6.Y 0.520706f
C3455 mux8_4.A0 mux8_4.NAND4F_4.B 1.5224f
C3456 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A 2.06e-19
C3457 mux8_5.NAND4F_4.B SEL2 0.734121f
C3458 V_FLAG_0.XOR2_0.Y SEL2 3.05e-19
C3459 OR8_0.S1 mux8_2.NAND4F_5.Y 2.34e-19
C3460 mux8_2.NAND4F_0.C VDD 1.40477f
C3461 mux8_6.NAND4F_6.Y Y7 1.95e-20
C3462 ZFLAG_0.nor4_0.Y Y5 1.07e-19
C3463 mux8_3.NAND4F_8.Y mux8_3.NAND4F_5.Y 0.001122f
C3464 mux8_6.NAND4F_9.Y Y7 0.012833f
C3465 MULT_0.4bit_ADDER_1.B0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A 5.19e-20
C3466 AND8_0.S4 OR8_0.NOT8_0.A7 1.82e-19
C3467 mux8_4.NAND4F_2.D SEL1 3.38954f
C3468 mux8_2.NAND4F_2.D SEL2 0.482633f
C3469 mux8_4.NAND4F_0.C mux8_4.NAND4F_5.Y 0.051024f
C3470 AND8_0.S0 mux8_4.A1 0.069391f
C3471 mux8_8.A0 MULT_0.S2 0.025236f
C3472 8bit_ADDER_0.S2 mux8_2.NAND4F_4.B 7.14e-21
C3473 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B VDD 1.82806f
C3474 NOT8_0.S3 SEL1 0.073664f
C3475 MULT_0.4bit_ADDER_1.A2 A1 0.003067f
C3476 mux8_6.A1 B4 0.055127f
C3477 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A 0.248956f
C3478 V_FLAG_0.XOR2_0.Y mux8_0.NAND4F_2.D 2.58e-19
C3479 mux8_4.NAND4F_0.C XOR8_0.S3 0.080897f
C3480 mux8_7.A0 XOR8_0.S2 0.024552f
C3481 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y mux8_5.A0 2.04e-19
C3482 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y A4 3.93e-19
C3483 mux8_3.NAND4F_3.Y mux8_3.NAND4F_1.Y 0.086984f
C3484 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y mux8_5.A0 2.04e-19
C3485 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 0.139263f
C3486 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A VDD 1.30816f
C3487 8bit_ADDER_0.S2 A1 0.441108f
C3488 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A A4 0.008956f
C3489 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A VDD 1.67078f
C3490 mux8_0.NAND4F_0.Y mux8_0.NAND4F_9.Y 2.96e-20
C3491 mux8_6.NAND4F_4.B XOR8_0.S7 0.96335f
C3492 A5 A3 0.027577f
C3493 mux8_1.NAND4F_2.D mux8_1.NAND4F_5.Y 9.34e-20
C3494 AND8_0.S0 XOR8_0.S0 0.025009f
C3495 mux8_0.NAND4F_3.Y mux8_0.NAND4F_5.Y 4.33e-19
C3496 OR8_0.S1 B1 0.013633f
C3497 mux8_4.NAND4F_0.C mux8_4.NAND4F_3.Y 0.399921f
C3498 AND8_0.S2 mux8_6.A1 0.044095f
C3499 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 6.28e-19
C3500 mux8_5.A0 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 0.005184f
C3501 mux8_7.A0 mux8_4.A0 0.010437f
C3502 AND8_0.S5 mux8_7.NAND4F_0.C 0.052524f
C3503 mux8_8.A0 8bit_ADDER_0.S2 1.01e-19
C3504 AND8_0.NOT8_0.A1 AND8_0.S4 2.87e-21
C3505 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y A1 2.72694f
C3506 mux8_4.A0 MULT_0.SO 0.02025f
C3507 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y A1 5.14e-19
C3508 mux8_2.NAND4F_7.Y mux8_3.NAND4F_0.Y 0.002061f
C3509 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y A1 5.14e-19
C3510 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A 0.001919f
C3511 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT mux8_4.A0 0.001724f
C3512 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B 0.005184f
C3513 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y A1 0.004073f
C3514 AND8_0.S1 XOR8_0.S2 8.16e-20
C3515 mux8_5.NAND4F_0.Y SEL2 2.97e-20
C3516 mux8_4.A1 mux8_4.NAND4F_2.D 0.107639f
C3517 mux8_1.NAND4F_8.Y mux8_1.NAND4F_6.Y 2.96e-20
C3518 A4 A1 0.025158f
C3519 mux8_2.NAND4F_2.Y mux8_2.NAND4F_5.Y 4.33e-19
C3520 mux8_2.NAND4F_8.Y mux8_2.NAND4F_9.Y 0.696806f
C3521 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y mux8_8.A0 1.08e-19
C3522 AND8_0.S5 B4 0.635157f
C3523 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y mux8_8.A0 1.08e-19
C3524 mux8_6.NAND4F_6.Y mux8_6.NAND4F_7.Y 0.14618f
C3525 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y mux8_8.A0 0.018985f
C3526 mux8_1.NAND4F_0.Y SEL2 2.97e-20
C3527 mux8_4.A1 NOT8_0.S3 0.009258f
C3528 mux8_8.NAND4F_2.Y mux8_8.NAND4F_6.Y 0.08709f
C3529 mux8_6.NAND4F_9.Y mux8_6.NAND4F_7.Y 0.248336f
C3530 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A mux8_8.A0 9.64e-19
C3531 mux8_7.A1 XOR8_0.S3 0.038314f
C3532 NOT8_0.S4 B6 0.030062f
C3533 mux8_4.A0 AND8_0.S1 0.015326f
C3534 mux8_4.NAND4F_7.Y SEL2 0.176544f
C3535 mux8_5.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B 0.028878f
C3536 MULT_0.inv_15.Y MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT 0.010334f
C3537 mux8_8.NAND4F_4.Y mux8_8.NAND4F_8.Y 0.404949f
C3538 mux8_2.NAND4F_3.Y SEL0 0.360934f
C3539 XOR8_0.S4 B5 0.018312f
C3540 B6 B2 0.018262f
C3541 AND8_0.S2 AND8_0.S5 7.95e-22
C3542 A2 A0 0.309221f
C3543 mux8_3.NAND4F_7.Y SEL2 0.176544f
C3544 mux8_6.NAND4F_2.D mux8_6.NAND4F_6.Y 2.96e-20
C3545 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT mux8_5.A1 0.177096f
C3546 mux8_1.NAND4F_4.B SEL0 1.61016f
C3547 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B VDD 1.97673f
C3548 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 0.132279f
C3549 mux8_5.A0 mux8_4.NAND4F_0.C 8.66e-21
C3550 NOT8_0.S2 SEL0 1.10234f
C3551 AND8_0.S1 OR8_0.NOT8_0.A0 0.001946f
C3552 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B A2 0.009827f
C3553 B7 SEL3 1.17333f
C3554 AND8_0.S0 AND8_0.NOT8_0.A2 2.98e-21
C3555 mux8_3.NAND4F_4.Y mux8_3.NAND4F_9.Y 5.28e-19
C3556 mux8_2.NAND4F_9.Y VDD 2.28332f
C3557 mux8_5.NAND4F_4.Y SEL1 0.30433f
C3558 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B 0.008371f
C3559 mux8_4.A0 mux8_2.NAND4F_0.C 2.46e-19
C3560 mux8_6.A1 B5 0.071925f
C3561 mux8_5.NAND4F_0.C SEL1 1.11989f
C3562 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B 0.00323f
C3563 mux8_1.NAND4F_4.Y SEL1 0.30433f
C3564 mux8_6.NAND4F_2.Y SEL2 3.61e-20
C3565 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT 0.003009f
C3566 SEL3 SEL0 4.24e-21
C3567 mux8_0.NAND4F_2.Y SEL2 3.61e-20
C3568 mux8_8.NAND4F_8.Y SEL0 4.08e-19
C3569 mux8_8.NAND4F_2.D mux8_8.NAND4F_7.Y 2.97e-20
C3570 mux8_1.NAND4F_1.Y SEL1 2.35e-20
C3571 mux8_4.A0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B 0.004182f
C3572 NOT8_0.S0 mux8_1.NAND4F_7.Y 0.431664f
C3573 mux8_3.NAND4F_0.Y SEL0 0.236427f
C3574 mux8_3.NAND4F_4.Y VDD 2.21728f
C3575 mux8_4.NAND4F_2.D mux8_4.NAND4F_4.B 1.27138f
C3576 mux8_7.A0 mux8_7.NAND4F_6.Y 2.97e-22
C3577 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A 0.186684f
C3578 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT SEL3 1.96e-19
C3579 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A VDD 1.66874f
C3580 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A mux8_4.A0 2.76e-19
C3581 mux8_7.A0 AND8_0.S0 0.013827f
C3582 NOT8_0.S1 mux8_2.NAND4F_6.Y 0.79864f
C3583 mux8_4.NAND4F_4.B NOT8_0.S3 0.105153f
C3584 MULT_0.S2 NOT8_0.S2 0.009258f
C3585 AND8_0.S0 MULT_0.SO 10.0202f
C3586 mux8_1.NAND4F_0.C mux8_1.NAND4F_2.Y 0.122872f
C3587 MULT_0.inv_15.Y A2 0.003977f
C3588 mux8_0.NAND4F_2.D mux8_0.NAND4F_2.Y 0.339934f
C3589 OR8_0.S1 AND8_0.S3 0.020288f
C3590 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT 0.094647f
C3591 mux8_3.NAND4F_0.C mux8_3.NAND4F_3.Y 0.399921f
C3592 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A VDD 1.35296f
C3593 mux8_1.NAND4F_0.C VDD 2.55839f
C3594 mux8_5.A0 NOT8_0.S0 0.012053f
C3595 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B VDD 1.85859f
C3596 mux8_3.NAND4F_2.D mux8_3.NAND4F_1.Y 2.96e-20
C3597 B1 A3 1.3619f
C3598 V_FLAG_0.XOR2_2.Y SEL2 0.010007f
C3599 XOR8_0.S1 mux8_5.A1 0.015837f
C3600 AND8_0.S5 B5 0.054593f
C3601 mux8_5.NAND4F_2.D mux8_5.NAND4F_1.Y 2.96e-20
C3602 mux8_6.NAND4F_6.Y SEL1 0.222305f
C3603 mux8_1.NAND4F_2.D SEL2 0.481923f
C3604 mux8_6.A0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 2.35e-19
C3605 mux8_4.NAND4F_2.Y SEL2 3.61e-20
C3606 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 0.792412f
C3607 mux8_5.A0 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A 0.002364f
C3608 8bit_ADDER_0.S2 mux8_1.NAND4F_4.B 5.66e-21
C3609 NOT8_0.S6 OR8_0.S7 1.48e-20
C3610 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B MULT_0.4bit_ADDER_1.B3 0.007216f
C3611 mux8_2.NAND4F_6.Y SEL2 0.419676f
C3612 8bit_ADDER_0.S2 NOT8_0.S2 1.33e-19
C3613 AND8_0.S0 AND8_0.S1 9.237309f
C3614 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 0.012283f
C3615 MULT_0.4bit_ADDER_2.B1 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A 0.002364f
C3616 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 0.00162f
C3617 mux8_4.NAND4F_0.Y mux8_4.NAND4F_9.Y 2.96e-20
C3618 XOR8_0.S4 B6 0.020637f
C3619 AND8_0.S4 B7 0.80678f
C3620 AND8_0.NOT8_0.A6 A4 0.022516f
C3621 mux8_8.A1 XOR8_0.S6 0.078168f
C3622 V_FLAG_0.XOR2_2.Y mux8_0.NAND4F_2.D 0.002215f
C3623 ZFLAG_0.nor4_0.Y ZFLAG_0.nor4_1.Y 0.845159f
C3624 OR8_0.NOT8_0.A6 B3 3.16e-21
C3625 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 1.58859f
C3626 mux8_5.NAND4F_5.Y SEL2 0.323263f
C3627 mux8_8.NAND4F_1.Y SEL1 2.35e-20
C3628 AND8_0.NOT8_0.A5 AND8_0.NOT8_0.A7 8.82e-20
C3629 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT A4 0.129004f
C3630 mux8_1.NAND4F_4.Y XOR8_0.S0 2.3e-19
C3631 mux8_1.NAND4F_7.Y mux8_2.NAND4F_2.D 9.03e-22
C3632 MULT_0.S2 mux8_3.NAND4F_0.Y 0.43187f
C3633 MULT_0.4bit_ADDER_0.B2 B1 0.002129f
C3634 mux8_7.A0 NOT8_0.S3 0.017532f
C3635 mux8_5.A0 mux8_5.NAND4F_4.B 1.52249f
C3636 8bit_ADDER_0.S0 mux8_1.NAND4F_3.Y 0.406267f
C3637 XOR8_0.S0 mux8_1.NAND4F_1.Y 0.404949f
C3638 mux8_8.NAND4F_2.Y mux8_8.NAND4F_9.Y 2.96e-20
C3639 mux8_6.A1 mux8_6.NAND4F_0.Y 0.43187f
C3640 mux8_4.NAND4F_6.Y mux8_4.NAND4F_1.Y 2.45057f
C3641 mux8_4.NAND4F_5.Y mux8_4.NAND4F_7.Y 0.235079f
C3642 AND8_0.S4 SEL0 0.128349f
C3643 mux8_5.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A 0.010664f
C3644 mux8_2.NAND4F_4.B mux8_2.NAND4F_3.Y 0.223331f
C3645 XOR8_0.S3 mux8_4.NAND4F_7.Y 9.74e-20
C3646 8bit_ADDER_0.S2 SEL3 1.72e-19
C3647 mux8_8.NAND4F_0.C mux8_8.NAND4F_3.Y 0.399921f
C3648 XOR8_0.S1 mux8_2.NAND4F_5.Y 0.602392f
C3649 mux8_5.A0 mux8_2.NAND4F_2.D 2.18e-19
C3650 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B 1.2618f
C3651 XOR8_0.S5 XOR8_0.S6 0.349358f
C3652 mux8_6.A1 B6 0.489863f
C3653 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A VDD 1.69389f
C3654 mux8_1.NAND4F_4.B mux8_2.NAND4F_4.B 0.001714f
C3655 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A 0.009184f
C3656 mux8_7.NAND4F_5.Y mux8_8.NAND4F_4.Y 0.002218f
C3657 mux8_7.NAND4F_4.Y SEL0 0.116645f
C3658 mux8_3.NAND4F_6.Y mux8_3.NAND4F_1.Y 2.45057f
C3659 mux8_3.NAND4F_5.Y mux8_3.NAND4F_7.Y 0.235079f
C3660 ZFLAG_0.nor4_1.Y Y0 8.73e-19
C3661 B0 A5 0.03332f
C3662 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A A2 0.001946f
C3663 mux8_6.NAND4F_0.Y mux8_6.NAND4F_4.Y 0.28646f
C3664 mux8_6.NAND4F_3.Y mux8_6.NAND4F_2.Y 1.63543f
C3665 ZFLAG_0.nor4_0.Y Y2 0.013348f
C3666 mux8_4.NAND4F_3.Y mux8_4.NAND4F_7.Y 5.28e-20
C3667 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT mux8_8.A0 0.015636f
C3668 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y SEL3 0.732287f
C3669 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y SEL3 0.732305f
C3670 mux8_3.NAND4F_4.Y XOR8_0.S2 2.3e-19
C3671 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y SEL3 0.735109f
C3672 XOR8_0.S5 A5 0.559514f
C3673 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y SEL3 0.571059f
C3674 mux8_8.A1 mux8_5.A1 0.001375f
C3675 mux8_0.NAND4F_0.Y mux8_0.NAND4F_4.Y 0.28646f
C3676 mux8_0.NAND4F_3.Y mux8_0.NAND4F_2.Y 1.63543f
C3677 MULT_0.4bit_ADDER_1.A2 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A 0.685441f
C3678 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A SEL3 7.01e-19
C3679 mux8_5.NAND4F_2.D SEL0 0.229145f
C3680 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B 0.007216f
C3681 MULT_0.4bit_ADDER_0.B2 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A 0.005938f
C3682 left_shifter_0.S7 mux8_6.NAND4F_0.C 0.052281f
C3683 SEL3 A4 0.253188f
C3684 mux8_7.NAND4F_3.Y mux8_7.NAND4F_7.Y 5.28e-20
C3685 NOT8_0.S5 B3 0.001682f
C3686 mux8_4.NAND4F_0.C mux8_5.NAND4F_4.B 0.002598f
C3687 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A 2.59e-19
C3688 mux8_8.A0 NOT8_0.S2 0.017307f
C3689 mux8_1.NAND4F_0.Y mux8_1.NAND4F_7.Y 0.08762f
C3690 XOR8_0.S1 B1 0.222819f
C3691 NOT8_0.S0 mux8_7.A1 0.012929f
C3692 OR8_0.S7 SEL2 0.029578f
C3693 mux8_8.A1 mux8_8.NAND4F_2.Y 1.16938f
C3694 mux8_5.A1 B0 0.00145f
C3695 mux8_7.NAND4F_3.Y mux8_7.NAND4F_8.Y 0.222524f
C3696 AND8_0.S5 B6 0.044545f
C3697 mux8_7.NAND4F_2.Y mux8_7.NAND4F_4.Y 2.04463f
C3698 mux8_4.A0 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A 2.76e-19
C3699 NOT8_0.S4 NOT8_0.S6 0.011385f
C3700 Y0 Y2 0.010733f
C3701 OR8_0.NOT8_0.A5 AND8_0.S6 0.069685f
C3702 SEL3 A1 0.300936f
C3703 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A 2.56e-19
C3704 mux8_7.NAND4F_5.Y SEL0 0.122766f
C3705 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B VDD 1.8288f
C3706 AND8_0.S3 A3 0.221398f
C3707 mux8_4.A0 mux8_1.NAND4F_0.C 2.46e-19
C3708 AND8_0.NOT8_0.A3 B3 0.174091f
C3709 VDD B3 8.45629f
C3710 mux8_6.NAND4F_0.C mux8_6.NAND4F_5.Y 0.051024f
C3711 AND8_0.NOT8_0.A0 A3 2.81e-19
C3712 A7 A5 0.112835f
C3713 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A A4 0.685441f
C3714 OR8_0.NOT8_0.A6 B4 0.06202f
C3715 B2 A0 1.48093f
C3716 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 0.008371f
C3717 XOR8_0.S3 A2 0.011125f
C3718 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A VDD 1.67113f
C3719 mux8_3.NAND4F_2.D mux8_3.NAND4F_0.C 1.55301f
C3720 mux8_7.NAND4F_4.B SEL0 1.61074f
C3721 mux8_4.NAND4F_2.Y mux8_4.NAND4F_5.Y 4.33e-19
C3722 mux8_7.A1 mux8_5.NAND4F_4.B 4.61e-21
C3723 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 0.001075f
C3724 mux8_7.NAND4F_4.B mux8_8.NAND4F_4.B 0.001581f
C3725 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT 0.127988f
C3726 XOR8_0.S7 VDD 0.797334f
C3727 mux8_4.NAND4F_2.Y XOR8_0.S3 1.49e-19
C3728 MULT_0.SO mux8_1.NAND4F_4.Y 0.157118f
C3729 mux8_0.NAND4F_9.Y SEL2 1.49e-20
C3730 MULT_0.4bit_ADDER_0.A2 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B 0.950228f
C3731 mux8_7.NAND4F_2.Y mux8_7.NAND4F_5.Y 4.33e-19
C3732 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT VDD 3.559f
C3733 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B 0.087175f
C3734 MULT_0.SO mux8_1.NAND4F_1.Y 8.98e-23
C3735 mux8_1.NAND4F_3.Y mux8_1.NAND4F_5.Y 4.33e-19
C3736 mux8_3.NAND4F_8.Y mux8_3.NAND4F_7.Y 9.84e-20
C3737 NOT8_0.S1 B2 6.75e-21
C3738 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A B0 0.009367f
C3739 mux8_4.NAND4F_0.Y mux8_4.NAND4F_4.Y 0.28646f
C3740 mux8_4.NAND4F_3.Y mux8_4.NAND4F_2.Y 1.63543f
C3741 AND8_0.S4 A4 0.007405f
C3742 mux8_1.NAND4F_8.Y mux8_1.NAND4F_9.Y 0.696806f
C3743 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A mux8_8.A0 1.08e-19
C3744 mux8_8.NAND4F_0.C mux8_8.NAND4F_1.Y 0.402437f
C3745 mux8_6.A0 XOR8_0.S7 0.009242f
C3746 NOT8_0.S5 mux8_7.NAND4F_0.C 0.054384f
C3747 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A 0.186684f
C3748 mux8_7.NAND4F_4.B mux8_7.NAND4F_2.Y 0.112019f
C3749 mux8_4.NAND4F_0.C mux8_4.NAND4F_7.Y 0.224691f
C3750 mux8_8.A1 B1 3.35e-19
C3751 B3 A6 0.022007f
C3752 mux8_5.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B 0.005184f
C3753 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y A2 2.72694f
C3754 mux8_6.NAND4F_2.Y mux8_6.NAND4F_1.Y 3.31e-22
C3755 NOT8_0.S4 SEL2 0.096656f
C3756 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A 0.127125f
C3757 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B VDD 1.97177f
C3758 AND8_0.S4 A1 8.6e-19
C3759 NOT8_0.S5 B4 0.584514f
C3760 B1 B0 1.16521f
C3761 mux8_5.NAND4F_4.Y mux8_5.NAND4F_6.Y 4.33e-19
C3762 mux8_1.NAND4F_2.D mux8_1.NAND4F_7.Y 2.97e-20
C3763 mux8_3.NAND4F_0.C mux8_3.NAND4F_6.Y 0.142729f
C3764 mux8_5.A0 A2 9.63e-20
C3765 XOR8_0.S7 A6 0.01001f
C3766 mux8_5.NAND4F_0.C mux8_5.NAND4F_6.Y 0.142729f
C3767 OR8_0.S7 mux8_6.NAND4F_3.Y 2.56e-19
C3768 mux8_7.NAND4F_0.C VDD 1.39513f
C3769 MULT_0.4bit_ADDER_2.B1 AND8_0.S2 1.18e-19
C3770 mux8_2.NAND4F_0.Y mux8_2.NAND4F_2.Y 0.170507f
C3771 mux8_8.A0 AND8_0.S4 0.019293f
C3772 AND8_0.NOT8_0.A1 A3 2.26e-19
C3773 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A 0.009055f
C3774 mux8_0.NAND4F_0.C mux8_0.NAND4F_6.Y 0.142729f
C3775 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT 1.58859f
C3776 XOR8_0.S1 AND8_0.S3 0.021609f
C3777 mux8_7.NAND4F_2.D SEL2 0.481921f
C3778 mux8_1.NAND4F_4.B mux8_2.NAND4F_3.Y 1.02e-21
C3779 NOT8_0.S6 XOR8_0.S4 0.04573f
C3780 mux8_5.A0 mux8_1.NAND4F_2.D 2.18e-19
C3781 AND8_0.NOT8_0.A3 B4 0.019626f
C3782 XOR8_0.S2 B3 0.008591f
C3783 mux8_7.NAND4F_2.D mux8_7.NAND4F_1.Y 2.96e-20
C3784 VDD B4 6.77754f
C3785 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B 0.003236f
C3786 mux8_1.NAND4F_0.C AND8_0.S0 0.037082f
C3787 mux8_7.NAND4F_3.Y XOR8_0.S5 5.23e-19
C3788 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A A7 0.685441f
C3789 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT mux8_7.A1 0.177264f
C3790 OR8_0.NOT8_0.A6 B5 0.031279f
C3791 mux8_1.NAND4F_0.Y NOT8_0.S0 5.24e-19
C3792 OR8_0.S2 mux8_5.A1 0.018541f
C3793 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A MULT_0.4bit_ADDER_1.B0 0.200037f
C3794 mux8_1.NAND4F_1.Y mux8_2.NAND4F_0.C 1.02e-21
C3795 XOR8_0.S6 SEL1 0.097094f
C3796 AND8_0.S6 XOR8_0.S6 8.01e-19
C3797 XOR8_0.S3 OR8_0.S7 0.004998f
C3798 mux8_5.A0 mux8_5.NAND4F_5.Y 2.08e-19
C3799 mux8_4.A0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B 0.004182f
C3800 mux8_4.NAND4F_1.Y SEL1 2.35e-20
C3801 mux8_4.A0 B3 5.02e-19
C3802 AND8_0.S2 AND8_0.NOT8_0.A3 2.48e-21
C3803 AND8_0.S7 B3 0.152005f
C3804 AND8_0.S2 VDD 1.91773f
C3805 MULT_0.4bit_ADDER_1.A2 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT 0.010334f
C3806 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT SEL3 1.95e-19
C3807 OR8_0.S1 SEL0 1.09979f
C3808 mux8_3.NAND4F_1.Y SEL1 2.35e-20
C3809 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A VDD 1.66874f
C3810 mux8_6.A1 NOT8_0.S6 0.047628f
C3811 mux8_3.NAND4F_4.B SEL2 0.734121f
C3812 AND8_0.S6 A5 0.008615f
C3813 A7 B1 0.050107f
C3814 mux8_3.NAND4F_2.Y mux8_3.NAND4F_1.Y 3.31e-22
C3815 mux8_5.NAND4F_9.Y mux8_7.NAND4F_8.Y 0.001427f
C3816 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A VDD 1.33873f
C3817 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A 0.005938f
C3818 mux8_4.NAND4F_9.Y SEL2 1.49e-20
C3819 AND8_0.S7 XOR8_0.S7 1.69e-19
C3820 mux8_6.A1 A0 0.036615f
C3821 mux8_6.A0 AND8_0.S2 0.016672f
C3822 mux8_4.NAND4F_0.C mux8_4.NAND4F_2.Y 0.122872f
C3823 mux8_0.NAND4F_2.Y mux8_0.NAND4F_5.Y 4.33e-19
C3824 left_shifter_0.S7 B7 0.888198f
C3825 8bit_ADDER_0.C A5 0.035357f
C3826 mux8_3.NAND4F_0.Y NOT8_0.S2 5.24e-19
C3827 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B 2.43e-19
C3828 mux8_8.NAND4F_5.Y mux8_6.NAND4F_4.Y 0.002218f
C3829 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 0.119902f
C3830 B4 A6 0.023842f
C3831 NOT8_0.S7 B3 4.65e-20
C3832 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B MULT_0.4bit_ADDER_1.B3 1.26434f
C3833 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A 0.186684f
C3834 mux8_5.A1 SEL1 0.070061f
C3835 mux8_4.A1 mux8_4.NAND4F_1.Y 8.98e-23
C3836 mux8_5.NAND4F_3.Y SEL2 2.96e-20
C3837 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT A4 0.010334f
C3838 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A 0.118063f
C3839 mux8_8.A1 AND8_0.S3 0.030155f
C3840 left_shifter_0.S7 SEL0 0.094947f
C3841 mux8_2.NAND4F_4.Y mux8_2.NAND4F_5.Y 0.087643f
C3842 NOT8_0.S5 B5 0.464495f
C3843 mux8_1.NAND4F_6.Y SEL0 0.353731f
C3844 XOR8_0.S4 SEL2 0.211868f
C3845 mux8_8.NAND4F_4.Y mux8_8.NAND4F_6.Y 4.33e-19
C3846 NOT8_0.S6 AND8_0.S5 0.01597f
C3847 mux8_1.NAND4F_3.Y SEL2 2.96e-20
C3848 NOT8_0.S7 XOR8_0.S7 7.91126f
C3849 OR8_0.S1 MULT_0.S2 0.023167f
C3850 MULT_0.4bit_ADDER_1.A2 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A 1.19e-19
C3851 mux8_8.NAND4F_2.Y SEL1 0.222331f
C3852 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A MULT_0.inv_9.Y 0.001139f
C3853 AND8_0.S6 mux8_8.NAND4F_2.Y 1.24e-19
C3854 mux8_2.NAND4F_2.Y SEL0 0.296541f
C3855 mux8_0.NAND4F_6.Y SEL1 0.222305f
C3856 AND8_0.S3 B0 0.779678f
C3857 mux8_5.A1 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A 0.002364f
C3858 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A mux8_5.A1 0.200037f
C3859 AND8_0.S4 AND8_0.NOT8_0.A6 3.43e-20
C3860 AND8_0.NOT8_0.A0 B0 0.188787f
C3861 XOR8_0.S2 B4 0.004643f
C3862 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B 0.209959f
C3863 mux8_3.NAND4F_0.C OR8_0.S2 0.051008f
C3864 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A VDD 1.69306f
C3865 OR8_0.S2 B1 0.021122f
C3866 XOR8_0.S3 NOT8_0.S4 0.944679f
C3867 VDD B5 5.77943f
C3868 mux8_6.NAND4F_0.Y mux8_6.NAND4F_8.Y 0.249057f
C3869 mux8_6.NAND4F_5.Y SEL0 0.117659f
C3870 VDD Y5 0.979029f
C3871 OR8_0.NOT8_0.A6 B6 0.03152f
C3872 MULT_0.inv_15.Y mux8_6.A1 0.668337f
C3873 mux8_6.A1 SEL2 0.021272f
C3874 XOR8_0.S3 B2 0.014797f
C3875 8bit_ADDER_0.C mux8_0.NAND4F_6.Y 2.97e-22
C3876 mux8_1.NAND4F_2.D NOT8_0.S0 4.43e-19
C3877 mux8_5.A1 mux8_4.A1 1.39356f
C3878 8bit_ADDER_0.S2 OR8_0.S1 0.038808f
C3879 mux8_2.NAND4F_5.Y SEL1 0.306449f
C3880 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A SEL3 7e-19
C3881 AND8_0.S7 B4 0.081945f
C3882 AND8_0.S2 XOR8_0.S2 4.15e-19
C3883 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B 1.2618f
C3884 mux8_4.NAND4F_7.Y mux8_5.NAND4F_0.Y 0.002217f
C3885 B7 A3 0.104369f
C3886 mux8_5.NAND4F_7.Y SEL2 0.176544f
C3887 mux8_8.NAND4F_6.Y SEL0 0.353713f
C3888 mux8_6.NAND4F_4.Y SEL2 8.74e-20
C3889 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A 3.28e-19
C3890 XOR8_0.S0 mux8_5.A1 0.018712f
C3891 mux8_0.NAND4F_4.Y SEL2 8.74e-20
C3892 mux8_4.A0 AND8_0.S2 0.019086f
C3893 mux8_8.NAND4F_4.B mux8_8.NAND4F_6.Y 0.187883f
C3894 mux8_3.NAND4F_3.Y SEL0 0.360934f
C3895 mux8_4.A0 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A 2.76e-19
C3896 MULT_0.4bit_ADDER_1.B3 B1 1.87e-19
C3897 mux8_4.NAND4F_4.B mux8_4.NAND4F_1.Y 0.222551f
C3898 mux8_8.NAND4F_0.C XOR8_0.S6 0.081857f
C3899 8bit_ADDER_0.C 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A 0.188141f
C3900 V_FLAG_0.XOR2_2.Y V_FLAG_0.XOR2_0.Y 0.767153f
C3901 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT 0.003012f
C3902 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A 0.248956f
C3903 AND8_0.S5 SEL2 0.180528f
C3904 XOR8_0.S1 mux8_2.NAND4F_7.Y 9.74e-20
C3905 B5 A6 0.054831f
C3906 mux8_3.NAND4F_0.C SEL1 1.11959f
C3907 NOT8_0.S7 B4 5.81e-20
C3908 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B VDD 1.82878f
C3909 mux8_2.NAND4F_4.B OR8_0.S1 0.079695f
C3910 mux8_1.NAND4F_0.C mux8_1.NAND4F_4.Y 0.049743f
C3911 mux8_0.NAND4F_2.D mux8_0.NAND4F_4.Y 0.349681f
C3912 AND8_0.S2 OR8_0.NOT8_0.A0 0.016829f
C3913 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y B2 0.202041f
C3914 mux8_3.NAND4F_0.C mux8_3.NAND4F_2.Y 0.122872f
C3915 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT A7 0.010334f
C3916 mux8_4.NAND4F_9.Y mux8_4.NAND4F_5.Y 0.402985f
C3917 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_1.B0 0.697503f
C3918 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B 0.139263f
C3919 OR8_0.S1 A1 0.015539f
C3920 mux8_1.NAND4F_0.C mux8_1.NAND4F_1.Y 0.402437f
C3921 mux8_3.NAND4F_4.B mux8_3.NAND4F_5.Y 0.248856f
C3922 mux8_5.A0 NOT8_0.S4 1.11e-19
C3923 NOT8_0.S5 B6 0.036298f
C3924 MULT_0.4bit_ADDER_2.B2 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A 2.56e-19
C3925 mux8_5.NAND4F_4.B mux8_5.NAND4F_5.Y 0.248856f
C3926 NOT8_0.S3 B3 0.511429f
C3927 mux8_2.NAND4F_2.D mux8_2.NAND4F_6.Y 2.96e-20
C3928 8bit_ADDER_0.C B1 0.008271f
C3929 AND8_0.NOT8_0.A1 B0 0.015331f
C3930 mux8_4.NAND4F_4.Y SEL2 8.74e-20
C3931 MULT_0.4bit_ADDER_1.B2 VDD 2.025f
C3932 mux8_8.A0 OR8_0.S1 0.024803f
C3933 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A B1 0.001945f
C3934 mux8_6.NAND4F_0.Y VDD 2.13487f
C3935 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A MULT_0.4bit_ADDER_1.B3 0.127125f
C3936 MULT_0.4bit_ADDER_0.A2 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B 0.00981f
C3937 mux8_0.NAND4F_0.Y VDD 2.13434f
C3938 mux8_0.NAND4F_6.Y mux8_0.NAND4F_1.Y 2.45057f
C3939 mux8_7.NAND4F_0.C mux8_7.NAND4F_6.Y 0.142729f
C3940 XOR8_0.S2 B5 0.003214f
C3941 mux8_6.NAND4F_4.B SEL2 0.734112f
C3942 OR8_0.NOT8_0.A7 A7 0.255162f
C3943 VDD B6 5.68514f
C3944 mux8_0.NAND4F_0.C mux8_0.NAND4F_4.B 2.13077f
C3945 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A mux8_8.A0 1.08e-19
C3946 MULT_0.S2 mux8_3.NAND4F_3.Y 0.541275f
C3947 XOR8_0.S3 XOR8_0.S4 2.40327f
C3948 mux8_8.NAND4F_4.Y mux8_8.NAND4F_9.Y 5.28e-19
C3949 8bit_ADDER_0.S0 mux8_1.NAND4F_2.Y 0.200461f
C3950 mux8_0.NAND4F_0.C mux8_0.NAND4F_7.Y 0.224691f
C3951 mux8_6.A1 mux8_6.NAND4F_3.Y 0.541275f
C3952 mux8_7.NAND4F_7.Y SEL0 0.234594f
C3953 AND8_0.NOT8_0.A5 AND8_0.S5 0.393093f
C3954 OR8_0.S2 AND8_0.S3 2.48365f
C3955 8bit_ADDER_0.S0 VDD 1.00337f
C3956 AND8_0.S7 B5 0.123533f
C3957 mux8_6.NAND4F_0.C mux8_6.NAND4F_7.Y 0.224691f
C3958 mux8_2.NAND4F_4.B mux8_2.NAND4F_2.Y 0.112019f
C3959 mux8_8.NAND4F_0.C mux8_8.NAND4F_2.Y 0.122872f
C3960 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT 0.132279f
C3961 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B 0.087175f
C3962 MULT_0.4bit_ADDER_1.A2 A3 0.006603f
C3963 mux8_0.NAND4F_9.Y mux8_0.NAND4F_5.Y 0.402985f
C3964 mux8_1.NAND4F_2.D mux8_1.NAND4F_0.Y 0.184536f
C3965 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A 8.33e-19
C3966 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A 1.01138f
C3967 mux8_7.NAND4F_8.Y SEL0 4.08e-19
C3968 8bit_ADDER_0.S2 mux8_3.NAND4F_3.Y 0.406267f
C3969 mux8_5.NAND4F_0.Y mux8_5.NAND4F_5.Y 4.32e-19
C3970 mux8_1.NAND4F_9.Y mux8_2.NAND4F_0.Y 1.02e-21
C3971 mux8_4.NAND4F_0.Y VDD 2.13487f
C3972 mux8_6.NAND4F_3.Y mux8_6.NAND4F_4.Y 0.102178f
C3973 mux8_6.A0 8bit_ADDER_0.S0 0.427226f
C3974 XOR8_0.S1 SEL0 0.167333f
C3975 mux8_6.NAND4F_2.D mux8_6.NAND4F_0.C 1.55388f
C3976 AND8_0.S0 AND8_0.S2 5.05e-19
C3977 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT MULT_0.inv_9.Y 0.034931f
C3978 mux8_6.A1 XOR8_0.S3 0.043557f
C3979 mux8_0.NAND4F_0.Y mux8_0.NAND4F_8.Y 0.249057f
C3980 mux8_7.A0 mux8_5.A1 0.022439f
C3981 mux8_0.NAND4F_3.Y mux8_0.NAND4F_4.Y 0.102178f
C3982 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT mux8_5.A1 0.742096f
C3983 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A 0.127125f
C3984 B6 A6 52.6843f
C3985 NOT8_0.S7 B5 6.31e-19
C3986 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y A3 2.7267f
C3987 AND8_0.S0 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A 2.06e-19
C3988 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y A3 8.66e-19
C3989 mux8_1.NAND4F_3.Y mux8_1.NAND4F_7.Y 5.28e-20
C3990 OR8_0.NOT8_0.A4 A4 0.256957f
C3991 mux8_8.NAND4F_9.Y SEL0 2.8e-19
C3992 mux8_8.A1 mux8_8.NAND4F_4.Y 0.157118f
C3993 A4 A3 0.068495f
C3994 mux8_7.A1 NOT8_0.S4 0.019866f
C3995 mux8_7.NAND4F_2.Y mux8_7.NAND4F_8.Y 0.222339f
C3996 mux8_5.A0 mux8_5.NAND4F_3.Y 0.406267f
C3997 AND8_0.S3 SEL1 0.110785f
C3998 mux8_5.NAND4F_2.D AND8_0.S4 0.076916f
C3999 AND8_0.NOT8_0.A4 A5 3.23e-20
C4000 AND8_0.S3 AND8_0.S6 1.86e-19
C4001 mux8_4.A0 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B 0.018146f
C4002 NOT8_0.S3 B4 0.206776f
C4003 left_shifter_0.S0 VDD 2.09067f
C4004 AND8_0.S1 mux8_5.A1 0.01438f
C4005 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT SEL3 1.92e-19
C4006 mux8_3.NAND4F_2.D SEL0 0.229749f
C4007 MULT_0.4bit_ADDER_0.A2 B1 0.001792f
C4008 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A mux8_5.A1 2.28e-19
C4009 mux8_5.A0 XOR8_0.S4 0.009216f
C4010 mux8_8.A0 mux8_8.NAND4F_6.Y 2.97e-22
C4011 mux8_1.NAND4F_5.Y mux8_2.NAND4F_8.Y 1.02e-21
C4012 mux8_3.NAND4F_0.C mux8_4.NAND4F_4.B 0.002598f
C4013 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A VDD 1.66874f
C4014 XOR8_0.S3 AND8_0.S5 0.031581f
C4015 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT 8bit_ADDER_0.S2 0.152789f
C4016 V_FLAG_0.XOR2_2.B VDD 0.92091f
C4017 A3 A1 0.676097f
C4018 mux8_4.NAND4F_0.C mux8_4.NAND4F_9.Y 4.79e-21
C4019 ZFLAG_0.nor4_1.Y VDD 0.228523f
C4020 mux8_7.A1 mux8_7.NAND4F_2.D 0.108116f
C4021 AND8_0.NOT8_0.A2 B1 0.013841f
C4022 XOR8_0.S2 B6 0.001548f
C4023 mux8_6.A0 left_shifter_0.S0 0.017859f
C4024 MULT_0.S2 XOR8_0.S1 0.029851f
C4025 mux8_0.NAND4F_4.B SEL1 4.35973f
C4026 S VSS 0.576747f
C4027 Y7 VSS 9.981952f
C4028 Y6 VSS 11.002562f
C4029 Y5 VSS 6.283913f
C4030 Y4 VSS 2.82598f
C4031 Z VSS 0.574471f
C4032 Y3 VSS 2.70484f
C4033 Y2 VSS 8.094442f
C4034 Y1 VSS 13.512403f
C4035 Y0 VSS 10.534714f
C4036 C VSS 0.636653f
C4037 A0 VSS 60.469715f
C4038 A1 VSS 60.198044f
C4039 A2 VSS 50.80682f
C4040 A3 VSS 47.31751f
C4041 A4 VSS 72.80435f
C4042 A5 VSS 68.22108f
C4043 A6 VSS 66.44732f
C4044 SEL0 VSS 65.05544f
C4045 SEL1 VSS 46.216084f
C4046 SEL2 VSS 55.184315f
C4047 B0 VSS 53.558285f
C4048 B1 VSS 49.44086f
C4049 B2 VSS 48.782375f
C4050 B3 VSS 48.467052f
C4051 B4 VSS 42.144352f
C4052 B5 VSS 48.35252f
C4053 B6 VSS 67.65343f
C4054 V VSS 0.584393f
C4055 SEL3 VSS 31.55541f
C4056 B7 VSS 71.146904f
C4057 A7 VSS 67.321236f
C4058 VDD VSS 1.477444p
C4059 mux8_6.NAND4F_7.Y VSS 2.530448f
C4060 mux8_6.NAND4F_1.Y VSS 3.905086f
C4061 mux8_6.NAND4F_6.Y VSS 2.459403f
C4062 mux8_6.NAND4F_5.Y VSS 3.571911f
C4063 mux8_6.NAND4F_9.Y VSS 2.63083f
C4064 mux8_6.NAND4F_8.Y VSS 2.630238f
C4065 XOR8_0.S7 VSS 17.756603f
C4066 mux8_6.NAND4F_4.Y VSS 3.953424f
C4067 mux8_6.NAND4F_2.Y VSS 2.515674f
C4068 mux8_6.NAND4F_3.Y VSS 2.678273f
C4069 mux8_6.NAND4F_0.Y VSS 2.620947f
C4070 mux8_6.NAND4F_4.B VSS 4.855343f
C4071 mux8_6.NAND4F_0.C VSS 6.4159f
C4072 mux8_6.NAND4F_2.D VSS 3.664538f
C4073 mux8_8.NAND4F_7.Y VSS 2.527498f
C4074 mux8_8.NAND4F_1.Y VSS 3.902316f
C4075 mux8_8.NAND4F_6.Y VSS 2.456373f
C4076 mux8_8.NAND4F_5.Y VSS 3.569941f
C4077 XOR8_0.S6 VSS 24.204159f
C4078 mux8_8.NAND4F_9.Y VSS 2.64868f
C4079 mux8_8.NAND4F_8.Y VSS 2.630278f
C4080 mux8_8.NAND4F_4.Y VSS 3.953424f
C4081 mux8_8.NAND4F_2.Y VSS 2.515674f
C4082 mux8_8.NAND4F_3.Y VSS 2.678273f
C4083 mux8_8.NAND4F_0.Y VSS 2.620947f
C4084 mux8_8.NAND4F_4.B VSS 4.854973f
C4085 mux8_8.NAND4F_0.C VSS 5.926896f
C4086 mux8_8.NAND4F_2.D VSS 3.635502f
C4087 mux8_7.NAND4F_7.Y VSS 2.527498f
C4088 mux8_7.NAND4F_1.Y VSS 3.902316f
C4089 mux8_7.NAND4F_6.Y VSS 2.456373f
C4090 mux8_7.NAND4F_5.Y VSS 3.569801f
C4091 XOR8_0.S5 VSS 30.5012f
C4092 mux8_7.NAND4F_9.Y VSS 2.64564f
C4093 mux8_7.NAND4F_8.Y VSS 2.630068f
C4094 mux8_7.NAND4F_4.Y VSS 3.953404f
C4095 mux8_7.NAND4F_2.Y VSS 2.515674f
C4096 mux8_7.NAND4F_3.Y VSS 2.678273f
C4097 mux8_7.NAND4F_0.Y VSS 2.620947f
C4098 mux8_7.NAND4F_4.B VSS 4.861272f
C4099 mux8_7.NAND4F_0.C VSS 5.929299f
C4100 mux8_7.NAND4F_2.D VSS 3.636972f
C4101 mux8_5.NAND4F_7.Y VSS 2.527498f
C4102 mux8_5.NAND4F_1.Y VSS 3.902316f
C4103 mux8_5.NAND4F_6.Y VSS 2.456373f
C4104 mux8_5.NAND4F_5.Y VSS 3.569891f
C4105 OR8_0.S7 VSS 33.60993f
C4106 AND8_0.S7 VSS 25.541004f
C4107 AND8_0.NOT8_0.A7 VSS 3.701097f
C4108 OR8_0.NOT8_0.A7 VSS 2.8824f
C4109 XOR8_0.S4 VSS 21.59798f
C4110 mux8_5.NAND4F_9.Y VSS 2.64865f
C4111 left_shifter_0.S7 VSS 23.236803f
C4112 OR8_0.NOT8_0.A6 VSS 1.84584f
C4113 AND8_0.S6 VSS 38.43716f
C4114 AND8_0.NOT8_0.A6 VSS 2.690751f
C4115 AND8_0.S5 VSS 36.90735f
C4116 AND8_0.NOT8_0.A5 VSS 2.202838f
C4117 OR8_0.NOT8_0.A5 VSS 1.65065f
C4118 OR8_0.NOT8_0.A4 VSS 1.40916f
C4119 mux8_5.NAND4F_8.Y VSS 2.630298f
C4120 mux8_5.NAND4F_4.Y VSS 3.953404f
C4121 mux8_5.NAND4F_2.Y VSS 2.515674f
C4122 mux8_5.NAND4F_3.Y VSS 2.678273f
C4123 mux8_5.NAND4F_0.Y VSS 2.620947f
C4124 AND8_0.S4 VSS 35.568565f
C4125 AND8_0.NOT8_0.A4 VSS 2.628171f
C4126 mux8_5.NAND4F_4.B VSS 4.854593f
C4127 mux8_5.NAND4F_0.C VSS 5.940899f
C4128 mux8_5.NAND4F_2.D VSS 3.627452f
C4129 NOT8_0.S7 VSS 26.57448f
C4130 OR8_0.NOT8_0.A3 VSS 1.79661f
C4131 ZFLAG_0.nor4_1.Y VSS 2.33398f
C4132 NOT8_0.S6 VSS 23.949272f
C4133 AND8_0.NOT8_0.A3 VSS 2.906079f
C4134 ZFLAG_0.nor4_0.Y VSS 2.36682f
C4135 NOT8_0.S5 VSS 22.13711f
C4136 mux8_4.NAND4F_7.Y VSS 2.527498f
C4137 mux8_4.NAND4F_1.Y VSS 3.902316f
C4138 mux8_4.NAND4F_6.Y VSS 2.456373f
C4139 mux8_4.NAND4F_5.Y VSS 3.570111f
C4140 NOT8_0.S4 VSS 21.5774f
C4141 AND8_0.NOT8_0.A2 VSS 3.048563f
C4142 OR8_0.NOT8_0.A2 VSS 1.87294f
C4143 NOT8_0.S3 VSS 15.62932f
C4144 XOR8_0.S3 VSS 19.727846f
C4145 mux8_4.NAND4F_9.Y VSS 2.64874f
C4146 AND8_0.NOT8_0.A1 VSS 3.367471f
C4147 OR8_0.NOT8_0.A1 VSS 1.84722f
C4148 mux8_4.NAND4F_8.Y VSS 2.630198f
C4149 mux8_4.NAND4F_4.Y VSS 3.953424f
C4150 mux8_4.NAND4F_2.Y VSS 2.515694f
C4151 mux8_4.NAND4F_3.Y VSS 2.678273f
C4152 mux8_4.NAND4F_0.Y VSS 2.620947f
C4153 AND8_0.S3 VSS 26.826406f
C4154 mux8_4.NAND4F_4.B VSS 4.860043f
C4155 mux8_4.NAND4F_0.C VSS 5.925688f
C4156 mux8_4.NAND4F_2.D VSS 3.633722f
C4157 AND8_0.NOT8_0.A0 VSS 4.447208f
C4158 OR8_0.NOT8_0.A0 VSS 2.79371f
C4159 mux8_3.NAND4F_7.Y VSS 2.527498f
C4160 mux8_3.NAND4F_1.Y VSS 3.902316f
C4161 mux8_3.NAND4F_6.Y VSS 2.456373f
C4162 mux8_3.NAND4F_5.Y VSS 3.569661f
C4163 mux8_6.A1 VSS 35.856014f
C4164 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.B VSS 2.06422f
C4165 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_2.A VSS 1.90576f
C4166 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.B VSS 1.83397f
C4167 MULT_0.4bit_ADDER_2.FULL_ADDER_2.NAND2_2.A VSS 0.884942f
C4168 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.B VSS 1.8542f
C4169 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_2.A VSS 0.892161f
C4170 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.B VSS 1.87674f
C4171 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_2.A VSS 0.90243f
C4172 NOT8_0.S2 VSS 26.022652f
C4173 XOR8_0.S2 VSS 27.056906f
C4174 mux8_3.NAND4F_9.Y VSS 2.64736f
C4175 mux8_3.NAND4F_8.Y VSS 2.630408f
C4176 mux8_4.A1 VSS 21.267946f
C4177 mux8_5.A1 VSS 27.873066f
C4178 mux8_7.A1 VSS 37.724857f
C4179 mux8_8.A1 VSS 34.382652f
C4180 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A VSS 5.371498f
C4181 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT VSS 6.520818f
C4182 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A VSS 3.763987f
C4183 MULT_0.inv_9.Y VSS 14.685481f
C4184 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT VSS 6.358377f
C4185 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A VSS 3.761637f
C4186 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT VSS 6.383528f
C4187 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A VSS 3.758327f
C4188 MULT_0.inv_15.Y VSS 4.057219f
C4189 mux8_3.NAND4F_4.Y VSS 3.953834f
C4190 mux8_3.NAND4F_2.Y VSS 2.516054f
C4191 mux8_3.NAND4F_3.Y VSS 2.678643f
C4192 mux8_3.NAND4F_0.Y VSS 2.621477f
C4193 OR8_0.S2 VSS 32.90203f
C4194 AND8_0.S2 VSS 49.60307f
C4195 mux8_3.NAND4F_4.B VSS 4.857792f
C4196 mux8_3.NAND4F_0.C VSS 5.962939f
C4197 mux8_3.NAND4F_2.D VSS 3.693452f
C4198 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.B VSS 1.94635f
C4199 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_2.A VSS 1.89752f
C4200 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.B VSS 1.67277f
C4201 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_2.A VSS 0.868503f
C4202 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.B VSS 1.66074f
C4203 MULT_0.4bit_ADDER_1.FULL_ADDER_1.NAND2_2.A VSS 0.868104f
C4204 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.B VSS 1.65744f
C4205 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_2.A VSS 0.867708f
C4206 mux8_2.NAND4F_7.Y VSS 2.528028f
C4207 mux8_2.NAND4F_1.Y VSS 3.902686f
C4208 mux8_2.NAND4F_6.Y VSS 2.456733f
C4209 mux8_2.NAND4F_5.Y VSS 3.570461f
C4210 NOT8_0.S1 VSS 41.80846f
C4211 XOR8_0.S1 VSS 39.509735f
C4212 mux8_2.NAND4F_9.Y VSS 2.64872f
C4213 MULT_0.S2 VSS 24.395802f
C4214 MULT_0.4bit_ADDER_2.B1 VSS 5.296375f
C4215 MULT_0.4bit_ADDER_2.B2 VSS 5.266288f
C4216 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A VSS 5.365667f
C4217 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT VSS 6.555182f
C4218 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A VSS 3.757387f
C4219 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT VSS 6.346919f
C4220 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A VSS 3.753927f
C4221 MULT_0.4bit_ADDER_1.A2 VSS 5.606205f
C4222 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT VSS 6.321439f
C4223 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A VSS 3.750067f
C4224 mux8_2.NAND4F_8.Y VSS 2.630008f
C4225 mux8_2.NAND4F_4.Y VSS 3.952874f
C4226 mux8_2.NAND4F_2.Y VSS 2.515194f
C4227 mux8_2.NAND4F_3.Y VSS 2.677063f
C4228 mux8_2.NAND4F_0.Y VSS 2.620177f
C4229 OR8_0.S1 VSS 52.68481f
C4230 AND8_0.S1 VSS 71.887505f
C4231 MULT_0.4bit_ADDER_1.B3 VSS 7.416202f
C4232 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.B VSS 1.94618f
C4233 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_2.A VSS 1.89748f
C4234 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.B VSS 1.67292f
C4235 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_2.A VSS 0.868522f
C4236 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.B VSS 1.6609f
C4237 MULT_0.4bit_ADDER_0.FULL_ADDER_1.NAND2_2.A VSS 0.868123f
C4238 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.B VSS 1.77269f
C4239 MULT_0.4bit_ADDER_0.FULL_ADDER_0.NAND2_2.A VSS 0.867727f
C4240 mux8_2.NAND4F_4.B VSS 4.857652f
C4241 mux8_2.NAND4F_0.C VSS 5.967943f
C4242 mux8_2.NAND4F_2.D VSS 3.639622f
C4243 MULT_0.4bit_ADDER_1.B0 VSS 5.332882f
C4244 MULT_0.4bit_ADDER_1.B1 VSS 5.251795f
C4245 MULT_0.4bit_ADDER_1.B2 VSS 6.013672f
C4246 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A VSS 5.369798f
C4247 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT VSS 6.555082f
C4248 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A VSS 3.761007f
C4249 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT VSS 6.346179f
C4250 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A VSS 3.755827f
C4251 MULT_0.4bit_ADDER_0.A2 VSS 5.692927f
C4252 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT VSS 6.32515f
C4253 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A VSS 3.997557f
C4254 mux8_1.NAND4F_7.Y VSS 2.526718f
C4255 mux8_1.NAND4F_1.Y VSS 3.901066f
C4256 mux8_1.NAND4F_6.Y VSS 2.455883f
C4257 mux8_1.NAND4F_5.Y VSS 3.569121f
C4258 NOT8_0.S0 VSS 39.935345f
C4259 XOR8_0.S0 VSS 40.661583f
C4260 left_shifter_0.S0 VSS 35.64056f
C4261 mux8_1.NAND4F_9.Y VSS 2.64807f
C4262 MULT_0.4bit_ADDER_0.B2 VSS 6.967605f
C4263 mux8_1.NAND4F_8.Y VSS 2.594868f
C4264 mux8_1.NAND4F_4.Y VSS 3.935111f
C4265 mux8_1.NAND4F_2.Y VSS 2.492794f
C4266 mux8_1.NAND4F_3.Y VSS 2.668517f
C4267 mux8_1.NAND4F_0.Y VSS 2.622518f
C4268 MULT_0.SO VSS 28.171358f
C4269 AND8_0.S0 VSS 57.08197f
C4270 mux8_1.NAND4F_4.B VSS 4.834332f
C4271 mux8_1.NAND4F_0.C VSS 5.957524f
C4272 mux8_1.NAND4F_2.D VSS 3.495212f
C4273 mux8_0.NAND4F_7.Y VSS 2.959778f
C4274 mux8_0.NAND4F_1.Y VSS 4.857377f
C4275 mux8_0.NAND4F_6.Y VSS 3.776243f
C4276 mux8_0.NAND4F_5.Y VSS 4.460581f
C4277 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.B VSS 1.83418f
C4278 8bit_ADDER_0.FULL_ADDER_XORED_7.NAND2_2.A VSS 0.88994f
C4279 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.B VSS 1.83571f
C4280 8bit_ADDER_0.FULL_ADDER_XORED_6.NAND2_2.A VSS 0.889051f
C4281 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.B VSS 1.84703f
C4282 8bit_ADDER_0.FULL_ADDER_XORED_5.NAND2_2.A VSS 0.891779f
C4283 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.B VSS 1.85539f
C4284 8bit_ADDER_0.FULL_ADDER_XORED_4.NAND2_2.A VSS 0.893631f
C4285 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.B VSS 1.86226f
C4286 8bit_ADDER_0.FULL_ADDER_XORED_3.NAND2_2.A VSS 0.895143f
C4287 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.B VSS 1.84179f
C4288 8bit_ADDER_0.FULL_ADDER_XORED_2.NAND2_2.A VSS 0.887789f
C4289 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.B VSS 1.83146f
C4290 8bit_ADDER_0.FULL_ADDER_XORED_1.NAND2_2.A VSS 0.890532f
C4291 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.B VSS 1.85572f
C4292 8bit_ADDER_0.FULL_ADDER_XORED_0.NAND2_2.A VSS 0.902927f
C4293 mux8_0.NAND4F_9.Y VSS 2.64857f
C4294 8bit_ADDER_0.S0 VSS 12.69156f
C4295 8bit_ADDER_0.S2 VSS 21.34066f
C4296 mux8_4.A0 VSS 28.319302f
C4297 mux8_5.A0 VSS 41.503902f
C4298 mux8_7.A0 VSS 43.662483f
C4299 mux8_8.A0 VSS 45.992508f
C4300 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A VSS 3.789287f
C4301 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT VSS 6.290631f
C4302 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A VSS 3.782427f
C4303 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT VSS 6.199451f
C4304 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A VSS 3.782707f
C4305 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT VSS 6.216218f
C4306 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A VSS 3.782947f
C4307 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT VSS 6.218491f
C4308 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A VSS 3.783167f
C4309 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT VSS 6.207281f
C4310 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A VSS 3.782947f
C4311 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT VSS 6.197631f
C4312 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A VSS 3.780097f
C4313 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT VSS 6.259958f
C4314 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A VSS 3.783517f
C4315 mux8_0.NAND4F_8.Y VSS 2.632418f
C4316 mux8_0.NAND4F_4.Y VSS 5.042604f
C4317 mux8_0.NAND4F_2.Y VSS 4.091314f
C4318 mux8_0.NAND4F_3.Y VSS 3.223563f
C4319 mux8_0.NAND4F_0.Y VSS 3.056837f
C4320 8bit_ADDER_0.C VSS 22.77708f
C4321 mux8_0.NAND4F_4.B VSS 7.152422f
C4322 mux8_0.NAND4F_0.C VSS 6.231926f
C4323 mux8_0.NAND4F_2.D VSS 3.916722f
C4324 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y VSS 5.366589f
C4325 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y VSS 5.364839f
C4326 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y VSS 5.364319f
C4327 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y VSS 5.364779f
C4328 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y VSS 5.364619f
C4329 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y VSS 5.364009f
C4330 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y VSS 5.363539f
C4331 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y VSS 5.567189f
C4332 V_FLAG_0.XOR2_0.Y VSS 2.405839f
C4333 mux8_6.A0 VSS 37.83299f
C4334 V_FLAG_0.XOR2_2.Y VSS 4.529007f
C4335 V_FLAG_0.XOR2_2.B VSS 2.661607f
C4336 right_shifter_0.S1.n0 VSS 8.33998f
C4337 mux8_2.NAND4F_6.A VSS 0.948172f
C4338 right_shifter_0.S1.t6 VSS 0.071826f
C4339 right_shifter_0.S1.t5 VSS 0.211621f
C4340 right_shifter_0.S1.t4 VSS 0.069882f
C4341 right_shifter_0.S1.n1 VSS 0.360292f
C4342 right_shifter_0.S1.t3 VSS 0.034431f
C4343 right_shifter_0.S1.t2 VSS 0.034431f
C4344 right_shifter_0.S1.n2 VSS 0.076728f
C4345 right_shifter_0.S1.t1 VSS 0.124883f
C4346 right_shifter_0.S1.t0 VSS 0.099312f
C4347 mux8_2.A7 VSS 8.92844f
C4348 left_shifter_0.S4.n0 VSS 7.10775f
C4349 mux8_5.NAND4F_5.A VSS 0.966515f
C4350 left_shifter_0.S4.t5 VSS 0.079776f
C4351 left_shifter_0.S4.t4 VSS 0.235044f
C4352 left_shifter_0.S4.t6 VSS 0.077617f
C4353 left_shifter_0.S4.n1 VSS 0.40017f
C4354 left_shifter_0.S4.t2 VSS 0.038243f
C4355 left_shifter_0.S4.t3 VSS 0.038243f
C4356 left_shifter_0.S4.n2 VSS 0.085311f
C4357 left_shifter_0.S4.t1 VSS 0.138805f
C4358 left_shifter_0.S4.t0 VSS 0.110304f
C4359 mux8_5.A6 VSS 6.62223f
C4360 left_shifter_0.S6.n0 VSS 8.84196f
C4361 mux8_8.NAND4F_5.A VSS 0.774942f
C4362 left_shifter_0.S6.t5 VSS 0.063797f
C4363 left_shifter_0.S6.t4 VSS 0.187963f
C4364 left_shifter_0.S6.t6 VSS 0.06207f
C4365 left_shifter_0.S6.n1 VSS 0.320013f
C4366 left_shifter_0.S6.t2 VSS 0.030582f
C4367 left_shifter_0.S6.t3 VSS 0.030582f
C4368 left_shifter_0.S6.n2 VSS 0.068223f
C4369 left_shifter_0.S6.t1 VSS 0.111001f
C4370 left_shifter_0.S6.t0 VSS 0.088209f
C4371 mux8_8.A6 VSS 8.62066f
C4372 mux8_4.NAND4F_8.Y.n0 VSS 0.539804f
C4373 mux8_4.NAND4F_8.Y.t9 VSS 0.026899f
C4374 mux8_4.NAND4F_8.Y.t10 VSS 0.028853f
C4375 mux8_4.NAND4F_8.Y.n1 VSS 0.042994f
C4376 mux8_4.NAND4F_8.Y.t11 VSS 0.026899f
C4377 mux8_4.NAND4F_8.Y.t13 VSS 0.026899f
C4378 mux8_4.NAND4F_8.Y.t12 VSS 0.026899f
C4379 mux8_4.NAND4F_8.Y.t14 VSS 0.033983f
C4380 mux8_4.NAND4F_8.Y.n2 VSS 0.072608f
C4381 mux8_4.NAND4F_8.Y.n3 VSS 0.045714f
C4382 mux8_4.NAND4F_8.Y.n4 VSS 0.037354f
C4383 mux8_4.NAND4F_8.Y.n5 VSS 0.018278f
C4384 mux8_4.NAND4F_8.Y.t4 VSS 0.026614f
C4385 mux8_4.NAND4F_8.Y.t5 VSS 0.026614f
C4386 mux8_4.NAND4F_8.Y.n6 VSS 0.0618f
C4387 mux8_4.NAND4F_8.Y.t1 VSS 0.026614f
C4388 mux8_4.NAND4F_8.Y.t0 VSS 0.026614f
C4389 mux8_4.NAND4F_8.Y.n7 VSS 0.061615f
C4390 mux8_4.NAND4F_8.Y.t3 VSS 0.026614f
C4391 mux8_4.NAND4F_8.Y.t2 VSS 0.026614f
C4392 mux8_4.NAND4F_8.Y.n8 VSS 0.061615f
C4393 mux8_4.NAND4F_8.Y.t8 VSS 0.026614f
C4394 mux8_4.NAND4F_8.Y.t7 VSS 0.026614f
C4395 mux8_4.NAND4F_8.Y.n9 VSS 0.061615f
C4396 mux8_4.NAND4F_8.Y.n10 VSS 0.268281f
C4397 mux8_4.NAND4F_8.Y.t6 VSS 0.21369f
C4398 OR8_0.S7.n0 VSS 1.76297f
C4399 OR8_0.S7.t4 VSS 0.085128f
C4400 OR8_0.S7.t6 VSS 0.082824f
C4401 OR8_0.S7.t5 VSS 0.250813f
C4402 OR8_0.S7.n1 VSS 0.427017f
C4403 OR8_0.S7.t2 VSS 0.040808f
C4404 OR8_0.S7.t3 VSS 0.040808f
C4405 OR8_0.S7.n2 VSS 0.090938f
C4406 OR8_0.S7.t1 VSS 0.14801f
C4407 OR8_0.S7.t0 VSS 0.117704f
C4408 mux8_3.NAND4F_6.Y.n0 VSS 0.599344f
C4409 mux8_3.NAND4F_6.Y.t2 VSS 0.244548f
C4410 mux8_3.NAND4F_6.Y.t10 VSS 0.038543f
C4411 mux8_3.NAND4F_6.Y.t11 VSS 0.118929f
C4412 mux8_3.NAND4F_6.Y.t9 VSS 0.044398f
C4413 mux8_3.NAND4F_6.Y.n1 VSS 0.149236f
C4414 mux8_3.NAND4F_6.Y.n2 VSS 0.032396f
C4415 mux8_3.NAND4F_6.Y.n3 VSS 1.72835f
C4416 mux8_3.NAND4F_6.Y.t1 VSS 0.029549f
C4417 mux8_3.NAND4F_6.Y.t0 VSS 0.029549f
C4418 mux8_3.NAND4F_6.Y.n4 VSS 0.068617f
C4419 mux8_3.NAND4F_6.Y.t5 VSS 0.029549f
C4420 mux8_3.NAND4F_6.Y.t6 VSS 0.029549f
C4421 mux8_3.NAND4F_6.Y.n5 VSS 0.068411f
C4422 mux8_3.NAND4F_6.Y.t8 VSS 0.029549f
C4423 mux8_3.NAND4F_6.Y.t7 VSS 0.029549f
C4424 mux8_3.NAND4F_6.Y.n6 VSS 0.068411f
C4425 mux8_3.NAND4F_6.Y.t4 VSS 0.029549f
C4426 mux8_3.NAND4F_6.Y.t3 VSS 0.029549f
C4427 mux8_3.NAND4F_6.Y.n7 VSS 0.068411f
C4428 mux8_3.NAND4F_6.Y.n8 VSS 0.281208f
C4429 mux8_4.NAND4F_2.Y.n0 VSS 0.530078f
C4430 mux8_4.NAND4F_2.Y.t1 VSS 0.026135f
C4431 mux8_4.NAND4F_2.Y.t0 VSS 0.026135f
C4432 mux8_4.NAND4F_2.Y.n1 VSS 0.060687f
C4433 mux8_4.NAND4F_2.Y.t6 VSS 0.026135f
C4434 mux8_4.NAND4F_2.Y.t5 VSS 0.026135f
C4435 mux8_4.NAND4F_2.Y.n2 VSS 0.060505f
C4436 mux8_4.NAND4F_2.Y.t7 VSS 0.026135f
C4437 mux8_4.NAND4F_2.Y.t8 VSS 0.026135f
C4438 mux8_4.NAND4F_2.Y.n3 VSS 0.060505f
C4439 mux8_4.NAND4F_2.Y.t4 VSS 0.026135f
C4440 mux8_4.NAND4F_2.Y.t3 VSS 0.026135f
C4441 mux8_4.NAND4F_2.Y.n4 VSS 0.060505f
C4442 mux8_4.NAND4F_2.Y.n5 VSS 0.263447f
C4443 mux8_4.NAND4F_2.Y.t2 VSS 0.213114f
C4444 mux8_4.NAND4F_2.Y.t11 VSS 0.034088f
C4445 mux8_4.NAND4F_2.Y.t9 VSS 0.105185f
C4446 mux8_4.NAND4F_2.Y.t10 VSS 0.039267f
C4447 mux8_4.NAND4F_2.Y.n6 VSS 0.131989f
C4448 mux8_4.NAND4F_2.Y.n7 VSS 0.028742f
C4449 mux8_4.NAND4F_2.Y.n8 VSS 1.53344f
C4450 a_n13975_n11063.n0 VSS 1.48365f
C4451 a_n13975_n11063.n1 VSS 1.48326f
C4452 a_n13975_n11063.t1 VSS 0.093341f
C4453 a_n13975_n11063.t3 VSS 0.093341f
C4454 a_n13975_n11063.t4 VSS 0.093341f
C4455 a_n13975_n11063.n2 VSS 0.202296f
C4456 a_n13975_n11063.t5 VSS 0.093341f
C4457 a_n13975_n11063.t9 VSS 0.093341f
C4458 a_n13975_n11063.n3 VSS 0.202001f
C4459 a_n13975_n11063.t10 VSS 0.093341f
C4460 a_n13975_n11063.t11 VSS 0.093341f
C4461 a_n13975_n11063.n4 VSS 0.202001f
C4462 a_n13975_n11063.t8 VSS 0.093341f
C4463 a_n13975_n11063.t7 VSS 0.093341f
C4464 a_n13975_n11063.n5 VSS 0.20269f
C4465 a_n13975_n11063.t0 VSS 0.093341f
C4466 a_n13975_n11063.t6 VSS 0.093341f
C4467 a_n13975_n11063.n6 VSS 0.202001f
C4468 a_n13975_n11063.n7 VSS 0.202001f
C4469 a_n13975_n11063.t2 VSS 0.093341f
C4470 mux8_6.NAND4F_2.Y.n0 VSS 0.530078f
C4471 mux8_6.NAND4F_2.Y.t1 VSS 0.026135f
C4472 mux8_6.NAND4F_2.Y.t0 VSS 0.026135f
C4473 mux8_6.NAND4F_2.Y.n1 VSS 0.060687f
C4474 mux8_6.NAND4F_2.Y.t5 VSS 0.026135f
C4475 mux8_6.NAND4F_2.Y.t6 VSS 0.026135f
C4476 mux8_6.NAND4F_2.Y.n2 VSS 0.060505f
C4477 mux8_6.NAND4F_2.Y.t8 VSS 0.026135f
C4478 mux8_6.NAND4F_2.Y.t7 VSS 0.026135f
C4479 mux8_6.NAND4F_2.Y.n3 VSS 0.060505f
C4480 mux8_6.NAND4F_2.Y.t2 VSS 0.026135f
C4481 mux8_6.NAND4F_2.Y.t4 VSS 0.026135f
C4482 mux8_6.NAND4F_2.Y.n4 VSS 0.060505f
C4483 mux8_6.NAND4F_2.Y.n5 VSS 0.263447f
C4484 mux8_6.NAND4F_2.Y.t3 VSS 0.213114f
C4485 mux8_6.NAND4F_2.Y.t11 VSS 0.034088f
C4486 mux8_6.NAND4F_2.Y.t9 VSS 0.105185f
C4487 mux8_6.NAND4F_2.Y.t10 VSS 0.039267f
C4488 mux8_6.NAND4F_2.Y.n6 VSS 0.131989f
C4489 mux8_6.NAND4F_2.Y.n7 VSS 0.028742f
C4490 mux8_6.NAND4F_2.Y.n8 VSS 1.53344f
C4491 right_shifter_0.S3.n0 VSS 1.94576f
C4492 mux8_4.NAND4F_6.A VSS 0.386792f
C4493 right_shifter_0.S3.t5 VSS 0.0293f
C4494 right_shifter_0.S3.t4 VSS 0.086328f
C4495 right_shifter_0.S3.t6 VSS 0.028507f
C4496 right_shifter_0.S3.n1 VSS 0.146976f
C4497 right_shifter_0.S3.t3 VSS 0.014046f
C4498 right_shifter_0.S3.t2 VSS 0.014046f
C4499 right_shifter_0.S3.n2 VSS 0.0313f
C4500 right_shifter_0.S3.t1 VSS 0.050944f
C4501 right_shifter_0.S3.t0 VSS 0.040513f
C4502 mux8_4.A7 VSS 1.82548f
C4503 right_shifter_0.S6.n0 VSS 4.06786f
C4504 mux8_8.NAND4F_6.A VSS 0.419174f
C4505 right_shifter_0.S6.t5 VSS 0.031753f
C4506 right_shifter_0.S6.t4 VSS 0.093555f
C4507 right_shifter_0.S6.t6 VSS 0.030894f
C4508 right_shifter_0.S6.n1 VSS 0.15928f
C4509 right_shifter_0.S6.t3 VSS 0.015222f
C4510 right_shifter_0.S6.t2 VSS 0.015222f
C4511 right_shifter_0.S6.n2 VSS 0.033921f
C4512 right_shifter_0.S6.t1 VSS 0.055209f
C4513 right_shifter_0.S6.t0 VSS 0.043904f
C4514 mux8_8.A7 VSS 3.834f
C4515 a_n9125_n11063.n0 VSS 1.48365f
C4516 a_n9125_n11063.n1 VSS 1.48326f
C4517 a_n9125_n11063.t3 VSS 0.093341f
C4518 a_n9125_n11063.t9 VSS 0.093341f
C4519 a_n9125_n11063.t10 VSS 0.093341f
C4520 a_n9125_n11063.n2 VSS 0.202296f
C4521 a_n9125_n11063.t11 VSS 0.093341f
C4522 a_n9125_n11063.t2 VSS 0.093341f
C4523 a_n9125_n11063.n3 VSS 0.202001f
C4524 a_n9125_n11063.t1 VSS 0.093341f
C4525 a_n9125_n11063.t0 VSS 0.093341f
C4526 a_n9125_n11063.n4 VSS 0.202001f
C4527 a_n9125_n11063.t7 VSS 0.093341f
C4528 a_n9125_n11063.t8 VSS 0.093341f
C4529 a_n9125_n11063.n5 VSS 0.202001f
C4530 a_n9125_n11063.t6 VSS 0.093341f
C4531 a_n9125_n11063.t4 VSS 0.093341f
C4532 a_n9125_n11063.n6 VSS 0.202001f
C4533 a_n9125_n11063.n7 VSS 0.20269f
C4534 a_n9125_n11063.t5 VSS 0.093341f
C4535 mux8_5.NAND4F_1.Y.n0 VSS 0.655599f
C4536 mux8_5.NAND4F_1.Y.t6 VSS 0.306614f
C4537 mux8_5.NAND4F_1.Y.t11 VSS 0.132168f
C4538 mux8_5.NAND4F_1.Y.t10 VSS 0.04216f
C4539 mux8_5.NAND4F_1.Y.t9 VSS 0.04216f
C4540 mux8_5.NAND4F_1.Y.n1 VSS 0.049498f
C4541 mux8_5.NAND4F_1.Y.n2 VSS 0.277534f
C4542 mux8_5.NAND4F_1.Y.t1 VSS 0.032323f
C4543 mux8_5.NAND4F_1.Y.t0 VSS 0.032323f
C4544 mux8_5.NAND4F_1.Y.n3 VSS 0.075057f
C4545 mux8_5.NAND4F_1.Y.t3 VSS 0.032323f
C4546 mux8_5.NAND4F_1.Y.t2 VSS 0.032323f
C4547 mux8_5.NAND4F_1.Y.n4 VSS 0.074832f
C4548 mux8_5.NAND4F_1.Y.t5 VSS 0.032323f
C4549 mux8_5.NAND4F_1.Y.t4 VSS 0.032323f
C4550 mux8_5.NAND4F_1.Y.n5 VSS 0.074832f
C4551 mux8_5.NAND4F_1.Y.t8 VSS 0.032323f
C4552 mux8_5.NAND4F_1.Y.t7 VSS 0.032323f
C4553 mux8_5.NAND4F_1.Y.n6 VSS 0.074832f
C4554 mux8_5.NAND4F_1.Y.n7 VSS 0.307603f
C4555 OR8_0.S6.n0 VSS 2.17413f
C4556 mux8_8.NAND4F_2.A VSS 1.67384f
C4557 OR8_0.S6.t4 VSS 0.104932f
C4558 OR8_0.S6.t5 VSS 0.102092f
C4559 OR8_0.S6.t6 VSS 0.309159f
C4560 OR8_0.S6.n1 VSS 0.526354f
C4561 mux8_8.A3 VSS 12.7354f
C4562 OR8_0.S6.t3 VSS 0.050301f
C4563 OR8_0.S6.t1 VSS 0.050301f
C4564 OR8_0.S6.n2 VSS 0.112093f
C4565 OR8_0.S6.t2 VSS 0.182442f
C4566 OR8_0.S6.t0 VSS 0.145085f
C4567 OR8_0.NOT8_0.S6 VSS 9.53386f
C4568 mux8_3.NAND4F_2.Y.n0 VSS 0.530078f
C4569 mux8_3.NAND4F_2.Y.t4 VSS 0.026135f
C4570 mux8_3.NAND4F_2.Y.t3 VSS 0.026135f
C4571 mux8_3.NAND4F_2.Y.n1 VSS 0.060687f
C4572 mux8_3.NAND4F_2.Y.t5 VSS 0.026135f
C4573 mux8_3.NAND4F_2.Y.t6 VSS 0.026135f
C4574 mux8_3.NAND4F_2.Y.n2 VSS 0.060505f
C4575 mux8_3.NAND4F_2.Y.t8 VSS 0.026135f
C4576 mux8_3.NAND4F_2.Y.t7 VSS 0.026135f
C4577 mux8_3.NAND4F_2.Y.n3 VSS 0.060505f
C4578 mux8_3.NAND4F_2.Y.t2 VSS 0.026135f
C4579 mux8_3.NAND4F_2.Y.t1 VSS 0.026135f
C4580 mux8_3.NAND4F_2.Y.n4 VSS 0.060505f
C4581 mux8_3.NAND4F_2.Y.n5 VSS 0.263447f
C4582 mux8_3.NAND4F_2.Y.t0 VSS 0.213114f
C4583 mux8_3.NAND4F_2.Y.t11 VSS 0.034088f
C4584 mux8_3.NAND4F_2.Y.t9 VSS 0.105185f
C4585 mux8_3.NAND4F_2.Y.t10 VSS 0.039267f
C4586 mux8_3.NAND4F_2.Y.n6 VSS 0.131989f
C4587 mux8_3.NAND4F_2.Y.n7 VSS 0.028742f
C4588 mux8_3.NAND4F_2.Y.n8 VSS 1.53344f
C4589 a_n17266_n11063.n0 VSS 1.48365f
C4590 a_n17266_n11063.n1 VSS 1.48326f
C4591 a_n17266_n11063.t1 VSS 0.093341f
C4592 a_n17266_n11063.t9 VSS 0.093341f
C4593 a_n17266_n11063.t10 VSS 0.093341f
C4594 a_n17266_n11063.n2 VSS 0.202296f
C4595 a_n17266_n11063.t11 VSS 0.093341f
C4596 a_n17266_n11063.t7 VSS 0.093341f
C4597 a_n17266_n11063.n3 VSS 0.202001f
C4598 a_n17266_n11063.t8 VSS 0.093341f
C4599 a_n17266_n11063.t6 VSS 0.093341f
C4600 a_n17266_n11063.n4 VSS 0.202001f
C4601 a_n17266_n11063.t3 VSS 0.093341f
C4602 a_n17266_n11063.t5 VSS 0.093341f
C4603 a_n17266_n11063.n5 VSS 0.202001f
C4604 a_n17266_n11063.t4 VSS 0.093341f
C4605 a_n17266_n11063.t0 VSS 0.093341f
C4606 a_n17266_n11063.n6 VSS 0.202001f
C4607 a_n17266_n11063.n7 VSS 0.20269f
C4608 a_n17266_n11063.t2 VSS 0.093341f
C4609 NOT8_0.S1.n0 VSS 3.61822f
C4610 NOT8_0.S1.t4 VSS 0.175296f
C4611 NOT8_0.S1.t5 VSS 0.516473f
C4612 NOT8_0.S1.t6 VSS 0.170551f
C4613 NOT8_0.S1.n1 VSS 0.879311f
C4614 NOT8_0.S1.t1 VSS 0.084032f
C4615 NOT8_0.S1.t3 VSS 0.084032f
C4616 NOT8_0.S1.n2 VSS 0.187259f
C4617 NOT8_0.S1.t2 VSS 0.304782f
C4618 NOT8_0.S1.t0 VSS 0.242375f
C4619 a_n15707_n7799.n0 VSS 1.48365f
C4620 a_n15707_n7799.n1 VSS 1.48326f
C4621 a_n15707_n7799.t5 VSS 0.093341f
C4622 a_n15707_n7799.t8 VSS 0.093341f
C4623 a_n15707_n7799.t7 VSS 0.093341f
C4624 a_n15707_n7799.n2 VSS 0.202296f
C4625 a_n15707_n7799.t6 VSS 0.093341f
C4626 a_n15707_n7799.t10 VSS 0.093341f
C4627 a_n15707_n7799.n3 VSS 0.202001f
C4628 a_n15707_n7799.t11 VSS 0.093341f
C4629 a_n15707_n7799.t9 VSS 0.093341f
C4630 a_n15707_n7799.n4 VSS 0.202001f
C4631 a_n15707_n7799.t4 VSS 0.093341f
C4632 a_n15707_n7799.t3 VSS 0.093341f
C4633 a_n15707_n7799.n5 VSS 0.202001f
C4634 a_n15707_n7799.t1 VSS 0.093341f
C4635 a_n15707_n7799.t0 VSS 0.093341f
C4636 a_n15707_n7799.n6 VSS 0.20269f
C4637 a_n15707_n7799.n7 VSS 0.202001f
C4638 a_n15707_n7799.t2 VSS 0.093341f
C4639 mux8_8.NAND4F_8.Y.n0 VSS 0.539804f
C4640 mux8_8.NAND4F_8.Y.t14 VSS 0.026899f
C4641 mux8_8.NAND4F_8.Y.t13 VSS 0.028853f
C4642 mux8_8.NAND4F_8.Y.n1 VSS 0.042994f
C4643 mux8_8.NAND4F_8.Y.t9 VSS 0.026899f
C4644 mux8_8.NAND4F_8.Y.t11 VSS 0.026899f
C4645 mux8_8.NAND4F_8.Y.t10 VSS 0.026899f
C4646 mux8_8.NAND4F_8.Y.t12 VSS 0.033983f
C4647 mux8_8.NAND4F_8.Y.n2 VSS 0.072608f
C4648 mux8_8.NAND4F_8.Y.n3 VSS 0.045714f
C4649 mux8_8.NAND4F_8.Y.n4 VSS 0.037354f
C4650 mux8_8.NAND4F_8.Y.n5 VSS 0.018278f
C4651 mux8_8.NAND4F_8.Y.t2 VSS 0.026614f
C4652 mux8_8.NAND4F_8.Y.t3 VSS 0.026614f
C4653 mux8_8.NAND4F_8.Y.n6 VSS 0.0618f
C4654 mux8_8.NAND4F_8.Y.t1 VSS 0.026614f
C4655 mux8_8.NAND4F_8.Y.t0 VSS 0.026614f
C4656 mux8_8.NAND4F_8.Y.n7 VSS 0.061615f
C4657 mux8_8.NAND4F_8.Y.t5 VSS 0.026614f
C4658 mux8_8.NAND4F_8.Y.t4 VSS 0.026614f
C4659 mux8_8.NAND4F_8.Y.n8 VSS 0.061615f
C4660 mux8_8.NAND4F_8.Y.t8 VSS 0.026614f
C4661 mux8_8.NAND4F_8.Y.t7 VSS 0.026614f
C4662 mux8_8.NAND4F_8.Y.n9 VSS 0.061615f
C4663 mux8_8.NAND4F_8.Y.n10 VSS 0.268281f
C4664 mux8_8.NAND4F_8.Y.t6 VSS 0.21369f
C4665 mux8_4.NAND4F_3.Y.n0 VSS 0.306333f
C4666 mux8_4.NAND4F_3.Y.t1 VSS 0.015103f
C4667 mux8_4.NAND4F_3.Y.t0 VSS 0.015103f
C4668 mux8_4.NAND4F_3.Y.n1 VSS 0.035071f
C4669 mux8_4.NAND4F_3.Y.t3 VSS 0.015103f
C4670 mux8_4.NAND4F_3.Y.t2 VSS 0.015103f
C4671 mux8_4.NAND4F_3.Y.n2 VSS 0.034966f
C4672 mux8_4.NAND4F_3.Y.t5 VSS 0.015103f
C4673 mux8_4.NAND4F_3.Y.t4 VSS 0.015103f
C4674 mux8_4.NAND4F_3.Y.n3 VSS 0.034966f
C4675 mux8_4.NAND4F_3.Y.t8 VSS 0.015103f
C4676 mux8_4.NAND4F_3.Y.t7 VSS 0.015103f
C4677 mux8_4.NAND4F_3.Y.n4 VSS 0.034966f
C4678 mux8_4.NAND4F_3.Y.n5 VSS 0.152246f
C4679 mux8_4.NAND4F_3.Y.t6 VSS 0.143521f
C4680 mux8_4.NAND4F_3.Y.t10 VSS 0.0197f
C4681 mux8_4.NAND4F_3.Y.t11 VSS 0.0197f
C4682 mux8_4.NAND4F_3.Y.n6 VSS 0.023128f
C4683 mux8_4.NAND4F_3.Y.t9 VSS 0.061756f
C4684 mux8_4.NAND4F_3.Y.n7 VSS 0.129679f
C4685 a_n17266_n4534.n0 VSS 1.48326f
C4686 a_n17266_n4534.n1 VSS 1.48365f
C4687 a_n17266_n4534.t1 VSS 0.093341f
C4688 a_n17266_n4534.t4 VSS 0.093341f
C4689 a_n17266_n4534.t3 VSS 0.093341f
C4690 a_n17266_n4534.n2 VSS 0.20269f
C4691 a_n17266_n4534.t6 VSS 0.093341f
C4692 a_n17266_n4534.t5 VSS 0.093341f
C4693 a_n17266_n4534.n3 VSS 0.202001f
C4694 a_n17266_n4534.t8 VSS 0.093341f
C4695 a_n17266_n4534.t7 VSS 0.093341f
C4696 a_n17266_n4534.n4 VSS 0.202001f
C4697 a_n17266_n4534.t11 VSS 0.093341f
C4698 a_n17266_n4534.t9 VSS 0.093341f
C4699 a_n17266_n4534.n5 VSS 0.202001f
C4700 a_n17266_n4534.t0 VSS 0.093341f
C4701 a_n17266_n4534.t10 VSS 0.093341f
C4702 a_n17266_n4534.n6 VSS 0.202001f
C4703 a_n17266_n4534.n7 VSS 0.202296f
C4704 a_n17266_n4534.t2 VSS 0.093341f
C4705 mux8_3.NAND4F_1.Y.n0 VSS 0.655599f
C4706 mux8_3.NAND4F_1.Y.t2 VSS 0.306614f
C4707 mux8_3.NAND4F_1.Y.t9 VSS 0.132168f
C4708 mux8_3.NAND4F_1.Y.t11 VSS 0.04216f
C4709 mux8_3.NAND4F_1.Y.t10 VSS 0.04216f
C4710 mux8_3.NAND4F_1.Y.n1 VSS 0.049498f
C4711 mux8_3.NAND4F_1.Y.n2 VSS 0.277534f
C4712 mux8_3.NAND4F_1.Y.t1 VSS 0.032323f
C4713 mux8_3.NAND4F_1.Y.t0 VSS 0.032323f
C4714 mux8_3.NAND4F_1.Y.n3 VSS 0.075057f
C4715 mux8_3.NAND4F_1.Y.t8 VSS 0.032323f
C4716 mux8_3.NAND4F_1.Y.t7 VSS 0.032323f
C4717 mux8_3.NAND4F_1.Y.n4 VSS 0.074832f
C4718 mux8_3.NAND4F_1.Y.t6 VSS 0.032323f
C4719 mux8_3.NAND4F_1.Y.t5 VSS 0.032323f
C4720 mux8_3.NAND4F_1.Y.n5 VSS 0.074832f
C4721 mux8_3.NAND4F_1.Y.t3 VSS 0.032323f
C4722 mux8_3.NAND4F_1.Y.t4 VSS 0.032323f
C4723 mux8_3.NAND4F_1.Y.n6 VSS 0.074832f
C4724 mux8_3.NAND4F_1.Y.n7 VSS 0.307603f
C4725 mux8_8.NAND4F_2.Y.n0 VSS 0.530078f
C4726 mux8_8.NAND4F_2.Y.t1 VSS 0.026135f
C4727 mux8_8.NAND4F_2.Y.t0 VSS 0.026135f
C4728 mux8_8.NAND4F_2.Y.n1 VSS 0.060687f
C4729 mux8_8.NAND4F_2.Y.t2 VSS 0.026135f
C4730 mux8_8.NAND4F_2.Y.t3 VSS 0.026135f
C4731 mux8_8.NAND4F_2.Y.n2 VSS 0.060505f
C4732 mux8_8.NAND4F_2.Y.t5 VSS 0.026135f
C4733 mux8_8.NAND4F_2.Y.t4 VSS 0.026135f
C4734 mux8_8.NAND4F_2.Y.n3 VSS 0.060505f
C4735 mux8_8.NAND4F_2.Y.t6 VSS 0.026135f
C4736 mux8_8.NAND4F_2.Y.t7 VSS 0.026135f
C4737 mux8_8.NAND4F_2.Y.n4 VSS 0.060505f
C4738 mux8_8.NAND4F_2.Y.n5 VSS 0.263447f
C4739 mux8_8.NAND4F_2.Y.t8 VSS 0.213114f
C4740 mux8_8.NAND4F_2.Y.t10 VSS 0.034088f
C4741 mux8_8.NAND4F_2.Y.t11 VSS 0.105185f
C4742 mux8_8.NAND4F_2.Y.t9 VSS 0.039267f
C4743 mux8_8.NAND4F_2.Y.n6 VSS 0.131989f
C4744 mux8_8.NAND4F_2.Y.n7 VSS 0.028742f
C4745 mux8_8.NAND4F_2.Y.n8 VSS 1.53344f
C4746 OR8_0.S2.n0 VSS 2.14487f
C4747 OR8_0.S2.t4 VSS 0.103766f
C4748 OR8_0.S2.t6 VSS 0.100957f
C4749 OR8_0.S2.t5 VSS 0.305724f
C4750 OR8_0.S2.n1 VSS 0.520505f
C4751 OR8_0.S2.t2 VSS 0.049742f
C4752 OR8_0.S2.t3 VSS 0.049742f
C4753 OR8_0.S2.n2 VSS 0.110847f
C4754 OR8_0.S2.t1 VSS 0.180415f
C4755 OR8_0.S2.t0 VSS 0.143473f
C4756 left_shifter_0.S2.n0 VSS 10.157599f
C4757 mux8_3.NAND4F_5.A VSS 1.26327f
C4758 left_shifter_0.S2.t4 VSS 0.103997f
C4759 left_shifter_0.S2.t6 VSS 0.306406f
C4760 left_shifter_0.S2.t5 VSS 0.101182f
C4761 left_shifter_0.S2.n1 VSS 0.521666f
C4762 left_shifter_0.S2.t2 VSS 0.049853f
C4763 left_shifter_0.S2.t3 VSS 0.049853f
C4764 left_shifter_0.S2.n2 VSS 0.111213f
C4765 left_shifter_0.S2.t1 VSS 0.180948f
C4766 left_shifter_0.S2.t0 VSS 0.143793f
C4767 mux8_3.A6 VSS 9.2102f
C4768 AND8_0.NOT8_0.A6.n0 VSS 0.749958f
C4769 AND8_0.NOT8_0.A6.t7 VSS 0.018598f
C4770 AND8_0.NOT8_0.A6.t8 VSS 0.025961f
C4771 AND8_0.NOT8_0.A6.t9 VSS 0.025961f
C4772 AND8_0.NOT8_0.A6.n1 VSS 0.084508f
C4773 AND8_0.NOT8_0.A6.t10 VSS 0.029791f
C4774 AND8_0.NOT8_0.A6.n2 VSS 0.258271f
C4775 AND8_0.NOT8_0.A6.t0 VSS 0.088073f
C4776 AND8_0.NOT8_0.A6.t2 VSS 0.014593f
C4777 AND8_0.NOT8_0.A6.t1 VSS 0.014593f
C4778 AND8_0.NOT8_0.A6.n3 VSS 0.032471f
C4779 AND8_0.NOT8_0.A6.t5 VSS 0.014593f
C4780 AND8_0.NOT8_0.A6.t4 VSS 0.014593f
C4781 AND8_0.NOT8_0.A6.n4 VSS 0.03256f
C4782 AND8_0.NOT8_0.A6.t3 VSS 0.014593f
C4783 AND8_0.NOT8_0.A6.t6 VSS 0.014593f
C4784 AND8_0.NOT8_0.A6.n5 VSS 0.032471f
C4785 MULT_0.4bit_ADDER_2.B1.t15 VSS 0.041628f
C4786 MULT_0.4bit_ADDER_2.B1.t14 VSS 0.013556f
C4787 MULT_0.4bit_ADDER_2.B1.t21 VSS 0.01872f
C4788 MULT_0.4bit_ADDER_2.B1.n0 VSS 0.020187f
C4789 MULT_0.4bit_ADDER_2.B1.t13 VSS 0.013936f
C4790 MULT_0.4bit_ADDER_2.B1.n1 VSS 0.035362f
C4791 MULT_0.4bit_ADDER_2.B1.n2 VSS 0.062031f
C4792 MULT_0.4bit_ADDER_2.B1.t16 VSS 0.019007f
C4793 MULT_0.4bit_ADDER_2.B1.t19 VSS 0.038242f
C4794 MULT_0.4bit_ADDER_2.B1.t22 VSS 0.037766f
C4795 MULT_0.4bit_ADDER_2.B1.t17 VSS 0.037766f
C4796 MULT_0.4bit_ADDER_2.B1.t23 VSS 0.037766f
C4797 MULT_0.4bit_ADDER_2.B1.t12 VSS 0.007848f
C4798 MULT_0.4bit_ADDER_2.B1.t20 VSS 0.007848f
C4799 MULT_0.4bit_ADDER_2.B1.t18 VSS 0.007848f
C4800 MULT_0.4bit_ADDER_2.B1.n3 VSS 0.232672f
C4801 MULT_0.4bit_ADDER_2.B1.n4 VSS 0.171374f
C4802 MULT_0.4bit_ADDER_2.B1.n5 VSS 0.093397f
C4803 MULT_0.4bit_ADDER_2.B1.n6 VSS 0.091755f
C4804 MULT_0.4bit_ADDER_2.B1.n7 VSS 0.05644f
C4805 MULT_0.4bit_ADDER_2.B1.n8 VSS 0.074039f
C4806 MULT_0.4bit_ADDER_2.B1.n9 VSS 0.814584f
C4807 MULT_0.4bit_ADDER_2.B1.t1 VSS 0.006802f
C4808 MULT_0.4bit_ADDER_2.B1.t2 VSS 0.006802f
C4809 MULT_0.4bit_ADDER_2.B1.n10 VSS 0.016451f
C4810 MULT_0.4bit_ADDER_2.B1.t4 VSS 0.006802f
C4811 MULT_0.4bit_ADDER_2.B1.t6 VSS 0.006802f
C4812 MULT_0.4bit_ADDER_2.B1.n11 VSS 0.016449f
C4813 MULT_0.4bit_ADDER_2.B1.n12 VSS 0.117953f
C4814 MULT_0.4bit_ADDER_2.B1.t0 VSS 0.006802f
C4815 MULT_0.4bit_ADDER_2.B1.t3 VSS 0.006802f
C4816 MULT_0.4bit_ADDER_2.B1.n13 VSS 0.013603f
C4817 MULT_0.4bit_ADDER_2.B1.n14 VSS 0.010686f
C4818 MULT_0.4bit_ADDER_2.B1.t9 VSS 0.028776f
C4819 MULT_0.4bit_ADDER_2.B1.t5 VSS 0.028776f
C4820 MULT_0.4bit_ADDER_2.B1.n15 VSS 0.057553f
C4821 MULT_0.4bit_ADDER_2.B1.n16 VSS 0.022884f
C4822 MULT_0.4bit_ADDER_2.B1.t10 VSS 0.028776f
C4823 MULT_0.4bit_ADDER_2.B1.t11 VSS 0.028776f
C4824 MULT_0.4bit_ADDER_2.B1.n17 VSS 0.057553f
C4825 MULT_0.4bit_ADDER_2.B1.n18 VSS 0.025313f
C4826 MULT_0.4bit_ADDER_2.B1.n19 VSS 0.260608f
C4827 MULT_0.4bit_ADDER_2.B1.t7 VSS 0.028776f
C4828 MULT_0.4bit_ADDER_2.B1.t8 VSS 0.028776f
C4829 MULT_0.4bit_ADDER_2.B1.n20 VSS 0.057553f
C4830 MULT_0.4bit_ADDER_2.B1.n21 VSS 0.025351f
C4831 MULT_0.4bit_ADDER_2.B1.n22 VSS 0.167143f
C4832 MULT_0.4bit_ADDER_2.B1.n23 VSS 0.037667f
C4833 MULT_0.4bit_ADDER_2.B1.n24 VSS 0.165331f
C4834 left_shifter_0.S3.n0 VSS 5.30967f
C4835 mux8_4.NAND4F_5.A VSS 0.806447f
C4836 left_shifter_0.S3.t5 VSS 0.06639f
C4837 left_shifter_0.S3.t4 VSS 0.195605f
C4838 left_shifter_0.S3.t6 VSS 0.064593f
C4839 left_shifter_0.S3.n1 VSS 0.333023f
C4840 left_shifter_0.S3.t1 VSS 0.031825f
C4841 left_shifter_0.S3.t2 VSS 0.031825f
C4842 left_shifter_0.S3.n2 VSS 0.070996f
C4843 left_shifter_0.S3.t3 VSS 0.115514f
C4844 left_shifter_0.S3.t0 VSS 0.091795f
C4845 mux8_4.A6 VSS 5.28232f
C4846 a_n12416_n11063.n0 VSS 1.48365f
C4847 a_n12416_n11063.n1 VSS 1.48326f
C4848 a_n12416_n11063.t8 VSS 0.093341f
C4849 a_n12416_n11063.t9 VSS 0.093341f
C4850 a_n12416_n11063.t10 VSS 0.093341f
C4851 a_n12416_n11063.n2 VSS 0.202296f
C4852 a_n12416_n11063.t11 VSS 0.093341f
C4853 a_n12416_n11063.t3 VSS 0.093341f
C4854 a_n12416_n11063.n3 VSS 0.202001f
C4855 a_n12416_n11063.t4 VSS 0.093341f
C4856 a_n12416_n11063.t5 VSS 0.093341f
C4857 a_n12416_n11063.n4 VSS 0.202001f
C4858 a_n12416_n11063.t1 VSS 0.093341f
C4859 a_n12416_n11063.t0 VSS 0.093341f
C4860 a_n12416_n11063.n5 VSS 0.202001f
C4861 a_n12416_n11063.t6 VSS 0.093341f
C4862 a_n12416_n11063.t7 VSS 0.093341f
C4863 a_n12416_n11063.n6 VSS 0.20269f
C4864 a_n12416_n11063.n7 VSS 0.202001f
C4865 a_n12416_n11063.t2 VSS 0.093341f
C4866 mux8_5.NAND4F_4.Y.n0 VSS 0.480308f
C4867 mux8_5.NAND4F_4.Y.t6 VSS 0.023681f
C4868 mux8_5.NAND4F_4.Y.t5 VSS 0.023681f
C4869 mux8_5.NAND4F_4.Y.n1 VSS 0.054989f
C4870 mux8_5.NAND4F_4.Y.t7 VSS 0.023681f
C4871 mux8_5.NAND4F_4.Y.t8 VSS 0.023681f
C4872 mux8_5.NAND4F_4.Y.n2 VSS 0.054824f
C4873 mux8_5.NAND4F_4.Y.t4 VSS 0.023681f
C4874 mux8_5.NAND4F_4.Y.t3 VSS 0.023681f
C4875 mux8_5.NAND4F_4.Y.n3 VSS 0.054824f
C4876 mux8_5.NAND4F_4.Y.t2 VSS 0.023681f
C4877 mux8_5.NAND4F_4.Y.t1 VSS 0.023681f
C4878 mux8_5.NAND4F_4.Y.n4 VSS 0.054824f
C4879 mux8_5.NAND4F_4.Y.n5 VSS 0.238711f
C4880 mux8_5.NAND4F_4.Y.t9 VSS 0.032831f
C4881 mux8_5.NAND4F_4.Y.t10 VSS 0.031942f
C4882 mux8_5.NAND4F_4.Y.t11 VSS 0.096729f
C4883 mux8_5.NAND4F_4.Y.n6 VSS 0.164667f
C4884 mux8_5.NAND4F_4.Y.t0 VSS 0.190137f
C4885 mux8_5.NAND4F_4.Y.n7 VSS 1.51729f
C4886 AND8_0.S7.n0 VSS 2.50819f
C4887 AND8_0.S7.t4 VSS 0.121112f
C4888 AND8_0.S7.t5 VSS 0.117834f
C4889 AND8_0.S7.t6 VSS 0.356832f
C4890 AND8_0.S7.n1 VSS 0.607468f
C4891 AND8_0.S7.n2 VSS 17.050098f
C4892 AND8_0.S7.t2 VSS 0.058058f
C4893 AND8_0.S7.t3 VSS 0.058058f
C4894 AND8_0.S7.n3 VSS 0.129378f
C4895 AND8_0.S7.t1 VSS 0.210575f
C4896 AND8_0.S7.t0 VSS 0.167458f
C4897 AND8_0.S5.n0 VSS 2.88069f
C4898 AND8_0.S5.t5 VSS 0.139371f
C4899 AND8_0.S5.t6 VSS 0.135599f
C4900 AND8_0.S5.t4 VSS 0.410627f
C4901 AND8_0.S5.n1 VSS 0.699049f
C4902 AND8_0.S5.t2 VSS 0.06681f
C4903 AND8_0.S5.t3 VSS 0.06681f
C4904 AND8_0.S5.n2 VSS 0.148883f
C4905 AND8_0.S5.t1 VSS 0.242321f
C4906 AND8_0.S5.t0 VSS 0.192703f
C4907 mux8_5.NAND4F_4.B.n0 VSS 0.921489f
C4908 mux8_5.NAND4F_4.B.t5 VSS 0.03989f
C4909 mux8_5.NAND4F_4.B.t9 VSS 0.123086f
C4910 mux8_5.NAND4F_4.B.t4 VSS 0.04595f
C4911 mux8_5.NAND4F_4.B.n1 VSS 0.154452f
C4912 mux8_5.NAND4F_4.B.n2 VSS 0.033769f
C4913 mux8_5.NAND4F_4.B.t14 VSS 0.03989f
C4914 mux8_5.NAND4F_4.B.t15 VSS 0.123086f
C4915 mux8_5.NAND4F_4.B.t12 VSS 0.04595f
C4916 mux8_5.NAND4F_4.B.n3 VSS 0.154452f
C4917 mux8_5.NAND4F_4.B.n4 VSS 0.032977f
C4918 mux8_5.NAND4F_4.B.t8 VSS 0.03989f
C4919 mux8_5.NAND4F_4.B.t10 VSS 0.123086f
C4920 mux8_5.NAND4F_4.B.t7 VSS 0.04595f
C4921 mux8_5.NAND4F_4.B.n5 VSS 0.154452f
C4922 mux8_5.NAND4F_4.B.n6 VSS 0.033699f
C4923 mux8_5.NAND4F_4.B.n7 VSS 0.612655f
C4924 mux8_5.NAND4F_4.B.t3 VSS 0.020325f
C4925 mux8_5.NAND4F_4.B.t2 VSS 0.020325f
C4926 mux8_5.NAND4F_4.B.n8 VSS 0.045293f
C4927 mux8_5.NAND4F_4.B.t1 VSS 0.073718f
C4928 mux8_5.NAND4F_4.B.t0 VSS 0.058624f
C4929 mux8_5.NAND4F_4.B.n9 VSS 0.607515f
C4930 mux8_5.NAND4F_4.B.t13 VSS 0.03989f
C4931 mux8_5.NAND4F_4.B.t6 VSS 0.123086f
C4932 mux8_5.NAND4F_4.B.t11 VSS 0.04595f
C4933 mux8_5.NAND4F_4.B.n10 VSS 0.154452f
C4934 mux8_5.NAND4F_4.B.n11 VSS 0.033659f
C4935 mux8_5.NAND4F_4.B.n12 VSS 0.776456f
C4936 a_n13975_n4534.n0 VSS 1.48326f
C4937 a_n13975_n4534.n1 VSS 1.48365f
C4938 a_n13975_n4534.t1 VSS 0.093341f
C4939 a_n13975_n4534.t9 VSS 0.093341f
C4940 a_n13975_n4534.t10 VSS 0.093341f
C4941 a_n13975_n4534.n2 VSS 0.20269f
C4942 a_n13975_n4534.t8 VSS 0.093341f
C4943 a_n13975_n4534.t11 VSS 0.093341f
C4944 a_n13975_n4534.n3 VSS 0.202001f
C4945 a_n13975_n4534.t7 VSS 0.093341f
C4946 a_n13975_n4534.t6 VSS 0.093341f
C4947 a_n13975_n4534.n4 VSS 0.202001f
C4948 a_n13975_n4534.t4 VSS 0.093341f
C4949 a_n13975_n4534.t3 VSS 0.093341f
C4950 a_n13975_n4534.n5 VSS 0.202001f
C4951 a_n13975_n4534.t0 VSS 0.093341f
C4952 a_n13975_n4534.t5 VSS 0.093341f
C4953 a_n13975_n4534.n6 VSS 0.202001f
C4954 a_n13975_n4534.n7 VSS 0.202296f
C4955 a_n13975_n4534.t2 VSS 0.093341f
C4956 MULT_0.inv_12.A.n0 VSS 1.18962f
C4957 MULT_0.inv_12.A.n1 VSS 0.18714f
C4958 MULT_0.inv_12.A.t3 VSS 0.138862f
C4959 MULT_0.inv_12.A.t6 VSS 0.023051f
C4960 MULT_0.inv_12.A.t5 VSS 0.023051f
C4961 MULT_0.inv_12.A.n2 VSS 0.051291f
C4962 MULT_0.inv_12.A.t1 VSS 0.023051f
C4963 MULT_0.inv_12.A.t0 VSS 0.023051f
C4964 MULT_0.inv_12.A.n3 VSS 0.051431f
C4965 MULT_0.inv_12.A.t4 VSS 0.023051f
C4966 MULT_0.inv_12.A.t2 VSS 0.023051f
C4967 MULT_0.inv_12.A.n4 VSS 0.051291f
C4968 MULT_0.inv_12.A.t9 VSS 0.029376f
C4969 MULT_0.inv_12.A.t8 VSS 0.041007f
C4970 MULT_0.inv_12.A.t10 VSS 0.041007f
C4971 MULT_0.inv_12.A.n5 VSS 0.133851f
C4972 MULT_0.inv_12.A.t7 VSS 0.04682f
C4973 left_shifter_0.C.n0 VSS 2.30077f
C4974 mux8_0.NAND4F_5.A VSS 0.146325f
C4975 left_shifter_0.C.t4 VSS 0.012046f
C4976 left_shifter_0.C.t6 VSS 0.035491f
C4977 left_shifter_0.C.t5 VSS 0.01172f
C4978 left_shifter_0.C.n1 VSS 0.060425f
C4979 left_shifter_0.C.t3 VSS 0.005775f
C4980 left_shifter_0.C.t2 VSS 0.005775f
C4981 left_shifter_0.C.n2 VSS 0.012882f
C4982 left_shifter_0.C.t0 VSS 0.020959f
C4983 left_shifter_0.C.t1 VSS 0.016656f
C4984 mux8_0.A6 VSS 2.47118f
C4985 MULT_0.S2.t12 VSS 0.065621f
C4986 MULT_0.S2.t14 VSS 0.063845f
C4987 MULT_0.S2.t13 VSS 0.193338f
C4988 MULT_0.S2.n0 VSS 0.329164f
C4989 MULT_0.S2.t11 VSS 0.019109f
C4990 MULT_0.S2.t10 VSS 0.019109f
C4991 MULT_0.S2.n1 VSS 0.046218f
C4992 MULT_0.S2.t8 VSS 0.019109f
C4993 MULT_0.S2.t4 VSS 0.019109f
C4994 MULT_0.S2.n2 VSS 0.046213f
C4995 MULT_0.S2.n3 VSS 0.331387f
C4996 MULT_0.S2.t9 VSS 0.019109f
C4997 MULT_0.S2.t7 VSS 0.019109f
C4998 MULT_0.S2.n4 VSS 0.038218f
C4999 MULT_0.S2.n5 VSS 0.030022f
C5000 MULT_0.S2.t2 VSS 0.080847f
C5001 MULT_0.S2.t3 VSS 0.080847f
C5002 MULT_0.S2.n6 VSS 0.161694f
C5003 MULT_0.S2.n7 VSS 0.064292f
C5004 MULT_0.S2.t1 VSS 0.080847f
C5005 MULT_0.S2.t0 VSS 0.080847f
C5006 MULT_0.S2.n8 VSS 0.161694f
C5007 MULT_0.S2.n9 VSS 0.071116f
C5008 MULT_0.S2.n10 VSS 0.732175f
C5009 MULT_0.S2.t5 VSS 0.080847f
C5010 MULT_0.S2.t6 VSS 0.080847f
C5011 MULT_0.S2.n11 VSS 0.161694f
C5012 MULT_0.S2.n12 VSS 0.071223f
C5013 MULT_0.S2.n13 VSS 0.469585f
C5014 MULT_0.S2.n14 VSS 0.105826f
C5015 MULT_0.S2.n15 VSS 0.464494f
C5016 a_n10684_n7799.n0 VSS 1.48326f
C5017 a_n10684_n7799.n1 VSS 1.48365f
C5018 a_n10684_n7799.t1 VSS 0.093341f
C5019 a_n10684_n7799.t10 VSS 0.093341f
C5020 a_n10684_n7799.t9 VSS 0.093341f
C5021 a_n10684_n7799.n2 VSS 0.202296f
C5022 a_n10684_n7799.t11 VSS 0.093341f
C5023 a_n10684_n7799.t2 VSS 0.093341f
C5024 a_n10684_n7799.n3 VSS 0.202001f
C5025 a_n10684_n7799.t6 VSS 0.093341f
C5026 a_n10684_n7799.t5 VSS 0.093341f
C5027 a_n10684_n7799.n4 VSS 0.20269f
C5028 a_n10684_n7799.t8 VSS 0.093341f
C5029 a_n10684_n7799.t4 VSS 0.093341f
C5030 a_n10684_n7799.n5 VSS 0.202001f
C5031 a_n10684_n7799.t0 VSS 0.093341f
C5032 a_n10684_n7799.t7 VSS 0.093341f
C5033 a_n10684_n7799.n6 VSS 0.202001f
C5034 a_n10684_n7799.n7 VSS 0.202001f
C5035 a_n10684_n7799.t3 VSS 0.093341f
C5036 a_n18998_n4534.n0 VSS 1.48365f
C5037 a_n18998_n4534.n1 VSS 1.48326f
C5038 a_n18998_n4534.t0 VSS 0.093341f
C5039 a_n18998_n4534.t6 VSS 0.093341f
C5040 a_n18998_n4534.t8 VSS 0.093341f
C5041 a_n18998_n4534.n2 VSS 0.202296f
C5042 a_n18998_n4534.t7 VSS 0.093341f
C5043 a_n18998_n4534.t9 VSS 0.093341f
C5044 a_n18998_n4534.n3 VSS 0.202001f
C5045 a_n18998_n4534.t10 VSS 0.093341f
C5046 a_n18998_n4534.t11 VSS 0.093341f
C5047 a_n18998_n4534.n4 VSS 0.202001f
C5048 a_n18998_n4534.t5 VSS 0.093341f
C5049 a_n18998_n4534.t4 VSS 0.093341f
C5050 a_n18998_n4534.n5 VSS 0.202001f
C5051 a_n18998_n4534.t3 VSS 0.093341f
C5052 a_n18998_n4534.t1 VSS 0.093341f
C5053 a_n18998_n4534.n6 VSS 0.202001f
C5054 a_n18998_n4534.n7 VSS 0.20269f
C5055 a_n18998_n4534.t2 VSS 0.093341f
C5056 mux8_6.NAND4F_0.Y.n0 VSS 0.350455f
C5057 mux8_6.NAND4F_0.Y.t10 VSS 0.022537f
C5058 mux8_6.NAND4F_0.Y.t9 VSS 0.079785f
C5059 mux8_6.NAND4F_0.Y.t11 VSS 0.024808f
C5060 mux8_6.NAND4F_0.Y.n1 VSS 0.070768f
C5061 mux8_6.NAND4F_0.Y.n2 VSS 0.020978f
C5062 mux8_6.NAND4F_0.Y.t1 VSS 0.017278f
C5063 mux8_6.NAND4F_0.Y.t0 VSS 0.017278f
C5064 mux8_6.NAND4F_0.Y.n3 VSS 0.040122f
C5065 mux8_6.NAND4F_0.Y.t3 VSS 0.017278f
C5066 mux8_6.NAND4F_0.Y.t2 VSS 0.017278f
C5067 mux8_6.NAND4F_0.Y.n4 VSS 0.040002f
C5068 mux8_6.NAND4F_0.Y.t8 VSS 0.017278f
C5069 mux8_6.NAND4F_0.Y.t7 VSS 0.017278f
C5070 mux8_6.NAND4F_0.Y.n5 VSS 0.040002f
C5071 mux8_6.NAND4F_0.Y.t6 VSS 0.017278f
C5072 mux8_6.NAND4F_0.Y.t5 VSS 0.017278f
C5073 mux8_6.NAND4F_0.Y.n6 VSS 0.040002f
C5074 mux8_6.NAND4F_0.Y.t4 VSS 0.166327f
C5075 Y2.t7 VSS 0.060228f
C5076 Y2.t5 VSS 0.129299f
C5077 Y2.t6 VSS 0.139704f
C5078 Y2.n0 VSS 0.110363f
C5079 Y2.t4 VSS 0.130039f
C5080 Y2.n1 VSS 0.062532f
C5081 Y2.n2 VSS 0.064234f
C5082 Y2.t3 VSS 0.024195f
C5083 Y2.t2 VSS 0.024195f
C5084 Y2.n3 VSS 0.053904f
C5085 Y2.t0 VSS 0.069885f
C5086 Y2.n4 VSS 0.292627f
C5087 Y2.t1 VSS 0.087754f
C5088 Y2.n5 VSS 0.12655f
C5089 MULT_0.NAND2_8.Y.n0 VSS 1.19272f
C5090 MULT_0.NAND2_8.Y.n1 VSS 0.186498f
C5091 MULT_0.NAND2_8.Y.t4 VSS 0.022972f
C5092 MULT_0.NAND2_8.Y.t6 VSS 0.022972f
C5093 MULT_0.NAND2_8.Y.n2 VSS 0.051117f
C5094 MULT_0.NAND2_8.Y.t1 VSS 0.022972f
C5095 MULT_0.NAND2_8.Y.t2 VSS 0.022972f
C5096 MULT_0.NAND2_8.Y.n3 VSS 0.051256f
C5097 MULT_0.NAND2_8.Y.t5 VSS 0.022972f
C5098 MULT_0.NAND2_8.Y.t0 VSS 0.022972f
C5099 MULT_0.NAND2_8.Y.n4 VSS 0.051117f
C5100 MULT_0.NAND2_8.Y.t3 VSS 0.13839f
C5101 MULT_0.NAND2_8.Y.t9 VSS 0.029277f
C5102 MULT_0.NAND2_8.Y.t7 VSS 0.040868f
C5103 MULT_0.NAND2_8.Y.t10 VSS 0.040868f
C5104 MULT_0.NAND2_8.Y.n5 VSS 0.133396f
C5105 MULT_0.NAND2_8.Y.t8 VSS 0.046661f
C5106 mux8_7.NAND4F_4.Y.n0 VSS 0.480308f
C5107 mux8_7.NAND4F_4.Y.t4 VSS 0.023681f
C5108 mux8_7.NAND4F_4.Y.t3 VSS 0.023681f
C5109 mux8_7.NAND4F_4.Y.n1 VSS 0.054989f
C5110 mux8_7.NAND4F_4.Y.t6 VSS 0.023681f
C5111 mux8_7.NAND4F_4.Y.t5 VSS 0.023681f
C5112 mux8_7.NAND4F_4.Y.n2 VSS 0.054824f
C5113 mux8_7.NAND4F_4.Y.t8 VSS 0.023681f
C5114 mux8_7.NAND4F_4.Y.t7 VSS 0.023681f
C5115 mux8_7.NAND4F_4.Y.n3 VSS 0.054824f
C5116 mux8_7.NAND4F_4.Y.t1 VSS 0.023681f
C5117 mux8_7.NAND4F_4.Y.t2 VSS 0.023681f
C5118 mux8_7.NAND4F_4.Y.n4 VSS 0.054824f
C5119 mux8_7.NAND4F_4.Y.n5 VSS 0.238711f
C5120 mux8_7.NAND4F_4.Y.t9 VSS 0.032831f
C5121 mux8_7.NAND4F_4.Y.t10 VSS 0.031942f
C5122 mux8_7.NAND4F_4.Y.t11 VSS 0.096729f
C5123 mux8_7.NAND4F_4.Y.n6 VSS 0.164667f
C5124 mux8_7.NAND4F_4.Y.t0 VSS 0.190137f
C5125 mux8_7.NAND4F_4.Y.n7 VSS 1.51729f
C5126 ZFLAG_0.NAND2_0.Y.n0 VSS 1.14261f
C5127 ZFLAG_0.NAND2_0.Y.n1 VSS 0.195221f
C5128 ZFLAG_0.NAND2_0.Y.t4 VSS 0.146393f
C5129 ZFLAG_0.NAND2_0.Y.t9 VSS 0.03097f
C5130 ZFLAG_0.NAND2_0.Y.t7 VSS 0.043231f
C5131 ZFLAG_0.NAND2_0.Y.t10 VSS 0.043231f
C5132 ZFLAG_0.NAND2_0.Y.n2 VSS 0.140768f
C5133 ZFLAG_0.NAND2_0.Y.t3 VSS 0.024301f
C5134 ZFLAG_0.NAND2_0.Y.t5 VSS 0.024301f
C5135 ZFLAG_0.NAND2_0.Y.n3 VSS 0.054073f
C5136 ZFLAG_0.NAND2_0.Y.t2 VSS 0.024301f
C5137 ZFLAG_0.NAND2_0.Y.t1 VSS 0.024301f
C5138 ZFLAG_0.NAND2_0.Y.n4 VSS 0.05422f
C5139 ZFLAG_0.NAND2_0.Y.t6 VSS 0.024301f
C5140 ZFLAG_0.NAND2_0.Y.t0 VSS 0.024301f
C5141 ZFLAG_0.NAND2_0.Y.n5 VSS 0.054073f
C5142 ZFLAG_0.NAND2_0.Y.t8 VSS 0.049404f
C5143 MULT_0.NAND2_0.Y.n0 VSS 1.19733f
C5144 MULT_0.NAND2_0.Y.n1 VSS 0.185543f
C5145 MULT_0.NAND2_0.Y.t5 VSS 0.022856f
C5146 MULT_0.NAND2_0.Y.t6 VSS 0.022856f
C5147 MULT_0.NAND2_0.Y.n2 VSS 0.050858f
C5148 MULT_0.NAND2_0.Y.t1 VSS 0.022856f
C5149 MULT_0.NAND2_0.Y.t0 VSS 0.022856f
C5150 MULT_0.NAND2_0.Y.n3 VSS 0.050996f
C5151 MULT_0.NAND2_0.Y.t4 VSS 0.022856f
C5152 MULT_0.NAND2_0.Y.t2 VSS 0.022856f
C5153 MULT_0.NAND2_0.Y.n4 VSS 0.050858f
C5154 MULT_0.NAND2_0.Y.t3 VSS 0.137689f
C5155 MULT_0.NAND2_0.Y.t10 VSS 0.029128f
C5156 MULT_0.NAND2_0.Y.t9 VSS 0.040661f
C5157 MULT_0.NAND2_0.Y.t7 VSS 0.040661f
C5158 MULT_0.NAND2_0.Y.n5 VSS 0.132719f
C5159 MULT_0.NAND2_0.Y.t8 VSS 0.046425f
C5160 mux8_6.NAND4F_3.Y.n0 VSS 0.306333f
C5161 mux8_6.NAND4F_3.Y.t1 VSS 0.015103f
C5162 mux8_6.NAND4F_3.Y.t0 VSS 0.015103f
C5163 mux8_6.NAND4F_3.Y.n1 VSS 0.035071f
C5164 mux8_6.NAND4F_3.Y.t3 VSS 0.015103f
C5165 mux8_6.NAND4F_3.Y.t2 VSS 0.015103f
C5166 mux8_6.NAND4F_3.Y.n2 VSS 0.034966f
C5167 mux8_6.NAND4F_3.Y.t5 VSS 0.015103f
C5168 mux8_6.NAND4F_3.Y.t4 VSS 0.015103f
C5169 mux8_6.NAND4F_3.Y.n3 VSS 0.034966f
C5170 mux8_6.NAND4F_3.Y.t7 VSS 0.015103f
C5171 mux8_6.NAND4F_3.Y.t8 VSS 0.015103f
C5172 mux8_6.NAND4F_3.Y.n4 VSS 0.034966f
C5173 mux8_6.NAND4F_3.Y.n5 VSS 0.152246f
C5174 mux8_6.NAND4F_3.Y.t6 VSS 0.143521f
C5175 mux8_6.NAND4F_3.Y.t10 VSS 0.0197f
C5176 mux8_6.NAND4F_3.Y.t11 VSS 0.0197f
C5177 mux8_6.NAND4F_3.Y.n6 VSS 0.023128f
C5178 mux8_6.NAND4F_3.Y.t9 VSS 0.061756f
C5179 mux8_6.NAND4F_3.Y.n7 VSS 0.129679f
C5180 mux8_3.NAND4F_0.Y.n0 VSS 0.350455f
C5181 mux8_3.NAND4F_0.Y.t10 VSS 0.022537f
C5182 mux8_3.NAND4F_0.Y.t9 VSS 0.079785f
C5183 mux8_3.NAND4F_0.Y.t11 VSS 0.024808f
C5184 mux8_3.NAND4F_0.Y.n1 VSS 0.070768f
C5185 mux8_3.NAND4F_0.Y.n2 VSS 0.020978f
C5186 mux8_3.NAND4F_0.Y.t4 VSS 0.017278f
C5187 mux8_3.NAND4F_0.Y.t3 VSS 0.017278f
C5188 mux8_3.NAND4F_0.Y.n3 VSS 0.040122f
C5189 mux8_3.NAND4F_0.Y.t6 VSS 0.017278f
C5190 mux8_3.NAND4F_0.Y.t5 VSS 0.017278f
C5191 mux8_3.NAND4F_0.Y.n4 VSS 0.040002f
C5192 mux8_3.NAND4F_0.Y.t8 VSS 0.017278f
C5193 mux8_3.NAND4F_0.Y.t7 VSS 0.017278f
C5194 mux8_3.NAND4F_0.Y.n5 VSS 0.040002f
C5195 mux8_3.NAND4F_0.Y.t0 VSS 0.017278f
C5196 mux8_3.NAND4F_0.Y.t2 VSS 0.017278f
C5197 mux8_3.NAND4F_0.Y.n6 VSS 0.040002f
C5198 mux8_3.NAND4F_0.Y.t1 VSS 0.166327f
C5199 AND8_0.S2.n0 VSS 3.01106f
C5200 AND8_0.S2.t4 VSS 0.14577f
C5201 AND8_0.S2.t5 VSS 0.141825f
C5202 AND8_0.S2.t6 VSS 0.429481f
C5203 AND8_0.S2.n1 VSS 0.731146f
C5204 AND8_0.S2.t2 VSS 0.069878f
C5205 AND8_0.S2.t3 VSS 0.069878f
C5206 AND8_0.S2.n2 VSS 0.155719f
C5207 AND8_0.S2.t1 VSS 0.253447f
C5208 AND8_0.S2.t0 VSS 0.201551f
C5209 MULT_0.NAND2_10.Y.n0 VSS 1.19348f
C5210 MULT_0.NAND2_10.Y.n1 VSS 0.186339f
C5211 MULT_0.NAND2_10.Y.t5 VSS 0.022953f
C5212 MULT_0.NAND2_10.Y.t4 VSS 0.022953f
C5213 MULT_0.NAND2_10.Y.n2 VSS 0.051074f
C5214 MULT_0.NAND2_10.Y.t1 VSS 0.022953f
C5215 MULT_0.NAND2_10.Y.t0 VSS 0.022953f
C5216 MULT_0.NAND2_10.Y.n3 VSS 0.051213f
C5217 MULT_0.NAND2_10.Y.t6 VSS 0.022953f
C5218 MULT_0.NAND2_10.Y.t2 VSS 0.022953f
C5219 MULT_0.NAND2_10.Y.n4 VSS 0.051074f
C5220 MULT_0.NAND2_10.Y.t3 VSS 0.138274f
C5221 MULT_0.NAND2_10.Y.t9 VSS 0.029252f
C5222 MULT_0.NAND2_10.Y.t8 VSS 0.040833f
C5223 MULT_0.NAND2_10.Y.t10 VSS 0.040833f
C5224 MULT_0.NAND2_10.Y.n5 VSS 0.133283f
C5225 MULT_0.NAND2_10.Y.t7 VSS 0.046622f
C5226 a_n12314_n21072.n0 VSS 1.48326f
C5227 a_n12314_n21072.n1 VSS 1.48365f
C5228 a_n12314_n21072.t1 VSS 0.093341f
C5229 a_n12314_n21072.t4 VSS 0.093341f
C5230 a_n12314_n21072.t3 VSS 0.093341f
C5231 a_n12314_n21072.n2 VSS 0.20269f
C5232 a_n12314_n21072.t11 VSS 0.093341f
C5233 a_n12314_n21072.t5 VSS 0.093341f
C5234 a_n12314_n21072.n3 VSS 0.202001f
C5235 a_n12314_n21072.t9 VSS 0.093341f
C5236 a_n12314_n21072.t10 VSS 0.093341f
C5237 a_n12314_n21072.n4 VSS 0.202001f
C5238 a_n12314_n21072.t7 VSS 0.093341f
C5239 a_n12314_n21072.t6 VSS 0.093341f
C5240 a_n12314_n21072.n5 VSS 0.202001f
C5241 a_n12314_n21072.t0 VSS 0.093341f
C5242 a_n12314_n21072.t8 VSS 0.093341f
C5243 a_n12314_n21072.n6 VSS 0.202001f
C5244 a_n12314_n21072.n7 VSS 0.202296f
C5245 a_n12314_n21072.t2 VSS 0.093341f
C5246 XOR8_0.S2.t14 VSS 0.069371f
C5247 XOR8_0.S2.t13 VSS 0.204388f
C5248 XOR8_0.S2.t12 VSS 0.067494f
C5249 XOR8_0.S2.n0 VSS 0.347956f
C5250 XOR8_0.S2.t0 VSS 0.020201f
C5251 XOR8_0.S2.t1 VSS 0.020201f
C5252 XOR8_0.S2.n1 VSS 0.04886f
C5253 XOR8_0.S2.t10 VSS 0.020201f
C5254 XOR8_0.S2.t11 VSS 0.020201f
C5255 XOR8_0.S2.n2 VSS 0.048854f
C5256 XOR8_0.S2.n3 VSS 0.350327f
C5257 XOR8_0.S2.t2 VSS 0.020201f
C5258 XOR8_0.S2.t9 VSS 0.020201f
C5259 XOR8_0.S2.n4 VSS 0.040403f
C5260 XOR8_0.S2.n5 VSS 0.031738f
C5261 XOR8_0.S2.t3 VSS 0.085467f
C5262 XOR8_0.S2.t6 VSS 0.085467f
C5263 XOR8_0.S2.n6 VSS 0.170935f
C5264 XOR8_0.S2.n7 VSS 0.067806f
C5265 XOR8_0.S2.t5 VSS 0.085467f
C5266 XOR8_0.S2.t4 VSS 0.085467f
C5267 XOR8_0.S2.n8 VSS 0.170935f
C5268 XOR8_0.S2.n9 VSS 0.07518f
C5269 XOR8_0.S2.n10 VSS 0.774021f
C5270 XOR8_0.S2.t7 VSS 0.085467f
C5271 XOR8_0.S2.t8 VSS 0.085467f
C5272 XOR8_0.S2.n11 VSS 0.170935f
C5273 XOR8_0.S2.n12 VSS 0.075294f
C5274 XOR8_0.S2.n13 VSS 0.496424f
C5275 XOR8_0.S2.n14 VSS 0.111738f
C5276 XOR8_0.S2.n15 VSS 0.491338f
C5277 XOR8_0.S5.t12 VSS 0.063165f
C5278 XOR8_0.S5.t14 VSS 0.186101f
C5279 XOR8_0.S5.t13 VSS 0.061455f
C5280 XOR8_0.S5.n0 VSS 0.316823f
C5281 XOR8_0.S5.t2 VSS 0.018394f
C5282 XOR8_0.S5.t1 VSS 0.018394f
C5283 XOR8_0.S5.n1 VSS 0.044488f
C5284 XOR8_0.S5.t0 VSS 0.018394f
C5285 XOR8_0.S5.t4 VSS 0.018394f
C5286 XOR8_0.S5.n2 VSS 0.044483f
C5287 XOR8_0.S5.n3 VSS 0.318983f
C5288 XOR8_0.S5.t3 VSS 0.018394f
C5289 XOR8_0.S5.t10 VSS 0.018394f
C5290 XOR8_0.S5.n4 VSS 0.036788f
C5291 XOR8_0.S5.n5 VSS 0.028898f
C5292 XOR8_0.S5.t6 VSS 0.077821f
C5293 XOR8_0.S5.t11 VSS 0.077821f
C5294 XOR8_0.S5.n6 VSS 0.155641f
C5295 XOR8_0.S5.n7 VSS 0.06174f
C5296 XOR8_0.S5.t8 VSS 0.077821f
C5297 XOR8_0.S5.t7 VSS 0.077821f
C5298 XOR8_0.S5.n8 VSS 0.155641f
C5299 XOR8_0.S5.n9 VSS 0.068454f
C5300 XOR8_0.S5.n10 VSS 0.704769f
C5301 XOR8_0.S5.t5 VSS 0.077821f
C5302 XOR8_0.S5.t9 VSS 0.077821f
C5303 XOR8_0.S5.n11 VSS 0.155641f
C5304 XOR8_0.S5.n12 VSS 0.068557f
C5305 XOR8_0.S5.n13 VSS 0.452008f
C5306 XOR8_0.S5.n14 VSS 0.10174f
C5307 XOR8_0.S5.n15 VSS 0.447377f
C5308 mux8_4.NAND4F_4.Y.n0 VSS 0.480308f
C5309 mux8_4.NAND4F_4.Y.t1 VSS 0.023681f
C5310 mux8_4.NAND4F_4.Y.t0 VSS 0.023681f
C5311 mux8_4.NAND4F_4.Y.n1 VSS 0.054989f
C5312 mux8_4.NAND4F_4.Y.t5 VSS 0.023681f
C5313 mux8_4.NAND4F_4.Y.t4 VSS 0.023681f
C5314 mux8_4.NAND4F_4.Y.n2 VSS 0.054824f
C5315 mux8_4.NAND4F_4.Y.t3 VSS 0.023681f
C5316 mux8_4.NAND4F_4.Y.t2 VSS 0.023681f
C5317 mux8_4.NAND4F_4.Y.n3 VSS 0.054824f
C5318 mux8_4.NAND4F_4.Y.t7 VSS 0.023681f
C5319 mux8_4.NAND4F_4.Y.t6 VSS 0.023681f
C5320 mux8_4.NAND4F_4.Y.n4 VSS 0.054824f
C5321 mux8_4.NAND4F_4.Y.n5 VSS 0.238711f
C5322 mux8_4.NAND4F_4.Y.t9 VSS 0.032831f
C5323 mux8_4.NAND4F_4.Y.t10 VSS 0.031942f
C5324 mux8_4.NAND4F_4.Y.t11 VSS 0.096729f
C5325 mux8_4.NAND4F_4.Y.n6 VSS 0.164667f
C5326 mux8_4.NAND4F_4.Y.t8 VSS 0.190137f
C5327 mux8_4.NAND4F_4.Y.n7 VSS 1.51729f
C5328 mux8_3.NAND4F_3.Y.n0 VSS 0.306333f
C5329 mux8_3.NAND4F_3.Y.t4 VSS 0.015103f
C5330 mux8_3.NAND4F_3.Y.t3 VSS 0.015103f
C5331 mux8_3.NAND4F_3.Y.n1 VSS 0.035071f
C5332 mux8_3.NAND4F_3.Y.t8 VSS 0.015103f
C5333 mux8_3.NAND4F_3.Y.t7 VSS 0.015103f
C5334 mux8_3.NAND4F_3.Y.n2 VSS 0.034966f
C5335 mux8_3.NAND4F_3.Y.t6 VSS 0.015103f
C5336 mux8_3.NAND4F_3.Y.t5 VSS 0.015103f
C5337 mux8_3.NAND4F_3.Y.n3 VSS 0.034966f
C5338 mux8_3.NAND4F_3.Y.t1 VSS 0.015103f
C5339 mux8_3.NAND4F_3.Y.t2 VSS 0.015103f
C5340 mux8_3.NAND4F_3.Y.n4 VSS 0.034966f
C5341 mux8_3.NAND4F_3.Y.n5 VSS 0.152246f
C5342 mux8_3.NAND4F_3.Y.t0 VSS 0.143521f
C5343 mux8_3.NAND4F_3.Y.t10 VSS 0.0197f
C5344 mux8_3.NAND4F_3.Y.t11 VSS 0.0197f
C5345 mux8_3.NAND4F_3.Y.n6 VSS 0.023128f
C5346 mux8_3.NAND4F_3.Y.t9 VSS 0.061756f
C5347 mux8_3.NAND4F_3.Y.n7 VSS 0.129679f
C5348 mux8_3.NAND4F_2.D.n0 VSS 0.664607f
C5349 mux8_3.NAND4F_2.D.t14 VSS 0.027742f
C5350 mux8_3.NAND4F_2.D.t5 VSS 0.098211f
C5351 mux8_3.NAND4F_2.D.t13 VSS 0.030538f
C5352 mux8_3.NAND4F_2.D.n1 VSS 0.087112f
C5353 mux8_3.NAND4F_2.D.n2 VSS 0.025808f
C5354 mux8_3.NAND4F_2.D.t3 VSS 0.014135f
C5355 mux8_3.NAND4F_2.D.t2 VSS 0.014135f
C5356 mux8_3.NAND4F_2.D.n3 VSS 0.031499f
C5357 mux8_3.NAND4F_2.D.t1 VSS 0.051268f
C5358 mux8_3.NAND4F_2.D.t0 VSS 0.040771f
C5359 mux8_3.NAND4F_2.D.t11 VSS 0.027742f
C5360 mux8_3.NAND4F_2.D.t15 VSS 0.098211f
C5361 mux8_3.NAND4F_2.D.t6 VSS 0.030538f
C5362 mux8_3.NAND4F_2.D.n4 VSS 0.087112f
C5363 mux8_3.NAND4F_2.D.n5 VSS 0.025813f
C5364 mux8_3.NAND4F_2.D.n6 VSS 0.620222f
C5365 mux8_3.NAND4F_2.D.t10 VSS 0.027742f
C5366 mux8_3.NAND4F_2.D.t8 VSS 0.098211f
C5367 mux8_3.NAND4F_2.D.t9 VSS 0.030538f
C5368 mux8_3.NAND4F_2.D.n7 VSS 0.087112f
C5369 mux8_3.NAND4F_2.D.n8 VSS 0.025807f
C5370 mux8_3.NAND4F_2.D.n9 VSS 0.261852f
C5371 mux8_3.NAND4F_2.D.t7 VSS 0.027742f
C5372 mux8_3.NAND4F_2.D.t12 VSS 0.098211f
C5373 mux8_3.NAND4F_2.D.t4 VSS 0.030538f
C5374 mux8_3.NAND4F_2.D.n10 VSS 0.087112f
C5375 mux8_3.NAND4F_2.D.n11 VSS 0.025808f
C5376 mux8_3.NAND4F_2.D.n12 VSS 0.407824f
C5377 AND8_0.S6.n0 VSS 2.48442f
C5378 AND8_0.S6.t4 VSS 0.119908f
C5379 AND8_0.S6.t5 VSS 0.116662f
C5380 AND8_0.S6.t6 VSS 0.353283f
C5381 AND8_0.S6.n1 VSS 0.601426f
C5382 AND8_0.S6.t0 VSS 0.05748f
C5383 AND8_0.S6.t2 VSS 0.05748f
C5384 AND8_0.S6.n2 VSS 0.128091f
C5385 AND8_0.S6.t1 VSS 0.20848f
C5386 AND8_0.S6.t3 VSS 0.165792f
C5387 mux8_2.NAND4F_6.Y.n0 VSS 0.599344f
C5388 mux8_2.NAND4F_6.Y.t3 VSS 0.244548f
C5389 mux8_2.NAND4F_6.Y.t9 VSS 0.038543f
C5390 mux8_2.NAND4F_6.Y.t11 VSS 0.118929f
C5391 mux8_2.NAND4F_6.Y.t10 VSS 0.044398f
C5392 mux8_2.NAND4F_6.Y.n1 VSS 0.149236f
C5393 mux8_2.NAND4F_6.Y.n2 VSS 0.032396f
C5394 mux8_2.NAND4F_6.Y.n3 VSS 1.72835f
C5395 mux8_2.NAND4F_6.Y.t0 VSS 0.029549f
C5396 mux8_2.NAND4F_6.Y.t1 VSS 0.029549f
C5397 mux8_2.NAND4F_6.Y.n4 VSS 0.068617f
C5398 mux8_2.NAND4F_6.Y.t6 VSS 0.029549f
C5399 mux8_2.NAND4F_6.Y.t5 VSS 0.029549f
C5400 mux8_2.NAND4F_6.Y.n5 VSS 0.068411f
C5401 mux8_2.NAND4F_6.Y.t7 VSS 0.029549f
C5402 mux8_2.NAND4F_6.Y.t8 VSS 0.029549f
C5403 mux8_2.NAND4F_6.Y.n6 VSS 0.068411f
C5404 mux8_2.NAND4F_6.Y.t4 VSS 0.029549f
C5405 mux8_2.NAND4F_6.Y.t2 VSS 0.029549f
C5406 mux8_2.NAND4F_6.Y.n7 VSS 0.068411f
C5407 mux8_2.NAND4F_6.Y.n8 VSS 0.281208f
C5408 NOT8_0.S2.n0 VSS 2.46464f
C5409 NOT8_0.S2.t6 VSS 0.119236f
C5410 NOT8_0.S2.t5 VSS 0.351304f
C5411 NOT8_0.S2.t4 VSS 0.116009f
C5412 NOT8_0.S2.n1 VSS 0.598106f
C5413 NOT8_0.S2.t1 VSS 0.057158f
C5414 NOT8_0.S2.t3 VSS 0.057158f
C5415 NOT8_0.S2.n2 VSS 0.127373f
C5416 NOT8_0.S2.t2 VSS 0.207312f
C5417 NOT8_0.S2.t0 VSS 0.164863f
C5418 a_n12314_n23651.n0 VSS 1.48365f
C5419 a_n12314_n23651.n1 VSS 1.48326f
C5420 a_n12314_n23651.t1 VSS 0.093341f
C5421 a_n12314_n23651.t3 VSS 0.093341f
C5422 a_n12314_n23651.t5 VSS 0.093341f
C5423 a_n12314_n23651.n2 VSS 0.202296f
C5424 a_n12314_n23651.t4 VSS 0.093341f
C5425 a_n12314_n23651.t11 VSS 0.093341f
C5426 a_n12314_n23651.n3 VSS 0.202001f
C5427 a_n12314_n23651.t10 VSS 0.093341f
C5428 a_n12314_n23651.t9 VSS 0.093341f
C5429 a_n12314_n23651.n4 VSS 0.202001f
C5430 a_n12314_n23651.t8 VSS 0.093341f
C5431 a_n12314_n23651.t7 VSS 0.093341f
C5432 a_n12314_n23651.n5 VSS 0.20269f
C5433 a_n12314_n23651.t0 VSS 0.093341f
C5434 a_n12314_n23651.t6 VSS 0.093341f
C5435 a_n12314_n23651.n6 VSS 0.202001f
C5436 a_n12314_n23651.n7 VSS 0.202001f
C5437 a_n12314_n23651.t2 VSS 0.093341f
C5438 mux8_8.NAND4F_1.Y.n0 VSS 0.655599f
C5439 mux8_8.NAND4F_1.Y.t2 VSS 0.306614f
C5440 mux8_8.NAND4F_1.Y.t11 VSS 0.132168f
C5441 mux8_8.NAND4F_1.Y.t10 VSS 0.04216f
C5442 mux8_8.NAND4F_1.Y.t9 VSS 0.04216f
C5443 mux8_8.NAND4F_1.Y.n1 VSS 0.049498f
C5444 mux8_8.NAND4F_1.Y.n2 VSS 0.277534f
C5445 mux8_8.NAND4F_1.Y.t1 VSS 0.032323f
C5446 mux8_8.NAND4F_1.Y.t0 VSS 0.032323f
C5447 mux8_8.NAND4F_1.Y.n3 VSS 0.075057f
C5448 mux8_8.NAND4F_1.Y.t8 VSS 0.032323f
C5449 mux8_8.NAND4F_1.Y.t7 VSS 0.032323f
C5450 mux8_8.NAND4F_1.Y.n4 VSS 0.074832f
C5451 mux8_8.NAND4F_1.Y.t6 VSS 0.032323f
C5452 mux8_8.NAND4F_1.Y.t5 VSS 0.032323f
C5453 mux8_8.NAND4F_1.Y.n5 VSS 0.074832f
C5454 mux8_8.NAND4F_1.Y.t4 VSS 0.032323f
C5455 mux8_8.NAND4F_1.Y.t3 VSS 0.032323f
C5456 mux8_8.NAND4F_1.Y.n6 VSS 0.074832f
C5457 mux8_8.NAND4F_1.Y.n7 VSS 0.307603f
C5458 left_shifter_0.S5.n0 VSS 7.45182f
C5459 mux8_7.NAND4F_5.A VSS 0.781467f
C5460 left_shifter_0.S5.t5 VSS 0.064334f
C5461 left_shifter_0.S5.t4 VSS 0.189546f
C5462 left_shifter_0.S5.t6 VSS 0.062592f
C5463 left_shifter_0.S5.n1 VSS 0.322708f
C5464 left_shifter_0.S5.t3 VSS 0.03084f
C5465 left_shifter_0.S5.t2 VSS 0.03084f
C5466 left_shifter_0.S5.n2 VSS 0.068797f
C5467 left_shifter_0.S5.t0 VSS 0.111936f
C5468 left_shifter_0.S5.t1 VSS 0.088952f
C5469 mux8_7.A6 VSS 6.99617f
C5470 a_n29_2026.n0 VSS 1.48326f
C5471 a_n29_2026.n1 VSS 1.48365f
C5472 a_n29_2026.t1 VSS 0.093341f
C5473 a_n29_2026.t10 VSS 0.093341f
C5474 a_n29_2026.t8 VSS 0.093341f
C5475 a_n29_2026.n2 VSS 0.20269f
C5476 a_n29_2026.t4 VSS 0.093341f
C5477 a_n29_2026.t9 VSS 0.093341f
C5478 a_n29_2026.n3 VSS 0.202001f
C5479 a_n29_2026.t3 VSS 0.093341f
C5480 a_n29_2026.t5 VSS 0.093341f
C5481 a_n29_2026.n4 VSS 0.202001f
C5482 a_n29_2026.t6 VSS 0.093341f
C5483 a_n29_2026.t11 VSS 0.093341f
C5484 a_n29_2026.n5 VSS 0.202001f
C5485 a_n29_2026.t0 VSS 0.093341f
C5486 a_n29_2026.t7 VSS 0.093341f
C5487 a_n29_2026.n6 VSS 0.202001f
C5488 a_n29_2026.n7 VSS 0.202296f
C5489 a_n29_2026.t2 VSS 0.093341f
C5490 mux8_4.NAND4F_0.Y.n0 VSS 0.350455f
C5491 mux8_4.NAND4F_0.Y.t10 VSS 0.022537f
C5492 mux8_4.NAND4F_0.Y.t9 VSS 0.079785f
C5493 mux8_4.NAND4F_0.Y.t11 VSS 0.024808f
C5494 mux8_4.NAND4F_0.Y.n1 VSS 0.070768f
C5495 mux8_4.NAND4F_0.Y.n2 VSS 0.020978f
C5496 mux8_4.NAND4F_0.Y.t1 VSS 0.017278f
C5497 mux8_4.NAND4F_0.Y.t0 VSS 0.017278f
C5498 mux8_4.NAND4F_0.Y.n3 VSS 0.040122f
C5499 mux8_4.NAND4F_0.Y.t3 VSS 0.017278f
C5500 mux8_4.NAND4F_0.Y.t2 VSS 0.017278f
C5501 mux8_4.NAND4F_0.Y.n4 VSS 0.040002f
C5502 mux8_4.NAND4F_0.Y.t8 VSS 0.017278f
C5503 mux8_4.NAND4F_0.Y.t7 VSS 0.017278f
C5504 mux8_4.NAND4F_0.Y.n5 VSS 0.040002f
C5505 mux8_4.NAND4F_0.Y.t5 VSS 0.017278f
C5506 mux8_4.NAND4F_0.Y.t6 VSS 0.017278f
C5507 mux8_4.NAND4F_0.Y.n6 VSS 0.040002f
C5508 mux8_4.NAND4F_0.Y.t4 VSS 0.166327f
C5509 a_n23065_2026.n0 VSS 1.48365f
C5510 a_n23065_2026.n1 VSS 1.48326f
C5511 a_n23065_2026.t1 VSS 0.093341f
C5512 a_n23065_2026.t4 VSS 0.093341f
C5513 a_n23065_2026.t5 VSS 0.093341f
C5514 a_n23065_2026.n2 VSS 0.202296f
C5515 a_n23065_2026.t3 VSS 0.093341f
C5516 a_n23065_2026.t7 VSS 0.093341f
C5517 a_n23065_2026.n3 VSS 0.202001f
C5518 a_n23065_2026.t8 VSS 0.093341f
C5519 a_n23065_2026.t6 VSS 0.093341f
C5520 a_n23065_2026.n4 VSS 0.202001f
C5521 a_n23065_2026.t10 VSS 0.093341f
C5522 a_n23065_2026.t11 VSS 0.093341f
C5523 a_n23065_2026.n5 VSS 0.202001f
C5524 a_n23065_2026.t9 VSS 0.093341f
C5525 a_n23065_2026.t0 VSS 0.093341f
C5526 a_n23065_2026.n6 VSS 0.202001f
C5527 a_n23065_2026.n7 VSS 0.20269f
C5528 a_n23065_2026.t2 VSS 0.093341f
C5529 mux8_2.NAND4F_2.D.n0 VSS 0.664607f
C5530 mux8_2.NAND4F_2.D.t7 VSS 0.027742f
C5531 mux8_2.NAND4F_2.D.t6 VSS 0.098211f
C5532 mux8_2.NAND4F_2.D.t8 VSS 0.030538f
C5533 mux8_2.NAND4F_2.D.n1 VSS 0.087112f
C5534 mux8_2.NAND4F_2.D.n2 VSS 0.025808f
C5535 mux8_2.NAND4F_2.D.t3 VSS 0.014135f
C5536 mux8_2.NAND4F_2.D.t2 VSS 0.014135f
C5537 mux8_2.NAND4F_2.D.n3 VSS 0.031499f
C5538 mux8_2.NAND4F_2.D.t1 VSS 0.051268f
C5539 mux8_2.NAND4F_2.D.t0 VSS 0.040771f
C5540 mux8_2.NAND4F_2.D.t13 VSS 0.027742f
C5541 mux8_2.NAND4F_2.D.t11 VSS 0.098211f
C5542 mux8_2.NAND4F_2.D.t14 VSS 0.030538f
C5543 mux8_2.NAND4F_2.D.n4 VSS 0.087112f
C5544 mux8_2.NAND4F_2.D.n5 VSS 0.025813f
C5545 mux8_2.NAND4F_2.D.n6 VSS 0.620222f
C5546 mux8_2.NAND4F_2.D.t9 VSS 0.027742f
C5547 mux8_2.NAND4F_2.D.t5 VSS 0.098211f
C5548 mux8_2.NAND4F_2.D.t10 VSS 0.030538f
C5549 mux8_2.NAND4F_2.D.n7 VSS 0.087112f
C5550 mux8_2.NAND4F_2.D.n8 VSS 0.025807f
C5551 mux8_2.NAND4F_2.D.n9 VSS 0.261852f
C5552 mux8_2.NAND4F_2.D.t12 VSS 0.027742f
C5553 mux8_2.NAND4F_2.D.t4 VSS 0.098211f
C5554 mux8_2.NAND4F_2.D.t15 VSS 0.030538f
C5555 mux8_2.NAND4F_2.D.n10 VSS 0.087112f
C5556 mux8_2.NAND4F_2.D.n11 VSS 0.025808f
C5557 mux8_2.NAND4F_2.D.n12 VSS 0.407824f
C5558 a_n15707_n4534.n0 VSS 1.48365f
C5559 a_n15707_n4534.n1 VSS 1.48326f
C5560 a_n15707_n4534.t5 VSS 0.093341f
C5561 a_n15707_n4534.t8 VSS 0.093341f
C5562 a_n15707_n4534.t7 VSS 0.093341f
C5563 a_n15707_n4534.n2 VSS 0.202296f
C5564 a_n15707_n4534.t6 VSS 0.093341f
C5565 a_n15707_n4534.t10 VSS 0.093341f
C5566 a_n15707_n4534.n3 VSS 0.202001f
C5567 a_n15707_n4534.t11 VSS 0.093341f
C5568 a_n15707_n4534.t9 VSS 0.093341f
C5569 a_n15707_n4534.n4 VSS 0.202001f
C5570 a_n15707_n4534.t4 VSS 0.093341f
C5571 a_n15707_n4534.t3 VSS 0.093341f
C5572 a_n15707_n4534.n5 VSS 0.202001f
C5573 a_n15707_n4534.t1 VSS 0.093341f
C5574 a_n15707_n4534.t0 VSS 0.093341f
C5575 a_n15707_n4534.n6 VSS 0.20269f
C5576 a_n15707_n4534.n7 VSS 0.202001f
C5577 a_n15707_n4534.t2 VSS 0.093341f
C5578 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n0 VSS 0.860417f
C5579 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t1 VSS 0.007445f
C5580 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t2 VSS 0.007445f
C5581 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n1 VSS 0.016566f
C5582 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t5 VSS 0.007445f
C5583 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t6 VSS 0.007445f
C5584 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n2 VSS 0.016611f
C5585 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t3 VSS 0.007445f
C5586 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t4 VSS 0.007445f
C5587 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n3 VSS 0.016566f
C5588 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t0 VSS 0.044951f
C5589 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t14 VSS 0.025427f
C5590 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t7 VSS 0.025111f
C5591 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t11 VSS 0.025111f
C5592 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t9 VSS 0.025111f
C5593 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n4 VSS 0.099949f
C5594 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t8 VSS 0.005218f
C5595 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t18 VSS 0.005218f
C5596 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t10 VSS 0.005218f
C5597 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t12 VSS 0.005218f
C5598 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n5 VSS 0.094423f
C5599 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n6 VSS 0.147672f
C5600 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t13 VSS 0.023482f
C5601 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t17 VSS 0.009013f
C5602 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t15 VSS 0.012447f
C5603 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n7 VSS 0.014327f
C5604 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.t16 VSS 0.009474f
C5605 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n8 VSS 0.014529f
C5606 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n9 VSS 0.049349f
C5607 8bit_ADDER_0.FULL_ADDER_XORED_6.COUT.n10 VSS 0.328172f
C5608 mux8_8.NAND4F_0.Y.n0 VSS 0.350455f
C5609 mux8_8.NAND4F_0.Y.t10 VSS 0.022537f
C5610 mux8_8.NAND4F_0.Y.t9 VSS 0.079785f
C5611 mux8_8.NAND4F_0.Y.t11 VSS 0.024808f
C5612 mux8_8.NAND4F_0.Y.n1 VSS 0.070768f
C5613 mux8_8.NAND4F_0.Y.n2 VSS 0.020978f
C5614 mux8_8.NAND4F_0.Y.t3 VSS 0.017278f
C5615 mux8_8.NAND4F_0.Y.t2 VSS 0.017278f
C5616 mux8_8.NAND4F_0.Y.n3 VSS 0.040122f
C5617 mux8_8.NAND4F_0.Y.t1 VSS 0.017278f
C5618 mux8_8.NAND4F_0.Y.t0 VSS 0.017278f
C5619 mux8_8.NAND4F_0.Y.n4 VSS 0.040002f
C5620 mux8_8.NAND4F_0.Y.t8 VSS 0.017278f
C5621 mux8_8.NAND4F_0.Y.t7 VSS 0.017278f
C5622 mux8_8.NAND4F_0.Y.n5 VSS 0.040002f
C5623 mux8_8.NAND4F_0.Y.t6 VSS 0.017278f
C5624 mux8_8.NAND4F_0.Y.t5 VSS 0.017278f
C5625 mux8_8.NAND4F_0.Y.n6 VSS 0.040002f
C5626 mux8_8.NAND4F_0.Y.t4 VSS 0.166327f
C5627 NOT8_0.S0.n0 VSS 3.50159f
C5628 NOT8_0.S0.t6 VSS 0.16986f
C5629 NOT8_0.S0.t5 VSS 0.500458f
C5630 NOT8_0.S0.t4 VSS 0.165263f
C5631 NOT8_0.S0.n1 VSS 0.852045f
C5632 NOT8_0.S0.t1 VSS 0.081426f
C5633 NOT8_0.S0.t3 VSS 0.081426f
C5634 NOT8_0.S0.n2 VSS 0.181453f
C5635 NOT8_0.S0.t2 VSS 0.295332f
C5636 NOT8_0.S0.t0 VSS 0.23486f
C5637 MULT_0.SO.n0 VSS 5.35653f
C5638 MULT_0.SO.t5 VSS 0.059065f
C5639 MULT_0.SO.t4 VSS 0.057466f
C5640 MULT_0.SO.t6 VSS 0.174023f
C5641 MULT_0.SO.n1 VSS 0.29628f
C5642 MULT_0.SO.t0 VSS 0.081804f
C5643 MULT_0.SO.t1 VSS 0.102695f
C5644 MULT_0.SO.t3 VSS 0.028314f
C5645 MULT_0.SO.t2 VSS 0.028314f
C5646 MULT_0.SO.n2 VSS 0.063082f
C5647 MULT_0.NAND2_3.Y.n0 VSS 0.294301f
C5648 MULT_0.NAND2_3.Y.n1 VSS 1.09643f
C5649 MULT_0.NAND2_3.Y.t9 VSS 0.028812f
C5650 MULT_0.NAND2_3.Y.t8 VSS 0.040219f
C5651 MULT_0.NAND2_3.Y.t10 VSS 0.040219f
C5652 MULT_0.NAND2_3.Y.n2 VSS 0.13121f
C5653 MULT_0.NAND2_3.Y.t7 VSS 0.045918f
C5654 MULT_0.NAND2_3.Y.t0 VSS 0.136194f
C5655 MULT_0.NAND2_3.Y.t5 VSS 0.022608f
C5656 MULT_0.NAND2_3.Y.t4 VSS 0.022608f
C5657 MULT_0.NAND2_3.Y.n3 VSS 0.050442f
C5658 MULT_0.NAND2_3.Y.t3 VSS 0.022608f
C5659 MULT_0.NAND2_3.Y.t6 VSS 0.022608f
C5660 MULT_0.NAND2_3.Y.n4 VSS 0.050306f
C5661 MULT_0.NAND2_3.Y.t2 VSS 0.022608f
C5662 MULT_0.NAND2_3.Y.t1 VSS 0.022608f
C5663 MULT_0.NAND2_3.Y.n5 VSS 0.050306f
C5664 a_n12314_n29052.n0 VSS 1.48365f
C5665 a_n12314_n29052.n1 VSS 1.48326f
C5666 a_n12314_n29052.t1 VSS 0.093341f
C5667 a_n12314_n29052.t3 VSS 0.093341f
C5668 a_n12314_n29052.t5 VSS 0.093341f
C5669 a_n12314_n29052.n2 VSS 0.202296f
C5670 a_n12314_n29052.t4 VSS 0.093341f
C5671 a_n12314_n29052.t9 VSS 0.093341f
C5672 a_n12314_n29052.n3 VSS 0.202001f
C5673 a_n12314_n29052.t8 VSS 0.093341f
C5674 a_n12314_n29052.t7 VSS 0.093341f
C5675 a_n12314_n29052.n4 VSS 0.202001f
C5676 a_n12314_n29052.t11 VSS 0.093341f
C5677 a_n12314_n29052.t6 VSS 0.093341f
C5678 a_n12314_n29052.n5 VSS 0.202001f
C5679 a_n12314_n29052.t10 VSS 0.093341f
C5680 a_n12314_n29052.t0 VSS 0.093341f
C5681 a_n12314_n29052.n6 VSS 0.202001f
C5682 a_n12314_n29052.n7 VSS 0.20269f
C5683 a_n12314_n29052.t2 VSS 0.093341f
C5684 OR8_0.S3.n0 VSS 1.08987f
C5685 mux8_4.NAND4F_2.A VSS 0.840041f
C5686 OR8_0.S3.t4 VSS 0.052718f
C5687 OR8_0.S3.t6 VSS 0.051291f
C5688 OR8_0.S3.t5 VSS 0.155322f
C5689 OR8_0.S3.n1 VSS 0.264441f
C5690 mux8_4.A3 VSS 5.5248f
C5691 OR8_0.S3.t1 VSS 0.025271f
C5692 OR8_0.S3.t2 VSS 0.025271f
C5693 OR8_0.S3.n2 VSS 0.056316f
C5694 OR8_0.S3.t3 VSS 0.091659f
C5695 OR8_0.S3.t0 VSS 0.072891f
C5696 OR8_0.NOT8_0.S3 VSS 3.95011f
C5697 MULT_0.inv_7.Y VSS 5.43413f
C5698 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_0.B VSS 0.867421f
C5699 MULT_0.4bit_ADDER_1.FULL_ADDER_2.A VSS 3.02874f
C5700 MULT_0.4bit_ADDER_1.A1.t14 VSS 0.066082f
C5701 MULT_0.4bit_ADDER_1.A1.t5 VSS 0.025365f
C5702 MULT_0.4bit_ADDER_1.A1.t4 VSS 0.035029f
C5703 MULT_0.4bit_ADDER_1.A1.n0 VSS 0.040318f
C5704 MULT_0.4bit_ADDER_1.A1.t6 VSS 0.026663f
C5705 MULT_0.4bit_ADDER_1.A1.n1 VSS 0.040888f
C5706 MULT_0.4bit_ADDER_1.A1.n2 VSS 0.169246f
C5707 MULT_0.4bit_ADDER_1.FULL_ADDER_2.NAND2_0.B VSS 0.653921f
C5708 MULT_0.4bit_ADDER_1.A1.t7 VSS 0.071557f
C5709 MULT_0.4bit_ADDER_1.A1.t12 VSS 0.070667f
C5710 MULT_0.4bit_ADDER_1.A1.t15 VSS 0.070667f
C5711 MULT_0.4bit_ADDER_1.A1.t13 VSS 0.070667f
C5712 MULT_0.4bit_ADDER_1.A1.n3 VSS 0.281275f
C5713 MULT_0.4bit_ADDER_1.A1.t10 VSS 0.014685f
C5714 MULT_0.4bit_ADDER_1.A1.t9 VSS 0.014685f
C5715 MULT_0.4bit_ADDER_1.A1.t11 VSS 0.014685f
C5716 MULT_0.4bit_ADDER_1.A1.t8 VSS 0.014685f
C5717 MULT_0.4bit_ADDER_1.A1.n4 VSS 0.265723f
C5718 MULT_0.4bit_ADDER_1.A1.n5 VSS 0.415645f
C5719 MULT_0.4bit_ADDER_1.A1.n6 VSS 0.982175f
C5720 MULT_0.4bit_ADDER_1.A1.t0 VSS 0.060568f
C5721 MULT_0.4bit_ADDER_1.A1.t2 VSS 0.075989f
C5722 MULT_0.4bit_ADDER_1.A1.t1 VSS 0.020951f
C5723 MULT_0.4bit_ADDER_1.A1.t3 VSS 0.020951f
C5724 MULT_0.4bit_ADDER_1.A1.n7 VSS 0.046618f
C5725 mux8_4.NAND4F_2.D.n0 VSS 0.664607f
C5726 mux8_4.NAND4F_2.D.t6 VSS 0.027742f
C5727 mux8_4.NAND4F_2.D.t9 VSS 0.098211f
C5728 mux8_4.NAND4F_2.D.t5 VSS 0.030538f
C5729 mux8_4.NAND4F_2.D.n1 VSS 0.087112f
C5730 mux8_4.NAND4F_2.D.n2 VSS 0.025808f
C5731 mux8_4.NAND4F_2.D.t3 VSS 0.014135f
C5732 mux8_4.NAND4F_2.D.t2 VSS 0.014135f
C5733 mux8_4.NAND4F_2.D.n3 VSS 0.031499f
C5734 mux8_4.NAND4F_2.D.t1 VSS 0.051268f
C5735 mux8_4.NAND4F_2.D.t0 VSS 0.040771f
C5736 mux8_4.NAND4F_2.D.t15 VSS 0.027742f
C5737 mux8_4.NAND4F_2.D.t7 VSS 0.098211f
C5738 mux8_4.NAND4F_2.D.t10 VSS 0.030538f
C5739 mux8_4.NAND4F_2.D.n4 VSS 0.087112f
C5740 mux8_4.NAND4F_2.D.n5 VSS 0.025813f
C5741 mux8_4.NAND4F_2.D.n6 VSS 0.620222f
C5742 mux8_4.NAND4F_2.D.t14 VSS 0.027742f
C5743 mux8_4.NAND4F_2.D.t12 VSS 0.098211f
C5744 mux8_4.NAND4F_2.D.t13 VSS 0.030538f
C5745 mux8_4.NAND4F_2.D.n7 VSS 0.087112f
C5746 mux8_4.NAND4F_2.D.n8 VSS 0.025807f
C5747 mux8_4.NAND4F_2.D.n9 VSS 0.261852f
C5748 mux8_4.NAND4F_2.D.t11 VSS 0.027742f
C5749 mux8_4.NAND4F_2.D.t4 VSS 0.098211f
C5750 mux8_4.NAND4F_2.D.t8 VSS 0.030538f
C5751 mux8_4.NAND4F_2.D.n10 VSS 0.087112f
C5752 mux8_4.NAND4F_2.D.n11 VSS 0.025808f
C5753 mux8_4.NAND4F_2.D.n12 VSS 0.407824f
C5754 a_n12416_n7799.n0 VSS 1.48365f
C5755 a_n12416_n7799.n1 VSS 1.48326f
C5756 a_n12416_n7799.t1 VSS 0.093341f
C5757 a_n12416_n7799.t8 VSS 0.093341f
C5758 a_n12416_n7799.t7 VSS 0.093341f
C5759 a_n12416_n7799.n2 VSS 0.202296f
C5760 a_n12416_n7799.t6 VSS 0.093341f
C5761 a_n12416_n7799.t10 VSS 0.093341f
C5762 a_n12416_n7799.n3 VSS 0.202001f
C5763 a_n12416_n7799.t11 VSS 0.093341f
C5764 a_n12416_n7799.t9 VSS 0.093341f
C5765 a_n12416_n7799.n4 VSS 0.202001f
C5766 a_n12416_n7799.t4 VSS 0.093341f
C5767 a_n12416_n7799.t3 VSS 0.093341f
C5768 a_n12416_n7799.n5 VSS 0.202001f
C5769 a_n12416_n7799.t5 VSS 0.093341f
C5770 a_n12416_n7799.t0 VSS 0.093341f
C5771 a_n12416_n7799.n6 VSS 0.202001f
C5772 a_n12416_n7799.n7 VSS 0.20269f
C5773 a_n12416_n7799.t2 VSS 0.093341f
C5774 mux8_4.NAND4F_1.Y.n0 VSS 0.655599f
C5775 mux8_4.NAND4F_1.Y.t4 VSS 0.306614f
C5776 mux8_4.NAND4F_1.Y.t11 VSS 0.132168f
C5777 mux8_4.NAND4F_1.Y.t10 VSS 0.04216f
C5778 mux8_4.NAND4F_1.Y.t9 VSS 0.04216f
C5779 mux8_4.NAND4F_1.Y.n1 VSS 0.049498f
C5780 mux8_4.NAND4F_1.Y.n2 VSS 0.277534f
C5781 mux8_4.NAND4F_1.Y.t1 VSS 0.032323f
C5782 mux8_4.NAND4F_1.Y.t0 VSS 0.032323f
C5783 mux8_4.NAND4F_1.Y.n3 VSS 0.075057f
C5784 mux8_4.NAND4F_1.Y.t3 VSS 0.032323f
C5785 mux8_4.NAND4F_1.Y.t2 VSS 0.032323f
C5786 mux8_4.NAND4F_1.Y.n4 VSS 0.074832f
C5787 mux8_4.NAND4F_1.Y.t8 VSS 0.032323f
C5788 mux8_4.NAND4F_1.Y.t7 VSS 0.032323f
C5789 mux8_4.NAND4F_1.Y.n5 VSS 0.074832f
C5790 mux8_4.NAND4F_1.Y.t6 VSS 0.032323f
C5791 mux8_4.NAND4F_1.Y.t5 VSS 0.032323f
C5792 mux8_4.NAND4F_1.Y.n6 VSS 0.074832f
C5793 mux8_4.NAND4F_1.Y.n7 VSS 0.307603f
C5794 MULT_0.4bit_ADDER_1.FULL_ADDER_2.OUT VSS 0.563979f
C5795 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_0.A VSS 0.1564f
C5796 MULT_0.4bit_ADDER_2.FULL_ADDER_3.B VSS 0.34251f
C5797 MULT_0.4bit_ADDER_2.B0.t23 VSS 0.041874f
C5798 MULT_0.4bit_ADDER_2.B0.t22 VSS 0.013636f
C5799 MULT_0.4bit_ADDER_2.B0.t14 VSS 0.018831f
C5800 MULT_0.4bit_ADDER_2.B0.n0 VSS 0.020307f
C5801 MULT_0.4bit_ADDER_2.B0.t21 VSS 0.014019f
C5802 MULT_0.4bit_ADDER_2.B0.n1 VSS 0.035571f
C5803 MULT_0.4bit_ADDER_2.B0.n2 VSS 0.062398f
C5804 MULT_0.4bit_ADDER_2.B0.t17 VSS 0.019119f
C5805 MULT_0.4bit_ADDER_2.B0.t19 VSS 0.038468f
C5806 MULT_0.4bit_ADDER_2.B0.t12 VSS 0.037989f
C5807 MULT_0.4bit_ADDER_2.B0.t13 VSS 0.037989f
C5808 MULT_0.4bit_ADDER_2.B0.t18 VSS 0.037989f
C5809 MULT_0.4bit_ADDER_2.B0.t20 VSS 0.007895f
C5810 MULT_0.4bit_ADDER_2.B0.t16 VSS 0.007895f
C5811 MULT_0.4bit_ADDER_2.B0.t15 VSS 0.007895f
C5812 MULT_0.4bit_ADDER_2.B0.n3 VSS 0.234048f
C5813 MULT_0.4bit_ADDER_2.B0.n4 VSS 0.172387f
C5814 MULT_0.4bit_ADDER_2.B0.n5 VSS 0.093949f
C5815 MULT_0.4bit_ADDER_2.B0.n6 VSS 0.092297f
C5816 MULT_0.4bit_ADDER_2.B0.n7 VSS 0.056773f
C5817 MULT_0.4bit_ADDER_2.B0.n8 VSS 0.074476f
C5818 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_0.A VSS 0.132446f
C5819 MULT_0.4bit_ADDER_2.B0.n9 VSS 0.822778f
C5820 MULT_0.4bit_ADDER_2.B0.t2 VSS 0.006842f
C5821 MULT_0.4bit_ADDER_2.B0.t0 VSS 0.006842f
C5822 MULT_0.4bit_ADDER_2.B0.n10 VSS 0.016548f
C5823 MULT_0.4bit_ADDER_2.B0.t7 VSS 0.006842f
C5824 MULT_0.4bit_ADDER_2.B0.t3 VSS 0.006842f
C5825 MULT_0.4bit_ADDER_2.B0.n11 VSS 0.016546f
C5826 MULT_0.4bit_ADDER_2.B0.n12 VSS 0.11865f
C5827 MULT_0.4bit_ADDER_2.B0.t1 VSS 0.006842f
C5828 MULT_0.4bit_ADDER_2.B0.t8 VSS 0.006842f
C5829 MULT_0.4bit_ADDER_2.B0.n13 VSS 0.013684f
C5830 MULT_0.4bit_ADDER_2.B0.n14 VSS 0.010749f
C5831 MULT_0.4bit_ADDER_2.B0.t9 VSS 0.028947f
C5832 MULT_0.4bit_ADDER_2.B0.t5 VSS 0.028947f
C5833 MULT_0.4bit_ADDER_2.B0.n15 VSS 0.057893f
C5834 MULT_0.4bit_ADDER_2.B0.n16 VSS 0.023019f
C5835 MULT_0.4bit_ADDER_2.B0.t10 VSS 0.028947f
C5836 MULT_0.4bit_ADDER_2.B0.t11 VSS 0.028947f
C5837 MULT_0.4bit_ADDER_2.B0.n17 VSS 0.057893f
C5838 MULT_0.4bit_ADDER_2.B0.n18 VSS 0.025462f
C5839 MULT_0.4bit_ADDER_2.B0.n19 VSS 0.262149f
C5840 MULT_0.4bit_ADDER_2.B0.t4 VSS 0.028947f
C5841 MULT_0.4bit_ADDER_2.B0.t6 VSS 0.028947f
C5842 MULT_0.4bit_ADDER_2.B0.n20 VSS 0.057893f
C5843 MULT_0.4bit_ADDER_2.B0.n21 VSS 0.025501f
C5844 MULT_0.4bit_ADDER_2.B0.n22 VSS 0.168131f
C5845 MULT_0.4bit_ADDER_2.B0.n23 VSS 0.03789f
C5846 MULT_0.4bit_ADDER_2.B0.n24 VSS 0.166308f
C5847 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.Y VSS 0.383036f
C5848 a_n12316_n34281.n0 VSS 1.48326f
C5849 a_n12316_n34281.n1 VSS 1.48365f
C5850 a_n12316_n34281.t0 VSS 0.093341f
C5851 a_n12316_n34281.t6 VSS 0.093341f
C5852 a_n12316_n34281.t8 VSS 0.093341f
C5853 a_n12316_n34281.n2 VSS 0.20269f
C5854 a_n12316_n34281.t3 VSS 0.093341f
C5855 a_n12316_n34281.t7 VSS 0.093341f
C5856 a_n12316_n34281.n3 VSS 0.202001f
C5857 a_n12316_n34281.t5 VSS 0.093341f
C5858 a_n12316_n34281.t4 VSS 0.093341f
C5859 a_n12316_n34281.n4 VSS 0.202001f
C5860 a_n12316_n34281.t10 VSS 0.093341f
C5861 a_n12316_n34281.t9 VSS 0.093341f
C5862 a_n12316_n34281.n5 VSS 0.202001f
C5863 a_n12316_n34281.t1 VSS 0.093341f
C5864 a_n12316_n34281.t11 VSS 0.093341f
C5865 a_n12316_n34281.n6 VSS 0.202001f
C5866 a_n12316_n34281.n7 VSS 0.202296f
C5867 a_n12316_n34281.t2 VSS 0.093341f
C5868 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t14 VSS 0.013766f
C5869 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t19 VSS 0.027698f
C5870 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t23 VSS 0.027354f
C5871 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t13 VSS 0.027354f
C5872 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t17 VSS 0.027354f
C5873 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t15 VSS 0.005684f
C5874 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t12 VSS 0.005684f
C5875 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t22 VSS 0.005684f
C5876 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n0 VSS 0.168523f
C5877 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n1 VSS 0.124125f
C5878 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n2 VSS 0.067647f
C5879 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n3 VSS 0.066457f
C5880 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n4 VSS 0.040879f
C5881 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n5 VSS 0.05311f
C5882 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t16 VSS 0.030151f
C5883 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t21 VSS 0.009818f
C5884 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t18 VSS 0.013559f
C5885 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n6 VSS 0.014622f
C5886 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t20 VSS 0.010094f
C5887 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n7 VSS 0.025612f
C5888 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n8 VSS 0.044927f
C5889 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t2 VSS 0.004926f
C5890 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t3 VSS 0.004926f
C5891 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n9 VSS 0.011915f
C5892 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t7 VSS 0.004926f
C5893 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t8 VSS 0.004926f
C5894 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n10 VSS 0.011914f
C5895 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n11 VSS 0.085433f
C5896 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t1 VSS 0.004926f
C5897 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t4 VSS 0.004926f
C5898 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n12 VSS 0.009853f
C5899 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n13 VSS 0.00774f
C5900 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t11 VSS 0.020843f
C5901 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t6 VSS 0.020843f
C5902 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n14 VSS 0.041685f
C5903 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n15 VSS 0.016575f
C5904 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t10 VSS 0.020843f
C5905 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t9 VSS 0.020843f
C5906 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n16 VSS 0.041685f
C5907 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n17 VSS 0.018334f
C5908 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n18 VSS 0.188757f
C5909 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t0 VSS 0.020843f
C5910 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.t5 VSS 0.020843f
C5911 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n19 VSS 0.041685f
C5912 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n20 VSS 0.018362f
C5913 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n21 VSS 0.12106f
C5914 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n22 VSS 0.027282f
C5915 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_1.A.n23 VSS 0.119748f
C5916 mux8_2.NAND4F_3.Y.n0 VSS 0.306333f
C5917 mux8_2.NAND4F_3.Y.t3 VSS 0.015103f
C5918 mux8_2.NAND4F_3.Y.t2 VSS 0.015103f
C5919 mux8_2.NAND4F_3.Y.n1 VSS 0.035071f
C5920 mux8_2.NAND4F_3.Y.t0 VSS 0.015103f
C5921 mux8_2.NAND4F_3.Y.t1 VSS 0.015103f
C5922 mux8_2.NAND4F_3.Y.n2 VSS 0.034966f
C5923 mux8_2.NAND4F_3.Y.t7 VSS 0.015103f
C5924 mux8_2.NAND4F_3.Y.t8 VSS 0.015103f
C5925 mux8_2.NAND4F_3.Y.n3 VSS 0.034966f
C5926 mux8_2.NAND4F_3.Y.t6 VSS 0.015103f
C5927 mux8_2.NAND4F_3.Y.t5 VSS 0.015103f
C5928 mux8_2.NAND4F_3.Y.n4 VSS 0.034966f
C5929 mux8_2.NAND4F_3.Y.n5 VSS 0.152246f
C5930 mux8_2.NAND4F_3.Y.t4 VSS 0.143521f
C5931 mux8_2.NAND4F_3.Y.t10 VSS 0.0197f
C5932 mux8_2.NAND4F_3.Y.t9 VSS 0.0197f
C5933 mux8_2.NAND4F_3.Y.n6 VSS 0.023128f
C5934 mux8_2.NAND4F_3.Y.t11 VSS 0.061756f
C5935 mux8_2.NAND4F_3.Y.n7 VSS 0.129679f
C5936 mux8_3.NAND4F_0.C.n0 VSS 1.72379f
C5937 mux8_3.NAND4F_0.C.t6 VSS 0.238621f
C5938 mux8_3.NAND4F_0.C.t10 VSS 0.076118f
C5939 mux8_3.NAND4F_0.C.t9 VSS 0.076118f
C5940 mux8_3.NAND4F_0.C.n1 VSS 0.089365f
C5941 mux8_3.NAND4F_0.C.n2 VSS 0.501052f
C5942 mux8_3.NAND4F_0.C.t5 VSS 0.076118f
C5943 mux8_3.NAND4F_0.C.t7 VSS 0.076118f
C5944 mux8_3.NAND4F_0.C.n3 VSS 0.089365f
C5945 mux8_3.NAND4F_0.C.t4 VSS 0.238621f
C5946 mux8_3.NAND4F_0.C.n4 VSS 0.501084f
C5947 mux8_3.NAND4F_0.C.t11 VSS 0.076118f
C5948 mux8_3.NAND4F_0.C.t12 VSS 0.076118f
C5949 mux8_3.NAND4F_0.C.n5 VSS 0.089365f
C5950 mux8_3.NAND4F_0.C.t8 VSS 0.238621f
C5951 mux8_3.NAND4F_0.C.n6 VSS 0.501098f
C5952 mux8_3.NAND4F_0.C.n7 VSS 1.82754f
C5953 mux8_3.NAND4F_0.C.t3 VSS 0.038784f
C5954 mux8_3.NAND4F_0.C.t2 VSS 0.038784f
C5955 mux8_3.NAND4F_0.C.n8 VSS 0.086427f
C5956 mux8_3.NAND4F_0.C.t1 VSS 0.140669f
C5957 mux8_3.NAND4F_0.C.t0 VSS 0.111866f
C5958 mux8_3.NAND4F_0.C.n9 VSS 3.19968f
C5959 mux8_3.NAND4F_0.C.t15 VSS 0.238621f
C5960 mux8_3.NAND4F_0.C.t14 VSS 0.076118f
C5961 mux8_3.NAND4F_0.C.t13 VSS 0.076118f
C5962 mux8_3.NAND4F_0.C.n10 VSS 0.089365f
C5963 mux8_3.NAND4F_0.C.n11 VSS 0.50107f
C5964 mux8_3.NAND4F_0.C.n12 VSS 2.56421f
C5965 mux8_8.NAND4F_2.D.n0 VSS 0.664607f
C5966 mux8_8.NAND4F_2.D.t14 VSS 0.027742f
C5967 mux8_8.NAND4F_2.D.t11 VSS 0.098211f
C5968 mux8_8.NAND4F_2.D.t13 VSS 0.030538f
C5969 mux8_8.NAND4F_2.D.n1 VSS 0.087112f
C5970 mux8_8.NAND4F_2.D.n2 VSS 0.025808f
C5971 mux8_8.NAND4F_2.D.t1 VSS 0.014135f
C5972 mux8_8.NAND4F_2.D.t3 VSS 0.014135f
C5973 mux8_8.NAND4F_2.D.n3 VSS 0.031499f
C5974 mux8_8.NAND4F_2.D.t2 VSS 0.051268f
C5975 mux8_8.NAND4F_2.D.t0 VSS 0.040771f
C5976 mux8_8.NAND4F_2.D.t10 VSS 0.027742f
C5977 mux8_8.NAND4F_2.D.t7 VSS 0.098211f
C5978 mux8_8.NAND4F_2.D.t5 VSS 0.030538f
C5979 mux8_8.NAND4F_2.D.n4 VSS 0.087112f
C5980 mux8_8.NAND4F_2.D.n5 VSS 0.025813f
C5981 mux8_8.NAND4F_2.D.n6 VSS 0.620222f
C5982 mux8_8.NAND4F_2.D.t9 VSS 0.027742f
C5983 mux8_8.NAND4F_2.D.t12 VSS 0.098211f
C5984 mux8_8.NAND4F_2.D.t8 VSS 0.030538f
C5985 mux8_8.NAND4F_2.D.n7 VSS 0.087112f
C5986 mux8_8.NAND4F_2.D.n8 VSS 0.025807f
C5987 mux8_8.NAND4F_2.D.n9 VSS 0.261852f
C5988 mux8_8.NAND4F_2.D.t6 VSS 0.027742f
C5989 mux8_8.NAND4F_2.D.t15 VSS 0.098211f
C5990 mux8_8.NAND4F_2.D.t4 VSS 0.030538f
C5991 mux8_8.NAND4F_2.D.n10 VSS 0.087112f
C5992 mux8_8.NAND4F_2.D.n11 VSS 0.025808f
C5993 mux8_8.NAND4F_2.D.n12 VSS 0.407824f
C5994 mux8_8.NAND4F_0.C.n0 VSS 1.66671f
C5995 mux8_8.NAND4F_0.C.t13 VSS 0.230719f
C5996 mux8_8.NAND4F_0.C.t10 VSS 0.073597f
C5997 mux8_8.NAND4F_0.C.t8 VSS 0.073597f
C5998 mux8_8.NAND4F_0.C.n1 VSS 0.086405f
C5999 mux8_8.NAND4F_0.C.n2 VSS 0.484461f
C6000 mux8_8.NAND4F_0.C.t4 VSS 0.073597f
C6001 mux8_8.NAND4F_0.C.t5 VSS 0.073597f
C6002 mux8_8.NAND4F_0.C.n3 VSS 0.086405f
C6003 mux8_8.NAND4F_0.C.t9 VSS 0.230719f
C6004 mux8_8.NAND4F_0.C.n4 VSS 0.484492f
C6005 mux8_8.NAND4F_0.C.t12 VSS 0.073597f
C6006 mux8_8.NAND4F_0.C.t14 VSS 0.073597f
C6007 mux8_8.NAND4F_0.C.n5 VSS 0.086405f
C6008 mux8_8.NAND4F_0.C.t15 VSS 0.230719f
C6009 mux8_8.NAND4F_0.C.n6 VSS 0.484506f
C6010 mux8_8.NAND4F_0.C.n7 VSS 1.76702f
C6011 mux8_8.NAND4F_0.C.t1 VSS 0.0375f
C6012 mux8_8.NAND4F_0.C.t3 VSS 0.0375f
C6013 mux8_8.NAND4F_0.C.n8 VSS 0.083565f
C6014 mux8_8.NAND4F_0.C.t2 VSS 0.136011f
C6015 mux8_8.NAND4F_0.C.t0 VSS 0.108161f
C6016 mux8_8.NAND4F_0.C.n9 VSS 3.09373f
C6017 mux8_8.NAND4F_0.C.t11 VSS 0.230719f
C6018 mux8_8.NAND4F_0.C.t7 VSS 0.073597f
C6019 mux8_8.NAND4F_0.C.t6 VSS 0.073597f
C6020 mux8_8.NAND4F_0.C.n10 VSS 0.086405f
C6021 mux8_8.NAND4F_0.C.n11 VSS 0.484478f
C6022 mux8_8.NAND4F_0.C.n12 VSS 2.47931f
C6023 mux8_2.NAND4F_3.A VSS 0.720312f
C6024 8bit_ADDER_0.FULL_ADDER_XORED_6.OUT VSS 3.66612f
C6025 8bit_ADDER_0.S1.t12 VSS 0.044741f
C6026 8bit_ADDER_0.S1.t14 VSS 0.04353f
C6027 8bit_ADDER_0.S1.t13 VSS 0.131821f
C6028 8bit_ADDER_0.S1.n0 VSS 0.224429f
C6029 mux8_2.A0 VSS 4.01562f
C6030 8bit_ADDER_0.S1.t1 VSS 0.013029f
C6031 8bit_ADDER_0.S1.t2 VSS 0.013029f
C6032 8bit_ADDER_0.S1.n1 VSS 0.031512f
C6033 8bit_ADDER_0.S1.t8 VSS 0.013029f
C6034 8bit_ADDER_0.S1.t7 VSS 0.013029f
C6035 8bit_ADDER_0.S1.n2 VSS 0.031509f
C6036 8bit_ADDER_0.S1.n3 VSS 0.225945f
C6037 8bit_ADDER_0.S1.t0 VSS 0.013029f
C6038 8bit_ADDER_0.S1.t6 VSS 0.013029f
C6039 8bit_ADDER_0.S1.n4 VSS 0.026058f
C6040 8bit_ADDER_0.S1.n5 VSS 0.020469f
C6041 8bit_ADDER_0.S1.t4 VSS 0.055123f
C6042 8bit_ADDER_0.S1.t10 VSS 0.055123f
C6043 8bit_ADDER_0.S1.n6 VSS 0.110245f
C6044 8bit_ADDER_0.S1.n7 VSS 0.043835f
C6045 8bit_ADDER_0.S1.t5 VSS 0.055123f
C6046 8bit_ADDER_0.S1.t3 VSS 0.055123f
C6047 8bit_ADDER_0.S1.n8 VSS 0.110245f
C6048 8bit_ADDER_0.S1.n9 VSS 0.048488f
C6049 8bit_ADDER_0.S1.n10 VSS 0.499209f
C6050 8bit_ADDER_0.S1.t9 VSS 0.055123f
C6051 8bit_ADDER_0.S1.t11 VSS 0.055123f
C6052 8bit_ADDER_0.S1.n11 VSS 0.110245f
C6053 8bit_ADDER_0.S1.n12 VSS 0.048561f
C6054 8bit_ADDER_0.S1.n13 VSS 0.320171f
C6055 8bit_ADDER_0.S1.n14 VSS 0.072154f
C6056 8bit_ADDER_0.S1.n15 VSS 0.316699f
C6057 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.Y VSS 0.729173f
C6058 a_n3320_2026.n0 VSS 1.48365f
C6059 a_n3320_2026.n1 VSS 1.48326f
C6060 a_n3320_2026.t0 VSS 0.093341f
C6061 a_n3320_2026.t8 VSS 0.093341f
C6062 a_n3320_2026.t6 VSS 0.093341f
C6063 a_n3320_2026.n2 VSS 0.202296f
C6064 a_n3320_2026.t7 VSS 0.093341f
C6065 a_n3320_2026.t5 VSS 0.093341f
C6066 a_n3320_2026.n3 VSS 0.202001f
C6067 a_n3320_2026.t3 VSS 0.093341f
C6068 a_n3320_2026.t4 VSS 0.093341f
C6069 a_n3320_2026.n4 VSS 0.202001f
C6070 a_n3320_2026.t10 VSS 0.093341f
C6071 a_n3320_2026.t9 VSS 0.093341f
C6072 a_n3320_2026.n5 VSS 0.202001f
C6073 a_n3320_2026.t11 VSS 0.093341f
C6074 a_n3320_2026.t1 VSS 0.093341f
C6075 a_n3320_2026.n6 VSS 0.202001f
C6076 a_n3320_2026.n7 VSS 0.20269f
C6077 a_n3320_2026.t2 VSS 0.093341f
C6078 mux8_8.A0.t14 VSS 0.060866f
C6079 mux8_8.A0.t12 VSS 0.059219f
C6080 mux8_8.A0.t13 VSS 0.179329f
C6081 mux8_8.A0.n0 VSS 0.305314f
C6082 mux8_8.A0.t0 VSS 0.017725f
C6083 mux8_8.A0.t5 VSS 0.017725f
C6084 mux8_8.A0.n1 VSS 0.042869f
C6085 mux8_8.A0.t10 VSS 0.017725f
C6086 mux8_8.A0.t11 VSS 0.017725f
C6087 mux8_8.A0.n2 VSS 0.042864f
C6088 mux8_8.A0.n3 VSS 0.307375f
C6089 mux8_8.A0.t4 VSS 0.017725f
C6090 mux8_8.A0.t6 VSS 0.017725f
C6091 mux8_8.A0.n4 VSS 0.035449f
C6092 mux8_8.A0.n5 VSS 0.027846f
C6093 mux8_8.A0.t3 VSS 0.074989f
C6094 mux8_8.A0.t8 VSS 0.074989f
C6095 mux8_8.A0.n6 VSS 0.149978f
C6096 mux8_8.A0.n7 VSS 0.059634f
C6097 mux8_8.A0.t2 VSS 0.074989f
C6098 mux8_8.A0.t1 VSS 0.074989f
C6099 mux8_8.A0.n8 VSS 0.149978f
C6100 mux8_8.A0.n9 VSS 0.065963f
C6101 mux8_8.A0.n10 VSS 0.679123f
C6102 mux8_8.A0.t9 VSS 0.074989f
C6103 mux8_8.A0.t7 VSS 0.074989f
C6104 mux8_8.A0.n11 VSS 0.149978f
C6105 mux8_8.A0.n12 VSS 0.066063f
C6106 mux8_8.A0.n13 VSS 0.43556f
C6107 mux8_8.A0.n14 VSS 0.098158f
C6108 mux8_8.A0.n15 VSS 0.430837f
C6109 Y5.t7 VSS 0.069463f
C6110 Y5.t4 VSS 0.075053f
C6111 Y5.n0 VSS 0.05929f
C6112 Y5.t6 VSS 0.069861f
C6113 Y5.n1 VSS 0.033594f
C6114 Y5.t5 VSS 0.032356f
C6115 Y5.n2 VSS 0.034509f
C6116 Y5.t3 VSS 0.012998f
C6117 Y5.t2 VSS 0.012998f
C6118 Y5.n3 VSS 0.028945f
C6119 Y5.t1 VSS 0.047144f
C6120 Y5.n4 VSS 0.056322f
C6121 Y5.t0 VSS 0.037543f
C6122 Y5.n5 VSS 0.147272f
C6123 a_n11460_2026.n0 VSS 1.48326f
C6124 a_n11460_2026.n1 VSS 1.48365f
C6125 a_n11460_2026.t1 VSS 0.093341f
C6126 a_n11460_2026.t3 VSS 0.093341f
C6127 a_n11460_2026.t4 VSS 0.093341f
C6128 a_n11460_2026.n2 VSS 0.202296f
C6129 a_n11460_2026.t5 VSS 0.093341f
C6130 a_n11460_2026.t0 VSS 0.093341f
C6131 a_n11460_2026.n3 VSS 0.202001f
C6132 a_n11460_2026.t8 VSS 0.093341f
C6133 a_n11460_2026.t6 VSS 0.093341f
C6134 a_n11460_2026.n4 VSS 0.20269f
C6135 a_n11460_2026.t10 VSS 0.093341f
C6136 a_n11460_2026.t7 VSS 0.093341f
C6137 a_n11460_2026.n5 VSS 0.202001f
C6138 a_n11460_2026.t11 VSS 0.093341f
C6139 a_n11460_2026.t9 VSS 0.093341f
C6140 a_n11460_2026.n6 VSS 0.202001f
C6141 a_n11460_2026.n7 VSS 0.202001f
C6142 a_n11460_2026.t2 VSS 0.093341f
C6143 a_n9125_n7799.n0 VSS 1.48365f
C6144 a_n9125_n7799.n1 VSS 1.48326f
C6145 a_n9125_n7799.t4 VSS 0.093341f
C6146 a_n9125_n7799.t11 VSS 0.093341f
C6147 a_n9125_n7799.t10 VSS 0.093341f
C6148 a_n9125_n7799.n2 VSS 0.202296f
C6149 a_n9125_n7799.t9 VSS 0.093341f
C6150 a_n9125_n7799.t7 VSS 0.093341f
C6151 a_n9125_n7799.n3 VSS 0.202001f
C6152 a_n9125_n7799.t8 VSS 0.093341f
C6153 a_n9125_n7799.t6 VSS 0.093341f
C6154 a_n9125_n7799.n4 VSS 0.202001f
C6155 a_n9125_n7799.t0 VSS 0.093341f
C6156 a_n9125_n7799.t1 VSS 0.093341f
C6157 a_n9125_n7799.n5 VSS 0.202001f
C6158 a_n9125_n7799.t2 VSS 0.093341f
C6159 a_n9125_n7799.t3 VSS 0.093341f
C6160 a_n9125_n7799.n6 VSS 0.202001f
C6161 a_n9125_n7799.n7 VSS 0.20269f
C6162 a_n9125_n7799.t5 VSS 0.093341f
C6163 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t16 VSS 0.013766f
C6164 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t20 VSS 0.027698f
C6165 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t13 VSS 0.027354f
C6166 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t12 VSS 0.027354f
C6167 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t22 VSS 0.027354f
C6168 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t19 VSS 0.005684f
C6169 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t14 VSS 0.005684f
C6170 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t17 VSS 0.005684f
C6171 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n0 VSS 0.168523f
C6172 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n1 VSS 0.124125f
C6173 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n2 VSS 0.067647f
C6174 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n3 VSS 0.066457f
C6175 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n4 VSS 0.040879f
C6176 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n5 VSS 0.05311f
C6177 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t15 VSS 0.030151f
C6178 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t21 VSS 0.009818f
C6179 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t18 VSS 0.013559f
C6180 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n6 VSS 0.014622f
C6181 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t23 VSS 0.010094f
C6182 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n7 VSS 0.025612f
C6183 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n8 VSS 0.044927f
C6184 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t2 VSS 0.004926f
C6185 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t4 VSS 0.004926f
C6186 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n9 VSS 0.011915f
C6187 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t0 VSS 0.004926f
C6188 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t8 VSS 0.004926f
C6189 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n10 VSS 0.011914f
C6190 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n11 VSS 0.085433f
C6191 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t3 VSS 0.004926f
C6192 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t11 VSS 0.004926f
C6193 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n12 VSS 0.009853f
C6194 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n13 VSS 0.00774f
C6195 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t7 VSS 0.020843f
C6196 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t1 VSS 0.020843f
C6197 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n14 VSS 0.041685f
C6198 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n15 VSS 0.016575f
C6199 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t5 VSS 0.020843f
C6200 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t6 VSS 0.020843f
C6201 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n16 VSS 0.041685f
C6202 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n17 VSS 0.018334f
C6203 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n18 VSS 0.188757f
C6204 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t9 VSS 0.020843f
C6205 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.t10 VSS 0.020843f
C6206 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n19 VSS 0.041685f
C6207 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n20 VSS 0.018362f
C6208 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n21 VSS 0.12106f
C6209 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n22 VSS 0.027282f
C6210 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_1.A.n23 VSS 0.119748f
C6211 mux8_6.NAND4F_2.D.n0 VSS 0.64506f
C6212 mux8_6.NAND4F_2.D.t14 VSS 0.026926f
C6213 mux8_6.NAND4F_2.D.t5 VSS 0.095322f
C6214 mux8_6.NAND4F_2.D.t13 VSS 0.029639f
C6215 mux8_6.NAND4F_2.D.n1 VSS 0.084549f
C6216 mux8_6.NAND4F_2.D.n2 VSS 0.025049f
C6217 mux8_6.NAND4F_2.D.t3 VSS 0.013719f
C6218 mux8_6.NAND4F_2.D.t2 VSS 0.013719f
C6219 mux8_6.NAND4F_2.D.n3 VSS 0.030573f
C6220 mux8_6.NAND4F_2.D.t1 VSS 0.04976f
C6221 mux8_6.NAND4F_2.D.t0 VSS 0.039572f
C6222 mux8_6.NAND4F_2.D.t11 VSS 0.026926f
C6223 mux8_6.NAND4F_2.D.t15 VSS 0.095322f
C6224 mux8_6.NAND4F_2.D.t6 VSS 0.029639f
C6225 mux8_6.NAND4F_2.D.n4 VSS 0.084549f
C6226 mux8_6.NAND4F_2.D.n5 VSS 0.025054f
C6227 mux8_6.NAND4F_2.D.n6 VSS 0.601981f
C6228 mux8_6.NAND4F_2.D.t10 VSS 0.026926f
C6229 mux8_6.NAND4F_2.D.t8 VSS 0.095322f
C6230 mux8_6.NAND4F_2.D.t9 VSS 0.029639f
C6231 mux8_6.NAND4F_2.D.n7 VSS 0.084549f
C6232 mux8_6.NAND4F_2.D.n8 VSS 0.025048f
C6233 mux8_6.NAND4F_2.D.n9 VSS 0.254151f
C6234 mux8_6.NAND4F_2.D.t7 VSS 0.026926f
C6235 mux8_6.NAND4F_2.D.t12 VSS 0.095322f
C6236 mux8_6.NAND4F_2.D.t4 VSS 0.029639f
C6237 mux8_6.NAND4F_2.D.n10 VSS 0.084549f
C6238 mux8_6.NAND4F_2.D.n11 VSS 0.025049f
C6239 mux8_6.NAND4F_2.D.n12 VSS 0.395829f
C6240 mux8_7.A1.t14 VSS 0.074864f
C6241 mux8_7.A1.t12 VSS 0.072838f
C6242 mux8_7.A1.t13 VSS 0.220572f
C6243 mux8_7.A1.n0 VSS 0.375531f
C6244 mux8_7.A1.t6 VSS 0.021801f
C6245 mux8_7.A1.t7 VSS 0.021801f
C6246 mux8_7.A1.n1 VSS 0.052729f
C6247 mux8_7.A1.t2 VSS 0.021801f
C6248 mux8_7.A1.t1 VSS 0.021801f
C6249 mux8_7.A1.n2 VSS 0.052722f
C6250 mux8_7.A1.n3 VSS 0.378067f
C6251 mux8_7.A1.t8 VSS 0.021801f
C6252 mux8_7.A1.t0 VSS 0.021801f
C6253 mux8_7.A1.n4 VSS 0.043602f
C6254 mux8_7.A1.n5 VSS 0.034251f
C6255 mux8_7.A1.t9 VSS 0.092235f
C6256 mux8_7.A1.t4 VSS 0.092235f
C6257 mux8_7.A1.n6 VSS 0.18447f
C6258 mux8_7.A1.n7 VSS 0.073348f
C6259 mux8_7.A1.t11 VSS 0.092235f
C6260 mux8_7.A1.t10 VSS 0.092235f
C6261 mux8_7.A1.n8 VSS 0.18447f
C6262 mux8_7.A1.n9 VSS 0.081133f
C6263 mux8_7.A1.n10 VSS 0.835311f
C6264 mux8_7.A1.t5 VSS 0.092235f
C6265 mux8_7.A1.t3 VSS 0.092235f
C6266 mux8_7.A1.n11 VSS 0.18447f
C6267 mux8_7.A1.n12 VSS 0.081256f
C6268 mux8_7.A1.n13 VSS 0.535732f
C6269 mux8_7.A1.n14 VSS 0.120733f
C6270 mux8_7.A1.n15 VSS 0.529923f
C6271 OR8_0.S4.n0 VSS 2.44222f
C6272 mux8_5.NAND4F_2.A VSS 1.88441f
C6273 OR8_0.S4.t4 VSS 0.118132f
C6274 OR8_0.S4.t5 VSS 0.114935f
C6275 OR8_0.S4.t6 VSS 0.348052f
C6276 OR8_0.S4.n1 VSS 0.59257f
C6277 mux8_5.A3 VSS 11.416901f
C6278 OR8_0.S4.t2 VSS 0.056629f
C6279 OR8_0.S4.t3 VSS 0.056629f
C6280 OR8_0.S4.n2 VSS 0.126195f
C6281 OR8_0.S4.t1 VSS 0.205394f
C6282 OR8_0.S4.t0 VSS 0.163338f
C6283 OR8_0.NOT8_0.S4 VSS 7.374629f
C6284 mux8_1.NAND4F_0.Y.n0 VSS 0.367143f
C6285 mux8_1.NAND4F_0.Y.t11 VSS 0.02361f
C6286 mux8_1.NAND4F_0.Y.t10 VSS 0.083584f
C6287 mux8_1.NAND4F_0.Y.t9 VSS 0.02599f
C6288 mux8_1.NAND4F_0.Y.n1 VSS 0.074138f
C6289 mux8_1.NAND4F_0.Y.n2 VSS 0.021976f
C6290 mux8_1.NAND4F_0.Y.t5 VSS 0.018101f
C6291 mux8_1.NAND4F_0.Y.t6 VSS 0.018101f
C6292 mux8_1.NAND4F_0.Y.n3 VSS 0.042033f
C6293 mux8_1.NAND4F_0.Y.t3 VSS 0.018101f
C6294 mux8_1.NAND4F_0.Y.t4 VSS 0.018101f
C6295 mux8_1.NAND4F_0.Y.n4 VSS 0.041907f
C6296 mux8_1.NAND4F_0.Y.t7 VSS 0.018101f
C6297 mux8_1.NAND4F_0.Y.t8 VSS 0.018101f
C6298 mux8_1.NAND4F_0.Y.n5 VSS 0.041907f
C6299 mux8_1.NAND4F_0.Y.t1 VSS 0.018101f
C6300 mux8_1.NAND4F_0.Y.t0 VSS 0.018101f
C6301 mux8_1.NAND4F_0.Y.n6 VSS 0.041907f
C6302 mux8_1.NAND4F_0.Y.t2 VSS 0.174248f
C6303 mux8_1.NAND4F_0.C.n0 VSS 2.02061f
C6304 mux8_1.NAND4F_0.C.t12 VSS 0.279708f
C6305 mux8_1.NAND4F_0.C.t13 VSS 0.089224f
C6306 mux8_1.NAND4F_0.C.t15 VSS 0.089224f
C6307 mux8_1.NAND4F_0.C.n1 VSS 0.104752f
C6308 mux8_1.NAND4F_0.C.n2 VSS 0.587326f
C6309 mux8_1.NAND4F_0.C.t6 VSS 0.089224f
C6310 mux8_1.NAND4F_0.C.t4 VSS 0.089224f
C6311 mux8_1.NAND4F_0.C.n3 VSS 0.104752f
C6312 mux8_1.NAND4F_0.C.t7 VSS 0.279708f
C6313 mux8_1.NAND4F_0.C.n4 VSS 0.587363f
C6314 mux8_1.NAND4F_0.C.t10 VSS 0.089224f
C6315 mux8_1.NAND4F_0.C.t8 VSS 0.089224f
C6316 mux8_1.NAND4F_0.C.n5 VSS 0.104752f
C6317 mux8_1.NAND4F_0.C.t5 VSS 0.279708f
C6318 mux8_1.NAND4F_0.C.n6 VSS 0.58738f
C6319 mux8_1.NAND4F_0.C.n7 VSS 2.14221f
C6320 mux8_1.NAND4F_0.C.t3 VSS 0.045462f
C6321 mux8_1.NAND4F_0.C.t2 VSS 0.045462f
C6322 mux8_1.NAND4F_0.C.n8 VSS 0.101309f
C6323 mux8_1.NAND4F_0.C.t1 VSS 0.16489f
C6324 mux8_1.NAND4F_0.C.t0 VSS 0.131127f
C6325 mux8_1.NAND4F_0.C.n9 VSS 3.75062f
C6326 mux8_1.NAND4F_0.C.t14 VSS 0.279708f
C6327 mux8_1.NAND4F_0.C.t9 VSS 0.089224f
C6328 mux8_1.NAND4F_0.C.t11 VSS 0.089224f
C6329 mux8_1.NAND4F_0.C.n10 VSS 0.104752f
C6330 mux8_1.NAND4F_0.C.n11 VSS 0.587347f
C6331 mux8_1.NAND4F_0.C.n12 VSS 3.00573f
C6332 mux8_0.NAND4F_7.Y.n0 VSS 0.11858f
C6333 mux8_0.NAND4F_7.Y.n1 VSS 0.350455f
C6334 mux8_0.NAND4F_7.Y.t4 VSS 0.168166f
C6335 mux8_0.NAND4F_7.Y.t11 VSS 0.022537f
C6336 mux8_0.NAND4F_7.Y.t9 VSS 0.079785f
C6337 mux8_0.NAND4F_7.Y.t10 VSS 0.024808f
C6338 mux8_0.NAND4F_7.Y.n2 VSS 0.070768f
C6339 mux8_0.NAND4F_7.Y.n3 VSS 0.020978f
C6340 mux8_0.NAND4F_7.Y.t1 VSS 0.017278f
C6341 mux8_0.NAND4F_7.Y.t0 VSS 0.017278f
C6342 mux8_0.NAND4F_7.Y.n4 VSS 0.040122f
C6343 mux8_0.NAND4F_7.Y.t3 VSS 0.017278f
C6344 mux8_0.NAND4F_7.Y.t2 VSS 0.017278f
C6345 mux8_0.NAND4F_7.Y.n5 VSS 0.040002f
C6346 mux8_0.NAND4F_7.Y.t7 VSS 0.017278f
C6347 mux8_0.NAND4F_7.Y.t8 VSS 0.017278f
C6348 mux8_0.NAND4F_7.Y.n6 VSS 0.040002f
C6349 mux8_0.NAND4F_7.Y.t6 VSS 0.017278f
C6350 mux8_0.NAND4F_7.Y.t5 VSS 0.017278f
C6351 mux8_0.NAND4F_7.Y.n7 VSS 0.040002f
C6352 a_n20557_n11063.n0 VSS 1.48365f
C6353 a_n20557_n11063.n1 VSS 1.48326f
C6354 a_n20557_n11063.t1 VSS 0.093341f
C6355 a_n20557_n11063.t9 VSS 0.093341f
C6356 a_n20557_n11063.t10 VSS 0.093341f
C6357 a_n20557_n11063.n2 VSS 0.202296f
C6358 a_n20557_n11063.t11 VSS 0.093341f
C6359 a_n20557_n11063.t8 VSS 0.093341f
C6360 a_n20557_n11063.n3 VSS 0.202001f
C6361 a_n20557_n11063.t7 VSS 0.093341f
C6362 a_n20557_n11063.t6 VSS 0.093341f
C6363 a_n20557_n11063.n4 VSS 0.202001f
C6364 a_n20557_n11063.t4 VSS 0.093341f
C6365 a_n20557_n11063.t5 VSS 0.093341f
C6366 a_n20557_n11063.n5 VSS 0.202001f
C6367 a_n20557_n11063.t3 VSS 0.093341f
C6368 a_n20557_n11063.t0 VSS 0.093341f
C6369 a_n20557_n11063.n6 VSS 0.202001f
C6370 a_n20557_n11063.n7 VSS 0.20269f
C6371 a_n20557_n11063.t2 VSS 0.093341f
C6372 MULT_0.inv_15.Y.n0 VSS 0.651777f
C6373 MULT_0.inv_15.Y.t14 VSS 0.020839f
C6374 MULT_0.inv_15.Y.t13 VSS 0.007999f
C6375 MULT_0.inv_15.Y.t15 VSS 0.011046f
C6376 MULT_0.inv_15.Y.n1 VSS 0.012714f
C6377 MULT_0.inv_15.Y.t8 VSS 0.008408f
C6378 MULT_0.inv_15.Y.n2 VSS 0.012894f
C6379 MULT_0.inv_15.Y.n3 VSS 0.053372f
C6380 MULT_0.inv_15.Y.t10 VSS 0.022566f
C6381 MULT_0.inv_15.Y.t5 VSS 0.022285f
C6382 MULT_0.inv_15.Y.t4 VSS 0.022285f
C6383 MULT_0.inv_15.Y.t9 VSS 0.022285f
C6384 MULT_0.inv_15.Y.n4 VSS 0.0887f
C6385 MULT_0.inv_15.Y.t11 VSS 0.004631f
C6386 MULT_0.inv_15.Y.t6 VSS 0.004631f
C6387 MULT_0.inv_15.Y.t7 VSS 0.004631f
C6388 MULT_0.inv_15.Y.t12 VSS 0.004631f
C6389 MULT_0.inv_15.Y.n5 VSS 0.083796f
C6390 MULT_0.inv_15.Y.n6 VSS 0.131073f
C6391 MULT_0.inv_15.Y.t0 VSS 0.019104f
C6392 MULT_0.inv_15.Y.t1 VSS 0.023963f
C6393 MULT_0.inv_15.Y.t3 VSS 0.006607f
C6394 MULT_0.inv_15.Y.t2 VSS 0.006607f
C6395 MULT_0.inv_15.Y.n7 VSS 0.014718f
C6396 MULT_0.4bit_ADDER_0.A0.n0 VSS 4.45631f
C6397 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_0.B VSS 0.77833f
C6398 MULT_0.4bit_ADDER_0.FULL_ADDER_3.A VSS 3.16142f
C6399 MULT_0.4bit_ADDER_0.A0.t4 VSS 0.059295f
C6400 MULT_0.4bit_ADDER_0.A0.t8 VSS 0.02276f
C6401 MULT_0.4bit_ADDER_0.A0.t7 VSS 0.031431f
C6402 MULT_0.4bit_ADDER_0.A0.n1 VSS 0.036177f
C6403 MULT_0.4bit_ADDER_0.A0.t12 VSS 0.023924f
C6404 MULT_0.4bit_ADDER_0.A0.n2 VSS 0.036689f
C6405 MULT_0.4bit_ADDER_0.A0.n3 VSS 0.151863f
C6406 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_0.B VSS 0.586758f
C6407 MULT_0.4bit_ADDER_0.A0.t5 VSS 0.064208f
C6408 MULT_0.4bit_ADDER_0.A0.t13 VSS 0.063409f
C6409 MULT_0.4bit_ADDER_0.A0.t6 VSS 0.063409f
C6410 MULT_0.4bit_ADDER_0.A0.t11 VSS 0.063409f
C6411 MULT_0.4bit_ADDER_0.A0.n4 VSS 0.252386f
C6412 MULT_0.4bit_ADDER_0.A0.t15 VSS 0.013177f
C6413 MULT_0.4bit_ADDER_0.A0.t9 VSS 0.013177f
C6414 MULT_0.4bit_ADDER_0.A0.t14 VSS 0.013177f
C6415 MULT_0.4bit_ADDER_0.A0.t10 VSS 0.013177f
C6416 MULT_0.4bit_ADDER_0.A0.n5 VSS 0.238431f
C6417 MULT_0.4bit_ADDER_0.A0.n6 VSS 0.372955f
C6418 MULT_0.4bit_ADDER_0.A0.n7 VSS 0.882102f
C6419 MULT_0.4bit_ADDER_0.A0.t3 VSS 0.018799f
C6420 MULT_0.4bit_ADDER_0.A0.t2 VSS 0.018799f
C6421 MULT_0.4bit_ADDER_0.A0.n8 VSS 0.041778f
C6422 MULT_0.4bit_ADDER_0.A0.t0 VSS 0.054468f
C6423 MULT_0.4bit_ADDER_0.A0.t1 VSS 0.068184f
C6424 a_n12316_n15299.n0 VSS 1.45527f
C6425 a_n12316_n15299.n1 VSS 1.45566f
C6426 a_n12316_n15299.t1 VSS 0.09158f
C6427 a_n12316_n15299.t11 VSS 0.09158f
C6428 a_n12316_n15299.t10 VSS 0.09158f
C6429 a_n12316_n15299.n2 VSS 0.198865f
C6430 a_n12316_n15299.t6 VSS 0.09158f
C6431 a_n12316_n15299.t9 VSS 0.09158f
C6432 a_n12316_n15299.n3 VSS 0.19819f
C6433 a_n12316_n15299.t8 VSS 0.09158f
C6434 a_n12316_n15299.t7 VSS 0.09158f
C6435 a_n12316_n15299.n4 VSS 0.19819f
C6436 a_n12316_n15299.t5 VSS 0.09158f
C6437 a_n12316_n15299.t3 VSS 0.09158f
C6438 a_n12316_n15299.n5 VSS 0.19819f
C6439 a_n12316_n15299.t0 VSS 0.09158f
C6440 a_n12316_n15299.t4 VSS 0.09158f
C6441 a_n12316_n15299.n6 VSS 0.19819f
C6442 a_n12316_n15299.n7 VSS 0.198479f
C6443 a_n12316_n15299.t2 VSS 0.09158f
C6444 Y6.t6 VSS 0.125015f
C6445 Y6.t5 VSS 0.135076f
C6446 Y6.n0 VSS 0.106706f
C6447 Y6.t7 VSS 0.125731f
C6448 Y6.n1 VSS 0.06046f
C6449 Y6.t4 VSS 0.058232f
C6450 Y6.n2 VSS 0.063129f
C6451 Y6.t2 VSS 0.023393f
C6452 Y6.t1 VSS 0.023393f
C6453 Y6.n3 VSS 0.0521f
C6454 Y6.t3 VSS 0.084846f
C6455 Y6.n4 VSS 0.117803f
C6456 Y6.t0 VSS 0.067568f
C6457 Y6.n5 VSS 0.291739f
C6458 mux8_8.NAND4F_3.Y.n0 VSS 0.306333f
C6459 mux8_8.NAND4F_3.Y.t0 VSS 0.015103f
C6460 mux8_8.NAND4F_3.Y.t6 VSS 0.015103f
C6461 mux8_8.NAND4F_3.Y.n1 VSS 0.035071f
C6462 mux8_8.NAND4F_3.Y.t7 VSS 0.015103f
C6463 mux8_8.NAND4F_3.Y.t8 VSS 0.015103f
C6464 mux8_8.NAND4F_3.Y.n2 VSS 0.034966f
C6465 mux8_8.NAND4F_3.Y.t2 VSS 0.015103f
C6466 mux8_8.NAND4F_3.Y.t1 VSS 0.015103f
C6467 mux8_8.NAND4F_3.Y.n3 VSS 0.034966f
C6468 mux8_8.NAND4F_3.Y.t5 VSS 0.015103f
C6469 mux8_8.NAND4F_3.Y.t3 VSS 0.015103f
C6470 mux8_8.NAND4F_3.Y.n4 VSS 0.034966f
C6471 mux8_8.NAND4F_3.Y.n5 VSS 0.152246f
C6472 mux8_8.NAND4F_3.Y.t4 VSS 0.143521f
C6473 mux8_8.NAND4F_3.Y.t10 VSS 0.0197f
C6474 mux8_8.NAND4F_3.Y.t11 VSS 0.0197f
C6475 mux8_8.NAND4F_3.Y.n6 VSS 0.023128f
C6476 mux8_8.NAND4F_3.Y.t9 VSS 0.061756f
C6477 mux8_8.NAND4F_3.Y.n7 VSS 0.129679f
C6478 mux8_1.NAND4F_5.Y.n0 VSS 0.25108f
C6479 mux8_1.NAND4F_5.Y.t10 VSS 0.017162f
C6480 mux8_1.NAND4F_5.Y.t11 VSS 0.050565f
C6481 mux8_1.NAND4F_5.Y.t9 VSS 0.016698f
C6482 mux8_1.NAND4F_5.Y.n1 VSS 0.086077f
C6483 mux8_1.NAND4F_5.Y.t2 VSS 0.099394f
C6484 mux8_1.NAND4F_5.Y.n2 VSS 0.798124f
C6485 mux8_1.NAND4F_5.Y.t0 VSS 0.012379f
C6486 mux8_1.NAND4F_5.Y.t1 VSS 0.012379f
C6487 mux8_1.NAND4F_5.Y.n3 VSS 0.028745f
C6488 mux8_1.NAND4F_5.Y.t5 VSS 0.012379f
C6489 mux8_1.NAND4F_5.Y.t6 VSS 0.012379f
C6490 mux8_1.NAND4F_5.Y.n4 VSS 0.028659f
C6491 mux8_1.NAND4F_5.Y.t7 VSS 0.012379f
C6492 mux8_1.NAND4F_5.Y.t8 VSS 0.012379f
C6493 mux8_1.NAND4F_5.Y.n5 VSS 0.028659f
C6494 mux8_1.NAND4F_5.Y.t3 VSS 0.012379f
C6495 mux8_1.NAND4F_5.Y.t4 VSS 0.012379f
C6496 mux8_1.NAND4F_5.Y.n6 VSS 0.028659f
C6497 mux8_1.NAND4F_5.Y.n7 VSS 0.117805f
C6498 8bit_ADDER_0.C.n0 VSS 0.2538f
C6499 8bit_ADDER_0.C.t6 VSS 0.002196f
C6500 8bit_ADDER_0.C.t5 VSS 0.002196f
C6501 8bit_ADDER_0.C.n1 VSS 0.0049f
C6502 8bit_ADDER_0.C.t2 VSS 0.002196f
C6503 8bit_ADDER_0.C.t4 VSS 0.002196f
C6504 8bit_ADDER_0.C.n2 VSS 0.004886f
C6505 8bit_ADDER_0.C.t1 VSS 0.002196f
C6506 8bit_ADDER_0.C.t3 VSS 0.002196f
C6507 8bit_ADDER_0.C.n3 VSS 0.004886f
C6508 8bit_ADDER_0.C.t0 VSS 0.013259f
C6509 8bit_ADDER_0.C.t8 VSS 0.004581f
C6510 8bit_ADDER_0.C.t7 VSS 0.004457f
C6511 8bit_ADDER_0.C.t9 VSS 0.013497f
C6512 8bit_ADDER_0.C.n4 VSS 0.022979f
C6513 mux8_2.NAND4F_4.B.n0 VSS 0.921489f
C6514 mux8_2.NAND4F_4.B.t7 VSS 0.03989f
C6515 mux8_2.NAND4F_4.B.t15 VSS 0.123086f
C6516 mux8_2.NAND4F_4.B.t9 VSS 0.04595f
C6517 mux8_2.NAND4F_4.B.n1 VSS 0.154452f
C6518 mux8_2.NAND4F_4.B.n2 VSS 0.033769f
C6519 mux8_2.NAND4F_4.B.t6 VSS 0.03989f
C6520 mux8_2.NAND4F_4.B.t5 VSS 0.123086f
C6521 mux8_2.NAND4F_4.B.t8 VSS 0.04595f
C6522 mux8_2.NAND4F_4.B.n3 VSS 0.154452f
C6523 mux8_2.NAND4F_4.B.n4 VSS 0.032977f
C6524 mux8_2.NAND4F_4.B.t10 VSS 0.03989f
C6525 mux8_2.NAND4F_4.B.t4 VSS 0.123086f
C6526 mux8_2.NAND4F_4.B.t12 VSS 0.04595f
C6527 mux8_2.NAND4F_4.B.n5 VSS 0.154452f
C6528 mux8_2.NAND4F_4.B.n6 VSS 0.033699f
C6529 mux8_2.NAND4F_4.B.n7 VSS 0.612655f
C6530 mux8_2.NAND4F_4.B.t1 VSS 0.020325f
C6531 mux8_2.NAND4F_4.B.t3 VSS 0.020325f
C6532 mux8_2.NAND4F_4.B.n8 VSS 0.045293f
C6533 mux8_2.NAND4F_4.B.t2 VSS 0.073718f
C6534 mux8_2.NAND4F_4.B.t0 VSS 0.058624f
C6535 mux8_2.NAND4F_4.B.n9 VSS 0.607515f
C6536 mux8_2.NAND4F_4.B.t11 VSS 0.03989f
C6537 mux8_2.NAND4F_4.B.t14 VSS 0.123086f
C6538 mux8_2.NAND4F_4.B.t13 VSS 0.04595f
C6539 mux8_2.NAND4F_4.B.n10 VSS 0.154452f
C6540 mux8_2.NAND4F_4.B.n11 VSS 0.033659f
C6541 mux8_2.NAND4F_4.B.n12 VSS 0.776456f
C6542 Y7.t10 VSS 0.052418f
C6543 Y7.t9 VSS 0.052418f
C6544 Y7.t8 VSS 0.056637f
C6545 Y7.n0 VSS 0.046867f
C6546 Y7.n1 VSS 0.035634f
C6547 Y7.t11 VSS 0.018926f
C6548 Y7.n2 VSS 0.035616f
C6549 Y7.n3 VSS 1.7678f
C6550 Y7.t3 VSS 0.009809f
C6551 Y7.t2 VSS 0.009809f
C6552 Y7.n4 VSS 0.021832f
C6553 Y7.n5 VSS 1.71363f
C6554 Y7.t1 VSS 0.035576f
C6555 Y7.n6 VSS 0.097717f
C6556 Y7.t0 VSS 0.028291f
C6557 Y7.n7 VSS 0.147694f
C6558 Y7.t6 VSS 0.019968f
C6559 Y7.t4 VSS 0.0125f
C6560 Y7.t7 VSS 0.017449f
C6561 Y7.t5 VSS 0.017449f
C6562 Y7.n8 VSS 0.056936f
C6563 Y7.n9 VSS 0.093853f
C6564 Y0.t7 VSS 0.029109f
C6565 Y0.t6 VSS 0.080619f
C6566 Y0.t5 VSS 0.080619f
C6567 Y0.t4 VSS 0.087106f
C6568 Y0.n0 VSS 0.07208f
C6569 Y0.n1 VSS 0.054804f
C6570 Y0.n2 VSS 0.054784f
C6571 Y0.t1 VSS 0.015086f
C6572 Y0.t3 VSS 0.015086f
C6573 Y0.n3 VSS 0.03361f
C6574 Y0.t0 VSS 0.043585f
C6575 Y0.t2 VSS 0.054715f
C6576 Y0.n4 VSS 0.226926f
C6577 Y0.n5 VSS 0.269464f
C6578 Y0.n6 VSS 2.67086f
C6579 mux8_2.NAND4F_0.C.n0 VSS 1.71238f
C6580 mux8_2.NAND4F_0.C.t12 VSS 0.23704f
C6581 mux8_2.NAND4F_0.C.t10 VSS 0.075614f
C6582 mux8_2.NAND4F_0.C.t11 VSS 0.075614f
C6583 mux8_2.NAND4F_0.C.n1 VSS 0.088773f
C6584 mux8_2.NAND4F_0.C.n2 VSS 0.497734f
C6585 mux8_2.NAND4F_0.C.t15 VSS 0.075614f
C6586 mux8_2.NAND4F_0.C.t13 VSS 0.075614f
C6587 mux8_2.NAND4F_0.C.n3 VSS 0.088773f
C6588 mux8_2.NAND4F_0.C.t9 VSS 0.23704f
C6589 mux8_2.NAND4F_0.C.n4 VSS 0.497766f
C6590 mux8_2.NAND4F_0.C.t7 VSS 0.075614f
C6591 mux8_2.NAND4F_0.C.t5 VSS 0.075614f
C6592 mux8_2.NAND4F_0.C.n5 VSS 0.088773f
C6593 mux8_2.NAND4F_0.C.t4 VSS 0.23704f
C6594 mux8_2.NAND4F_0.C.n6 VSS 0.49778f
C6595 mux8_2.NAND4F_0.C.n7 VSS 1.81543f
C6596 mux8_2.NAND4F_0.C.t1 VSS 0.038527f
C6597 mux8_2.NAND4F_0.C.t3 VSS 0.038527f
C6598 mux8_2.NAND4F_0.C.n8 VSS 0.085855f
C6599 mux8_2.NAND4F_0.C.t2 VSS 0.139737f
C6600 mux8_2.NAND4F_0.C.t0 VSS 0.111125f
C6601 mux8_2.NAND4F_0.C.n9 VSS 3.17849f
C6602 mux8_2.NAND4F_0.C.t14 VSS 0.23704f
C6603 mux8_2.NAND4F_0.C.t6 VSS 0.075614f
C6604 mux8_2.NAND4F_0.C.t8 VSS 0.075614f
C6605 mux8_2.NAND4F_0.C.n10 VSS 0.088773f
C6606 mux8_2.NAND4F_0.C.n11 VSS 0.497751f
C6607 mux8_2.NAND4F_0.C.n12 VSS 2.54723f
C6608 mux8_0.NAND4F_9.Y.n0 VSS 0.358256f
C6609 mux8_0.NAND4F_9.Y.t13 VSS 0.017853f
C6610 mux8_0.NAND4F_9.Y.t11 VSS 0.017853f
C6611 mux8_0.NAND4F_9.Y.t9 VSS 0.017853f
C6612 mux8_0.NAND4F_9.Y.t14 VSS 0.017853f
C6613 mux8_0.NAND4F_9.Y.t12 VSS 0.022554f
C6614 mux8_0.NAND4F_9.Y.n1 VSS 0.048188f
C6615 mux8_0.NAND4F_9.Y.n2 VSS 0.030339f
C6616 mux8_0.NAND4F_9.Y.n3 VSS 0.030339f
C6617 mux8_0.NAND4F_9.Y.n4 VSS 0.026149f
C6618 mux8_0.NAND4F_9.Y.t10 VSS 0.014813f
C6619 mux8_0.NAND4F_9.Y.n5 VSS 0.021261f
C6620 mux8_0.NAND4F_9.Y.t0 VSS 0.141821f
C6621 mux8_0.NAND4F_9.Y.t7 VSS 0.017663f
C6622 mux8_0.NAND4F_9.Y.t8 VSS 0.017663f
C6623 mux8_0.NAND4F_9.Y.n6 VSS 0.041015f
C6624 mux8_0.NAND4F_9.Y.t3 VSS 0.017663f
C6625 mux8_0.NAND4F_9.Y.t4 VSS 0.017663f
C6626 mux8_0.NAND4F_9.Y.n7 VSS 0.040893f
C6627 mux8_0.NAND4F_9.Y.t6 VSS 0.017663f
C6628 mux8_0.NAND4F_9.Y.t5 VSS 0.017663f
C6629 mux8_0.NAND4F_9.Y.n8 VSS 0.040893f
C6630 mux8_0.NAND4F_9.Y.t2 VSS 0.017663f
C6631 mux8_0.NAND4F_9.Y.t1 VSS 0.017663f
C6632 mux8_0.NAND4F_9.Y.n9 VSS 0.040893f
C6633 mux8_0.NAND4F_9.Y.n10 VSS 0.168091f
C6634 mux8_8.NAND4F_4.B.n0 VSS 0.921489f
C6635 mux8_8.NAND4F_4.B.t7 VSS 0.03989f
C6636 mux8_8.NAND4F_4.B.t9 VSS 0.123086f
C6637 mux8_8.NAND4F_4.B.t5 VSS 0.04595f
C6638 mux8_8.NAND4F_4.B.n1 VSS 0.154452f
C6639 mux8_8.NAND4F_4.B.n2 VSS 0.033769f
C6640 mux8_8.NAND4F_4.B.t12 VSS 0.03989f
C6641 mux8_8.NAND4F_4.B.t13 VSS 0.123086f
C6642 mux8_8.NAND4F_4.B.t11 VSS 0.04595f
C6643 mux8_8.NAND4F_4.B.n3 VSS 0.154452f
C6644 mux8_8.NAND4F_4.B.n4 VSS 0.032977f
C6645 mux8_8.NAND4F_4.B.t8 VSS 0.03989f
C6646 mux8_8.NAND4F_4.B.t10 VSS 0.123086f
C6647 mux8_8.NAND4F_4.B.t6 VSS 0.04595f
C6648 mux8_8.NAND4F_4.B.n5 VSS 0.154452f
C6649 mux8_8.NAND4F_4.B.n6 VSS 0.033699f
C6650 mux8_8.NAND4F_4.B.n7 VSS 0.612655f
C6651 mux8_8.NAND4F_4.B.t3 VSS 0.020325f
C6652 mux8_8.NAND4F_4.B.t2 VSS 0.020325f
C6653 mux8_8.NAND4F_4.B.n8 VSS 0.045293f
C6654 mux8_8.NAND4F_4.B.t1 VSS 0.073718f
C6655 mux8_8.NAND4F_4.B.t0 VSS 0.058624f
C6656 mux8_8.NAND4F_4.B.n9 VSS 0.607515f
C6657 mux8_8.NAND4F_4.B.t15 VSS 0.03989f
C6658 mux8_8.NAND4F_4.B.t4 VSS 0.123086f
C6659 mux8_8.NAND4F_4.B.t14 VSS 0.04595f
C6660 mux8_8.NAND4F_4.B.n10 VSS 0.154452f
C6661 mux8_8.NAND4F_4.B.n11 VSS 0.033659f
C6662 mux8_8.NAND4F_4.B.n12 VSS 0.776456f
C6663 mux8_7.NAND4F_2.D.n0 VSS 0.664607f
C6664 mux8_7.NAND4F_2.D.t6 VSS 0.027742f
C6665 mux8_7.NAND4F_2.D.t7 VSS 0.098211f
C6666 mux8_7.NAND4F_2.D.t4 VSS 0.030538f
C6667 mux8_7.NAND4F_2.D.n1 VSS 0.087112f
C6668 mux8_7.NAND4F_2.D.n2 VSS 0.025808f
C6669 mux8_7.NAND4F_2.D.t3 VSS 0.014135f
C6670 mux8_7.NAND4F_2.D.t2 VSS 0.014135f
C6671 mux8_7.NAND4F_2.D.n3 VSS 0.031499f
C6672 mux8_7.NAND4F_2.D.t1 VSS 0.051268f
C6673 mux8_7.NAND4F_2.D.t0 VSS 0.040771f
C6674 mux8_7.NAND4F_2.D.t15 VSS 0.027742f
C6675 mux8_7.NAND4F_2.D.t5 VSS 0.098211f
C6676 mux8_7.NAND4F_2.D.t10 VSS 0.030538f
C6677 mux8_7.NAND4F_2.D.n4 VSS 0.087112f
C6678 mux8_7.NAND4F_2.D.n5 VSS 0.025813f
C6679 mux8_7.NAND4F_2.D.n6 VSS 0.620222f
C6680 mux8_7.NAND4F_2.D.t14 VSS 0.027742f
C6681 mux8_7.NAND4F_2.D.t8 VSS 0.098211f
C6682 mux8_7.NAND4F_2.D.t13 VSS 0.030538f
C6683 mux8_7.NAND4F_2.D.n7 VSS 0.087112f
C6684 mux8_7.NAND4F_2.D.n8 VSS 0.025807f
C6685 mux8_7.NAND4F_2.D.n9 VSS 0.261852f
C6686 mux8_7.NAND4F_2.D.t11 VSS 0.027742f
C6687 mux8_7.NAND4F_2.D.t12 VSS 0.098211f
C6688 mux8_7.NAND4F_2.D.t9 VSS 0.030538f
C6689 mux8_7.NAND4F_2.D.n10 VSS 0.087112f
C6690 mux8_7.NAND4F_2.D.n11 VSS 0.025808f
C6691 mux8_7.NAND4F_2.D.n12 VSS 0.407824f
C6692 mux8_0.NAND4F_1.Y.n0 VSS 0.655599f
C6693 mux8_0.NAND4F_1.Y.t6 VSS 0.306614f
C6694 mux8_0.NAND4F_1.Y.t9 VSS 0.132168f
C6695 mux8_0.NAND4F_1.Y.t10 VSS 0.04216f
C6696 mux8_0.NAND4F_1.Y.t11 VSS 0.04216f
C6697 mux8_0.NAND4F_1.Y.n1 VSS 0.049498f
C6698 mux8_0.NAND4F_1.Y.n2 VSS 0.277534f
C6699 mux8_0.NAND4F_1.Y.t1 VSS 0.032323f
C6700 mux8_0.NAND4F_1.Y.t0 VSS 0.032323f
C6701 mux8_0.NAND4F_1.Y.n3 VSS 0.075057f
C6702 mux8_0.NAND4F_1.Y.t5 VSS 0.032323f
C6703 mux8_0.NAND4F_1.Y.t4 VSS 0.032323f
C6704 mux8_0.NAND4F_1.Y.n4 VSS 0.074832f
C6705 mux8_0.NAND4F_1.Y.t3 VSS 0.032323f
C6706 mux8_0.NAND4F_1.Y.t2 VSS 0.032323f
C6707 mux8_0.NAND4F_1.Y.n5 VSS 0.074832f
C6708 mux8_0.NAND4F_1.Y.t8 VSS 0.032323f
C6709 mux8_0.NAND4F_1.Y.t7 VSS 0.032323f
C6710 mux8_0.NAND4F_1.Y.n6 VSS 0.074832f
C6711 mux8_0.NAND4F_1.Y.n7 VSS 0.307603f
C6712 a_n12314_n31661.n0 VSS 1.48326f
C6713 a_n12314_n31661.n1 VSS 1.48365f
C6714 a_n12314_n31661.t0 VSS 0.093341f
C6715 a_n12314_n31661.t5 VSS 0.093341f
C6716 a_n12314_n31661.t4 VSS 0.093341f
C6717 a_n12314_n31661.n2 VSS 0.20269f
C6718 a_n12314_n31661.t9 VSS 0.093341f
C6719 a_n12314_n31661.t3 VSS 0.093341f
C6720 a_n12314_n31661.n3 VSS 0.202001f
C6721 a_n12314_n31661.t11 VSS 0.093341f
C6722 a_n12314_n31661.t10 VSS 0.093341f
C6723 a_n12314_n31661.n4 VSS 0.202001f
C6724 a_n12314_n31661.t7 VSS 0.093341f
C6725 a_n12314_n31661.t6 VSS 0.093341f
C6726 a_n12314_n31661.n5 VSS 0.202001f
C6727 a_n12314_n31661.t1 VSS 0.093341f
C6728 a_n12314_n31661.t8 VSS 0.093341f
C6729 a_n12314_n31661.n6 VSS 0.202001f
C6730 a_n12314_n31661.n7 VSS 0.202296f
C6731 a_n12314_n31661.t2 VSS 0.093341f
C6732 mux8_7.NAND4F_0.Y.n0 VSS 0.350455f
C6733 mux8_7.NAND4F_0.Y.t10 VSS 0.022537f
C6734 mux8_7.NAND4F_0.Y.t9 VSS 0.079785f
C6735 mux8_7.NAND4F_0.Y.t11 VSS 0.024808f
C6736 mux8_7.NAND4F_0.Y.n1 VSS 0.070768f
C6737 mux8_7.NAND4F_0.Y.n2 VSS 0.020978f
C6738 mux8_7.NAND4F_0.Y.t7 VSS 0.017278f
C6739 mux8_7.NAND4F_0.Y.t8 VSS 0.017278f
C6740 mux8_7.NAND4F_0.Y.n3 VSS 0.040122f
C6741 mux8_7.NAND4F_0.Y.t1 VSS 0.017278f
C6742 mux8_7.NAND4F_0.Y.t0 VSS 0.017278f
C6743 mux8_7.NAND4F_0.Y.n4 VSS 0.040002f
C6744 mux8_7.NAND4F_0.Y.t6 VSS 0.017278f
C6745 mux8_7.NAND4F_0.Y.t5 VSS 0.017278f
C6746 mux8_7.NAND4F_0.Y.n5 VSS 0.040002f
C6747 mux8_7.NAND4F_0.Y.t4 VSS 0.017278f
C6748 mux8_7.NAND4F_0.Y.t2 VSS 0.017278f
C6749 mux8_7.NAND4F_0.Y.n6 VSS 0.040002f
C6750 mux8_7.NAND4F_0.Y.t3 VSS 0.166327f
C6751 a_n7496_3810.n0 VSS 1.45527f
C6752 a_n7496_3810.n1 VSS 1.45566f
C6753 a_n7496_3810.t4 VSS 0.09158f
C6754 a_n7496_3810.t9 VSS 0.09158f
C6755 a_n7496_3810.t10 VSS 0.09158f
C6756 a_n7496_3810.n2 VSS 0.198865f
C6757 a_n7496_3810.t11 VSS 0.09158f
C6758 a_n7496_3810.t7 VSS 0.09158f
C6759 a_n7496_3810.n3 VSS 0.19819f
C6760 a_n7496_3810.t8 VSS 0.09158f
C6761 a_n7496_3810.t6 VSS 0.09158f
C6762 a_n7496_3810.n4 VSS 0.19819f
C6763 a_n7496_3810.t5 VSS 0.09158f
C6764 a_n7496_3810.t3 VSS 0.09158f
C6765 a_n7496_3810.n5 VSS 0.19819f
C6766 a_n7496_3810.t0 VSS 0.09158f
C6767 a_n7496_3810.t1 VSS 0.09158f
C6768 a_n7496_3810.n6 VSS 0.198479f
C6769 a_n7496_3810.n7 VSS 0.19819f
C6770 a_n7496_3810.t2 VSS 0.09158f
C6771 a_n19774_2026.n0 VSS 1.48326f
C6772 a_n19774_2026.n1 VSS 1.48365f
C6773 a_n19774_2026.t1 VSS 0.093341f
C6774 a_n19774_2026.t0 VSS 0.093341f
C6775 a_n19774_2026.t10 VSS 0.093341f
C6776 a_n19774_2026.n2 VSS 0.20269f
C6777 a_n19774_2026.t7 VSS 0.093341f
C6778 a_n19774_2026.t9 VSS 0.093341f
C6779 a_n19774_2026.n3 VSS 0.202001f
C6780 a_n19774_2026.t11 VSS 0.093341f
C6781 a_n19774_2026.t8 VSS 0.093341f
C6782 a_n19774_2026.n4 VSS 0.202001f
C6783 a_n19774_2026.t4 VSS 0.093341f
C6784 a_n19774_2026.t6 VSS 0.093341f
C6785 a_n19774_2026.n5 VSS 0.202001f
C6786 a_n19774_2026.t2 VSS 0.093341f
C6787 a_n19774_2026.t5 VSS 0.093341f
C6788 a_n19774_2026.n6 VSS 0.202001f
C6789 a_n19774_2026.n7 VSS 0.202296f
C6790 a_n19774_2026.t3 VSS 0.093341f
C6791 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n0 VSS 0.860417f
C6792 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t1 VSS 0.007445f
C6793 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t0 VSS 0.007445f
C6794 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n1 VSS 0.016611f
C6795 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t5 VSS 0.007445f
C6796 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t2 VSS 0.007445f
C6797 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n2 VSS 0.016566f
C6798 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t4 VSS 0.007445f
C6799 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t6 VSS 0.007445f
C6800 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n3 VSS 0.016566f
C6801 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t3 VSS 0.044951f
C6802 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t11 VSS 0.025427f
C6803 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t17 VSS 0.025111f
C6804 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t9 VSS 0.025111f
C6805 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t7 VSS 0.025111f
C6806 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n4 VSS 0.099949f
C6807 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t18 VSS 0.005218f
C6808 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t15 VSS 0.005218f
C6809 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t8 VSS 0.005218f
C6810 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t10 VSS 0.005218f
C6811 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n5 VSS 0.094423f
C6812 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n6 VSS 0.147672f
C6813 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t12 VSS 0.023482f
C6814 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t13 VSS 0.009013f
C6815 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t14 VSS 0.012447f
C6816 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n7 VSS 0.014327f
C6817 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.t16 VSS 0.009474f
C6818 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n8 VSS 0.014529f
C6819 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n9 VSS 0.049349f
C6820 8bit_ADDER_0.FULL_ADDER_XORED_2.COUT.n10 VSS 0.328172f
C6821 MULT_0.NAND2_4.Y.n0 VSS 1.19194f
C6822 MULT_0.NAND2_4.Y.n1 VSS 0.186659f
C6823 MULT_0.NAND2_4.Y.t6 VSS 0.022992f
C6824 MULT_0.NAND2_4.Y.t5 VSS 0.022992f
C6825 MULT_0.NAND2_4.Y.n2 VSS 0.0513f
C6826 MULT_0.NAND2_4.Y.t2 VSS 0.022992f
C6827 MULT_0.NAND2_4.Y.t4 VSS 0.022992f
C6828 MULT_0.NAND2_4.Y.n3 VSS 0.051161f
C6829 MULT_0.NAND2_4.Y.t3 VSS 0.022992f
C6830 MULT_0.NAND2_4.Y.t1 VSS 0.022992f
C6831 MULT_0.NAND2_4.Y.n4 VSS 0.051161f
C6832 MULT_0.NAND2_4.Y.t0 VSS 0.138509f
C6833 MULT_0.NAND2_4.Y.t9 VSS 0.029302f
C6834 MULT_0.NAND2_4.Y.t8 VSS 0.040903f
C6835 MULT_0.NAND2_4.Y.t10 VSS 0.040903f
C6836 MULT_0.NAND2_4.Y.n5 VSS 0.13351f
C6837 MULT_0.NAND2_4.Y.t7 VSS 0.046701f
C6838 mux8_8.NAND4F_4.Y.n0 VSS 0.480308f
C6839 mux8_8.NAND4F_4.Y.t3 VSS 0.023681f
C6840 mux8_8.NAND4F_4.Y.t4 VSS 0.023681f
C6841 mux8_8.NAND4F_4.Y.n1 VSS 0.054989f
C6842 mux8_8.NAND4F_4.Y.t5 VSS 0.023681f
C6843 mux8_8.NAND4F_4.Y.t6 VSS 0.023681f
C6844 mux8_8.NAND4F_4.Y.n2 VSS 0.054824f
C6845 mux8_8.NAND4F_4.Y.t7 VSS 0.023681f
C6846 mux8_8.NAND4F_4.Y.t8 VSS 0.023681f
C6847 mux8_8.NAND4F_4.Y.n3 VSS 0.054824f
C6848 mux8_8.NAND4F_4.Y.t0 VSS 0.023681f
C6849 mux8_8.NAND4F_4.Y.t1 VSS 0.023681f
C6850 mux8_8.NAND4F_4.Y.n4 VSS 0.054824f
C6851 mux8_8.NAND4F_4.Y.n5 VSS 0.238711f
C6852 mux8_8.NAND4F_4.Y.t10 VSS 0.032831f
C6853 mux8_8.NAND4F_4.Y.t11 VSS 0.031942f
C6854 mux8_8.NAND4F_4.Y.t9 VSS 0.096729f
C6855 mux8_8.NAND4F_4.Y.n6 VSS 0.164667f
C6856 mux8_8.NAND4F_4.Y.t2 VSS 0.190137f
C6857 mux8_8.NAND4F_4.Y.n7 VSS 1.51729f
C6858 mux8_4.A1.t14 VSS 0.046446f
C6859 mux8_4.A1.t13 VSS 0.045189f
C6860 mux8_4.A1.t12 VSS 0.136842f
C6861 mux8_4.A1.n0 VSS 0.232979f
C6862 mux8_4.A1.t3 VSS 0.013525f
C6863 mux8_4.A1.t4 VSS 0.013525f
C6864 mux8_4.A1.n1 VSS 0.032713f
C6865 mux8_4.A1.t11 VSS 0.013525f
C6866 mux8_4.A1.t9 VSS 0.013525f
C6867 mux8_4.A1.n2 VSS 0.032709f
C6868 mux8_4.A1.n3 VSS 0.234552f
C6869 mux8_4.A1.t5 VSS 0.013525f
C6870 mux8_4.A1.t10 VSS 0.013525f
C6871 mux8_4.A1.n4 VSS 0.027051f
C6872 mux8_4.A1.n5 VSS 0.021249f
C6873 mux8_4.A1.t0 VSS 0.057222f
C6874 mux8_4.A1.t7 VSS 0.057222f
C6875 mux8_4.A1.n6 VSS 0.114445f
C6876 mux8_4.A1.n7 VSS 0.045505f
C6877 mux8_4.A1.t2 VSS 0.057222f
C6878 mux8_4.A1.t1 VSS 0.057222f
C6879 mux8_4.A1.n8 VSS 0.114445f
C6880 mux8_4.A1.n9 VSS 0.050335f
C6881 mux8_4.A1.n10 VSS 0.518225f
C6882 mux8_4.A1.t8 VSS 0.057222f
C6883 mux8_4.A1.t6 VSS 0.057222f
C6884 mux8_4.A1.n11 VSS 0.114445f
C6885 mux8_4.A1.n12 VSS 0.050411f
C6886 mux8_4.A1.n13 VSS 0.332367f
C6887 mux8_4.A1.n14 VSS 0.074903f
C6888 mux8_4.A1.n15 VSS 0.328763f
C6889 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n0 VSS 0.887305f
C6890 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t6 VSS 0.007677f
C6891 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t5 VSS 0.007677f
C6892 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n1 VSS 0.01713f
C6893 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t2 VSS 0.007677f
C6894 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t4 VSS 0.007677f
C6895 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n2 VSS 0.017083f
C6896 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t3 VSS 0.007677f
C6897 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t1 VSS 0.007677f
C6898 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n3 VSS 0.017083f
C6899 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t0 VSS 0.046356f
C6900 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t10 VSS 0.026222f
C6901 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t8 VSS 0.025896f
C6902 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t17 VSS 0.025896f
C6903 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t9 VSS 0.025896f
C6904 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n4 VSS 0.103072f
C6905 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t12 VSS 0.005381f
C6906 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t18 VSS 0.005381f
C6907 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t7 VSS 0.005381f
C6908 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t15 VSS 0.005381f
C6909 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n5 VSS 0.097373f
C6910 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n6 VSS 0.152286f
C6911 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t11 VSS 0.024216f
C6912 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t13 VSS 0.009295f
C6913 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t16 VSS 0.012836f
C6914 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n7 VSS 0.014774f
C6915 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.t14 VSS 0.00977f
C6916 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n8 VSS 0.014983f
C6917 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n9 VSS 0.050891f
C6918 8bit_ADDER_0.FULL_ADDER_XORED_1.COUT.n10 VSS 0.338427f
C6919 right_shifter_0.S4.n0 VSS 3.45602f
C6920 mux8_5.NAND4F_6.A VSS 0.508231f
C6921 right_shifter_0.S4.t5 VSS 0.038847f
C6922 right_shifter_0.S4.t4 VSS 0.114454f
C6923 right_shifter_0.S4.t6 VSS 0.037795f
C6924 right_shifter_0.S4.n1 VSS 0.194861f
C6925 right_shifter_0.S4.t3 VSS 0.018622f
C6926 right_shifter_0.S4.t2 VSS 0.018622f
C6927 right_shifter_0.S4.n2 VSS 0.041498f
C6928 right_shifter_0.S4.t1 VSS 0.067542f
C6929 right_shifter_0.S4.t0 VSS 0.053712f
C6930 mux8_5.A7 VSS 3.1498f
C6931 MULT_0.inv_7.A.n0 VSS 1.19272f
C6932 MULT_0.inv_7.A.n1 VSS 0.186498f
C6933 MULT_0.inv_7.A.t3 VSS 0.13839f
C6934 MULT_0.inv_7.A.t4 VSS 0.022972f
C6935 MULT_0.inv_7.A.t5 VSS 0.022972f
C6936 MULT_0.inv_7.A.n2 VSS 0.051117f
C6937 MULT_0.inv_7.A.t1 VSS 0.022972f
C6938 MULT_0.inv_7.A.t0 VSS 0.022972f
C6939 MULT_0.inv_7.A.n3 VSS 0.051256f
C6940 MULT_0.inv_7.A.t6 VSS 0.022972f
C6941 MULT_0.inv_7.A.t2 VSS 0.022972f
C6942 MULT_0.inv_7.A.n4 VSS 0.051117f
C6943 MULT_0.inv_7.A.t7 VSS 0.029277f
C6944 MULT_0.inv_7.A.t10 VSS 0.040868f
C6945 MULT_0.inv_7.A.t8 VSS 0.040868f
C6946 MULT_0.inv_7.A.n5 VSS 0.133396f
C6947 MULT_0.inv_7.A.t9 VSS 0.046661f
C6948 mux8_5.A0.t12 VSS 0.077554f
C6949 mux8_5.A0.t13 VSS 0.075455f
C6950 mux8_5.A0.t14 VSS 0.228497f
C6951 mux8_5.A0.n0 VSS 0.389023f
C6952 mux8_5.A0.t2 VSS 0.022584f
C6953 mux8_5.A0.t0 VSS 0.022584f
C6954 mux8_5.A0.n1 VSS 0.054623f
C6955 mux8_5.A0.t4 VSS 0.022584f
C6956 mux8_5.A0.t5 VSS 0.022584f
C6957 mux8_5.A0.n2 VSS 0.054617f
C6958 mux8_5.A0.n3 VSS 0.39165f
C6959 mux8_5.A0.t1 VSS 0.022584f
C6960 mux8_5.A0.t3 VSS 0.022584f
C6961 mux8_5.A0.n4 VSS 0.045168f
C6962 mux8_5.A0.n5 VSS 0.035481f
C6963 mux8_5.A0.t10 VSS 0.095549f
C6964 mux8_5.A0.t8 VSS 0.095549f
C6965 mux8_5.A0.n6 VSS 0.191098f
C6966 mux8_5.A0.n7 VSS 0.075984f
C6967 mux8_5.A0.t11 VSS 0.095549f
C6968 mux8_5.A0.t9 VSS 0.095549f
C6969 mux8_5.A0.n8 VSS 0.191098f
C6970 mux8_5.A0.n9 VSS 0.084048f
C6971 mux8_5.A0.n10 VSS 0.865322f
C6972 mux8_5.A0.t6 VSS 0.095549f
C6973 mux8_5.A0.t7 VSS 0.095549f
C6974 mux8_5.A0.n11 VSS 0.191098f
C6975 mux8_5.A0.n12 VSS 0.084175f
C6976 mux8_5.A0.n13 VSS 0.55498f
C6977 mux8_5.A0.n14 VSS 0.125071f
C6978 mux8_5.A0.n15 VSS 0.548962f
C6979 MULT_0.inv_6.A.n0 VSS 1.19194f
C6980 MULT_0.inv_6.A.n1 VSS 0.186659f
C6981 MULT_0.inv_6.A.t3 VSS 0.138509f
C6982 MULT_0.inv_6.A.t6 VSS 0.022992f
C6983 MULT_0.inv_6.A.t5 VSS 0.022992f
C6984 MULT_0.inv_6.A.n2 VSS 0.0513f
C6985 MULT_0.inv_6.A.t1 VSS 0.022992f
C6986 MULT_0.inv_6.A.t4 VSS 0.022992f
C6987 MULT_0.inv_6.A.n3 VSS 0.051161f
C6988 MULT_0.inv_6.A.t2 VSS 0.022992f
C6989 MULT_0.inv_6.A.t0 VSS 0.022992f
C6990 MULT_0.inv_6.A.n4 VSS 0.051161f
C6991 MULT_0.inv_6.A.t9 VSS 0.029302f
C6992 MULT_0.inv_6.A.t8 VSS 0.040903f
C6993 MULT_0.inv_6.A.t10 VSS 0.040903f
C6994 MULT_0.inv_6.A.n5 VSS 0.13351f
C6995 MULT_0.inv_6.A.t7 VSS 0.046701f
C6996 mux8_3.NAND4F_4.B.n0 VSS 0.921489f
C6997 mux8_3.NAND4F_4.B.t14 VSS 0.03989f
C6998 mux8_3.NAND4F_4.B.t15 VSS 0.123086f
C6999 mux8_3.NAND4F_4.B.t13 VSS 0.04595f
C7000 mux8_3.NAND4F_4.B.n1 VSS 0.154452f
C7001 mux8_3.NAND4F_4.B.n2 VSS 0.033769f
C7002 mux8_3.NAND4F_4.B.t11 VSS 0.03989f
C7003 mux8_3.NAND4F_4.B.t9 VSS 0.123086f
C7004 mux8_3.NAND4F_4.B.t10 VSS 0.04595f
C7005 mux8_3.NAND4F_4.B.n3 VSS 0.154452f
C7006 mux8_3.NAND4F_4.B.n4 VSS 0.032977f
C7007 mux8_3.NAND4F_4.B.t6 VSS 0.03989f
C7008 mux8_3.NAND4F_4.B.t4 VSS 0.123086f
C7009 mux8_3.NAND4F_4.B.t5 VSS 0.04595f
C7010 mux8_3.NAND4F_4.B.n5 VSS 0.154452f
C7011 mux8_3.NAND4F_4.B.n6 VSS 0.033699f
C7012 mux8_3.NAND4F_4.B.n7 VSS 0.612655f
C7013 mux8_3.NAND4F_4.B.t3 VSS 0.020325f
C7014 mux8_3.NAND4F_4.B.t2 VSS 0.020325f
C7015 mux8_3.NAND4F_4.B.n8 VSS 0.045293f
C7016 mux8_3.NAND4F_4.B.t1 VSS 0.073718f
C7017 mux8_3.NAND4F_4.B.t0 VSS 0.058624f
C7018 mux8_3.NAND4F_4.B.n9 VSS 0.607515f
C7019 mux8_3.NAND4F_4.B.t8 VSS 0.03989f
C7020 mux8_3.NAND4F_4.B.t12 VSS 0.123086f
C7021 mux8_3.NAND4F_4.B.t7 VSS 0.04595f
C7022 mux8_3.NAND4F_4.B.n10 VSS 0.154452f
C7023 mux8_3.NAND4F_4.B.n11 VSS 0.033659f
C7024 mux8_3.NAND4F_4.B.n12 VSS 0.776456f
C7025 right_shifter_0.C.n0 VSS 3.26408f
C7026 mux8_0.NAND4F_6.A VSS 0.322623f
C7027 right_shifter_0.C.t4 VSS 0.02444f
C7028 right_shifter_0.C.t6 VSS 0.072006f
C7029 right_shifter_0.C.t5 VSS 0.023778f
C7030 right_shifter_0.C.n1 VSS 0.122592f
C7031 right_shifter_0.C.t1 VSS 0.011716f
C7032 right_shifter_0.C.t2 VSS 0.011716f
C7033 right_shifter_0.C.n2 VSS 0.026107f
C7034 right_shifter_0.C.t3 VSS 0.042492f
C7035 right_shifter_0.C.t0 VSS 0.033792f
C7036 mux8_0.A7 VSS 3.74466f
C7037 mux8_6.NAND4F_6.Y.n0 VSS 0.599344f
C7038 mux8_6.NAND4F_6.Y.t2 VSS 0.244548f
C7039 mux8_6.NAND4F_6.Y.t11 VSS 0.038543f
C7040 mux8_6.NAND4F_6.Y.t9 VSS 0.118929f
C7041 mux8_6.NAND4F_6.Y.t10 VSS 0.044398f
C7042 mux8_6.NAND4F_6.Y.n1 VSS 0.149236f
C7043 mux8_6.NAND4F_6.Y.n2 VSS 0.032396f
C7044 mux8_6.NAND4F_6.Y.n3 VSS 1.72835f
C7045 mux8_6.NAND4F_6.Y.t1 VSS 0.029549f
C7046 mux8_6.NAND4F_6.Y.t0 VSS 0.029549f
C7047 mux8_6.NAND4F_6.Y.n4 VSS 0.068617f
C7048 mux8_6.NAND4F_6.Y.t6 VSS 0.029549f
C7049 mux8_6.NAND4F_6.Y.t5 VSS 0.029549f
C7050 mux8_6.NAND4F_6.Y.n5 VSS 0.068411f
C7051 mux8_6.NAND4F_6.Y.t7 VSS 0.029549f
C7052 mux8_6.NAND4F_6.Y.t8 VSS 0.029549f
C7053 mux8_6.NAND4F_6.Y.n6 VSS 0.068411f
C7054 mux8_6.NAND4F_6.Y.t4 VSS 0.029549f
C7055 mux8_6.NAND4F_6.Y.t3 VSS 0.029549f
C7056 mux8_6.NAND4F_6.Y.n7 VSS 0.068411f
C7057 mux8_6.NAND4F_6.Y.n8 VSS 0.281208f
C7058 right_shifter_0.S7.n0 VSS 3.57377f
C7059 mux8_6.NAND4F_6.A VSS 0.300721f
C7060 right_shifter_0.S7.t5 VSS 0.02278f
C7061 right_shifter_0.S7.t4 VSS 0.067118f
C7062 right_shifter_0.S7.t6 VSS 0.022164f
C7063 right_shifter_0.S7.n1 VSS 0.11427f
C7064 right_shifter_0.S7.t3 VSS 0.01092f
C7065 right_shifter_0.S7.t2 VSS 0.01092f
C7066 right_shifter_0.S7.n2 VSS 0.024335f
C7067 right_shifter_0.S7.t1 VSS 0.039608f
C7068 right_shifter_0.S7.t0 VSS 0.031498f
C7069 mux8_6.A7 VSS 2.9819f
C7070 mux8_6.A1.n0 VSS 1.56671f
C7071 mux8_6.A1.t7 VSS 0.028292f
C7072 mux8_6.A1.t9 VSS 0.027526f
C7073 mux8_6.A1.t8 VSS 0.083357f
C7074 mux8_6.A1.n1 VSS 0.141918f
C7075 mux8_6.A1.t5 VSS 0.013562f
C7076 mux8_6.A1.t6 VSS 0.013562f
C7077 mux8_6.A1.n2 VSS 0.030261f
C7078 mux8_6.A1.t2 VSS 0.013562f
C7079 mux8_6.A1.t4 VSS 0.013562f
C7080 mux8_6.A1.n3 VSS 0.030179f
C7081 mux8_6.A1.t1 VSS 0.013562f
C7082 mux8_6.A1.t3 VSS 0.013562f
C7083 mux8_6.A1.n4 VSS 0.030179f
C7084 mux8_6.A1.t0 VSS 0.08189f
C7085 XOR8_0.S7.t12 VSS 0.030249f
C7086 XOR8_0.S7.t14 VSS 0.089121f
C7087 XOR8_0.S7.t13 VSS 0.02943f
C7088 XOR8_0.S7.n0 VSS 0.151723f
C7089 XOR8_0.S7.t10 VSS 0.008809f
C7090 XOR8_0.S7.t9 VSS 0.008809f
C7091 XOR8_0.S7.n1 VSS 0.021305f
C7092 XOR8_0.S7.t6 VSS 0.008809f
C7093 XOR8_0.S7.t8 VSS 0.008809f
C7094 XOR8_0.S7.n2 VSS 0.021302f
C7095 XOR8_0.S7.n3 VSS 0.152757f
C7096 XOR8_0.S7.t11 VSS 0.008809f
C7097 XOR8_0.S7.t7 VSS 0.008809f
C7098 XOR8_0.S7.n4 VSS 0.017617f
C7099 XOR8_0.S7.n5 VSS 0.013839f
C7100 XOR8_0.S7.t2 VSS 0.037267f
C7101 XOR8_0.S7.t5 VSS 0.037267f
C7102 XOR8_0.S7.n6 VSS 0.074534f
C7103 XOR8_0.S7.n7 VSS 0.029566f
C7104 XOR8_0.S7.t0 VSS 0.037267f
C7105 XOR8_0.S7.t1 VSS 0.037267f
C7106 XOR8_0.S7.n8 VSS 0.074534f
C7107 XOR8_0.S7.n9 VSS 0.032782f
C7108 XOR8_0.S7.n10 VSS 0.337505f
C7109 XOR8_0.S7.t4 VSS 0.037267f
C7110 XOR8_0.S7.t3 VSS 0.037267f
C7111 XOR8_0.S7.n11 VSS 0.074534f
C7112 XOR8_0.S7.n12 VSS 0.032831f
C7113 XOR8_0.S7.n13 VSS 0.216461f
C7114 XOR8_0.S7.n14 VSS 0.048722f
C7115 XOR8_0.S7.n15 VSS 0.214243f
C7116 mux8_5.NAND4F_2.D.n0 VSS 0.664607f
C7117 mux8_5.NAND4F_2.D.t15 VSS 0.027742f
C7118 mux8_5.NAND4F_2.D.t11 VSS 0.098211f
C7119 mux8_5.NAND4F_2.D.t14 VSS 0.030538f
C7120 mux8_5.NAND4F_2.D.n1 VSS 0.087112f
C7121 mux8_5.NAND4F_2.D.n2 VSS 0.025808f
C7122 mux8_5.NAND4F_2.D.t1 VSS 0.014135f
C7123 mux8_5.NAND4F_2.D.t3 VSS 0.014135f
C7124 mux8_5.NAND4F_2.D.n3 VSS 0.031499f
C7125 mux8_5.NAND4F_2.D.t2 VSS 0.051268f
C7126 mux8_5.NAND4F_2.D.t0 VSS 0.040771f
C7127 mux8_5.NAND4F_2.D.t13 VSS 0.027742f
C7128 mux8_5.NAND4F_2.D.t7 VSS 0.098211f
C7129 mux8_5.NAND4F_2.D.t6 VSS 0.030538f
C7130 mux8_5.NAND4F_2.D.n4 VSS 0.087112f
C7131 mux8_5.NAND4F_2.D.n5 VSS 0.025813f
C7132 mux8_5.NAND4F_2.D.n6 VSS 0.620222f
C7133 mux8_5.NAND4F_2.D.t10 VSS 0.027742f
C7134 mux8_5.NAND4F_2.D.t12 VSS 0.098211f
C7135 mux8_5.NAND4F_2.D.t9 VSS 0.030538f
C7136 mux8_5.NAND4F_2.D.n7 VSS 0.087112f
C7137 mux8_5.NAND4F_2.D.n8 VSS 0.025807f
C7138 mux8_5.NAND4F_2.D.n9 VSS 0.261852f
C7139 mux8_5.NAND4F_2.D.t8 VSS 0.027742f
C7140 mux8_5.NAND4F_2.D.t4 VSS 0.098211f
C7141 mux8_5.NAND4F_2.D.t5 VSS 0.030538f
C7142 mux8_5.NAND4F_2.D.n10 VSS 0.087112f
C7143 mux8_5.NAND4F_2.D.n11 VSS 0.025808f
C7144 mux8_5.NAND4F_2.D.n12 VSS 0.407824f
C7145 a_1887_5534.n0 VSS 1.45566f
C7146 a_1887_5534.n1 VSS 1.45527f
C7147 a_1887_5534.t0 VSS 0.09158f
C7148 a_1887_5534.t7 VSS 0.09158f
C7149 a_1887_5534.t6 VSS 0.09158f
C7150 a_1887_5534.n2 VSS 0.198479f
C7151 a_1887_5534.t8 VSS 0.09158f
C7152 a_1887_5534.t9 VSS 0.09158f
C7153 a_1887_5534.n3 VSS 0.19819f
C7154 a_1887_5534.t10 VSS 0.09158f
C7155 a_1887_5534.t11 VSS 0.09158f
C7156 a_1887_5534.n4 VSS 0.19819f
C7157 a_1887_5534.t4 VSS 0.09158f
C7158 a_1887_5534.t5 VSS 0.09158f
C7159 a_1887_5534.n5 VSS 0.19819f
C7160 a_1887_5534.t2 VSS 0.09158f
C7161 a_1887_5534.t1 VSS 0.09158f
C7162 a_1887_5534.n6 VSS 0.198865f
C7163 a_1887_5534.n7 VSS 0.19819f
C7164 a_1887_5534.t3 VSS 0.09158f
C7165 B7.t30 VSS 0.044159f
C7166 B7.t40 VSS 0.088849f
C7167 B7.t19 VSS 0.087744f
C7168 B7.t14 VSS 0.087744f
C7169 B7.t1 VSS 0.087744f
C7170 B7.t18 VSS 0.018234f
C7171 B7.t35 VSS 0.018234f
C7172 B7.t26 VSS 0.018234f
C7173 B7.n0 VSS 0.540583f
C7174 B7.n1 VSS 0.398164f
C7175 B7.n2 VSS 0.216996f
C7176 B7.n3 VSS 0.21318f
C7177 B7.n4 VSS 0.13113f
C7178 B7.n5 VSS 0.149122f
C7179 B7.n6 VSS 0.227034f
C7180 B7.t6 VSS 0.088849f
C7181 B7.t21 VSS 0.087744f
C7182 B7.t0 VSS 0.087744f
C7183 B7.t15 VSS 0.087744f
C7184 B7.n7 VSS 0.349246f
C7185 B7.t25 VSS 0.018234f
C7186 B7.t43 VSS 0.018234f
C7187 B7.t29 VSS 0.018234f
C7188 B7.t3 VSS 0.018234f
C7189 B7.n8 VSS 0.329937f
C7190 B7.n9 VSS 0.516456f
C7191 B7.n10 VSS 19.1576f
C7192 B7.t16 VSS 0.096828f
C7193 B7.t23 VSS 0.041469f
C7194 B7.t42 VSS 0.033153f
C7195 B7.n11 VSS 0.048928f
C7196 B7.t13 VSS 0.03238f
C7197 B7.n12 VSS 0.080772f
C7198 B7.n13 VSS 0.144104f
C7199 B7.n14 VSS 0.226206f
C7200 B7.n15 VSS 2.26575f
C7201 B7.t36 VSS 0.039562f
C7202 B7.t31 VSS 0.042436f
C7203 B7.n16 VSS 0.063233f
C7204 B7.t38 VSS 0.039562f
C7205 B7.t11 VSS 0.039562f
C7206 B7.t12 VSS 0.039562f
C7207 B7.t27 VSS 0.049981f
C7208 B7.n17 VSS 0.106788f
C7209 B7.n18 VSS 0.067234f
C7210 B7.n19 VSS 0.054938f
C7211 B7.n20 VSS 0.026883f
C7212 B7.n21 VSS 0.172162f
C7213 B7.n22 VSS 6.06138f
C7214 B7.t17 VSS 0.044159f
C7215 B7.t44 VSS 0.088849f
C7216 B7.t9 VSS 0.087744f
C7217 B7.t41 VSS 0.087744f
C7218 B7.t22 VSS 0.087744f
C7219 B7.t39 VSS 0.018234f
C7220 B7.t10 VSS 0.018234f
C7221 B7.t45 VSS 0.018234f
C7222 B7.n23 VSS 0.540447f
C7223 B7.n24 VSS 0.3983f
C7224 B7.n25 VSS 0.216996f
C7225 B7.n26 VSS 0.21318f
C7226 B7.n27 VSS 0.13113f
C7227 B7.n28 VSS 0.168739f
C7228 B7.n29 VSS 0.696577f
C7229 B7.n30 VSS 9.0305f
C7230 B7.t7 VSS 0.033153f
C7231 B7.t33 VSS 0.046278f
C7232 B7.t32 VSS 0.046278f
C7233 B7.n31 VSS 0.150647f
C7234 B7.t24 VSS 0.053107f
C7235 B7.n32 VSS 0.449659f
C7236 B7.n33 VSS 0.240952f
C7237 B7.n34 VSS 6.33584f
C7238 B7.t34 VSS 0.033153f
C7239 B7.t8 VSS 0.046278f
C7240 B7.t28 VSS 0.046278f
C7241 B7.n35 VSS 0.150647f
C7242 B7.t20 VSS 0.053107f
C7243 B7.n36 VSS 0.395441f
C7244 B7.n37 VSS 2.62905f
C7245 B7.t2 VSS 0.033153f
C7246 B7.t5 VSS 0.046278f
C7247 B7.t4 VSS 0.046278f
C7248 B7.n38 VSS 0.150647f
C7249 B7.t37 VSS 0.053107f
C7250 B7.n39 VSS 0.394907f
C7251 B7.n40 VSS 0.533757f
C7252 mux8_5.NAND4F_2.Y.n0 VSS 0.530078f
C7253 mux8_5.NAND4F_2.Y.t0 VSS 0.026135f
C7254 mux8_5.NAND4F_2.Y.t1 VSS 0.026135f
C7255 mux8_5.NAND4F_2.Y.n1 VSS 0.060687f
C7256 mux8_5.NAND4F_2.Y.t6 VSS 0.026135f
C7257 mux8_5.NAND4F_2.Y.t5 VSS 0.026135f
C7258 mux8_5.NAND4F_2.Y.n2 VSS 0.060505f
C7259 mux8_5.NAND4F_2.Y.t7 VSS 0.026135f
C7260 mux8_5.NAND4F_2.Y.t8 VSS 0.026135f
C7261 mux8_5.NAND4F_2.Y.n3 VSS 0.060505f
C7262 mux8_5.NAND4F_2.Y.t2 VSS 0.026135f
C7263 mux8_5.NAND4F_2.Y.t3 VSS 0.026135f
C7264 mux8_5.NAND4F_2.Y.n4 VSS 0.060505f
C7265 mux8_5.NAND4F_2.Y.n5 VSS 0.263447f
C7266 mux8_5.NAND4F_2.Y.t4 VSS 0.213114f
C7267 mux8_5.NAND4F_2.Y.t10 VSS 0.034088f
C7268 mux8_5.NAND4F_2.Y.t11 VSS 0.105185f
C7269 mux8_5.NAND4F_2.Y.t9 VSS 0.039267f
C7270 mux8_5.NAND4F_2.Y.n6 VSS 0.131989f
C7271 mux8_5.NAND4F_2.Y.n7 VSS 0.028742f
C7272 mux8_5.NAND4F_2.Y.n8 VSS 1.53344f
C7273 mux8_4.NAND4F_0.C.n0 VSS 1.68955f
C7274 mux8_4.NAND4F_0.C.t13 VSS 0.23388f
C7275 mux8_4.NAND4F_0.C.t10 VSS 0.074606f
C7276 mux8_4.NAND4F_0.C.t9 VSS 0.074606f
C7277 mux8_4.NAND4F_0.C.n1 VSS 0.087589f
C7278 mux8_4.NAND4F_0.C.n2 VSS 0.491098f
C7279 mux8_4.NAND4F_0.C.t14 VSS 0.074606f
C7280 mux8_4.NAND4F_0.C.t15 VSS 0.074606f
C7281 mux8_4.NAND4F_0.C.n3 VSS 0.087589f
C7282 mux8_4.NAND4F_0.C.t12 VSS 0.23388f
C7283 mux8_4.NAND4F_0.C.n4 VSS 0.491129f
C7284 mux8_4.NAND4F_0.C.t5 VSS 0.074606f
C7285 mux8_4.NAND4F_0.C.t7 VSS 0.074606f
C7286 mux8_4.NAND4F_0.C.n5 VSS 0.087589f
C7287 mux8_4.NAND4F_0.C.t4 VSS 0.23388f
C7288 mux8_4.NAND4F_0.C.n6 VSS 0.491143f
C7289 mux8_4.NAND4F_0.C.n7 VSS 1.79123f
C7290 mux8_4.NAND4F_0.C.t3 VSS 0.038013f
C7291 mux8_4.NAND4F_0.C.t2 VSS 0.038013f
C7292 mux8_4.NAND4F_0.C.n8 VSS 0.08471f
C7293 mux8_4.NAND4F_0.C.t1 VSS 0.137874f
C7294 mux8_4.NAND4F_0.C.t0 VSS 0.109643f
C7295 mux8_4.NAND4F_0.C.n9 VSS 3.13611f
C7296 mux8_4.NAND4F_0.C.t11 VSS 0.23388f
C7297 mux8_4.NAND4F_0.C.t8 VSS 0.074606f
C7298 mux8_4.NAND4F_0.C.t6 VSS 0.074606f
C7299 mux8_4.NAND4F_0.C.n10 VSS 0.087589f
C7300 mux8_4.NAND4F_0.C.n11 VSS 0.491115f
C7301 mux8_4.NAND4F_0.C.n12 VSS 2.51327f
C7302 a_n6611_2026.n0 VSS 1.48365f
C7303 a_n6611_2026.n1 VSS 1.48326f
C7304 a_n6611_2026.t4 VSS 0.093341f
C7305 a_n6611_2026.t1 VSS 0.093341f
C7306 a_n6611_2026.t0 VSS 0.093341f
C7307 a_n6611_2026.n2 VSS 0.202296f
C7308 a_n6611_2026.t2 VSS 0.093341f
C7309 a_n6611_2026.t9 VSS 0.093341f
C7310 a_n6611_2026.n3 VSS 0.202001f
C7311 a_n6611_2026.t8 VSS 0.093341f
C7312 a_n6611_2026.t10 VSS 0.093341f
C7313 a_n6611_2026.n4 VSS 0.202001f
C7314 a_n6611_2026.t7 VSS 0.093341f
C7315 a_n6611_2026.t11 VSS 0.093341f
C7316 a_n6611_2026.n5 VSS 0.202001f
C7317 a_n6611_2026.t6 VSS 0.093341f
C7318 a_n6611_2026.t3 VSS 0.093341f
C7319 a_n6611_2026.n6 VSS 0.202001f
C7320 a_n6611_2026.n7 VSS 0.20269f
C7321 a_n6611_2026.t5 VSS 0.093341f
C7322 mux8_0.NAND4F_5.Y.n0 VSS 0.25108f
C7323 mux8_0.NAND4F_5.Y.t10 VSS 0.017162f
C7324 mux8_0.NAND4F_5.Y.t9 VSS 0.050565f
C7325 mux8_0.NAND4F_5.Y.t11 VSS 0.016698f
C7326 mux8_0.NAND4F_5.Y.n1 VSS 0.086077f
C7327 mux8_0.NAND4F_5.Y.t6 VSS 0.099394f
C7328 mux8_0.NAND4F_5.Y.n2 VSS 0.798124f
C7329 mux8_0.NAND4F_5.Y.t0 VSS 0.012379f
C7330 mux8_0.NAND4F_5.Y.t1 VSS 0.012379f
C7331 mux8_0.NAND4F_5.Y.n3 VSS 0.028745f
C7332 mux8_0.NAND4F_5.Y.t8 VSS 0.012379f
C7333 mux8_0.NAND4F_5.Y.t7 VSS 0.012379f
C7334 mux8_0.NAND4F_5.Y.n4 VSS 0.028659f
C7335 mux8_0.NAND4F_5.Y.t2 VSS 0.012379f
C7336 mux8_0.NAND4F_5.Y.t3 VSS 0.012379f
C7337 mux8_0.NAND4F_5.Y.n5 VSS 0.028659f
C7338 mux8_0.NAND4F_5.Y.t4 VSS 0.012379f
C7339 mux8_0.NAND4F_5.Y.t5 VSS 0.012379f
C7340 mux8_0.NAND4F_5.Y.n6 VSS 0.028659f
C7341 mux8_0.NAND4F_5.Y.n7 VSS 0.117805f
C7342 mux8_0.NAND4F_4.B.n0 VSS 0.921489f
C7343 mux8_0.NAND4F_4.B.t4 VSS 0.03989f
C7344 mux8_0.NAND4F_4.B.t13 VSS 0.123086f
C7345 mux8_0.NAND4F_4.B.t15 VSS 0.04595f
C7346 mux8_0.NAND4F_4.B.n1 VSS 0.154452f
C7347 mux8_0.NAND4F_4.B.n2 VSS 0.033769f
C7348 mux8_0.NAND4F_4.B.t14 VSS 0.03989f
C7349 mux8_0.NAND4F_4.B.t7 VSS 0.123086f
C7350 mux8_0.NAND4F_4.B.t12 VSS 0.04595f
C7351 mux8_0.NAND4F_4.B.n3 VSS 0.154452f
C7352 mux8_0.NAND4F_4.B.n4 VSS 0.032977f
C7353 mux8_0.NAND4F_4.B.t10 VSS 0.03989f
C7354 mux8_0.NAND4F_4.B.t5 VSS 0.123086f
C7355 mux8_0.NAND4F_4.B.t9 VSS 0.04595f
C7356 mux8_0.NAND4F_4.B.n5 VSS 0.154452f
C7357 mux8_0.NAND4F_4.B.n6 VSS 0.033699f
C7358 mux8_0.NAND4F_4.B.n7 VSS 0.612655f
C7359 mux8_0.NAND4F_4.B.t3 VSS 0.020325f
C7360 mux8_0.NAND4F_4.B.t1 VSS 0.020325f
C7361 mux8_0.NAND4F_4.B.n8 VSS 0.045293f
C7362 mux8_0.NAND4F_4.B.t2 VSS 0.073718f
C7363 mux8_0.NAND4F_4.B.t0 VSS 0.058624f
C7364 mux8_0.NAND4F_4.B.n9 VSS 0.607515f
C7365 mux8_0.NAND4F_4.B.t8 VSS 0.03989f
C7366 mux8_0.NAND4F_4.B.t11 VSS 0.123086f
C7367 mux8_0.NAND4F_4.B.t6 VSS 0.04595f
C7368 mux8_0.NAND4F_4.B.n10 VSS 0.154452f
C7369 mux8_0.NAND4F_4.B.n11 VSS 0.033659f
C7370 mux8_0.NAND4F_4.B.n12 VSS 0.776456f
C7371 MULT_0.4bit_ADDER_1.B0.t19 VSS 0.042561f
C7372 MULT_0.4bit_ADDER_1.B0.t13 VSS 0.01386f
C7373 MULT_0.4bit_ADDER_1.B0.t12 VSS 0.01914f
C7374 MULT_0.4bit_ADDER_1.B0.n0 VSS 0.02064f
C7375 MULT_0.4bit_ADDER_1.B0.t15 VSS 0.014249f
C7376 MULT_0.4bit_ADDER_1.B0.n1 VSS 0.036155f
C7377 MULT_0.4bit_ADDER_1.B0.n2 VSS 0.063422f
C7378 MULT_0.4bit_ADDER_1.B0.t18 VSS 0.019433f
C7379 MULT_0.4bit_ADDER_1.B0.t22 VSS 0.039099f
C7380 MULT_0.4bit_ADDER_1.B0.t16 VSS 0.038613f
C7381 MULT_0.4bit_ADDER_1.B0.t14 VSS 0.038613f
C7382 MULT_0.4bit_ADDER_1.B0.t21 VSS 0.038613f
C7383 MULT_0.4bit_ADDER_1.B0.t20 VSS 0.008024f
C7384 MULT_0.4bit_ADDER_1.B0.t23 VSS 0.008024f
C7385 MULT_0.4bit_ADDER_1.B0.t17 VSS 0.008024f
C7386 MULT_0.4bit_ADDER_1.B0.n3 VSS 0.237888f
C7387 MULT_0.4bit_ADDER_1.B0.n4 VSS 0.175215f
C7388 MULT_0.4bit_ADDER_1.B0.n5 VSS 0.095491f
C7389 MULT_0.4bit_ADDER_1.B0.n6 VSS 0.093811f
C7390 MULT_0.4bit_ADDER_1.B0.n7 VSS 0.057705f
C7391 MULT_0.4bit_ADDER_1.B0.n8 VSS 0.075698f
C7392 MULT_0.4bit_ADDER_1.B0.n9 VSS 0.836755f
C7393 MULT_0.4bit_ADDER_1.B0.t11 VSS 0.006954f
C7394 MULT_0.4bit_ADDER_1.B0.t10 VSS 0.006954f
C7395 MULT_0.4bit_ADDER_1.B0.n10 VSS 0.016819f
C7396 MULT_0.4bit_ADDER_1.B0.t1 VSS 0.006954f
C7397 MULT_0.4bit_ADDER_1.B0.t8 VSS 0.006954f
C7398 MULT_0.4bit_ADDER_1.B0.n11 VSS 0.016818f
C7399 MULT_0.4bit_ADDER_1.B0.n12 VSS 0.120597f
C7400 MULT_0.4bit_ADDER_1.B0.t9 VSS 0.006954f
C7401 MULT_0.4bit_ADDER_1.B0.t2 VSS 0.006954f
C7402 MULT_0.4bit_ADDER_1.B0.n13 VSS 0.013908f
C7403 MULT_0.4bit_ADDER_1.B0.n14 VSS 0.010925f
C7404 MULT_0.4bit_ADDER_1.B0.t5 VSS 0.029422f
C7405 MULT_0.4bit_ADDER_1.B0.t7 VSS 0.029422f
C7406 MULT_0.4bit_ADDER_1.B0.n15 VSS 0.058843f
C7407 MULT_0.4bit_ADDER_1.B0.n16 VSS 0.023397f
C7408 MULT_0.4bit_ADDER_1.B0.t4 VSS 0.029422f
C7409 MULT_0.4bit_ADDER_1.B0.t3 VSS 0.029422f
C7410 MULT_0.4bit_ADDER_1.B0.n17 VSS 0.058843f
C7411 MULT_0.4bit_ADDER_1.B0.n18 VSS 0.02588f
C7412 MULT_0.4bit_ADDER_1.B0.n19 VSS 0.26645f
C7413 MULT_0.4bit_ADDER_1.B0.t6 VSS 0.029422f
C7414 MULT_0.4bit_ADDER_1.B0.t0 VSS 0.029422f
C7415 MULT_0.4bit_ADDER_1.B0.n20 VSS 0.058843f
C7416 MULT_0.4bit_ADDER_1.B0.n21 VSS 0.025919f
C7417 MULT_0.4bit_ADDER_1.B0.n22 VSS 0.17089f
C7418 MULT_0.4bit_ADDER_1.B0.n23 VSS 0.038512f
C7419 MULT_0.4bit_ADDER_1.B0.n24 VSS 0.169037f
C7420 A4.t13 VSS 0.030079f
C7421 A4.t11 VSS 0.030079f
C7422 A4.t19 VSS 0.030079f
C7423 A4.t8 VSS 0.030079f
C7424 A4.n0 VSS 0.54618f
C7425 A4.t4 VSS 0.144745f
C7426 A4.t21 VSS 0.144745f
C7427 A4.t25 VSS 0.146568f
C7428 A4.t23 VSS 0.144745f
C7429 A4.n1 VSS 0.574218f
C7430 A4.n2 VSS 0.851995f
C7431 A4.t0 VSS 0.135354f
C7432 A4.t3 VSS 0.051955f
C7433 A4.t1 VSS 0.071749f
C7434 A4.n3 VSS 0.082582f
C7435 A4.t2 VSS 0.054612f
C7436 A4.n4 VSS 0.08375f
C7437 A4.n5 VSS 0.34666f
C7438 A4.t14 VSS 0.146568f
C7439 A4.t20 VSS 0.144745f
C7440 A4.t6 VSS 0.144745f
C7441 A4.t26 VSS 0.144745f
C7442 A4.n6 VSS 0.576126f
C7443 A4.t22 VSS 0.030079f
C7444 A4.t16 VSS 0.030079f
C7445 A4.t28 VSS 0.030079f
C7446 A4.t9 VSS 0.030079f
C7447 A4.n7 VSS 0.544272f
C7448 A4.n8 VSS 0.851351f
C7449 A4.n9 VSS 1.69243f
C7450 A4.n10 VSS 2.16974f
C7451 A4.t7 VSS 0.13535f
C7452 A4.t5 VSS 0.068408f
C7453 A4.t15 VSS 0.05469f
C7454 A4.n11 VSS 0.086848f
C7455 A4.t24 VSS 0.054612f
C7456 A4.n12 VSS 0.080093f
C7457 A4.n13 VSS 0.347696f
C7458 A4.n14 VSS 0.636684f
C7459 A4.n15 VSS 4.47315f
C7460 A4.t10 VSS 0.054151f
C7461 A4.t12 VSS 0.065263f
C7462 A4.t29 VSS 0.065263f
C7463 A4.t27 VSS 0.065263f
C7464 A4.t18 VSS 0.065263f
C7465 A4.t17 VSS 0.08245f
C7466 A4.n16 VSS 0.17616f
C7467 A4.n17 VSS 0.110911f
C7468 A4.n18 VSS 0.110911f
C7469 A4.n19 VSS 0.09559f
C7470 A4.n20 VSS 0.078126f
C7471 A4.n21 VSS 0.41925f
C7472 A4.n22 VSS 10.801f
C7473 mux8_1.NAND4F_4.Y.n0 VSS 0.491744f
C7474 mux8_1.NAND4F_4.Y.t3 VSS 0.024245f
C7475 mux8_1.NAND4F_4.Y.t4 VSS 0.024245f
C7476 mux8_1.NAND4F_4.Y.n1 VSS 0.056298f
C7477 mux8_1.NAND4F_4.Y.t5 VSS 0.024245f
C7478 mux8_1.NAND4F_4.Y.t6 VSS 0.024245f
C7479 mux8_1.NAND4F_4.Y.n2 VSS 0.056129f
C7480 mux8_1.NAND4F_4.Y.t7 VSS 0.024245f
C7481 mux8_1.NAND4F_4.Y.t8 VSS 0.024245f
C7482 mux8_1.NAND4F_4.Y.n3 VSS 0.056129f
C7483 mux8_1.NAND4F_4.Y.t1 VSS 0.024245f
C7484 mux8_1.NAND4F_4.Y.t2 VSS 0.024245f
C7485 mux8_1.NAND4F_4.Y.n4 VSS 0.056129f
C7486 mux8_1.NAND4F_4.Y.n5 VSS 0.244395f
C7487 mux8_1.NAND4F_4.Y.t11 VSS 0.033612f
C7488 mux8_1.NAND4F_4.Y.t10 VSS 0.032702f
C7489 mux8_1.NAND4F_4.Y.t9 VSS 0.099032f
C7490 mux8_1.NAND4F_4.Y.n6 VSS 0.168587f
C7491 mux8_1.NAND4F_4.Y.t0 VSS 0.194665f
C7492 mux8_1.NAND4F_4.Y.n7 VSS 1.55341f
C7493 AND8_0.S3.n0 VSS 1.53099f
C7494 AND8_0.S3.t4 VSS 0.074075f
C7495 AND8_0.S3.t5 VSS 0.07207f
C7496 AND8_0.S3.t6 VSS 0.218246f
C7497 AND8_0.S3.n1 VSS 0.37154f
C7498 AND8_0.S3.t1 VSS 0.035509f
C7499 AND8_0.S3.t2 VSS 0.035509f
C7500 AND8_0.S3.n2 VSS 0.07913f
C7501 AND8_0.S3.t3 VSS 0.128792f
C7502 AND8_0.S3.t0 VSS 0.102421f
C7503 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t16 VSS 0.013766f
C7504 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t20 VSS 0.027698f
C7505 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t12 VSS 0.027354f
C7506 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t23 VSS 0.027354f
C7507 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t22 VSS 0.027354f
C7508 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t19 VSS 0.005684f
C7509 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t15 VSS 0.005684f
C7510 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t17 VSS 0.005684f
C7511 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n0 VSS 0.168523f
C7512 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n1 VSS 0.124125f
C7513 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n2 VSS 0.067647f
C7514 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n3 VSS 0.066457f
C7515 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n4 VSS 0.040879f
C7516 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n5 VSS 0.05311f
C7517 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t18 VSS 0.030151f
C7518 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t14 VSS 0.009818f
C7519 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t13 VSS 0.013559f
C7520 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n6 VSS 0.014622f
C7521 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t21 VSS 0.010094f
C7522 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n7 VSS 0.025612f
C7523 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n8 VSS 0.044927f
C7524 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t11 VSS 0.004926f
C7525 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t10 VSS 0.004926f
C7526 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n9 VSS 0.011915f
C7527 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t1 VSS 0.004926f
C7528 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t0 VSS 0.004926f
C7529 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n10 VSS 0.011914f
C7530 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n11 VSS 0.085433f
C7531 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t9 VSS 0.004926f
C7532 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t2 VSS 0.004926f
C7533 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n12 VSS 0.009853f
C7534 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n13 VSS 0.00774f
C7535 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t6 VSS 0.020843f
C7536 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t5 VSS 0.020843f
C7537 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n14 VSS 0.041685f
C7538 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n15 VSS 0.016575f
C7539 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t8 VSS 0.020843f
C7540 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t7 VSS 0.020843f
C7541 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n16 VSS 0.041685f
C7542 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n17 VSS 0.018334f
C7543 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n18 VSS 0.188757f
C7544 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t4 VSS 0.020843f
C7545 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.t3 VSS 0.020843f
C7546 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n19 VSS 0.041685f
C7547 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n20 VSS 0.018362f
C7548 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n21 VSS 0.12106f
C7549 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n22 VSS 0.027282f
C7550 MULT_0.4bit_ADDER_0.FULL_ADDER_0.XOR2_1.A.n23 VSS 0.119748f
C7551 a_n9901_2026.n0 VSS 1.48326f
C7552 a_n9901_2026.n1 VSS 1.48365f
C7553 a_n9901_2026.t5 VSS 0.093341f
C7554 a_n9901_2026.t3 VSS 0.093341f
C7555 a_n9901_2026.t4 VSS 0.093341f
C7556 a_n9901_2026.n2 VSS 0.202296f
C7557 a_n9901_2026.t7 VSS 0.093341f
C7558 a_n9901_2026.t8 VSS 0.093341f
C7559 a_n9901_2026.n3 VSS 0.20269f
C7560 a_n9901_2026.t10 VSS 0.093341f
C7561 a_n9901_2026.t6 VSS 0.093341f
C7562 a_n9901_2026.n4 VSS 0.202001f
C7563 a_n9901_2026.t11 VSS 0.093341f
C7564 a_n9901_2026.t9 VSS 0.093341f
C7565 a_n9901_2026.n5 VSS 0.202001f
C7566 a_n9901_2026.t0 VSS 0.093341f
C7567 a_n9901_2026.t1 VSS 0.093341f
C7568 a_n9901_2026.n6 VSS 0.202001f
C7569 a_n9901_2026.n7 VSS 0.202001f
C7570 a_n9901_2026.t2 VSS 0.093341f
C7571 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t3 VSS 0.007073f
C7572 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t4 VSS 0.007073f
C7573 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n0 VSS 0.017105f
C7574 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t10 VSS 0.007073f
C7575 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t11 VSS 0.007073f
C7576 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n1 VSS 0.017107f
C7577 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n2 VSS 0.122656f
C7578 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t5 VSS 0.007073f
C7579 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t9 VSS 0.007073f
C7580 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n3 VSS 0.014146f
C7581 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n4 VSS 0.011112f
C7582 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t8 VSS 0.029924f
C7583 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t2 VSS 0.029924f
C7584 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n5 VSS 0.059848f
C7585 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n6 VSS 0.023796f
C7586 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t6 VSS 0.029924f
C7587 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t7 VSS 0.029924f
C7588 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n7 VSS 0.059848f
C7589 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n8 VSS 0.026362f
C7590 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n9 VSS 0.271f
C7591 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t1 VSS 0.029924f
C7592 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t0 VSS 0.029924f
C7593 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n10 VSS 0.059848f
C7594 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n11 VSS 0.026322f
C7595 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n12 VSS 0.173808f
C7596 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n13 VSS 0.03917f
C7597 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n14 VSS 0.172104f
C7598 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t15 VSS 0.043288f
C7599 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t18 VSS 0.014096f
C7600 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t19 VSS 0.019467f
C7601 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n15 VSS 0.020992f
C7602 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t13 VSS 0.014492f
C7603 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n16 VSS 0.036772f
C7604 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n17 VSS 0.064505f
C7605 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t23 VSS 0.019764f
C7606 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t14 VSS 0.039767f
C7607 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t21 VSS 0.039272f
C7608 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t12 VSS 0.039272f
C7609 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t16 VSS 0.039272f
C7610 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t17 VSS 0.008161f
C7611 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t22 VSS 0.008161f
C7612 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.t20 VSS 0.008161f
C7613 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n18 VSS 0.24195f
C7614 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n19 VSS 0.178207f
C7615 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n20 VSS 0.097121f
C7616 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n21 VSS 0.095413f
C7617 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n22 VSS 0.05869f
C7618 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n23 VSS 0.076991f
C7619 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_2.Y.n24 VSS 1.26966f
C7620 mux8_2.NAND4F_2.Y.n0 VSS 0.530078f
C7621 mux8_2.NAND4F_2.Y.t5 VSS 0.026135f
C7622 mux8_2.NAND4F_2.Y.t4 VSS 0.026135f
C7623 mux8_2.NAND4F_2.Y.n1 VSS 0.060687f
C7624 mux8_2.NAND4F_2.Y.t1 VSS 0.026135f
C7625 mux8_2.NAND4F_2.Y.t0 VSS 0.026135f
C7626 mux8_2.NAND4F_2.Y.n2 VSS 0.060505f
C7627 mux8_2.NAND4F_2.Y.t2 VSS 0.026135f
C7628 mux8_2.NAND4F_2.Y.t3 VSS 0.026135f
C7629 mux8_2.NAND4F_2.Y.n3 VSS 0.060505f
C7630 mux8_2.NAND4F_2.Y.t7 VSS 0.026135f
C7631 mux8_2.NAND4F_2.Y.t8 VSS 0.026135f
C7632 mux8_2.NAND4F_2.Y.n4 VSS 0.060505f
C7633 mux8_2.NAND4F_2.Y.n5 VSS 0.263447f
C7634 mux8_2.NAND4F_2.Y.t6 VSS 0.213114f
C7635 mux8_2.NAND4F_2.Y.t10 VSS 0.034088f
C7636 mux8_2.NAND4F_2.Y.t9 VSS 0.105185f
C7637 mux8_2.NAND4F_2.Y.t11 VSS 0.039267f
C7638 mux8_2.NAND4F_2.Y.n6 VSS 0.131989f
C7639 mux8_2.NAND4F_2.Y.n7 VSS 0.028742f
C7640 mux8_2.NAND4F_2.Y.n8 VSS 1.53344f
C7641 OR8_0.S1.n0 VSS 3.45178f
C7642 OR8_0.S1.t6 VSS 0.167204f
C7643 OR8_0.S1.t5 VSS 0.162679f
C7644 OR8_0.S1.t4 VSS 0.492633f
C7645 OR8_0.S1.n1 VSS 0.838723f
C7646 OR8_0.S1.t1 VSS 0.080153f
C7647 OR8_0.S1.t0 VSS 0.080153f
C7648 OR8_0.S1.n2 VSS 0.178616f
C7649 OR8_0.S1.t2 VSS 0.290714f
C7650 OR8_0.S1.t3 VSS 0.231188f
C7651 mux8_1.NAND4F_3.Y.n0 VSS 0.320257f
C7652 mux8_1.NAND4F_3.Y.t5 VSS 0.01579f
C7653 mux8_1.NAND4F_3.Y.t6 VSS 0.01579f
C7654 mux8_1.NAND4F_3.Y.n1 VSS 0.036665f
C7655 mux8_1.NAND4F_3.Y.t1 VSS 0.01579f
C7656 mux8_1.NAND4F_3.Y.t0 VSS 0.01579f
C7657 mux8_1.NAND4F_3.Y.n2 VSS 0.036555f
C7658 mux8_1.NAND4F_3.Y.t8 VSS 0.01579f
C7659 mux8_1.NAND4F_3.Y.t7 VSS 0.01579f
C7660 mux8_1.NAND4F_3.Y.n3 VSS 0.036555f
C7661 mux8_1.NAND4F_3.Y.t3 VSS 0.01579f
C7662 mux8_1.NAND4F_3.Y.t4 VSS 0.01579f
C7663 mux8_1.NAND4F_3.Y.n4 VSS 0.036555f
C7664 mux8_1.NAND4F_3.Y.n5 VSS 0.159167f
C7665 mux8_1.NAND4F_3.Y.t2 VSS 0.150045f
C7666 mux8_1.NAND4F_3.Y.t10 VSS 0.020595f
C7667 mux8_1.NAND4F_3.Y.t9 VSS 0.020595f
C7668 mux8_1.NAND4F_3.Y.n6 VSS 0.024179f
C7669 mux8_1.NAND4F_3.Y.t11 VSS 0.064563f
C7670 mux8_1.NAND4F_3.Y.n7 VSS 0.135573f
C7671 a_n20557_n7799.n0 VSS 1.48326f
C7672 a_n20557_n7799.n1 VSS 1.48365f
C7673 a_n20557_n7799.t0 VSS 0.093341f
C7674 a_n20557_n7799.t6 VSS 0.093341f
C7675 a_n20557_n7799.t8 VSS 0.093341f
C7676 a_n20557_n7799.n2 VSS 0.202296f
C7677 a_n20557_n7799.t7 VSS 0.093341f
C7678 a_n20557_n7799.t1 VSS 0.093341f
C7679 a_n20557_n7799.n3 VSS 0.202001f
C7680 a_n20557_n7799.t3 VSS 0.093341f
C7681 a_n20557_n7799.t5 VSS 0.093341f
C7682 a_n20557_n7799.n4 VSS 0.20269f
C7683 a_n20557_n7799.t11 VSS 0.093341f
C7684 a_n20557_n7799.t4 VSS 0.093341f
C7685 a_n20557_n7799.n5 VSS 0.202001f
C7686 a_n20557_n7799.t9 VSS 0.093341f
C7687 a_n20557_n7799.t10 VSS 0.093341f
C7688 a_n20557_n7799.n6 VSS 0.202001f
C7689 a_n20557_n7799.n7 VSS 0.202001f
C7690 a_n20557_n7799.t2 VSS 0.093341f
C7691 mux8_0.NAND4F_6.Y.n0 VSS 0.599344f
C7692 mux8_0.NAND4F_6.Y.t6 VSS 0.244548f
C7693 mux8_0.NAND4F_6.Y.t11 VSS 0.038543f
C7694 mux8_0.NAND4F_6.Y.t9 VSS 0.118929f
C7695 mux8_0.NAND4F_6.Y.t10 VSS 0.044398f
C7696 mux8_0.NAND4F_6.Y.n1 VSS 0.149236f
C7697 mux8_0.NAND4F_6.Y.n2 VSS 0.032396f
C7698 mux8_0.NAND4F_6.Y.n3 VSS 1.72835f
C7699 mux8_0.NAND4F_6.Y.t1 VSS 0.029549f
C7700 mux8_0.NAND4F_6.Y.t0 VSS 0.029549f
C7701 mux8_0.NAND4F_6.Y.n4 VSS 0.068617f
C7702 mux8_0.NAND4F_6.Y.t3 VSS 0.029549f
C7703 mux8_0.NAND4F_6.Y.t2 VSS 0.029549f
C7704 mux8_0.NAND4F_6.Y.n5 VSS 0.068411f
C7705 mux8_0.NAND4F_6.Y.t8 VSS 0.029549f
C7706 mux8_0.NAND4F_6.Y.t7 VSS 0.029549f
C7707 mux8_0.NAND4F_6.Y.n6 VSS 0.068411f
C7708 mux8_0.NAND4F_6.Y.t4 VSS 0.029549f
C7709 mux8_0.NAND4F_6.Y.t5 VSS 0.029549f
C7710 mux8_0.NAND4F_6.Y.n7 VSS 0.068411f
C7711 mux8_0.NAND4F_6.Y.n8 VSS 0.281208f
C7712 a_n17368_3810.n0 VSS 1.45527f
C7713 a_n17368_3810.n1 VSS 1.45566f
C7714 a_n17368_3810.t1 VSS 0.09158f
C7715 a_n17368_3810.t7 VSS 0.09158f
C7716 a_n17368_3810.t8 VSS 0.09158f
C7717 a_n17368_3810.n2 VSS 0.198865f
C7718 a_n17368_3810.t6 VSS 0.09158f
C7719 a_n17368_3810.t4 VSS 0.09158f
C7720 a_n17368_3810.n3 VSS 0.19819f
C7721 a_n17368_3810.t5 VSS 0.09158f
C7722 a_n17368_3810.t3 VSS 0.09158f
C7723 a_n17368_3810.n4 VSS 0.19819f
C7724 a_n17368_3810.t9 VSS 0.09158f
C7725 a_n17368_3810.t10 VSS 0.09158f
C7726 a_n17368_3810.n5 VSS 0.19819f
C7727 a_n17368_3810.t11 VSS 0.09158f
C7728 a_n17368_3810.t0 VSS 0.09158f
C7729 a_n17368_3810.n6 VSS 0.19819f
C7730 a_n17368_3810.n7 VSS 0.198479f
C7731 a_n17368_3810.t2 VSS 0.09158f
C7732 right_shifter_0.S2.n0 VSS 2.26828f
C7733 mux8_3.NAND4F_6.A VSS 0.36191f
C7734 right_shifter_0.S2.t4 VSS 0.027483f
C7735 right_shifter_0.S2.t6 VSS 0.080973f
C7736 right_shifter_0.S2.t5 VSS 0.026739f
C7737 right_shifter_0.S2.n1 VSS 0.137859f
C7738 right_shifter_0.S2.t3 VSS 0.013175f
C7739 right_shifter_0.S2.t2 VSS 0.013175f
C7740 right_shifter_0.S2.n2 VSS 0.029358f
C7741 right_shifter_0.S2.t1 VSS 0.047784f
C7742 right_shifter_0.S2.t0 VSS 0.038f
C7743 mux8_3.A7 VSS 2.35526f
C7744 a_n10786_3810.n0 VSS 1.45527f
C7745 a_n10786_3810.n1 VSS 1.45566f
C7746 a_n10786_3810.t11 VSS 0.09158f
C7747 a_n10786_3810.t8 VSS 0.09158f
C7748 a_n10786_3810.t9 VSS 0.09158f
C7749 a_n10786_3810.n2 VSS 0.198865f
C7750 a_n10786_3810.t10 VSS 0.09158f
C7751 a_n10786_3810.t4 VSS 0.09158f
C7752 a_n10786_3810.n3 VSS 0.19819f
C7753 a_n10786_3810.t5 VSS 0.09158f
C7754 a_n10786_3810.t3 VSS 0.09158f
C7755 a_n10786_3810.n4 VSS 0.19819f
C7756 a_n10786_3810.t7 VSS 0.09158f
C7757 a_n10786_3810.t6 VSS 0.09158f
C7758 a_n10786_3810.n5 VSS 0.19819f
C7759 a_n10786_3810.t0 VSS 0.09158f
C7760 a_n10786_3810.t1 VSS 0.09158f
C7761 a_n10786_3810.n6 VSS 0.198479f
C7762 a_n10786_3810.n7 VSS 0.19819f
C7763 a_n10786_3810.t2 VSS 0.09158f
C7764 mux8_7.NAND4F_6.Y.n0 VSS 0.599344f
C7765 mux8_7.NAND4F_6.Y.t2 VSS 0.244548f
C7766 mux8_7.NAND4F_6.Y.t11 VSS 0.038543f
C7767 mux8_7.NAND4F_6.Y.t9 VSS 0.118929f
C7768 mux8_7.NAND4F_6.Y.t10 VSS 0.044398f
C7769 mux8_7.NAND4F_6.Y.n1 VSS 0.149236f
C7770 mux8_7.NAND4F_6.Y.n2 VSS 0.032396f
C7771 mux8_7.NAND4F_6.Y.n3 VSS 1.72835f
C7772 mux8_7.NAND4F_6.Y.t1 VSS 0.029549f
C7773 mux8_7.NAND4F_6.Y.t0 VSS 0.029549f
C7774 mux8_7.NAND4F_6.Y.n4 VSS 0.068617f
C7775 mux8_7.NAND4F_6.Y.t6 VSS 0.029549f
C7776 mux8_7.NAND4F_6.Y.t5 VSS 0.029549f
C7777 mux8_7.NAND4F_6.Y.n5 VSS 0.068411f
C7778 mux8_7.NAND4F_6.Y.t7 VSS 0.029549f
C7779 mux8_7.NAND4F_6.Y.t8 VSS 0.029549f
C7780 mux8_7.NAND4F_6.Y.n6 VSS 0.068411f
C7781 mux8_7.NAND4F_6.Y.t4 VSS 0.029549f
C7782 mux8_7.NAND4F_6.Y.t3 VSS 0.029549f
C7783 mux8_7.NAND4F_6.Y.n7 VSS 0.068411f
C7784 mux8_7.NAND4F_6.Y.n8 VSS 0.281208f
C7785 right_shifter_0.S5.n0 VSS 2.71757f
C7786 mux8_7.NAND4F_6.A VSS 0.341619f
C7787 right_shifter_0.S5.t5 VSS 0.025879f
C7788 right_shifter_0.S5.t4 VSS 0.076246f
C7789 right_shifter_0.S5.t6 VSS 0.025178f
C7790 right_shifter_0.S5.n1 VSS 0.129811f
C7791 right_shifter_0.S5.t3 VSS 0.012405f
C7792 right_shifter_0.S5.t2 VSS 0.012405f
C7793 right_shifter_0.S5.n2 VSS 0.027645f
C7794 right_shifter_0.S5.t1 VSS 0.044994f
C7795 right_shifter_0.S5.t0 VSS 0.035781f
C7796 mux8_7.A7 VSS 2.45047f
C7797 AND8_0.S1.n0 VSS 4.55957f
C7798 AND8_0.S1.t2 VSS 0.1059f
C7799 AND8_0.S1.t3 VSS 0.1059f
C7800 AND8_0.S1.n1 VSS 0.235991f
C7801 AND8_0.S1.t1 VSS 0.384099f
C7802 AND8_0.S1.t0 VSS 0.305451f
C7803 AND8_0.S1.t6 VSS 0.220915f
C7804 AND8_0.S1.t5 VSS 0.214935f
C7805 AND8_0.S1.t4 VSS 0.650879f
C7806 AND8_0.S1.n2 VSS 1.10805f
C7807 mux8_4.A0.t12 VSS 0.05837f
C7808 mux8_4.A0.t14 VSS 0.05679f
C7809 mux8_4.A0.t13 VSS 0.171976f
C7810 mux8_4.A0.n0 VSS 0.292794f
C7811 mux8_4.A0.t2 VSS 0.016998f
C7812 mux8_4.A0.t3 VSS 0.016998f
C7813 mux8_4.A0.n1 VSS 0.041111f
C7814 mux8_4.A0.t5 VSS 0.016998f
C7815 mux8_4.A0.t6 VSS 0.016998f
C7816 mux8_4.A0.n2 VSS 0.041107f
C7817 mux8_4.A0.n3 VSS 0.294772f
C7818 mux8_4.A0.t1 VSS 0.016998f
C7819 mux8_4.A0.t4 VSS 0.016998f
C7820 mux8_4.A0.n4 VSS 0.033996f
C7821 mux8_4.A0.n5 VSS 0.026705f
C7822 mux8_4.A0.t11 VSS 0.071914f
C7823 mux8_4.A0.t9 VSS 0.071914f
C7824 mux8_4.A0.n6 VSS 0.143828f
C7825 mux8_4.A0.n7 VSS 0.057188f
C7826 mux8_4.A0.t10 VSS 0.071914f
C7827 mux8_4.A0.t0 VSS 0.071914f
C7828 mux8_4.A0.n8 VSS 0.143828f
C7829 mux8_4.A0.n9 VSS 0.063258f
C7830 mux8_4.A0.n10 VSS 0.651276f
C7831 mux8_4.A0.t7 VSS 0.071914f
C7832 mux8_4.A0.t8 VSS 0.071914f
C7833 mux8_4.A0.n11 VSS 0.143828f
C7834 mux8_4.A0.n12 VSS 0.063354f
C7835 mux8_4.A0.n13 VSS 0.4177f
C7836 mux8_4.A0.n14 VSS 0.094133f
C7837 mux8_4.A0.n15 VSS 0.413171f
C7838 mux8_3.NAND4F_5.Y.n0 VSS 0.25108f
C7839 mux8_3.NAND4F_5.Y.t9 VSS 0.017162f
C7840 mux8_3.NAND4F_5.Y.t11 VSS 0.050565f
C7841 mux8_3.NAND4F_5.Y.t10 VSS 0.016698f
C7842 mux8_3.NAND4F_5.Y.n1 VSS 0.086077f
C7843 mux8_3.NAND4F_5.Y.t8 VSS 0.099394f
C7844 mux8_3.NAND4F_5.Y.n2 VSS 0.798124f
C7845 mux8_3.NAND4F_5.Y.t1 VSS 0.012379f
C7846 mux8_3.NAND4F_5.Y.t0 VSS 0.012379f
C7847 mux8_3.NAND4F_5.Y.n3 VSS 0.028745f
C7848 mux8_3.NAND4F_5.Y.t2 VSS 0.012379f
C7849 mux8_3.NAND4F_5.Y.t3 VSS 0.012379f
C7850 mux8_3.NAND4F_5.Y.n4 VSS 0.028659f
C7851 mux8_3.NAND4F_5.Y.t4 VSS 0.012379f
C7852 mux8_3.NAND4F_5.Y.t5 VSS 0.012379f
C7853 mux8_3.NAND4F_5.Y.n5 VSS 0.028659f
C7854 mux8_3.NAND4F_5.Y.t6 VSS 0.012379f
C7855 mux8_3.NAND4F_5.Y.t7 VSS 0.012379f
C7856 mux8_3.NAND4F_5.Y.n6 VSS 0.028659f
C7857 mux8_3.NAND4F_5.Y.n7 VSS 0.117805f
C7858 mux8_6.NAND4F_1.Y.n0 VSS 0.655599f
C7859 mux8_6.NAND4F_1.Y.t8 VSS 0.306614f
C7860 mux8_6.NAND4F_1.Y.t11 VSS 0.132168f
C7861 mux8_6.NAND4F_1.Y.t10 VSS 0.04216f
C7862 mux8_6.NAND4F_1.Y.t9 VSS 0.04216f
C7863 mux8_6.NAND4F_1.Y.n1 VSS 0.049498f
C7864 mux8_6.NAND4F_1.Y.n2 VSS 0.277534f
C7865 mux8_6.NAND4F_1.Y.t1 VSS 0.032323f
C7866 mux8_6.NAND4F_1.Y.t0 VSS 0.032323f
C7867 mux8_6.NAND4F_1.Y.n3 VSS 0.075057f
C7868 mux8_6.NAND4F_1.Y.t3 VSS 0.032323f
C7869 mux8_6.NAND4F_1.Y.t2 VSS 0.032323f
C7870 mux8_6.NAND4F_1.Y.n4 VSS 0.074832f
C7871 mux8_6.NAND4F_1.Y.t5 VSS 0.032323f
C7872 mux8_6.NAND4F_1.Y.t4 VSS 0.032323f
C7873 mux8_6.NAND4F_1.Y.n5 VSS 0.074832f
C7874 mux8_6.NAND4F_1.Y.t6 VSS 0.032323f
C7875 mux8_6.NAND4F_1.Y.t7 VSS 0.032323f
C7876 mux8_6.NAND4F_1.Y.n6 VSS 0.074832f
C7877 mux8_6.NAND4F_1.Y.n7 VSS 0.307603f
C7878 mux8_6.NAND4F_0.C.n0 VSS 1.44981f
C7879 mux8_6.NAND4F_0.C.t10 VSS 0.200694f
C7880 mux8_6.NAND4F_0.C.t15 VSS 0.06402f
C7881 mux8_6.NAND4F_0.C.t14 VSS 0.06402f
C7882 mux8_6.NAND4F_0.C.n1 VSS 0.075161f
C7883 mux8_6.NAND4F_0.C.n2 VSS 0.421415f
C7884 mux8_6.NAND4F_0.C.t7 VSS 0.06402f
C7885 mux8_6.NAND4F_0.C.t9 VSS 0.06402f
C7886 mux8_6.NAND4F_0.C.n3 VSS 0.075161f
C7887 mux8_6.NAND4F_0.C.t6 VSS 0.200694f
C7888 mux8_6.NAND4F_0.C.n4 VSS 0.421442f
C7889 mux8_6.NAND4F_0.C.t12 VSS 0.06402f
C7890 mux8_6.NAND4F_0.C.t13 VSS 0.06402f
C7891 mux8_6.NAND4F_0.C.n5 VSS 0.075161f
C7892 mux8_6.NAND4F_0.C.t11 VSS 0.200694f
C7893 mux8_6.NAND4F_0.C.n6 VSS 0.421454f
C7894 mux8_6.NAND4F_0.C.n7 VSS 1.53707f
C7895 mux8_6.NAND4F_0.C.t3 VSS 0.03262f
C7896 mux8_6.NAND4F_0.C.t2 VSS 0.03262f
C7897 mux8_6.NAND4F_0.C.n8 VSS 0.072691f
C7898 mux8_6.NAND4F_0.C.t1 VSS 0.118311f
C7899 mux8_6.NAND4F_0.C.t0 VSS 0.094086f
C7900 mux8_6.NAND4F_0.C.n9 VSS 2.69112f
C7901 mux8_6.NAND4F_0.C.t8 VSS 0.200694f
C7902 mux8_6.NAND4F_0.C.t5 VSS 0.06402f
C7903 mux8_6.NAND4F_0.C.t4 VSS 0.06402f
C7904 mux8_6.NAND4F_0.C.n10 VSS 0.075161f
C7905 mux8_6.NAND4F_0.C.n11 VSS 0.42143f
C7906 mux8_6.NAND4F_0.C.n12 VSS 2.15666f
C7907 a_n10684_n4534.n0 VSS 1.48326f
C7908 a_n10684_n4534.n1 VSS 1.48365f
C7909 a_n10684_n4534.t0 VSS 0.093341f
C7910 a_n10684_n4534.t4 VSS 0.093341f
C7911 a_n10684_n4534.t5 VSS 0.093341f
C7912 a_n10684_n4534.n2 VSS 0.202296f
C7913 a_n10684_n4534.t3 VSS 0.093341f
C7914 a_n10684_n4534.t1 VSS 0.093341f
C7915 a_n10684_n4534.n3 VSS 0.202001f
C7916 a_n10684_n4534.t8 VSS 0.093341f
C7917 a_n10684_n4534.t7 VSS 0.093341f
C7918 a_n10684_n4534.n4 VSS 0.20269f
C7919 a_n10684_n4534.t11 VSS 0.093341f
C7920 a_n10684_n4534.t6 VSS 0.093341f
C7921 a_n10684_n4534.n5 VSS 0.202001f
C7922 a_n10684_n4534.t9 VSS 0.093341f
C7923 a_n10684_n4534.t10 VSS 0.093341f
C7924 a_n10684_n4534.n6 VSS 0.202001f
C7925 a_n10684_n4534.n7 VSS 0.202001f
C7926 a_n10684_n4534.t2 VSS 0.093341f
C7927 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t15 VSS 0.013766f
C7928 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t18 VSS 0.027698f
C7929 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t12 VSS 0.027354f
C7930 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t23 VSS 0.027354f
C7931 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t20 VSS 0.027354f
C7932 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t21 VSS 0.005684f
C7933 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t14 VSS 0.005684f
C7934 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t16 VSS 0.005684f
C7935 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n0 VSS 0.168523f
C7936 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n1 VSS 0.124125f
C7937 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n2 VSS 0.067647f
C7938 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n3 VSS 0.066457f
C7939 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n4 VSS 0.040879f
C7940 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n5 VSS 0.05311f
C7941 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t22 VSS 0.030151f
C7942 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t17 VSS 0.009818f
C7943 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t13 VSS 0.013559f
C7944 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n6 VSS 0.014622f
C7945 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t19 VSS 0.010094f
C7946 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n7 VSS 0.025612f
C7947 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n8 VSS 0.044927f
C7948 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t8 VSS 0.004926f
C7949 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t7 VSS 0.004926f
C7950 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n9 VSS 0.011915f
C7951 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t1 VSS 0.004926f
C7952 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t2 VSS 0.004926f
C7953 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n10 VSS 0.011914f
C7954 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n11 VSS 0.085433f
C7955 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t6 VSS 0.004926f
C7956 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t0 VSS 0.004926f
C7957 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n12 VSS 0.009853f
C7958 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n13 VSS 0.00774f
C7959 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t5 VSS 0.020843f
C7960 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t9 VSS 0.020843f
C7961 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n14 VSS 0.041685f
C7962 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n15 VSS 0.016575f
C7963 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t4 VSS 0.020843f
C7964 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t3 VSS 0.020843f
C7965 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n16 VSS 0.041685f
C7966 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n17 VSS 0.018334f
C7967 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n18 VSS 0.188757f
C7968 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t10 VSS 0.020843f
C7969 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.t11 VSS 0.020843f
C7970 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n19 VSS 0.041685f
C7971 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n20 VSS 0.018362f
C7972 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n21 VSS 0.12106f
C7973 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n22 VSS 0.027282f
C7974 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.A.n23 VSS 0.119748f
C7975 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_0.A VSS 0.361534f
C7976 MULT_0.4bit_ADDER_0.B1.n0 VSS 2.7934f
C7977 MULT_0.4bit_ADDER_0.FULL_ADDER_2.B VSS 5.46099f
C7978 MULT_0.4bit_ADDER_0.B1.t0 VSS 0.07522f
C7979 MULT_0.4bit_ADDER_0.B1.t1 VSS 0.094429f
C7980 MULT_0.4bit_ADDER_0.B1.t3 VSS 0.026035f
C7981 MULT_0.4bit_ADDER_0.B1.t2 VSS 0.026035f
C7982 MULT_0.4bit_ADDER_0.B1.n1 VSS 0.058005f
C7983 MULT_0.4bit_ADDER_0.B1.t13 VSS 0.096796f
C7984 MULT_0.4bit_ADDER_0.B1.t8 VSS 0.031521f
C7985 MULT_0.4bit_ADDER_0.B1.t5 VSS 0.043529f
C7986 MULT_0.4bit_ADDER_0.B1.n2 VSS 0.046941f
C7987 MULT_0.4bit_ADDER_0.B1.t9 VSS 0.032406f
C7988 MULT_0.4bit_ADDER_0.B1.n3 VSS 0.082226f
C7989 MULT_0.4bit_ADDER_0.B1.n4 VSS 0.144239f
C7990 MULT_0.4bit_ADDER_0.B1.t10 VSS 0.044195f
C7991 MULT_0.4bit_ADDER_0.B1.t14 VSS 0.088922f
C7992 MULT_0.4bit_ADDER_0.B1.t11 VSS 0.087816f
C7993 MULT_0.4bit_ADDER_0.B1.t12 VSS 0.087816f
C7994 MULT_0.4bit_ADDER_0.B1.t6 VSS 0.087816f
C7995 MULT_0.4bit_ADDER_0.B1.t7 VSS 0.018249f
C7996 MULT_0.4bit_ADDER_0.B1.t15 VSS 0.018249f
C7997 MULT_0.4bit_ADDER_0.B1.t4 VSS 0.018249f
C7998 MULT_0.4bit_ADDER_0.B1.n5 VSS 0.541024f
C7999 MULT_0.4bit_ADDER_0.B1.n6 VSS 0.398489f
C8000 MULT_0.4bit_ADDER_0.B1.n7 VSS 0.217173f
C8001 MULT_0.4bit_ADDER_0.B1.n8 VSS 0.213354f
C8002 MULT_0.4bit_ADDER_0.B1.n9 VSS 0.131237f
C8003 MULT_0.4bit_ADDER_0.B1.n10 VSS 0.17216f
C8004 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_0.A VSS 0.306162f
C8005 MULT_0.4bit_ADDER_0.B1.n11 VSS 1.89578f
C8006 MULT_0.NAND2_1.Y.n0 VSS 1.24053f
C8007 MULT_0.NAND2_1.Y.n1 VSS 0.197241f
C8008 MULT_0.NAND2_1.Y.t5 VSS 0.024293f
C8009 MULT_0.NAND2_1.Y.t4 VSS 0.024293f
C8010 MULT_0.NAND2_1.Y.n2 VSS 0.054203f
C8011 MULT_0.NAND2_1.Y.t2 VSS 0.024293f
C8012 MULT_0.NAND2_1.Y.t6 VSS 0.024293f
C8013 MULT_0.NAND2_1.Y.n3 VSS 0.054056f
C8014 MULT_0.NAND2_1.Y.t1 VSS 0.024293f
C8015 MULT_0.NAND2_1.Y.t3 VSS 0.024293f
C8016 MULT_0.NAND2_1.Y.n4 VSS 0.054056f
C8017 MULT_0.NAND2_1.Y.t0 VSS 0.146348f
C8018 MULT_0.NAND2_1.Y.t8 VSS 0.03096f
C8019 MULT_0.NAND2_1.Y.t7 VSS 0.043218f
C8020 MULT_0.NAND2_1.Y.t9 VSS 0.043218f
C8021 MULT_0.NAND2_1.Y.n5 VSS 0.141069f
C8022 MULT_0.NAND2_1.Y.t10 VSS 0.049344f
C8023 a_n8170_2026.n0 VSS 1.48365f
C8024 a_n8170_2026.n1 VSS 1.48326f
C8025 a_n8170_2026.t1 VSS 0.093341f
C8026 a_n8170_2026.t4 VSS 0.093341f
C8027 a_n8170_2026.t5 VSS 0.093341f
C8028 a_n8170_2026.n2 VSS 0.202296f
C8029 a_n8170_2026.t3 VSS 0.093341f
C8030 a_n8170_2026.t10 VSS 0.093341f
C8031 a_n8170_2026.n3 VSS 0.202001f
C8032 a_n8170_2026.t11 VSS 0.093341f
C8033 a_n8170_2026.t9 VSS 0.093341f
C8034 a_n8170_2026.n4 VSS 0.202001f
C8035 a_n8170_2026.t6 VSS 0.093341f
C8036 a_n8170_2026.t7 VSS 0.093341f
C8037 a_n8170_2026.n5 VSS 0.202001f
C8038 a_n8170_2026.t8 VSS 0.093341f
C8039 a_n8170_2026.t0 VSS 0.093341f
C8040 a_n8170_2026.n6 VSS 0.202001f
C8041 a_n8170_2026.n7 VSS 0.20269f
C8042 a_n8170_2026.t2 VSS 0.093341f
C8043 mux8_1.NAND4F_2.D.n0 VSS 0.664607f
C8044 mux8_1.NAND4F_2.D.t11 VSS 0.027742f
C8045 mux8_1.NAND4F_2.D.t10 VSS 0.098211f
C8046 mux8_1.NAND4F_2.D.t13 VSS 0.030538f
C8047 mux8_1.NAND4F_2.D.n1 VSS 0.087112f
C8048 mux8_1.NAND4F_2.D.n2 VSS 0.025808f
C8049 mux8_1.NAND4F_2.D.t3 VSS 0.014135f
C8050 mux8_1.NAND4F_2.D.t2 VSS 0.014135f
C8051 mux8_1.NAND4F_2.D.n3 VSS 0.031499f
C8052 mux8_1.NAND4F_2.D.t1 VSS 0.051268f
C8053 mux8_1.NAND4F_2.D.t0 VSS 0.040771f
C8054 mux8_1.NAND4F_2.D.t6 VSS 0.027742f
C8055 mux8_1.NAND4F_2.D.t12 VSS 0.098211f
C8056 mux8_1.NAND4F_2.D.t7 VSS 0.030538f
C8057 mux8_1.NAND4F_2.D.n4 VSS 0.087112f
C8058 mux8_1.NAND4F_2.D.n5 VSS 0.025813f
C8059 mux8_1.NAND4F_2.D.n6 VSS 0.620222f
C8060 mux8_1.NAND4F_2.D.t14 VSS 0.027742f
C8061 mux8_1.NAND4F_2.D.t9 VSS 0.098211f
C8062 mux8_1.NAND4F_2.D.t15 VSS 0.030538f
C8063 mux8_1.NAND4F_2.D.n7 VSS 0.087112f
C8064 mux8_1.NAND4F_2.D.n8 VSS 0.025807f
C8065 mux8_1.NAND4F_2.D.n9 VSS 0.261852f
C8066 mux8_1.NAND4F_2.D.t5 VSS 0.027742f
C8067 mux8_1.NAND4F_2.D.t4 VSS 0.098211f
C8068 mux8_1.NAND4F_2.D.t8 VSS 0.030538f
C8069 mux8_1.NAND4F_2.D.n10 VSS 0.087112f
C8070 mux8_1.NAND4F_2.D.n11 VSS 0.025808f
C8071 mux8_1.NAND4F_2.D.n12 VSS 0.407824f
C8072 a_n1588_2026.n0 VSS 1.48326f
C8073 a_n1588_2026.n1 VSS 1.48365f
C8074 a_n1588_2026.t0 VSS 0.093341f
C8075 a_n1588_2026.t9 VSS 0.093341f
C8076 a_n1588_2026.t11 VSS 0.093341f
C8077 a_n1588_2026.n2 VSS 0.20269f
C8078 a_n1588_2026.t3 VSS 0.093341f
C8079 a_n1588_2026.t10 VSS 0.093341f
C8080 a_n1588_2026.n3 VSS 0.202001f
C8081 a_n1588_2026.t4 VSS 0.093341f
C8082 a_n1588_2026.t5 VSS 0.093341f
C8083 a_n1588_2026.n4 VSS 0.202001f
C8084 a_n1588_2026.t8 VSS 0.093341f
C8085 a_n1588_2026.t6 VSS 0.093341f
C8086 a_n1588_2026.n5 VSS 0.202001f
C8087 a_n1588_2026.t1 VSS 0.093341f
C8088 a_n1588_2026.t7 VSS 0.093341f
C8089 a_n1588_2026.n6 VSS 0.202001f
C8090 a_n1588_2026.n7 VSS 0.202296f
C8091 a_n1588_2026.t2 VSS 0.093341f
C8092 a_n21333_2026.n0 VSS 1.48365f
C8093 a_n21333_2026.n1 VSS 1.48326f
C8094 a_n21333_2026.t7 VSS 0.093341f
C8095 a_n21333_2026.t6 VSS 0.093341f
C8096 a_n21333_2026.t4 VSS 0.093341f
C8097 a_n21333_2026.n2 VSS 0.202296f
C8098 a_n21333_2026.t5 VSS 0.093341f
C8099 a_n21333_2026.t10 VSS 0.093341f
C8100 a_n21333_2026.n3 VSS 0.202001f
C8101 a_n21333_2026.t9 VSS 0.093341f
C8102 a_n21333_2026.t11 VSS 0.093341f
C8103 a_n21333_2026.n4 VSS 0.202001f
C8104 a_n21333_2026.t8 VSS 0.093341f
C8105 a_n21333_2026.t0 VSS 0.093341f
C8106 a_n21333_2026.n5 VSS 0.202001f
C8107 a_n21333_2026.t1 VSS 0.093341f
C8108 a_n21333_2026.t2 VSS 0.093341f
C8109 a_n21333_2026.n6 VSS 0.20269f
C8110 a_n21333_2026.n7 VSS 0.202001f
C8111 a_n21333_2026.t3 VSS 0.093341f
C8112 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t9 VSS 0.007073f
C8113 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t10 VSS 0.007073f
C8114 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n0 VSS 0.017105f
C8115 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t1 VSS 0.007073f
C8116 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t0 VSS 0.007073f
C8117 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n1 VSS 0.017107f
C8118 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n2 VSS 0.122656f
C8119 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t11 VSS 0.007073f
C8120 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t2 VSS 0.007073f
C8121 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n3 VSS 0.014146f
C8122 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n4 VSS 0.011112f
C8123 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t8 VSS 0.029924f
C8124 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t3 VSS 0.029924f
C8125 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n5 VSS 0.059848f
C8126 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n6 VSS 0.023796f
C8127 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t6 VSS 0.029924f
C8128 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t7 VSS 0.029924f
C8129 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n7 VSS 0.059848f
C8130 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n8 VSS 0.026362f
C8131 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n9 VSS 0.271f
C8132 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t4 VSS 0.029924f
C8133 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t5 VSS 0.029924f
C8134 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n10 VSS 0.059848f
C8135 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n11 VSS 0.026322f
C8136 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n12 VSS 0.173808f
C8137 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n13 VSS 0.03917f
C8138 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n14 VSS 0.172104f
C8139 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t18 VSS 0.043288f
C8140 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t21 VSS 0.014096f
C8141 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t19 VSS 0.019467f
C8142 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n15 VSS 0.020992f
C8143 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t20 VSS 0.014492f
C8144 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n16 VSS 0.036772f
C8145 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n17 VSS 0.064505f
C8146 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t16 VSS 0.019764f
C8147 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t22 VSS 0.039767f
C8148 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t14 VSS 0.039272f
C8149 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t17 VSS 0.039272f
C8150 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t12 VSS 0.039272f
C8151 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t15 VSS 0.008161f
C8152 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t13 VSS 0.008161f
C8153 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.t23 VSS 0.008161f
C8154 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n18 VSS 0.24195f
C8155 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n19 VSS 0.178207f
C8156 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n20 VSS 0.097121f
C8157 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n21 VSS 0.095413f
C8158 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n22 VSS 0.05869f
C8159 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n23 VSS 0.076991f
C8160 8bit_ADDER_0.FULL_ADDER_XORED_1.XOR2_2.Y.n24 VSS 1.26966f
C8161 AND8_0.NOT8_0.A5.n0 VSS 0.826718f
C8162 AND8_0.NOT8_0.A5.t8 VSS 0.020493f
C8163 AND8_0.NOT8_0.A5.t9 VSS 0.028606f
C8164 AND8_0.NOT8_0.A5.t7 VSS 0.028606f
C8165 AND8_0.NOT8_0.A5.n1 VSS 0.09312f
C8166 AND8_0.NOT8_0.A5.t10 VSS 0.032827f
C8167 AND8_0.NOT8_0.A5.n2 VSS 0.286655f
C8168 AND8_0.NOT8_0.A5.t3 VSS 0.097059f
C8169 AND8_0.NOT8_0.A5.t4 VSS 0.01608f
C8170 AND8_0.NOT8_0.A5.t6 VSS 0.01608f
C8171 AND8_0.NOT8_0.A5.n3 VSS 0.03578f
C8172 AND8_0.NOT8_0.A5.t0 VSS 0.01608f
C8173 AND8_0.NOT8_0.A5.t2 VSS 0.01608f
C8174 AND8_0.NOT8_0.A5.n4 VSS 0.035878f
C8175 AND8_0.NOT8_0.A5.t5 VSS 0.01608f
C8176 AND8_0.NOT8_0.A5.t1 VSS 0.01608f
C8177 AND8_0.NOT8_0.A5.n5 VSS 0.03578f
C8178 MULT_0.NAND2_15.Y.n0 VSS 1.243f
C8179 MULT_0.NAND2_15.Y.n1 VSS 0.196728f
C8180 MULT_0.NAND2_15.Y.t1 VSS 0.024231f
C8181 MULT_0.NAND2_15.Y.t2 VSS 0.024231f
C8182 MULT_0.NAND2_15.Y.n2 VSS 0.053917f
C8183 MULT_0.NAND2_15.Y.t6 VSS 0.024231f
C8184 MULT_0.NAND2_15.Y.t4 VSS 0.024231f
C8185 MULT_0.NAND2_15.Y.n3 VSS 0.054064f
C8186 MULT_0.NAND2_15.Y.t3 VSS 0.024231f
C8187 MULT_0.NAND2_15.Y.t5 VSS 0.024231f
C8188 MULT_0.NAND2_15.Y.n4 VSS 0.053917f
C8189 MULT_0.NAND2_15.Y.t0 VSS 0.145972f
C8190 MULT_0.NAND2_15.Y.t8 VSS 0.030881f
C8191 MULT_0.NAND2_15.Y.t7 VSS 0.043107f
C8192 MULT_0.NAND2_15.Y.t9 VSS 0.043107f
C8193 MULT_0.NAND2_15.Y.n5 VSS 0.140705f
C8194 MULT_0.NAND2_15.Y.t10 VSS 0.049217f
C8195 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t16 VSS 0.013766f
C8196 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t22 VSS 0.027698f
C8197 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t12 VSS 0.027354f
C8198 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t17 VSS 0.027354f
C8199 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t18 VSS 0.027354f
C8200 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t13 VSS 0.005684f
C8201 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t23 VSS 0.005684f
C8202 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t14 VSS 0.005684f
C8203 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n0 VSS 0.168523f
C8204 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n1 VSS 0.124125f
C8205 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n2 VSS 0.067647f
C8206 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n3 VSS 0.066457f
C8207 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n4 VSS 0.040879f
C8208 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n5 VSS 0.05311f
C8209 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t15 VSS 0.030151f
C8210 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t19 VSS 0.009818f
C8211 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t21 VSS 0.013559f
C8212 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n6 VSS 0.014622f
C8213 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t20 VSS 0.010094f
C8214 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n7 VSS 0.025612f
C8215 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n8 VSS 0.044927f
C8216 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t2 VSS 0.004926f
C8217 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t0 VSS 0.004926f
C8218 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n9 VSS 0.011915f
C8219 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t7 VSS 0.004926f
C8220 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t3 VSS 0.004926f
C8221 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n10 VSS 0.011914f
C8222 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n11 VSS 0.085433f
C8223 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t1 VSS 0.004926f
C8224 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t8 VSS 0.004926f
C8225 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n12 VSS 0.009853f
C8226 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n13 VSS 0.00774f
C8227 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t11 VSS 0.020843f
C8228 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t4 VSS 0.020843f
C8229 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n14 VSS 0.041685f
C8230 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n15 VSS 0.016575f
C8231 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t10 VSS 0.020843f
C8232 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t9 VSS 0.020843f
C8233 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n16 VSS 0.041685f
C8234 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n17 VSS 0.018334f
C8235 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n18 VSS 0.188757f
C8236 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t6 VSS 0.020843f
C8237 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.t5 VSS 0.020843f
C8238 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n19 VSS 0.041685f
C8239 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n20 VSS 0.018362f
C8240 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n21 VSS 0.12106f
C8241 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n22 VSS 0.027282f
C8242 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_1.A.n23 VSS 0.119748f
C8243 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t7 VSS 0.007073f
C8244 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t8 VSS 0.007073f
C8245 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n0 VSS 0.017105f
C8246 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t10 VSS 0.007073f
C8247 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t11 VSS 0.007073f
C8248 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n1 VSS 0.017107f
C8249 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n2 VSS 0.122656f
C8250 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t6 VSS 0.007073f
C8251 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t9 VSS 0.007073f
C8252 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n3 VSS 0.014146f
C8253 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n4 VSS 0.011112f
C8254 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t3 VSS 0.029924f
C8255 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t2 VSS 0.029924f
C8256 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n5 VSS 0.059848f
C8257 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n6 VSS 0.023796f
C8258 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t4 VSS 0.029924f
C8259 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t5 VSS 0.029924f
C8260 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n7 VSS 0.059848f
C8261 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n8 VSS 0.026362f
C8262 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n9 VSS 0.271f
C8263 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t0 VSS 0.029924f
C8264 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t1 VSS 0.029924f
C8265 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n10 VSS 0.059848f
C8266 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n11 VSS 0.026322f
C8267 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n12 VSS 0.173808f
C8268 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n13 VSS 0.03917f
C8269 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n14 VSS 0.172104f
C8270 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t12 VSS 0.043288f
C8271 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t20 VSS 0.014096f
C8272 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t22 VSS 0.019467f
C8273 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n15 VSS 0.020992f
C8274 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t17 VSS 0.014492f
C8275 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n16 VSS 0.036772f
C8276 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n17 VSS 0.064505f
C8277 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t21 VSS 0.019764f
C8278 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t13 VSS 0.039767f
C8279 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t15 VSS 0.039272f
C8280 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t18 VSS 0.039272f
C8281 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t23 VSS 0.039272f
C8282 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t16 VSS 0.008161f
C8283 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t14 VSS 0.008161f
C8284 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.t19 VSS 0.008161f
C8285 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n18 VSS 0.24195f
C8286 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n19 VSS 0.178207f
C8287 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n20 VSS 0.097121f
C8288 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n21 VSS 0.095413f
C8289 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n22 VSS 0.05869f
C8290 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n23 VSS 0.076991f
C8291 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_2.Y.n24 VSS 1.26966f
C8292 AND8_0.S4.n0 VSS 2.29868f
C8293 AND8_0.S4.t4 VSS 0.111189f
C8294 AND8_0.S4.t5 VSS 0.10818f
C8295 AND8_0.S4.t6 VSS 0.327596f
C8296 AND8_0.S4.n1 VSS 0.557696f
C8297 AND8_0.S4.t2 VSS 0.053301f
C8298 AND8_0.S4.t3 VSS 0.053301f
C8299 AND8_0.S4.n2 VSS 0.118777f
C8300 AND8_0.S4.t1 VSS 0.193322f
C8301 AND8_0.S4.t0 VSS 0.153737f
C8302 AND8_0.NOT8_0.A4.n0 VSS 0.752308f
C8303 AND8_0.NOT8_0.A4.t9 VSS 0.018579f
C8304 AND8_0.NOT8_0.A4.t10 VSS 0.025934f
C8305 AND8_0.NOT8_0.A4.t8 VSS 0.025934f
C8306 AND8_0.NOT8_0.A4.n1 VSS 0.084422f
C8307 AND8_0.NOT8_0.A4.t7 VSS 0.029761f
C8308 AND8_0.NOT8_0.A4.n2 VSS 0.26005f
C8309 AND8_0.NOT8_0.A4.t4 VSS 0.087948f
C8310 AND8_0.NOT8_0.A4.t3 VSS 0.014578f
C8311 AND8_0.NOT8_0.A4.t5 VSS 0.014578f
C8312 AND8_0.NOT8_0.A4.n3 VSS 0.032438f
C8313 AND8_0.NOT8_0.A4.t0 VSS 0.014578f
C8314 AND8_0.NOT8_0.A4.t2 VSS 0.014578f
C8315 AND8_0.NOT8_0.A4.n4 VSS 0.032527f
C8316 AND8_0.NOT8_0.A4.t6 VSS 0.014578f
C8317 AND8_0.NOT8_0.A4.t1 VSS 0.014578f
C8318 AND8_0.NOT8_0.A4.n5 VSS 0.032438f
C8319 a_n20557_n4534.n0 VSS 1.48326f
C8320 a_n20557_n4534.n1 VSS 1.48365f
C8321 a_n20557_n4534.t9 VSS 0.093341f
C8322 a_n20557_n4534.t1 VSS 0.093341f
C8323 a_n20557_n4534.t0 VSS 0.093341f
C8324 a_n20557_n4534.n2 VSS 0.202296f
C8325 a_n20557_n4534.t7 VSS 0.093341f
C8326 a_n20557_n4534.t6 VSS 0.093341f
C8327 a_n20557_n4534.n3 VSS 0.20269f
C8328 a_n20557_n4534.t5 VSS 0.093341f
C8329 a_n20557_n4534.t8 VSS 0.093341f
C8330 a_n20557_n4534.n4 VSS 0.202001f
C8331 a_n20557_n4534.t3 VSS 0.093341f
C8332 a_n20557_n4534.t4 VSS 0.093341f
C8333 a_n20557_n4534.n5 VSS 0.202001f
C8334 a_n20557_n4534.t10 VSS 0.093341f
C8335 a_n20557_n4534.t11 VSS 0.093341f
C8336 a_n20557_n4534.n6 VSS 0.202001f
C8337 a_n20557_n4534.n7 VSS 0.202001f
C8338 a_n20557_n4534.t2 VSS 0.093341f
C8339 MULT_0.4bit_ADDER_0.S0 VSS 4.31108f
C8340 mux8_2.NAND4F_0.A VSS 1.42478f
C8341 MULT_0.S1.t13 VSS 0.072645f
C8342 MULT_0.S1.t12 VSS 0.070679f
C8343 MULT_0.S1.t14 VSS 0.214032f
C8344 MULT_0.S1.n0 VSS 0.364397f
C8345 mux8_2.A1 VSS 8.13292f
C8346 MULT_0.S1.t3 VSS 0.021155f
C8347 MULT_0.S1.t4 VSS 0.021155f
C8348 MULT_0.S1.n1 VSS 0.051165f
C8349 MULT_0.S1.t6 VSS 0.021155f
C8350 MULT_0.S1.t7 VSS 0.021155f
C8351 MULT_0.S1.n2 VSS 0.051159f
C8352 MULT_0.S1.n3 VSS 0.366858f
C8353 MULT_0.S1.t5 VSS 0.021155f
C8354 MULT_0.S1.t8 VSS 0.021155f
C8355 MULT_0.S1.n4 VSS 0.042309f
C8356 MULT_0.S1.n5 VSS 0.033235f
C8357 MULT_0.S1.t0 VSS 0.0895f
C8358 MULT_0.S1.t11 VSS 0.0895f
C8359 MULT_0.S1.n6 VSS 0.179001f
C8360 MULT_0.S1.n7 VSS 0.071173f
C8361 MULT_0.S1.t1 VSS 0.0895f
C8362 MULT_0.S1.t2 VSS 0.0895f
C8363 MULT_0.S1.n8 VSS 0.179001f
C8364 MULT_0.S1.n9 VSS 0.078728f
C8365 MULT_0.S1.n10 VSS 0.810545f
C8366 MULT_0.S1.t10 VSS 0.0895f
C8367 MULT_0.S1.t9 VSS 0.0895f
C8368 MULT_0.S1.n11 VSS 0.179001f
C8369 MULT_0.S1.n12 VSS 0.078847f
C8370 MULT_0.S1.n13 VSS 0.519848f
C8371 MULT_0.S1.n14 VSS 0.117154f
C8372 MULT_0.S1.n15 VSS 0.514212f
C8373 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_1.Y VSS 1.1733f
C8374 a_n15707_n11063.n0 VSS 1.48326f
C8375 a_n15707_n11063.n1 VSS 1.48365f
C8376 a_n15707_n11063.t3 VSS 0.093341f
C8377 a_n15707_n11063.t8 VSS 0.093341f
C8378 a_n15707_n11063.t7 VSS 0.093341f
C8379 a_n15707_n11063.n2 VSS 0.20269f
C8380 a_n15707_n11063.t11 VSS 0.093341f
C8381 a_n15707_n11063.t9 VSS 0.093341f
C8382 a_n15707_n11063.n3 VSS 0.202001f
C8383 a_n15707_n11063.t10 VSS 0.093341f
C8384 a_n15707_n11063.t6 VSS 0.093341f
C8385 a_n15707_n11063.n4 VSS 0.202001f
C8386 a_n15707_n11063.t1 VSS 0.093341f
C8387 a_n15707_n11063.t0 VSS 0.093341f
C8388 a_n15707_n11063.n5 VSS 0.202001f
C8389 a_n15707_n11063.t4 VSS 0.093341f
C8390 a_n15707_n11063.t2 VSS 0.093341f
C8391 a_n15707_n11063.n6 VSS 0.202001f
C8392 a_n15707_n11063.n7 VSS 0.202296f
C8393 a_n15707_n11063.t5 VSS 0.093341f
C8394 mux8_6.NAND4F_9.Y.n0 VSS 0.358256f
C8395 mux8_6.NAND4F_9.Y.t10 VSS 0.017853f
C8396 mux8_6.NAND4F_9.Y.t9 VSS 0.017853f
C8397 mux8_6.NAND4F_9.Y.t13 VSS 0.017853f
C8398 mux8_6.NAND4F_9.Y.t12 VSS 0.017853f
C8399 mux8_6.NAND4F_9.Y.t11 VSS 0.022554f
C8400 mux8_6.NAND4F_9.Y.n1 VSS 0.048188f
C8401 mux8_6.NAND4F_9.Y.n2 VSS 0.030339f
C8402 mux8_6.NAND4F_9.Y.n3 VSS 0.030339f
C8403 mux8_6.NAND4F_9.Y.n4 VSS 0.026149f
C8404 mux8_6.NAND4F_9.Y.t14 VSS 0.014813f
C8405 mux8_6.NAND4F_9.Y.n5 VSS 0.021261f
C8406 mux8_6.NAND4F_9.Y.t2 VSS 0.141821f
C8407 mux8_6.NAND4F_9.Y.t7 VSS 0.017663f
C8408 mux8_6.NAND4F_9.Y.t8 VSS 0.017663f
C8409 mux8_6.NAND4F_9.Y.n6 VSS 0.041015f
C8410 mux8_6.NAND4F_9.Y.t5 VSS 0.017663f
C8411 mux8_6.NAND4F_9.Y.t6 VSS 0.017663f
C8412 mux8_6.NAND4F_9.Y.n7 VSS 0.040893f
C8413 mux8_6.NAND4F_9.Y.t0 VSS 0.017663f
C8414 mux8_6.NAND4F_9.Y.t1 VSS 0.017663f
C8415 mux8_6.NAND4F_9.Y.n8 VSS 0.040893f
C8416 mux8_6.NAND4F_9.Y.t4 VSS 0.017663f
C8417 mux8_6.NAND4F_9.Y.t3 VSS 0.017663f
C8418 mux8_6.NAND4F_9.Y.n9 VSS 0.040893f
C8419 mux8_6.NAND4F_9.Y.n10 VSS 0.168091f
C8420 a_n18998_n7799.n0 VSS 1.48365f
C8421 a_n18998_n7799.n1 VSS 1.48326f
C8422 a_n18998_n7799.t4 VSS 0.093341f
C8423 a_n18998_n7799.t11 VSS 0.093341f
C8424 a_n18998_n7799.t10 VSS 0.093341f
C8425 a_n18998_n7799.n2 VSS 0.202296f
C8426 a_n18998_n7799.t9 VSS 0.093341f
C8427 a_n18998_n7799.t7 VSS 0.093341f
C8428 a_n18998_n7799.n3 VSS 0.202001f
C8429 a_n18998_n7799.t6 VSS 0.093341f
C8430 a_n18998_n7799.t8 VSS 0.093341f
C8431 a_n18998_n7799.n4 VSS 0.202001f
C8432 a_n18998_n7799.t0 VSS 0.093341f
C8433 a_n18998_n7799.t1 VSS 0.093341f
C8434 a_n18998_n7799.n5 VSS 0.202001f
C8435 a_n18998_n7799.t2 VSS 0.093341f
C8436 a_n18998_n7799.t3 VSS 0.093341f
C8437 a_n18998_n7799.n6 VSS 0.202001f
C8438 a_n18998_n7799.n7 VSS 0.20269f
C8439 a_n18998_n7799.t5 VSS 0.093341f
C8440 A6.t15 VSS 0.027744f
C8441 A6.t16 VSS 0.027744f
C8442 A6.t17 VSS 0.027744f
C8443 A6.t10 VSS 0.027744f
C8444 A6.n0 VSS 0.503784f
C8445 A6.t6 VSS 0.13351f
C8446 A6.t22 VSS 0.13351f
C8447 A6.t4 VSS 0.135191f
C8448 A6.t5 VSS 0.13351f
C8449 A6.n1 VSS 0.529645f
C8450 A6.n2 VSS 0.785861f
C8451 A6.t21 VSS 0.124847f
C8452 A6.t3 VSS 0.047922f
C8453 A6.t0 VSS 0.066179f
C8454 A6.n3 VSS 0.076172f
C8455 A6.t2 VSS 0.050373f
C8456 A6.n4 VSS 0.077249f
C8457 A6.n5 VSS 0.319752f
C8458 A6.t20 VSS 0.135191f
C8459 A6.t29 VSS 0.13351f
C8460 A6.t23 VSS 0.13351f
C8461 A6.t8 VSS 0.13351f
C8462 A6.n6 VSS 0.531405f
C8463 A6.t12 VSS 0.027744f
C8464 A6.t25 VSS 0.027744f
C8465 A6.t11 VSS 0.027744f
C8466 A6.t18 VSS 0.027744f
C8467 A6.n7 VSS 0.502024f
C8468 A6.n8 VSS 0.785267f
C8469 A6.n9 VSS 1.56105f
C8470 A6.n10 VSS 2.00131f
C8471 A6.t19 VSS 0.124844f
C8472 A6.t27 VSS 0.063098f
C8473 A6.t28 VSS 0.050445f
C8474 A6.n11 VSS 0.080106f
C8475 A6.t9 VSS 0.050373f
C8476 A6.n12 VSS 0.073876f
C8477 A6.n13 VSS 0.320707f
C8478 A6.n14 VSS 0.586335f
C8479 A6.n15 VSS 4.14521f
C8480 A6.t24 VSS 0.049947f
C8481 A6.t26 VSS 0.060197f
C8482 A6.t14 VSS 0.060197f
C8483 A6.t13 VSS 0.060197f
C8484 A6.t7 VSS 0.060197f
C8485 A6.t1 VSS 0.07605f
C8486 A6.n16 VSS 0.162486f
C8487 A6.n17 VSS 0.102302f
C8488 A6.n18 VSS 0.102302f
C8489 A6.n19 VSS 0.08817f
C8490 A6.n20 VSS 0.072061f
C8491 A6.n21 VSS 15.259001f
C8492 a_n20659_3810.n0 VSS 1.45527f
C8493 a_n20659_3810.n1 VSS 1.45566f
C8494 a_n20659_3810.t8 VSS 0.09158f
C8495 a_n20659_3810.t4 VSS 0.09158f
C8496 a_n20659_3810.t5 VSS 0.09158f
C8497 a_n20659_3810.n2 VSS 0.198865f
C8498 a_n20659_3810.t3 VSS 0.09158f
C8499 a_n20659_3810.t9 VSS 0.09158f
C8500 a_n20659_3810.n3 VSS 0.19819f
C8501 a_n20659_3810.t10 VSS 0.09158f
C8502 a_n20659_3810.t11 VSS 0.09158f
C8503 a_n20659_3810.n4 VSS 0.19819f
C8504 a_n20659_3810.t6 VSS 0.09158f
C8505 a_n20659_3810.t7 VSS 0.09158f
C8506 a_n20659_3810.n5 VSS 0.19819f
C8507 a_n20659_3810.t0 VSS 0.09158f
C8508 a_n20659_3810.t1 VSS 0.09158f
C8509 a_n20659_3810.n6 VSS 0.198479f
C8510 a_n20659_3810.n7 VSS 0.19819f
C8511 a_n20659_3810.t2 VSS 0.09158f
C8512 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n0 VSS 0.887305f
C8513 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t6 VSS 0.007677f
C8514 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t4 VSS 0.007677f
C8515 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n1 VSS 0.017083f
C8516 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t0 VSS 0.007677f
C8517 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t1 VSS 0.007677f
C8518 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n2 VSS 0.01713f
C8519 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t3 VSS 0.007677f
C8520 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t2 VSS 0.007677f
C8521 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n3 VSS 0.017083f
C8522 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t5 VSS 0.046356f
C8523 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t14 VSS 0.026222f
C8524 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t9 VSS 0.025896f
C8525 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t8 VSS 0.025896f
C8526 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t10 VSS 0.025896f
C8527 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n4 VSS 0.103072f
C8528 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t17 VSS 0.005381f
C8529 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t7 VSS 0.005381f
C8530 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t12 VSS 0.005381f
C8531 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t18 VSS 0.005381f
C8532 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n5 VSS 0.097373f
C8533 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n6 VSS 0.152286f
C8534 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t13 VSS 0.024216f
C8535 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t15 VSS 0.009295f
C8536 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t16 VSS 0.012836f
C8537 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n7 VSS 0.014774f
C8538 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.t11 VSS 0.00977f
C8539 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n8 VSS 0.014983f
C8540 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n9 VSS 0.050891f
C8541 MULT_0.4bit_ADDER_2.FULL_ADDER_3.COUT.n10 VSS 0.338427f
C8542 a_n16483_2026.n0 VSS 1.48326f
C8543 a_n16483_2026.n1 VSS 1.48365f
C8544 a_n16483_2026.t3 VSS 0.093341f
C8545 a_n16483_2026.t11 VSS 0.093341f
C8546 a_n16483_2026.t9 VSS 0.093341f
C8547 a_n16483_2026.n2 VSS 0.20269f
C8548 a_n16483_2026.t2 VSS 0.093341f
C8549 a_n16483_2026.t10 VSS 0.093341f
C8550 a_n16483_2026.n3 VSS 0.202001f
C8551 a_n16483_2026.t1 VSS 0.093341f
C8552 a_n16483_2026.t0 VSS 0.093341f
C8553 a_n16483_2026.n4 VSS 0.202001f
C8554 a_n16483_2026.t8 VSS 0.093341f
C8555 a_n16483_2026.t7 VSS 0.093341f
C8556 a_n16483_2026.n5 VSS 0.202001f
C8557 a_n16483_2026.t4 VSS 0.093341f
C8558 a_n16483_2026.t6 VSS 0.093341f
C8559 a_n16483_2026.n6 VSS 0.202001f
C8560 a_n16483_2026.n7 VSS 0.202296f
C8561 a_n16483_2026.t5 VSS 0.093341f
C8562 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n0 VSS 0.860417f
C8563 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t1 VSS 0.007445f
C8564 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t6 VSS 0.007445f
C8565 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n1 VSS 0.016566f
C8566 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t3 VSS 0.007445f
C8567 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t4 VSS 0.007445f
C8568 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n2 VSS 0.016611f
C8569 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t5 VSS 0.007445f
C8570 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t2 VSS 0.007445f
C8571 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n3 VSS 0.016566f
C8572 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t0 VSS 0.044951f
C8573 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t11 VSS 0.025427f
C8574 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t14 VSS 0.025111f
C8575 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t9 VSS 0.025111f
C8576 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t7 VSS 0.025111f
C8577 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n4 VSS 0.099949f
C8578 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t18 VSS 0.005218f
C8579 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t12 VSS 0.005218f
C8580 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t8 VSS 0.005218f
C8581 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t10 VSS 0.005218f
C8582 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n5 VSS 0.094423f
C8583 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n6 VSS 0.147672f
C8584 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t13 VSS 0.023482f
C8585 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t17 VSS 0.009013f
C8586 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t15 VSS 0.012447f
C8587 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n7 VSS 0.014327f
C8588 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.t16 VSS 0.009474f
C8589 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n8 VSS 0.014529f
C8590 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n9 VSS 0.049349f
C8591 8bit_ADDER_0.FULL_ADDER_XORED_3.COUT.n10 VSS 0.328172f
C8592 mux8_2.NAND4F_9.Y.n0 VSS 0.358256f
C8593 mux8_2.NAND4F_9.Y.t13 VSS 0.017853f
C8594 mux8_2.NAND4F_9.Y.t9 VSS 0.017853f
C8595 mux8_2.NAND4F_9.Y.t10 VSS 0.017853f
C8596 mux8_2.NAND4F_9.Y.t11 VSS 0.017853f
C8597 mux8_2.NAND4F_9.Y.t12 VSS 0.022554f
C8598 mux8_2.NAND4F_9.Y.n1 VSS 0.048188f
C8599 mux8_2.NAND4F_9.Y.n2 VSS 0.030339f
C8600 mux8_2.NAND4F_9.Y.n3 VSS 0.030339f
C8601 mux8_2.NAND4F_9.Y.n4 VSS 0.026149f
C8602 mux8_2.NAND4F_9.Y.t14 VSS 0.014813f
C8603 mux8_2.NAND4F_9.Y.n5 VSS 0.021261f
C8604 mux8_2.NAND4F_9.Y.t5 VSS 0.141821f
C8605 mux8_2.NAND4F_9.Y.t1 VSS 0.017663f
C8606 mux8_2.NAND4F_9.Y.t0 VSS 0.017663f
C8607 mux8_2.NAND4F_9.Y.n6 VSS 0.041015f
C8608 mux8_2.NAND4F_9.Y.t3 VSS 0.017663f
C8609 mux8_2.NAND4F_9.Y.t4 VSS 0.017663f
C8610 mux8_2.NAND4F_9.Y.n7 VSS 0.040893f
C8611 mux8_2.NAND4F_9.Y.t2 VSS 0.017663f
C8612 mux8_2.NAND4F_9.Y.t8 VSS 0.017663f
C8613 mux8_2.NAND4F_9.Y.n8 VSS 0.040893f
C8614 mux8_2.NAND4F_9.Y.t6 VSS 0.017663f
C8615 mux8_2.NAND4F_9.Y.t7 VSS 0.017663f
C8616 mux8_2.NAND4F_9.Y.n9 VSS 0.040893f
C8617 mux8_2.NAND4F_9.Y.n10 VSS 0.168091f
C8618 mux8_2.NAND4F_7.Y.n0 VSS 0.11858f
C8619 mux8_2.NAND4F_7.Y.n1 VSS 0.350455f
C8620 mux8_2.NAND4F_7.Y.t3 VSS 0.168166f
C8621 mux8_2.NAND4F_7.Y.t11 VSS 0.022537f
C8622 mux8_2.NAND4F_7.Y.t10 VSS 0.079785f
C8623 mux8_2.NAND4F_7.Y.t9 VSS 0.024808f
C8624 mux8_2.NAND4F_7.Y.n2 VSS 0.070768f
C8625 mux8_2.NAND4F_7.Y.n3 VSS 0.020978f
C8626 mux8_2.NAND4F_7.Y.t0 VSS 0.017278f
C8627 mux8_2.NAND4F_7.Y.t1 VSS 0.017278f
C8628 mux8_2.NAND4F_7.Y.n4 VSS 0.040122f
C8629 mux8_2.NAND4F_7.Y.t8 VSS 0.017278f
C8630 mux8_2.NAND4F_7.Y.t7 VSS 0.017278f
C8631 mux8_2.NAND4F_7.Y.n5 VSS 0.040002f
C8632 mux8_2.NAND4F_7.Y.t5 VSS 0.017278f
C8633 mux8_2.NAND4F_7.Y.t6 VSS 0.017278f
C8634 mux8_2.NAND4F_7.Y.n6 VSS 0.040002f
C8635 mux8_2.NAND4F_7.Y.t2 VSS 0.017278f
C8636 mux8_2.NAND4F_7.Y.t4 VSS 0.017278f
C8637 mux8_2.NAND4F_7.Y.n7 VSS 0.040002f
C8638 a_n14751_2026.n0 VSS 1.48365f
C8639 a_n14751_2026.n1 VSS 1.48326f
C8640 a_n14751_2026.t4 VSS 0.093341f
C8641 a_n14751_2026.t11 VSS 0.093341f
C8642 a_n14751_2026.t10 VSS 0.093341f
C8643 a_n14751_2026.n2 VSS 0.202296f
C8644 a_n14751_2026.t9 VSS 0.093341f
C8645 a_n14751_2026.t0 VSS 0.093341f
C8646 a_n14751_2026.n3 VSS 0.202001f
C8647 a_n14751_2026.t2 VSS 0.093341f
C8648 a_n14751_2026.t1 VSS 0.093341f
C8649 a_n14751_2026.n4 VSS 0.202001f
C8650 a_n14751_2026.t7 VSS 0.093341f
C8651 a_n14751_2026.t8 VSS 0.093341f
C8652 a_n14751_2026.n5 VSS 0.20269f
C8653 a_n14751_2026.t3 VSS 0.093341f
C8654 a_n14751_2026.t6 VSS 0.093341f
C8655 a_n14751_2026.n6 VSS 0.202001f
C8656 a_n14751_2026.n7 VSS 0.202001f
C8657 a_n14751_2026.t5 VSS 0.093341f
C8658 mux8_0.NAND4F_4.Y.n0 VSS 0.480308f
C8659 mux8_0.NAND4F_4.Y.t2 VSS 0.023681f
C8660 mux8_0.NAND4F_4.Y.t3 VSS 0.023681f
C8661 mux8_0.NAND4F_4.Y.n1 VSS 0.054989f
C8662 mux8_0.NAND4F_4.Y.t8 VSS 0.023681f
C8663 mux8_0.NAND4F_4.Y.t7 VSS 0.023681f
C8664 mux8_0.NAND4F_4.Y.n2 VSS 0.054824f
C8665 mux8_0.NAND4F_4.Y.t0 VSS 0.023681f
C8666 mux8_0.NAND4F_4.Y.t1 VSS 0.023681f
C8667 mux8_0.NAND4F_4.Y.n3 VSS 0.054824f
C8668 mux8_0.NAND4F_4.Y.t4 VSS 0.023681f
C8669 mux8_0.NAND4F_4.Y.t5 VSS 0.023681f
C8670 mux8_0.NAND4F_4.Y.n4 VSS 0.054824f
C8671 mux8_0.NAND4F_4.Y.n5 VSS 0.238711f
C8672 mux8_0.NAND4F_4.Y.t9 VSS 0.032831f
C8673 mux8_0.NAND4F_4.Y.t10 VSS 0.031942f
C8674 mux8_0.NAND4F_4.Y.t11 VSS 0.096729f
C8675 mux8_0.NAND4F_4.Y.n6 VSS 0.164667f
C8676 mux8_0.NAND4F_4.Y.t6 VSS 0.190137f
C8677 mux8_0.NAND4F_4.Y.n7 VSS 1.51729f
C8678 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t1 VSS 0.007073f
C8679 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t2 VSS 0.007073f
C8680 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n0 VSS 0.017105f
C8681 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t7 VSS 0.007073f
C8682 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t6 VSS 0.007073f
C8683 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n1 VSS 0.017107f
C8684 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n2 VSS 0.122656f
C8685 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t0 VSS 0.007073f
C8686 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t8 VSS 0.007073f
C8687 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n3 VSS 0.014146f
C8688 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n4 VSS 0.011112f
C8689 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t3 VSS 0.029924f
C8690 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t9 VSS 0.029924f
C8691 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n5 VSS 0.059848f
C8692 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n6 VSS 0.023796f
C8693 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t4 VSS 0.029924f
C8694 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t5 VSS 0.029924f
C8695 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n7 VSS 0.059848f
C8696 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n8 VSS 0.026362f
C8697 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n9 VSS 0.271f
C8698 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t10 VSS 0.029924f
C8699 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t11 VSS 0.029924f
C8700 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n10 VSS 0.059848f
C8701 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n11 VSS 0.026322f
C8702 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n12 VSS 0.173808f
C8703 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n13 VSS 0.03917f
C8704 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n14 VSS 0.172104f
C8705 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t18 VSS 0.043288f
C8706 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t21 VSS 0.014096f
C8707 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t19 VSS 0.019467f
C8708 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n15 VSS 0.020992f
C8709 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t20 VSS 0.014492f
C8710 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n16 VSS 0.036772f
C8711 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n17 VSS 0.064505f
C8712 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t16 VSS 0.019764f
C8713 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t22 VSS 0.039767f
C8714 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t13 VSS 0.039272f
C8715 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t12 VSS 0.039272f
C8716 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t14 VSS 0.039272f
C8717 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t15 VSS 0.008161f
C8718 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t23 VSS 0.008161f
C8719 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.t17 VSS 0.008161f
C8720 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n18 VSS 0.24195f
C8721 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n19 VSS 0.178207f
C8722 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n20 VSS 0.097121f
C8723 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n21 VSS 0.095413f
C8724 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n22 VSS 0.05869f
C8725 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n23 VSS 0.076991f
C8726 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_2.Y.n24 VSS 1.26966f
C8727 MULT_0.4bit_ADDER_0.B2.t1 VSS 0.050264f
C8728 MULT_0.4bit_ADDER_0.B2.t0 VSS 0.0631f
C8729 MULT_0.4bit_ADDER_0.B2.n0 VSS 0.261702f
C8730 MULT_0.4bit_ADDER_0.B2.t2 VSS 0.017397f
C8731 MULT_0.4bit_ADDER_0.B2.t3 VSS 0.017397f
C8732 MULT_0.4bit_ADDER_0.B2.n1 VSS 0.03876f
C8733 MULT_0.4bit_ADDER_0.B2.n2 VSS 2.46335f
C8734 MULT_0.4bit_ADDER_0.B2.t10 VSS 0.012194f
C8735 MULT_0.4bit_ADDER_0.B2.t9 VSS 0.012194f
C8736 MULT_0.4bit_ADDER_0.B2.t4 VSS 0.012194f
C8737 MULT_0.4bit_ADDER_0.B2.n3 VSS 0.361527f
C8738 MULT_0.4bit_ADDER_0.B2.t13 VSS 0.058681f
C8739 MULT_0.4bit_ADDER_0.B2.n4 VSS 0.266281f
C8740 MULT_0.4bit_ADDER_0.B2.t14 VSS 0.058681f
C8741 MULT_0.4bit_ADDER_0.B2.n5 VSS 0.145121f
C8742 MULT_0.4bit_ADDER_0.B2.t15 VSS 0.058681f
C8743 MULT_0.4bit_ADDER_0.B2.n6 VSS 0.142569f
C8744 MULT_0.4bit_ADDER_0.B2.t8 VSS 0.05942f
C8745 MULT_0.4bit_ADDER_0.B2.n7 VSS 0.087696f
C8746 MULT_0.4bit_ADDER_0.B2.t6 VSS 0.029532f
C8747 MULT_0.4bit_ADDER_0.B2.n8 VSS 0.115042f
C8748 MULT_0.4bit_ADDER_0.B2.n9 VSS 1.26771f
C8749 MULT_0.4bit_ADDER_0.B2.n10 VSS 0.096385f
C8750 MULT_0.4bit_ADDER_0.B2.t7 VSS 0.064682f
C8751 MULT_0.4bit_ADDER_0.B2.t12 VSS 0.029087f
C8752 MULT_0.4bit_ADDER_0.B2.t11 VSS 0.021063f
C8753 MULT_0.4bit_ADDER_0.B2.n11 VSS 0.031367f
C8754 MULT_0.4bit_ADDER_0.B2.n12 VSS 0.054945f
C8755 MULT_0.4bit_ADDER_0.B2.t5 VSS 0.021654f
C8756 MULT_0.4bit_ADDER_0.B2.n13 VSS 0.214651f
C8757 MULT_0.4bit_ADDER_0.B2.n14 VSS 0.014422f
C8758 mux8_7.NAND4F_1.Y.n0 VSS 0.655599f
C8759 mux8_7.NAND4F_1.Y.t6 VSS 0.306614f
C8760 mux8_7.NAND4F_1.Y.t11 VSS 0.132168f
C8761 mux8_7.NAND4F_1.Y.t10 VSS 0.04216f
C8762 mux8_7.NAND4F_1.Y.t9 VSS 0.04216f
C8763 mux8_7.NAND4F_1.Y.n1 VSS 0.049498f
C8764 mux8_7.NAND4F_1.Y.n2 VSS 0.277534f
C8765 mux8_7.NAND4F_1.Y.t1 VSS 0.032323f
C8766 mux8_7.NAND4F_1.Y.t0 VSS 0.032323f
C8767 mux8_7.NAND4F_1.Y.n3 VSS 0.075057f
C8768 mux8_7.NAND4F_1.Y.t3 VSS 0.032323f
C8769 mux8_7.NAND4F_1.Y.t2 VSS 0.032323f
C8770 mux8_7.NAND4F_1.Y.n4 VSS 0.074832f
C8771 mux8_7.NAND4F_1.Y.t8 VSS 0.032323f
C8772 mux8_7.NAND4F_1.Y.t7 VSS 0.032323f
C8773 mux8_7.NAND4F_1.Y.n5 VSS 0.074832f
C8774 mux8_7.NAND4F_1.Y.t4 VSS 0.032323f
C8775 mux8_7.NAND4F_1.Y.t5 VSS 0.032323f
C8776 mux8_7.NAND4F_1.Y.n6 VSS 0.074832f
C8777 mux8_7.NAND4F_1.Y.n7 VSS 0.307603f
C8778 mux8_7.NAND4F_0.C.n0 VSS 1.68955f
C8779 mux8_7.NAND4F_0.C.t12 VSS 0.23388f
C8780 mux8_7.NAND4F_0.C.t7 VSS 0.074606f
C8781 mux8_7.NAND4F_0.C.t6 VSS 0.074606f
C8782 mux8_7.NAND4F_0.C.n1 VSS 0.087589f
C8783 mux8_7.NAND4F_0.C.n2 VSS 0.491098f
C8784 mux8_7.NAND4F_0.C.t13 VSS 0.074606f
C8785 mux8_7.NAND4F_0.C.t14 VSS 0.074606f
C8786 mux8_7.NAND4F_0.C.n3 VSS 0.087589f
C8787 mux8_7.NAND4F_0.C.t11 VSS 0.23388f
C8788 mux8_7.NAND4F_0.C.n4 VSS 0.491129f
C8789 mux8_7.NAND4F_0.C.t9 VSS 0.074606f
C8790 mux8_7.NAND4F_0.C.t10 VSS 0.074606f
C8791 mux8_7.NAND4F_0.C.n5 VSS 0.087589f
C8792 mux8_7.NAND4F_0.C.t15 VSS 0.23388f
C8793 mux8_7.NAND4F_0.C.n6 VSS 0.491143f
C8794 mux8_7.NAND4F_0.C.n7 VSS 1.79123f
C8795 mux8_7.NAND4F_0.C.t3 VSS 0.038013f
C8796 mux8_7.NAND4F_0.C.t2 VSS 0.038013f
C8797 mux8_7.NAND4F_0.C.n8 VSS 0.08471f
C8798 mux8_7.NAND4F_0.C.t1 VSS 0.137874f
C8799 mux8_7.NAND4F_0.C.t0 VSS 0.109643f
C8800 mux8_7.NAND4F_0.C.n9 VSS 3.13611f
C8801 mux8_7.NAND4F_0.C.t8 VSS 0.23388f
C8802 mux8_7.NAND4F_0.C.t5 VSS 0.074606f
C8803 mux8_7.NAND4F_0.C.t4 VSS 0.074606f
C8804 mux8_7.NAND4F_0.C.n10 VSS 0.087589f
C8805 mux8_7.NAND4F_0.C.n11 VSS 0.491115f
C8806 mux8_7.NAND4F_0.C.n12 VSS 2.51327f
C8807 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t1 VSS 0.007073f
C8808 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t5 VSS 0.007073f
C8809 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n0 VSS 0.017105f
C8810 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t9 VSS 0.007073f
C8811 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t8 VSS 0.007073f
C8812 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n1 VSS 0.017107f
C8813 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n2 VSS 0.122656f
C8814 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t3 VSS 0.007073f
C8815 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t10 VSS 0.007073f
C8816 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n3 VSS 0.014146f
C8817 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n4 VSS 0.011112f
C8818 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t4 VSS 0.029924f
C8819 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t7 VSS 0.029924f
C8820 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n5 VSS 0.059848f
C8821 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n6 VSS 0.023796f
C8822 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t2 VSS 0.029924f
C8823 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t0 VSS 0.029924f
C8824 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n7 VSS 0.059848f
C8825 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n8 VSS 0.026362f
C8826 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n9 VSS 0.271f
C8827 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t6 VSS 0.029924f
C8828 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t11 VSS 0.029924f
C8829 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n10 VSS 0.059848f
C8830 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n11 VSS 0.026322f
C8831 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n12 VSS 0.173808f
C8832 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n13 VSS 0.03917f
C8833 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n14 VSS 0.172104f
C8834 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t15 VSS 0.043288f
C8835 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t17 VSS 0.014096f
C8836 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t18 VSS 0.019467f
C8837 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n15 VSS 0.020992f
C8838 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t16 VSS 0.014492f
C8839 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n16 VSS 0.036772f
C8840 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n17 VSS 0.064505f
C8841 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t13 VSS 0.019764f
C8842 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t20 VSS 0.039767f
C8843 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t22 VSS 0.039272f
C8844 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t14 VSS 0.039272f
C8845 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t19 VSS 0.039272f
C8846 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t23 VSS 0.008161f
C8847 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t21 VSS 0.008161f
C8848 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.t12 VSS 0.008161f
C8849 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n18 VSS 0.24195f
C8850 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n19 VSS 0.178207f
C8851 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n20 VSS 0.097121f
C8852 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n21 VSS 0.095413f
C8853 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n22 VSS 0.05869f
C8854 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n23 VSS 0.076991f
C8855 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_2.Y.n24 VSS 1.26966f
C8856 B3.t21 VSS 0.055789f
C8857 B3.t16 VSS 0.05984f
C8858 B3.n0 VSS 0.089168f
C8859 B3.t25 VSS 0.055789f
C8860 B3.t42 VSS 0.055789f
C8861 B3.t46 VSS 0.055789f
C8862 B3.t8 VSS 0.07048f
C8863 B3.n1 VSS 0.150586f
C8864 B3.n2 VSS 0.094809f
C8865 B3.n3 VSS 0.07747f
C8866 B3.n4 VSS 0.037908f
C8867 B3.t19 VSS 0.04675f
C8868 B3.t24 VSS 0.065259f
C8869 B3.t23 VSS 0.065259f
C8870 B3.n5 VSS 0.212434f
C8871 B3.t6 VSS 0.074888f
C8872 B3.n6 VSS 0.528106f
C8873 B3.n7 VSS 0.603493f
C8874 B3.t10 VSS 0.04675f
C8875 B3.t36 VSS 0.065259f
C8876 B3.t9 VSS 0.065259f
C8877 B3.n8 VSS 0.212434f
C8878 B3.t45 VSS 0.074888f
C8879 B3.n9 VSS 0.525484f
C8880 B3.n10 VSS 0.466549f
C8881 B3.n11 VSS 3.02523f
C8882 B3.t1 VSS 0.04675f
C8883 B3.t39 VSS 0.065259f
C8884 B3.t37 VSS 0.065259f
C8885 B3.n12 VSS 0.212434f
C8886 B3.t27 VSS 0.074888f
C8887 B3.n13 VSS 0.640608f
C8888 B3.n14 VSS 0.461903f
C8889 B3.n15 VSS 4.88433f
C8890 B3.t40 VSS 0.062271f
C8891 B3.t13 VSS 0.12529f
C8892 B3.t35 VSS 0.123732f
C8893 B3.t12 VSS 0.123732f
C8894 B3.t49 VSS 0.123732f
C8895 B3.t53 VSS 0.025713f
C8896 B3.t20 VSS 0.025713f
C8897 B3.t3 VSS 0.025713f
C8898 B3.n16 VSS 0.762107f
C8899 B3.n17 VSS 0.56166f
C8900 B3.n18 VSS 0.305995f
C8901 B3.n19 VSS 0.300614f
C8902 B3.n20 VSS 0.184913f
C8903 B3.n21 VSS 0.237946f
C8904 B3.n22 VSS 6.69274f
C8905 B3.n23 VSS 6.05689f
C8906 B3.t11 VSS 0.062271f
C8907 B3.t15 VSS 0.12529f
C8908 B3.t47 VSS 0.123732f
C8909 B3.t38 VSS 0.123732f
C8910 B3.t26 VSS 0.123732f
C8911 B3.t34 VSS 0.025713f
C8912 B3.t14 VSS 0.025713f
C8913 B3.t0 VSS 0.025713f
C8914 B3.n24 VSS 0.762299f
C8915 B3.n25 VSS 0.561468f
C8916 B3.n26 VSS 0.305995f
C8917 B3.n27 VSS 0.300614f
C8918 B3.n28 VSS 0.184913f
C8919 B3.n29 VSS 0.210283f
C8920 B3.t31 VSS 0.115704f
C8921 B3.t28 VSS 0.044413f
C8922 B3.t30 VSS 0.061333f
C8923 B3.n30 VSS 0.070593f
C8924 B3.t4 VSS 0.046684f
C8925 B3.n31 VSS 0.071592f
C8926 B3.n32 VSS 0.297073f
C8927 B3.t48 VSS 0.136385f
C8928 B3.t2 VSS 0.044413f
C8929 B3.t5 VSS 0.061333f
C8930 B3.n33 VSS 0.06614f
C8931 B3.t43 VSS 0.04566f
C8932 B3.n34 VSS 0.115855f
C8933 B3.n35 VSS 0.203599f
C8934 B3.n36 VSS 2.80972f
C8935 B3.t17 VSS 0.115704f
C8936 B3.t32 VSS 0.044413f
C8937 B3.t51 VSS 0.061333f
C8938 B3.n37 VSS 0.070593f
C8939 B3.t50 VSS 0.046684f
C8940 B3.n38 VSS 0.071592f
C8941 B3.n39 VSS 0.297073f
C8942 B3.t41 VSS 0.136385f
C8943 B3.t33 VSS 0.044413f
C8944 B3.t52 VSS 0.061333f
C8945 B3.n40 VSS 0.06614f
C8946 B3.t29 VSS 0.04566f
C8947 B3.n41 VSS 0.115855f
C8948 B3.n42 VSS 0.203599f
C8949 B3.n43 VSS 3.26772f
C8950 B3.n44 VSS 21.271599f
C8951 B3.t7 VSS 0.136542f
C8952 B3.t18 VSS 0.058477f
C8953 B3.t22 VSS 0.04675f
C8954 B3.n45 VSS 0.068995f
C8955 B3.t44 VSS 0.04566f
C8956 B3.n46 VSS 0.113899f
C8957 B3.n47 VSS 0.203207f
C8958 B3.n48 VSS 0.306442f
C8959 B3.n49 VSS 0.078154f
C8960 B3.n50 VSS 3.00916f
C8961 B5.t11 VSS 0.057388f
C8962 B5.t18 VSS 0.080109f
C8963 B5.t14 VSS 0.080109f
C8964 B5.n0 VSS 0.260773f
C8965 B5.t3 VSS 0.091928f
C8966 B5.n1 VSS 0.647349f
C8967 B5.t23 VSS 0.07644f
C8968 B5.t27 VSS 0.1538f
C8969 B5.t21 VSS 0.151887f
C8970 B5.t2 VSS 0.151887f
C8971 B5.t33 VSS 0.151887f
C8972 B5.t36 VSS 0.031563f
C8973 B5.t9 VSS 0.031563f
C8974 B5.t19 VSS 0.031563f
C8975 B5.n2 VSS 0.935756f
C8976 B5.n3 VSS 0.689227f
C8977 B5.n4 VSS 0.375623f
C8978 B5.n5 VSS 0.369017f
C8979 B5.n6 VSS 0.226988f
C8980 B5.n7 VSS 0.258132f
C8981 B5.t6 VSS 0.167611f
C8982 B5.t15 VSS 0.071783f
C8983 B5.t29 VSS 0.057388f
C8984 B5.n8 VSS 0.084695f
C8985 B5.t1 VSS 0.056049f
C8986 B5.n9 VSS 0.139817f
C8987 B5.n10 VSS 0.249446f
C8988 B5.n11 VSS 0.411813f
C8989 B5.n12 VSS 25.6608f
C8990 B5.t17 VSS 0.068483f
C8991 B5.t13 VSS 0.073456f
C8992 B5.n13 VSS 0.109458f
C8993 B5.t20 VSS 0.068483f
C8994 B5.t31 VSS 0.068483f
C8995 B5.t34 VSS 0.068483f
C8996 B5.t5 VSS 0.086517f
C8997 B5.n14 VSS 0.184851f
C8998 B5.n15 VSS 0.116383f
C8999 B5.n16 VSS 0.095098f
C9000 B5.n17 VSS 0.046534f
C9001 B5.n18 VSS 9.30811f
C9002 B5.t26 VSS 0.07644f
C9003 B5.t7 VSS 0.1538f
C9004 B5.t22 VSS 0.151887f
C9005 B5.t4 VSS 0.151887f
C9006 B5.t32 VSS 0.151887f
C9007 B5.t35 VSS 0.031563f
C9008 B5.t8 VSS 0.031563f
C9009 B5.t37 VSS 0.031563f
C9010 B5.n19 VSS 0.93552f
C9011 B5.n20 VSS 0.689463f
C9012 B5.n21 VSS 0.375623f
C9013 B5.n22 VSS 0.369017f
C9014 B5.n23 VSS 0.226988f
C9015 B5.n24 VSS 0.29209f
C9016 B5.n25 VSS 12.767599f
C9017 B5.t0 VSS 0.057388f
C9018 B5.t25 VSS 0.080109f
C9019 B5.t24 VSS 0.080109f
C9020 B5.n26 VSS 0.260773f
C9021 B5.t16 VSS 0.091928f
C9022 B5.n27 VSS 0.789037f
C9023 B5.n28 VSS 0.485593f
C9024 B5.n29 VSS 9.02913f
C9025 B5.t12 VSS 0.057388f
C9026 B5.t30 VSS 0.080109f
C9027 B5.t10 VSS 0.080109f
C9028 B5.n30 VSS 0.260773f
C9029 B5.t28 VSS 0.091928f
C9030 B5.n31 VSS 0.645512f
C9031 B5.n32 VSS 0.573311f
C9032 B5.n33 VSS 4.386509f
C9033 B5.n34 VSS 0.745263f
C9034 right_shifter_0.S0.n0 VSS 11.7812f
C9035 mux8_1.NAND4F_6.A VSS 0.917785f
C9036 right_shifter_0.S0.t4 VSS 0.069524f
C9037 right_shifter_0.S0.t5 VSS 0.204839f
C9038 right_shifter_0.S0.t6 VSS 0.067643f
C9039 right_shifter_0.S0.n1 VSS 0.348745f
C9040 right_shifter_0.S0.t1 VSS 0.033328f
C9041 right_shifter_0.S0.t2 VSS 0.033328f
C9042 right_shifter_0.S0.n2 VSS 0.074269f
C9043 right_shifter_0.S0.t3 VSS 0.12088f
C9044 right_shifter_0.S0.t0 VSS 0.096129f
C9045 mux8_1.A7 VSS 11.0523f
C9046 A0.t41 VSS 0.025817f
C9047 A0.t31 VSS 0.025817f
C9048 A0.t44 VSS 0.025817f
C9049 A0.t29 VSS 0.025817f
C9050 A0.n0 VSS 0.468783f
C9051 A0.t21 VSS 0.124234f
C9052 A0.t4 VSS 0.124234f
C9053 A0.t16 VSS 0.125799f
C9054 A0.t5 VSS 0.124234f
C9055 A0.n1 VSS 0.492848f
C9056 A0.n2 VSS 0.731262f
C9057 A0.t22 VSS 0.116174f
C9058 A0.t25 VSS 0.044593f
C9059 A0.t26 VSS 0.061581f
C9060 A0.n3 VSS 0.07088f
C9061 A0.t24 VSS 0.046873f
C9062 A0.n4 VSS 0.071882f
C9063 A0.n5 VSS 0.297536f
C9064 A0.t32 VSS 0.125799f
C9065 A0.t45 VSS 0.124234f
C9066 A0.t36 VSS 0.124234f
C9067 A0.t19 VSS 0.124234f
C9068 A0.n6 VSS 0.494485f
C9069 A0.t12 VSS 0.025817f
C9070 A0.t1 VSS 0.025817f
C9071 A0.t9 VSS 0.025817f
C9072 A0.t30 VSS 0.025817f
C9073 A0.n7 VSS 0.467145f
C9074 A0.n8 VSS 0.730709f
C9075 A0.n9 VSS 1.4526f
C9076 A0.n10 VSS 1.86227f
C9077 A0.t20 VSS 0.136939f
C9078 A0.t11 VSS 0.044593f
C9079 A0.t43 VSS 0.061581f
C9080 A0.n11 VSS 0.066408f
C9081 A0.t14 VSS 0.045845f
C9082 A0.n12 VSS 0.116326f
C9083 A0.n13 VSS 0.204425f
C9084 A0.t8 VSS 0.136939f
C9085 A0.t3 VSS 0.044593f
C9086 A0.t34 VSS 0.061581f
C9087 A0.n14 VSS 0.066408f
C9088 A0.t7 VSS 0.045845f
C9089 A0.n15 VSS 0.116326f
C9090 A0.n16 VSS 0.204425f
C9091 A0.t27 VSS 0.116174f
C9092 A0.t42 VSS 0.044593f
C9093 A0.t38 VSS 0.061581f
C9094 A0.n17 VSS 0.07088f
C9095 A0.t10 VSS 0.046873f
C9096 A0.n18 VSS 0.071882f
C9097 A0.n19 VSS 0.298279f
C9098 A0.n20 VSS 11.620099f
C9099 A0.n21 VSS 5.75284f
C9100 A0.t33 VSS 0.136939f
C9101 A0.t23 VSS 0.044593f
C9102 A0.t39 VSS 0.061581f
C9103 A0.n22 VSS 0.066408f
C9104 A0.t17 VSS 0.045845f
C9105 A0.n23 VSS 0.116326f
C9106 A0.n24 VSS 0.204425f
C9107 A0.n25 VSS 3.29156f
C9108 A0.n26 VSS 28.1041f
C9109 A0.t13 VSS 0.11617f
C9110 A0.t28 VSS 0.058714f
C9111 A0.t40 VSS 0.04694f
C9112 A0.n27 VSS 0.074541f
C9113 A0.t6 VSS 0.046873f
C9114 A0.n28 VSS 0.068743f
C9115 A0.n29 VSS 0.298425f
C9116 A0.n30 VSS 0.521869f
C9117 A0.n31 VSS 3.25728f
C9118 A0.t35 VSS 0.046477f
C9119 A0.t37 VSS 0.056015f
C9120 A0.t18 VSS 0.056015f
C9121 A0.t15 VSS 0.056015f
C9122 A0.t2 VSS 0.056015f
C9123 A0.t0 VSS 0.070766f
C9124 A0.n32 VSS 0.151197f
C9125 A0.n33 VSS 0.095194f
C9126 A0.n34 VSS 0.095194f
C9127 A0.n35 VSS 0.082044f
C9128 A0.n36 VSS 0.067055f
C9129 A0.n37 VSS 6.80143f
C9130 A0.n38 VSS 1.02699f
C9131 A0.n39 VSS 0.076387f
C9132 mux8_2.NAND4F_4.Y.n0 VSS 0.480308f
C9133 mux8_2.NAND4F_4.Y.t6 VSS 0.023681f
C9134 mux8_2.NAND4F_4.Y.t5 VSS 0.023681f
C9135 mux8_2.NAND4F_4.Y.n1 VSS 0.054989f
C9136 mux8_2.NAND4F_4.Y.t4 VSS 0.023681f
C9137 mux8_2.NAND4F_4.Y.t3 VSS 0.023681f
C9138 mux8_2.NAND4F_4.Y.n2 VSS 0.054824f
C9139 mux8_2.NAND4F_4.Y.t8 VSS 0.023681f
C9140 mux8_2.NAND4F_4.Y.t7 VSS 0.023681f
C9141 mux8_2.NAND4F_4.Y.n3 VSS 0.054824f
C9142 mux8_2.NAND4F_4.Y.t2 VSS 0.023681f
C9143 mux8_2.NAND4F_4.Y.t1 VSS 0.023681f
C9144 mux8_2.NAND4F_4.Y.n4 VSS 0.054824f
C9145 mux8_2.NAND4F_4.Y.n5 VSS 0.238711f
C9146 mux8_2.NAND4F_4.Y.t10 VSS 0.032831f
C9147 mux8_2.NAND4F_4.Y.t9 VSS 0.031942f
C9148 mux8_2.NAND4F_4.Y.t11 VSS 0.096729f
C9149 mux8_2.NAND4F_4.Y.n6 VSS 0.164667f
C9150 mux8_2.NAND4F_4.Y.t0 VSS 0.190137f
C9151 mux8_2.NAND4F_4.Y.n7 VSS 1.51729f
C9152 mux8_0.NAND4F_2.D.n0 VSS 0.664607f
C9153 mux8_0.NAND4F_2.D.t8 VSS 0.027742f
C9154 mux8_0.NAND4F_2.D.t7 VSS 0.098211f
C9155 mux8_0.NAND4F_2.D.t6 VSS 0.030538f
C9156 mux8_0.NAND4F_2.D.n1 VSS 0.087112f
C9157 mux8_0.NAND4F_2.D.n2 VSS 0.025808f
C9158 mux8_0.NAND4F_2.D.t2 VSS 0.014135f
C9159 mux8_0.NAND4F_2.D.t3 VSS 0.014135f
C9160 mux8_0.NAND4F_2.D.n3 VSS 0.031499f
C9161 mux8_0.NAND4F_2.D.t1 VSS 0.051268f
C9162 mux8_0.NAND4F_2.D.t0 VSS 0.040771f
C9163 mux8_0.NAND4F_2.D.t4 VSS 0.027742f
C9164 mux8_0.NAND4F_2.D.t13 VSS 0.098211f
C9165 mux8_0.NAND4F_2.D.t12 VSS 0.030538f
C9166 mux8_0.NAND4F_2.D.n4 VSS 0.087112f
C9167 mux8_0.NAND4F_2.D.n5 VSS 0.025813f
C9168 mux8_0.NAND4F_2.D.n6 VSS 0.620222f
C9169 mux8_0.NAND4F_2.D.t15 VSS 0.027742f
C9170 mux8_0.NAND4F_2.D.t5 VSS 0.098211f
C9171 mux8_0.NAND4F_2.D.t11 VSS 0.030538f
C9172 mux8_0.NAND4F_2.D.n7 VSS 0.087112f
C9173 mux8_0.NAND4F_2.D.n8 VSS 0.025807f
C9174 mux8_0.NAND4F_2.D.n9 VSS 0.261852f
C9175 mux8_0.NAND4F_2.D.t14 VSS 0.027742f
C9176 mux8_0.NAND4F_2.D.t9 VSS 0.098211f
C9177 mux8_0.NAND4F_2.D.t10 VSS 0.030538f
C9178 mux8_0.NAND4F_2.D.n10 VSS 0.087112f
C9179 mux8_0.NAND4F_2.D.n11 VSS 0.025808f
C9180 mux8_0.NAND4F_2.D.n12 VSS 0.407824f
C9181 V_FLAG_0.XOR2_2.B.t16 VSS 0.035749f
C9182 V_FLAG_0.XOR2_2.B.t13 VSS 0.035304f
C9183 V_FLAG_0.XOR2_2.B.t15 VSS 0.035304f
C9184 V_FLAG_0.XOR2_2.B.t17 VSS 0.035304f
C9185 V_FLAG_0.XOR2_2.B.n0 VSS 0.14052f
C9186 V_FLAG_0.XOR2_2.B.t19 VSS 0.007337f
C9187 V_FLAG_0.XOR2_2.B.t14 VSS 0.007337f
C9188 V_FLAG_0.XOR2_2.B.t12 VSS 0.007337f
C9189 V_FLAG_0.XOR2_2.B.t18 VSS 0.007337f
C9190 V_FLAG_0.XOR2_2.B.n1 VSS 0.132751f
C9191 V_FLAG_0.XOR2_2.B.n2 VSS 0.207798f
C9192 V_FLAG_0.XOR2_2.B.t3 VSS 0.006358f
C9193 V_FLAG_0.XOR2_2.B.t1 VSS 0.006358f
C9194 V_FLAG_0.XOR2_2.B.n3 VSS 0.015378f
C9195 V_FLAG_0.XOR2_2.B.t6 VSS 0.006358f
C9196 V_FLAG_0.XOR2_2.B.t11 VSS 0.006358f
C9197 V_FLAG_0.XOR2_2.B.n4 VSS 0.015377f
C9198 V_FLAG_0.XOR2_2.B.n5 VSS 0.110264f
C9199 V_FLAG_0.XOR2_2.B.t2 VSS 0.006358f
C9200 V_FLAG_0.XOR2_2.B.t4 VSS 0.006358f
C9201 V_FLAG_0.XOR2_2.B.n6 VSS 0.012717f
C9202 V_FLAG_0.XOR2_2.B.n7 VSS 0.009989f
C9203 V_FLAG_0.XOR2_2.B.t10 VSS 0.026901f
C9204 V_FLAG_0.XOR2_2.B.t5 VSS 0.026901f
C9205 V_FLAG_0.XOR2_2.B.n8 VSS 0.053801f
C9206 V_FLAG_0.XOR2_2.B.n9 VSS 0.021392f
C9207 V_FLAG_0.XOR2_2.B.t8 VSS 0.026901f
C9208 V_FLAG_0.XOR2_2.B.t9 VSS 0.026901f
C9209 V_FLAG_0.XOR2_2.B.n10 VSS 0.053801f
C9210 V_FLAG_0.XOR2_2.B.n11 VSS 0.023663f
C9211 V_FLAG_0.XOR2_2.B.n12 VSS 0.24362f
C9212 V_FLAG_0.XOR2_2.B.t7 VSS 0.026901f
C9213 V_FLAG_0.XOR2_2.B.t0 VSS 0.026901f
C9214 V_FLAG_0.XOR2_2.B.n13 VSS 0.053801f
C9215 V_FLAG_0.XOR2_2.B.n14 VSS 0.023698f
C9216 V_FLAG_0.XOR2_2.B.n15 VSS 0.156247f
C9217 V_FLAG_0.XOR2_2.B.n16 VSS 0.035212f
C9218 V_FLAG_0.XOR2_2.B.n17 VSS 0.154552f
C9219 mux8_6.NAND4F_8.Y.n0 VSS 0.539804f
C9220 mux8_6.NAND4F_8.Y.t9 VSS 0.026899f
C9221 mux8_6.NAND4F_8.Y.t14 VSS 0.028853f
C9222 mux8_6.NAND4F_8.Y.n1 VSS 0.042994f
C9223 mux8_6.NAND4F_8.Y.t10 VSS 0.026899f
C9224 mux8_6.NAND4F_8.Y.t12 VSS 0.026899f
C9225 mux8_6.NAND4F_8.Y.t11 VSS 0.026899f
C9226 mux8_6.NAND4F_8.Y.t13 VSS 0.033983f
C9227 mux8_6.NAND4F_8.Y.n2 VSS 0.072608f
C9228 mux8_6.NAND4F_8.Y.n3 VSS 0.045714f
C9229 mux8_6.NAND4F_8.Y.n4 VSS 0.037354f
C9230 mux8_6.NAND4F_8.Y.n5 VSS 0.018278f
C9231 mux8_6.NAND4F_8.Y.t1 VSS 0.026614f
C9232 mux8_6.NAND4F_8.Y.t0 VSS 0.026614f
C9233 mux8_6.NAND4F_8.Y.n6 VSS 0.0618f
C9234 mux8_6.NAND4F_8.Y.t5 VSS 0.026614f
C9235 mux8_6.NAND4F_8.Y.t6 VSS 0.026614f
C9236 mux8_6.NAND4F_8.Y.n7 VSS 0.061615f
C9237 mux8_6.NAND4F_8.Y.t7 VSS 0.026614f
C9238 mux8_6.NAND4F_8.Y.t8 VSS 0.026614f
C9239 mux8_6.NAND4F_8.Y.n8 VSS 0.061615f
C9240 mux8_6.NAND4F_8.Y.t3 VSS 0.026614f
C9241 mux8_6.NAND4F_8.Y.t4 VSS 0.026614f
C9242 mux8_6.NAND4F_8.Y.n9 VSS 0.061615f
C9243 mux8_6.NAND4F_8.Y.n10 VSS 0.268281f
C9244 mux8_6.NAND4F_8.Y.t2 VSS 0.21369f
C9245 mux8_6.NAND4F_4.Y.n0 VSS 0.480308f
C9246 mux8_6.NAND4F_4.Y.t0 VSS 0.023681f
C9247 mux8_6.NAND4F_4.Y.t1 VSS 0.023681f
C9248 mux8_6.NAND4F_4.Y.n1 VSS 0.054989f
C9249 mux8_6.NAND4F_4.Y.t5 VSS 0.023681f
C9250 mux8_6.NAND4F_4.Y.t6 VSS 0.023681f
C9251 mux8_6.NAND4F_4.Y.n2 VSS 0.054824f
C9252 mux8_6.NAND4F_4.Y.t8 VSS 0.023681f
C9253 mux8_6.NAND4F_4.Y.t7 VSS 0.023681f
C9254 mux8_6.NAND4F_4.Y.n3 VSS 0.054824f
C9255 mux8_6.NAND4F_4.Y.t2 VSS 0.023681f
C9256 mux8_6.NAND4F_4.Y.t3 VSS 0.023681f
C9257 mux8_6.NAND4F_4.Y.n4 VSS 0.054824f
C9258 mux8_6.NAND4F_4.Y.n5 VSS 0.238711f
C9259 mux8_6.NAND4F_4.Y.t11 VSS 0.032831f
C9260 mux8_6.NAND4F_4.Y.t9 VSS 0.031942f
C9261 mux8_6.NAND4F_4.Y.t10 VSS 0.096729f
C9262 mux8_6.NAND4F_4.Y.n6 VSS 0.164667f
C9263 mux8_6.NAND4F_4.Y.t4 VSS 0.190137f
C9264 mux8_6.NAND4F_4.Y.n7 VSS 1.51729f
C9265 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n0 VSS 0.967969f
C9266 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t1 VSS 0.008375f
C9267 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t2 VSS 0.008375f
C9268 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n1 VSS 0.018687f
C9269 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t4 VSS 0.008375f
C9270 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t0 VSS 0.008375f
C9271 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n2 VSS 0.018636f
C9272 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t6 VSS 0.008375f
C9273 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t5 VSS 0.008375f
C9274 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n3 VSS 0.018636f
C9275 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t3 VSS 0.05057f
C9276 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t7 VSS 0.028606f
C9277 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t16 VSS 0.02825f
C9278 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t17 VSS 0.02825f
C9279 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t12 VSS 0.02825f
C9280 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n4 VSS 0.112442f
C9281 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t14 VSS 0.005871f
C9282 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t9 VSS 0.005871f
C9283 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t18 VSS 0.005871f
C9284 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t13 VSS 0.005871f
C9285 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n5 VSS 0.106225f
C9286 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n6 VSS 0.166131f
C9287 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t8 VSS 0.026417f
C9288 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t11 VSS 0.01014f
C9289 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t10 VSS 0.014003f
C9290 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n7 VSS 0.016118f
C9291 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.t15 VSS 0.010659f
C9292 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n8 VSS 0.016345f
C9293 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n9 VSS 0.055518f
C9294 MULT_0.4bit_ADDER_0.FULL_ADDER_2.COUT.n10 VSS 0.369194f
C9295 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t22 VSS 0.013766f
C9296 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t15 VSS 0.027698f
C9297 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t19 VSS 0.027354f
C9298 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t17 VSS 0.027354f
C9299 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t14 VSS 0.027354f
C9300 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t23 VSS 0.005684f
C9301 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t21 VSS 0.005684f
C9302 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t20 VSS 0.005684f
C9303 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n0 VSS 0.168523f
C9304 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n1 VSS 0.124125f
C9305 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n2 VSS 0.067647f
C9306 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n3 VSS 0.066457f
C9307 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n4 VSS 0.040879f
C9308 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n5 VSS 0.05311f
C9309 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t18 VSS 0.030151f
C9310 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t13 VSS 0.009818f
C9311 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t12 VSS 0.013559f
C9312 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n6 VSS 0.014622f
C9313 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t16 VSS 0.010094f
C9314 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n7 VSS 0.025612f
C9315 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n8 VSS 0.044927f
C9316 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t10 VSS 0.004926f
C9317 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t9 VSS 0.004926f
C9318 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n9 VSS 0.011915f
C9319 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t4 VSS 0.004926f
C9320 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t5 VSS 0.004926f
C9321 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n10 VSS 0.011914f
C9322 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n11 VSS 0.085433f
C9323 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t8 VSS 0.004926f
C9324 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t3 VSS 0.004926f
C9325 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n12 VSS 0.009853f
C9326 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n13 VSS 0.00774f
C9327 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t1 VSS 0.020843f
C9328 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t6 VSS 0.020843f
C9329 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n14 VSS 0.041685f
C9330 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n15 VSS 0.016575f
C9331 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t0 VSS 0.020843f
C9332 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t2 VSS 0.020843f
C9333 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n16 VSS 0.041685f
C9334 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n17 VSS 0.018334f
C9335 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n18 VSS 0.188757f
C9336 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t7 VSS 0.020843f
C9337 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.t11 VSS 0.020843f
C9338 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n19 VSS 0.041685f
C9339 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n20 VSS 0.018362f
C9340 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n21 VSS 0.12106f
C9341 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n22 VSS 0.027282f
C9342 MULT_0.4bit_ADDER_1.FULL_ADDER_1.XOR2_1.A.n23 VSS 0.119748f
C9343 a_n17266_n7799.n0 VSS 1.48365f
C9344 a_n17266_n7799.n1 VSS 1.48326f
C9345 a_n17266_n7799.t5 VSS 0.093341f
C9346 a_n17266_n7799.t11 VSS 0.093341f
C9347 a_n17266_n7799.t10 VSS 0.093341f
C9348 a_n17266_n7799.n2 VSS 0.202296f
C9349 a_n17266_n7799.t9 VSS 0.093341f
C9350 a_n17266_n7799.t0 VSS 0.093341f
C9351 a_n17266_n7799.n3 VSS 0.202001f
C9352 a_n17266_n7799.t2 VSS 0.093341f
C9353 a_n17266_n7799.t1 VSS 0.093341f
C9354 a_n17266_n7799.n4 VSS 0.202001f
C9355 a_n17266_n7799.t3 VSS 0.093341f
C9356 a_n17266_n7799.t4 VSS 0.093341f
C9357 a_n17266_n7799.n5 VSS 0.202001f
C9358 a_n17266_n7799.t8 VSS 0.093341f
C9359 a_n17266_n7799.t6 VSS 0.093341f
C9360 a_n17266_n7799.n6 VSS 0.202001f
C9361 a_n17266_n7799.n7 VSS 0.20269f
C9362 a_n17266_n7799.t7 VSS 0.093341f
C9363 8bit_ADDER_0.S2.t14 VSS 0.052755f
C9364 8bit_ADDER_0.S2.t13 VSS 0.051327f
C9365 8bit_ADDER_0.S2.t12 VSS 0.155431f
C9366 8bit_ADDER_0.S2.n0 VSS 0.264627f
C9367 8bit_ADDER_0.S2.t6 VSS 0.015363f
C9368 8bit_ADDER_0.S2.t5 VSS 0.015363f
C9369 8bit_ADDER_0.S2.n1 VSS 0.037156f
C9370 8bit_ADDER_0.S2.t0 VSS 0.015363f
C9371 8bit_ADDER_0.S2.t9 VSS 0.015363f
C9372 8bit_ADDER_0.S2.n2 VSS 0.037152f
C9373 8bit_ADDER_0.S2.n3 VSS 0.266414f
C9374 8bit_ADDER_0.S2.t4 VSS 0.015363f
C9375 8bit_ADDER_0.S2.t11 VSS 0.015363f
C9376 8bit_ADDER_0.S2.n4 VSS 0.030725f
C9377 8bit_ADDER_0.S2.n5 VSS 0.024136f
C9378 8bit_ADDER_0.S2.t1 VSS 0.064996f
C9379 8bit_ADDER_0.S2.t8 VSS 0.064996f
C9380 8bit_ADDER_0.S2.n6 VSS 0.129991f
C9381 8bit_ADDER_0.S2.n7 VSS 0.051686f
C9382 8bit_ADDER_0.S2.t2 VSS 0.064996f
C9383 8bit_ADDER_0.S2.t3 VSS 0.064996f
C9384 8bit_ADDER_0.S2.n8 VSS 0.129991f
C9385 8bit_ADDER_0.S2.n9 VSS 0.057172f
C9386 8bit_ADDER_0.S2.n10 VSS 0.588621f
C9387 8bit_ADDER_0.S2.t10 VSS 0.064996f
C9388 8bit_ADDER_0.S2.t7 VSS 0.064996f
C9389 8bit_ADDER_0.S2.n11 VSS 0.129991f
C9390 8bit_ADDER_0.S2.n12 VSS 0.057259f
C9391 8bit_ADDER_0.S2.n13 VSS 0.377516f
C9392 8bit_ADDER_0.S2.n14 VSS 0.085077f
C9393 8bit_ADDER_0.S2.n15 VSS 0.373423f
C9394 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t14 VSS 0.013766f
C9395 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t20 VSS 0.027698f
C9396 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t13 VSS 0.027354f
C9397 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t15 VSS 0.027354f
C9398 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t17 VSS 0.027354f
C9399 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t18 VSS 0.005684f
C9400 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t12 VSS 0.005684f
C9401 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t16 VSS 0.005684f
C9402 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n0 VSS 0.168523f
C9403 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n1 VSS 0.124125f
C9404 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n2 VSS 0.067647f
C9405 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n3 VSS 0.066457f
C9406 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n4 VSS 0.040879f
C9407 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n5 VSS 0.05311f
C9408 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t19 VSS 0.030151f
C9409 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t22 VSS 0.009818f
C9410 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t23 VSS 0.013559f
C9411 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n6 VSS 0.014622f
C9412 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t21 VSS 0.010094f
C9413 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n7 VSS 0.025612f
C9414 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n8 VSS 0.044927f
C9415 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t6 VSS 0.004926f
C9416 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t5 VSS 0.004926f
C9417 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n9 VSS 0.011915f
C9418 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t11 VSS 0.004926f
C9419 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t10 VSS 0.004926f
C9420 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n10 VSS 0.011914f
C9421 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n11 VSS 0.085433f
C9422 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t7 VSS 0.004926f
C9423 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t1 VSS 0.004926f
C9424 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n12 VSS 0.009853f
C9425 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n13 VSS 0.00774f
C9426 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t4 VSS 0.020843f
C9427 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t9 VSS 0.020843f
C9428 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n14 VSS 0.041685f
C9429 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n15 VSS 0.016575f
C9430 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t3 VSS 0.020843f
C9431 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t2 VSS 0.020843f
C9432 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n16 VSS 0.041685f
C9433 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n17 VSS 0.018334f
C9434 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n18 VSS 0.188757f
C9435 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t8 VSS 0.020843f
C9436 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.t0 VSS 0.020843f
C9437 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n19 VSS 0.041685f
C9438 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n20 VSS 0.018362f
C9439 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n21 VSS 0.12106f
C9440 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n22 VSS 0.027282f
C9441 8bit_ADDER_0.FULL_ADDER_XORED_5.XOR2_1.A.n23 VSS 0.119748f
C9442 mux8_6.A0.t20 VSS 0.036758f
C9443 mux8_6.A0.t14 VSS 0.035764f
C9444 mux8_6.A0.t13 VSS 0.108301f
C9445 mux8_6.A0.n0 VSS 0.184386f
C9446 mux8_6.A0.t15 VSS 0.060184f
C9447 mux8_6.A0.t22 VSS 0.059435f
C9448 mux8_6.A0.t17 VSS 0.059435f
C9449 mux8_6.A0.t19 VSS 0.059435f
C9450 mux8_6.A0.n1 VSS 0.236568f
C9451 mux8_6.A0.t12 VSS 0.012351f
C9452 mux8_6.A0.t16 VSS 0.012351f
C9453 mux8_6.A0.t21 VSS 0.012351f
C9454 mux8_6.A0.t18 VSS 0.012351f
C9455 mux8_6.A0.n2 VSS 0.223488f
C9456 mux8_6.A0.n3 VSS 0.349758f
C9457 mux8_6.A0.n4 VSS 1.81464f
C9458 mux8_6.A0.n5 VSS 13.1639f
C9459 mux8_6.A0.t1 VSS 0.010704f
C9460 mux8_6.A0.t2 VSS 0.010704f
C9461 mux8_6.A0.n6 VSS 0.02589f
C9462 mux8_6.A0.t6 VSS 0.010704f
C9463 mux8_6.A0.t7 VSS 0.010704f
C9464 mux8_6.A0.n7 VSS 0.025887f
C9465 mux8_6.A0.n8 VSS 0.185631f
C9466 mux8_6.A0.t0 VSS 0.010704f
C9467 mux8_6.A0.t11 VSS 0.010704f
C9468 mux8_6.A0.n9 VSS 0.021409f
C9469 mux8_6.A0.n10 VSS 0.016817f
C9470 mux8_6.A0.t5 VSS 0.045288f
C9471 mux8_6.A0.t10 VSS 0.045288f
C9472 mux8_6.A0.n11 VSS 0.090575f
C9473 mux8_6.A0.n12 VSS 0.036014f
C9474 mux8_6.A0.t4 VSS 0.045288f
C9475 mux8_6.A0.t3 VSS 0.045288f
C9476 mux8_6.A0.n13 VSS 0.090575f
C9477 mux8_6.A0.n14 VSS 0.039836f
C9478 mux8_6.A0.n15 VSS 0.410138f
C9479 mux8_6.A0.t8 VSS 0.045288f
C9480 mux8_6.A0.t9 VSS 0.045288f
C9481 mux8_6.A0.n16 VSS 0.090575f
C9482 mux8_6.A0.n17 VSS 0.039897f
C9483 mux8_6.A0.n18 VSS 0.263045f
C9484 mux8_6.A0.n19 VSS 0.05928f
C9485 mux8_6.A0.n20 VSS 0.260193f
C9486 mux8_3.NAND4F_9.Y.n0 VSS 0.358256f
C9487 mux8_3.NAND4F_9.Y.t13 VSS 0.017853f
C9488 mux8_3.NAND4F_9.Y.t12 VSS 0.017853f
C9489 mux8_3.NAND4F_9.Y.t11 VSS 0.017853f
C9490 mux8_3.NAND4F_9.Y.t10 VSS 0.017853f
C9491 mux8_3.NAND4F_9.Y.t9 VSS 0.022554f
C9492 mux8_3.NAND4F_9.Y.n1 VSS 0.048188f
C9493 mux8_3.NAND4F_9.Y.n2 VSS 0.030339f
C9494 mux8_3.NAND4F_9.Y.n3 VSS 0.030339f
C9495 mux8_3.NAND4F_9.Y.n4 VSS 0.026149f
C9496 mux8_3.NAND4F_9.Y.t14 VSS 0.014813f
C9497 mux8_3.NAND4F_9.Y.n5 VSS 0.021261f
C9498 mux8_3.NAND4F_9.Y.t2 VSS 0.141821f
C9499 mux8_3.NAND4F_9.Y.t6 VSS 0.017663f
C9500 mux8_3.NAND4F_9.Y.t5 VSS 0.017663f
C9501 mux8_3.NAND4F_9.Y.n6 VSS 0.041015f
C9502 mux8_3.NAND4F_9.Y.t7 VSS 0.017663f
C9503 mux8_3.NAND4F_9.Y.t8 VSS 0.017663f
C9504 mux8_3.NAND4F_9.Y.n7 VSS 0.040893f
C9505 mux8_3.NAND4F_9.Y.t3 VSS 0.017663f
C9506 mux8_3.NAND4F_9.Y.t4 VSS 0.017663f
C9507 mux8_3.NAND4F_9.Y.n8 VSS 0.040893f
C9508 mux8_3.NAND4F_9.Y.t0 VSS 0.017663f
C9509 mux8_3.NAND4F_9.Y.t1 VSS 0.017663f
C9510 mux8_3.NAND4F_9.Y.n9 VSS 0.040893f
C9511 mux8_3.NAND4F_9.Y.n10 VSS 0.168091f
C9512 mux8_3.NAND4F_7.Y.n0 VSS 0.11858f
C9513 mux8_3.NAND4F_7.Y.n1 VSS 0.350455f
C9514 mux8_3.NAND4F_7.Y.t3 VSS 0.168166f
C9515 mux8_3.NAND4F_7.Y.t11 VSS 0.022537f
C9516 mux8_3.NAND4F_7.Y.t10 VSS 0.079785f
C9517 mux8_3.NAND4F_7.Y.t9 VSS 0.024808f
C9518 mux8_3.NAND4F_7.Y.n2 VSS 0.070768f
C9519 mux8_3.NAND4F_7.Y.n3 VSS 0.020978f
C9520 mux8_3.NAND4F_7.Y.t1 VSS 0.017278f
C9521 mux8_3.NAND4F_7.Y.t0 VSS 0.017278f
C9522 mux8_3.NAND4F_7.Y.n4 VSS 0.040122f
C9523 mux8_3.NAND4F_7.Y.t5 VSS 0.017278f
C9524 mux8_3.NAND4F_7.Y.t6 VSS 0.017278f
C9525 mux8_3.NAND4F_7.Y.n5 VSS 0.040002f
C9526 mux8_3.NAND4F_7.Y.t8 VSS 0.017278f
C9527 mux8_3.NAND4F_7.Y.t7 VSS 0.017278f
C9528 mux8_3.NAND4F_7.Y.n6 VSS 0.040002f
C9529 mux8_3.NAND4F_7.Y.t4 VSS 0.017278f
C9530 mux8_3.NAND4F_7.Y.t2 VSS 0.017278f
C9531 mux8_3.NAND4F_7.Y.n7 VSS 0.040002f
C9532 a_n12416_n4534.n0 VSS 1.48326f
C9533 a_n12416_n4534.n1 VSS 1.48365f
C9534 a_n12416_n4534.t2 VSS 0.093341f
C9535 a_n12416_n4534.t6 VSS 0.093341f
C9536 a_n12416_n4534.t8 VSS 0.093341f
C9537 a_n12416_n4534.n2 VSS 0.20269f
C9538 a_n12416_n4534.t0 VSS 0.093341f
C9539 a_n12416_n4534.t7 VSS 0.093341f
C9540 a_n12416_n4534.n3 VSS 0.202001f
C9541 a_n12416_n4534.t5 VSS 0.093341f
C9542 a_n12416_n4534.t4 VSS 0.093341f
C9543 a_n12416_n4534.n4 VSS 0.202001f
C9544 a_n12416_n4534.t10 VSS 0.093341f
C9545 a_n12416_n4534.t11 VSS 0.093341f
C9546 a_n12416_n4534.n5 VSS 0.202001f
C9547 a_n12416_n4534.t1 VSS 0.093341f
C9548 a_n12416_n4534.t9 VSS 0.093341f
C9549 a_n12416_n4534.n6 VSS 0.202001f
C9550 a_n12416_n4534.n7 VSS 0.202296f
C9551 a_n12416_n4534.t3 VSS 0.093341f
C9552 MULT_0.4bit_ADDER_2.FULL_ADDER_1.XOR2_0.B VSS 0.752862f
C9553 MULT_0.4bit_ADDER_2.A2 VSS 1.05688f
C9554 MULT_0.inv_14.Y.n0 VSS 2.79153f
C9555 MULT_0.inv_14.Y.t3 VSS 0.065961f
C9556 MULT_0.inv_14.Y.t2 VSS 0.018184f
C9557 MULT_0.inv_14.Y.t1 VSS 0.018184f
C9558 MULT_0.inv_14.Y.n1 VSS 0.040543f
C9559 MULT_0.inv_14.Y.t0 VSS 0.052505f
C9560 MULT_0.inv_14.Y.t14 VSS 0.057355f
C9561 MULT_0.inv_14.Y.t8 VSS 0.022015f
C9562 MULT_0.inv_14.Y.t10 VSS 0.030403f
C9563 MULT_0.inv_14.Y.n2 VSS 0.034993f
C9564 MULT_0.inv_14.Y.t4 VSS 0.023141f
C9565 MULT_0.inv_14.Y.n3 VSS 0.035488f
C9566 MULT_0.inv_14.Y.n4 VSS 0.146894f
C9567 MULT_0.4bit_ADDER_2.FULL_ADDER_1.NAND2_0.B VSS 0.567559f
C9568 MULT_0.inv_14.Y.t5 VSS 0.062107f
C9569 MULT_0.inv_14.Y.t12 VSS 0.061334f
C9570 MULT_0.inv_14.Y.t11 VSS 0.061334f
C9571 MULT_0.inv_14.Y.t13 VSS 0.061334f
C9572 MULT_0.inv_14.Y.n5 VSS 0.244128f
C9573 MULT_0.inv_14.Y.t6 VSS 0.012746f
C9574 MULT_0.inv_14.Y.t9 VSS 0.012746f
C9575 MULT_0.inv_14.Y.t15 VSS 0.012746f
C9576 MULT_0.inv_14.Y.t7 VSS 0.012746f
C9577 MULT_0.inv_14.Y.n6 VSS 0.23063f
C9578 MULT_0.inv_14.Y.n7 VSS 0.360752f
C9579 MULT_0.inv_14.Y.n8 VSS 0.852904f
C9580 MULT_0.4bit_ADDER_1.FULL_ADDER_3.NAND2_0.B VSS 0.687724f
C9581 MULT_0.4bit_ADDER_1.A0.n0 VSS 4.14855f
C9582 MULT_0.4bit_ADDER_1.FULL_ADDER_3.XOR2_0.B VSS 0.724697f
C9583 MULT_0.4bit_ADDER_1.FULL_ADDER_3.A VSS 2.94359f
C9584 MULT_0.4bit_ADDER_1.A0.t5 VSS 0.055209f
C9585 MULT_0.4bit_ADDER_1.A0.t11 VSS 0.021192f
C9586 MULT_0.4bit_ADDER_1.A0.t10 VSS 0.029265f
C9587 MULT_0.4bit_ADDER_1.A0.n1 VSS 0.033684f
C9588 MULT_0.4bit_ADDER_1.A0.t4 VSS 0.022275f
C9589 MULT_0.4bit_ADDER_1.A0.n2 VSS 0.03416f
C9590 MULT_0.4bit_ADDER_1.A0.t6 VSS 0.059783f
C9591 MULT_0.4bit_ADDER_1.A0.t15 VSS 0.05904f
C9592 MULT_0.4bit_ADDER_1.A0.t7 VSS 0.05904f
C9593 MULT_0.4bit_ADDER_1.A0.t13 VSS 0.05904f
C9594 MULT_0.4bit_ADDER_1.A0.n3 VSS 0.234994f
C9595 MULT_0.4bit_ADDER_1.A0.t14 VSS 0.012269f
C9596 MULT_0.4bit_ADDER_1.A0.t8 VSS 0.012269f
C9597 MULT_0.4bit_ADDER_1.A0.t12 VSS 0.012269f
C9598 MULT_0.4bit_ADDER_1.A0.t9 VSS 0.012269f
C9599 MULT_0.4bit_ADDER_1.A0.n4 VSS 0.222002f
C9600 MULT_0.4bit_ADDER_1.A0.n5 VSS 0.347255f
C9601 MULT_0.4bit_ADDER_1.A0.n6 VSS 0.821319f
C9602 MULT_0.4bit_ADDER_1.A0.t1 VSS 0.017504f
C9603 MULT_0.4bit_ADDER_1.A0.t2 VSS 0.017504f
C9604 MULT_0.4bit_ADDER_1.A0.n7 VSS 0.038899f
C9605 MULT_0.4bit_ADDER_1.A0.t0 VSS 0.050712f
C9606 MULT_0.4bit_ADDER_1.A0.t3 VSS 0.063486f
C9607 mux8_7.NAND4F_3.Y.n0 VSS 0.306333f
C9608 mux8_7.NAND4F_3.Y.t7 VSS 0.015103f
C9609 mux8_7.NAND4F_3.Y.t8 VSS 0.015103f
C9610 mux8_7.NAND4F_3.Y.n1 VSS 0.035071f
C9611 mux8_7.NAND4F_3.Y.t0 VSS 0.015103f
C9612 mux8_7.NAND4F_3.Y.t1 VSS 0.015103f
C9613 mux8_7.NAND4F_3.Y.n2 VSS 0.034966f
C9614 mux8_7.NAND4F_3.Y.t6 VSS 0.015103f
C9615 mux8_7.NAND4F_3.Y.t5 VSS 0.015103f
C9616 mux8_7.NAND4F_3.Y.n3 VSS 0.034966f
C9617 mux8_7.NAND4F_3.Y.t4 VSS 0.015103f
C9618 mux8_7.NAND4F_3.Y.t3 VSS 0.015103f
C9619 mux8_7.NAND4F_3.Y.n4 VSS 0.034966f
C9620 mux8_7.NAND4F_3.Y.n5 VSS 0.152246f
C9621 mux8_7.NAND4F_3.Y.t2 VSS 0.143521f
C9622 mux8_7.NAND4F_3.Y.t10 VSS 0.0197f
C9623 mux8_7.NAND4F_3.Y.t11 VSS 0.0197f
C9624 mux8_7.NAND4F_3.Y.n6 VSS 0.023128f
C9625 mux8_7.NAND4F_3.Y.t9 VSS 0.061756f
C9626 mux8_7.NAND4F_3.Y.n7 VSS 0.129679f
C9627 mux8_7.A0.t12 VSS 0.067168f
C9628 mux8_7.A0.t14 VSS 0.06535f
C9629 mux8_7.A0.t13 VSS 0.197897f
C9630 mux8_7.A0.n0 VSS 0.336925f
C9631 mux8_7.A0.t9 VSS 0.01956f
C9632 mux8_7.A0.t11 VSS 0.01956f
C9633 mux8_7.A0.n1 VSS 0.047308f
C9634 mux8_7.A0.t4 VSS 0.01956f
C9635 mux8_7.A0.t2 VSS 0.01956f
C9636 mux8_7.A0.n2 VSS 0.047302f
C9637 mux8_7.A0.n3 VSS 0.3392f
C9638 mux8_7.A0.t10 VSS 0.01956f
C9639 mux8_7.A0.t1 VSS 0.01956f
C9640 mux8_7.A0.n4 VSS 0.03912f
C9641 mux8_7.A0.n5 VSS 0.03073f
C9642 mux8_7.A0.t7 VSS 0.082753f
C9643 mux8_7.A0.t3 VSS 0.082753f
C9644 mux8_7.A0.n6 VSS 0.165506f
C9645 mux8_7.A0.n7 VSS 0.065808f
C9646 mux8_7.A0.t6 VSS 0.082753f
C9647 mux8_7.A0.t8 VSS 0.082753f
C9648 mux8_7.A0.n8 VSS 0.165506f
C9649 mux8_7.A0.n9 VSS 0.072792f
C9650 mux8_7.A0.n10 VSS 0.749438f
C9651 mux8_7.A0.t0 VSS 0.082753f
C9652 mux8_7.A0.t5 VSS 0.082753f
C9653 mux8_7.A0.n11 VSS 0.165506f
C9654 mux8_7.A0.n12 VSS 0.072903f
C9655 mux8_7.A0.n13 VSS 0.480657f
C9656 mux8_7.A0.n14 VSS 0.108322f
C9657 mux8_7.A0.n15 VSS 0.475445f
C9658 MULT_0.4bit_ADDER_1.B3.n0 VSS 1.29534f
C9659 MULT_0.4bit_ADDER_1.B3.t13 VSS 0.04169f
C9660 MULT_0.4bit_ADDER_1.B3.t7 VSS 0.013576f
C9661 MULT_0.4bit_ADDER_1.B3.t18 VSS 0.018748f
C9662 MULT_0.4bit_ADDER_1.B3.n1 VSS 0.020218f
C9663 MULT_0.4bit_ADDER_1.B3.t12 VSS 0.013957f
C9664 MULT_0.4bit_ADDER_1.B3.n2 VSS 0.035415f
C9665 MULT_0.4bit_ADDER_1.B3.n3 VSS 0.062124f
C9666 MULT_0.4bit_ADDER_1.B3.t11 VSS 0.019035f
C9667 MULT_0.4bit_ADDER_1.B3.t16 VSS 0.038299f
C9668 MULT_0.4bit_ADDER_1.B3.t9 VSS 0.037822f
C9669 MULT_0.4bit_ADDER_1.B3.t17 VSS 0.037822f
C9670 MULT_0.4bit_ADDER_1.B3.t15 VSS 0.037822f
C9671 MULT_0.4bit_ADDER_1.B3.t14 VSS 0.00786f
C9672 MULT_0.4bit_ADDER_1.B3.t8 VSS 0.00786f
C9673 MULT_0.4bit_ADDER_1.B3.t10 VSS 0.00786f
C9674 MULT_0.4bit_ADDER_1.B3.n4 VSS 0.233019f
C9675 MULT_0.4bit_ADDER_1.B3.n5 VSS 0.171629f
C9676 MULT_0.4bit_ADDER_1.B3.n6 VSS 0.093536f
C9677 MULT_0.4bit_ADDER_1.B3.n7 VSS 0.091891f
C9678 MULT_0.4bit_ADDER_1.B3.n8 VSS 0.056524f
C9679 MULT_0.4bit_ADDER_1.B3.n9 VSS 0.074149f
C9680 MULT_0.4bit_ADDER_1.B3.n10 VSS 0.820717f
C9681 MULT_0.4bit_ADDER_1.B3.t2 VSS 0.011213f
C9682 MULT_0.4bit_ADDER_1.B3.t1 VSS 0.011213f
C9683 MULT_0.4bit_ADDER_1.B3.n11 VSS 0.024951f
C9684 MULT_0.4bit_ADDER_1.B3.t5 VSS 0.011213f
C9685 MULT_0.4bit_ADDER_1.B3.t4 VSS 0.011213f
C9686 MULT_0.4bit_ADDER_1.B3.n12 VSS 0.025019f
C9687 MULT_0.4bit_ADDER_1.B3.t0 VSS 0.011213f
C9688 MULT_0.4bit_ADDER_1.B3.t6 VSS 0.011213f
C9689 MULT_0.4bit_ADDER_1.B3.n13 VSS 0.024951f
C9690 MULT_0.4bit_ADDER_1.B3.t3 VSS 0.067706f
C9691 mux8_8.A1.t12 VSS 0.045589f
C9692 mux8_8.A1.t13 VSS 0.044355f
C9693 mux8_8.A1.t14 VSS 0.134319f
C9694 mux8_8.A1.n0 VSS 0.228683f
C9695 mux8_8.A1.t5 VSS 0.013276f
C9696 mux8_8.A1.t6 VSS 0.013276f
C9697 mux8_8.A1.n1 VSS 0.032109f
C9698 mux8_8.A1.t11 VSS 0.013276f
C9699 mux8_8.A1.t3 VSS 0.013276f
C9700 mux8_8.A1.n2 VSS 0.032106f
C9701 mux8_8.A1.n3 VSS 0.230227f
C9702 mux8_8.A1.t4 VSS 0.013276f
C9703 mux8_8.A1.t0 VSS 0.013276f
C9704 mux8_8.A1.n4 VSS 0.026552f
C9705 mux8_8.A1.n5 VSS 0.020857f
C9706 mux8_8.A1.t8 VSS 0.056167f
C9707 mux8_8.A1.t2 VSS 0.056167f
C9708 mux8_8.A1.n6 VSS 0.112335f
C9709 mux8_8.A1.n7 VSS 0.044666f
C9710 mux8_8.A1.t9 VSS 0.056167f
C9711 mux8_8.A1.t7 VSS 0.056167f
C9712 mux8_8.A1.n8 VSS 0.112335f
C9713 mux8_8.A1.n9 VSS 0.049407f
C9714 mux8_8.A1.n10 VSS 0.50867f
C9715 mux8_8.A1.t1 VSS 0.056167f
C9716 mux8_8.A1.t10 VSS 0.056167f
C9717 mux8_8.A1.n11 VSS 0.112335f
C9718 mux8_8.A1.n12 VSS 0.049481f
C9719 mux8_8.A1.n13 VSS 0.326239f
C9720 mux8_8.A1.n14 VSS 0.073522f
C9721 mux8_8.A1.n15 VSS 0.322701f
C9722 mux8_8.NAND4F_9.Y.n0 VSS 0.358256f
C9723 mux8_8.NAND4F_9.Y.t14 VSS 0.017853f
C9724 mux8_8.NAND4F_9.Y.t13 VSS 0.017853f
C9725 mux8_8.NAND4F_9.Y.t11 VSS 0.017853f
C9726 mux8_8.NAND4F_9.Y.t10 VSS 0.017853f
C9727 mux8_8.NAND4F_9.Y.t9 VSS 0.022554f
C9728 mux8_8.NAND4F_9.Y.n1 VSS 0.048188f
C9729 mux8_8.NAND4F_9.Y.n2 VSS 0.030339f
C9730 mux8_8.NAND4F_9.Y.n3 VSS 0.030339f
C9731 mux8_8.NAND4F_9.Y.n4 VSS 0.026149f
C9732 mux8_8.NAND4F_9.Y.t12 VSS 0.014813f
C9733 mux8_8.NAND4F_9.Y.n5 VSS 0.021261f
C9734 mux8_8.NAND4F_9.Y.t0 VSS 0.141821f
C9735 mux8_8.NAND4F_9.Y.t7 VSS 0.017663f
C9736 mux8_8.NAND4F_9.Y.t8 VSS 0.017663f
C9737 mux8_8.NAND4F_9.Y.n6 VSS 0.041015f
C9738 mux8_8.NAND4F_9.Y.t5 VSS 0.017663f
C9739 mux8_8.NAND4F_9.Y.t6 VSS 0.017663f
C9740 mux8_8.NAND4F_9.Y.n7 VSS 0.040893f
C9741 mux8_8.NAND4F_9.Y.t3 VSS 0.017663f
C9742 mux8_8.NAND4F_9.Y.t4 VSS 0.017663f
C9743 mux8_8.NAND4F_9.Y.n8 VSS 0.040893f
C9744 mux8_8.NAND4F_9.Y.t2 VSS 0.017663f
C9745 mux8_8.NAND4F_9.Y.t1 VSS 0.017663f
C9746 mux8_8.NAND4F_9.Y.n9 VSS 0.040893f
C9747 mux8_8.NAND4F_9.Y.n10 VSS 0.168091f
C9748 Y1.t7 VSS 0.091566f
C9749 Y1.t5 VSS 0.196577f
C9750 Y1.t4 VSS 0.212396f
C9751 Y1.n0 VSS 0.167788f
C9752 Y1.t6 VSS 0.197703f
C9753 Y1.n1 VSS 0.095069f
C9754 Y1.n2 VSS 0.099249f
C9755 Y1.t2 VSS 0.036784f
C9756 Y1.t3 VSS 0.036784f
C9757 Y1.n3 VSS 0.081952f
C9758 Y1.t1 VSS 0.106275f
C9759 Y1.t0 VSS 0.133415f
C9760 Y1.n4 VSS 0.553327f
C9761 Y1.n5 VSS 0.707877f
C9762 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n0 VSS 0.860468f
C9763 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t5 VSS 0.007445f
C9764 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t4 VSS 0.007445f
C9765 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n1 VSS 0.016612f
C9766 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t1 VSS 0.007445f
C9767 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t6 VSS 0.007445f
C9768 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n2 VSS 0.016567f
C9769 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t3 VSS 0.007445f
C9770 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t2 VSS 0.007445f
C9771 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n3 VSS 0.016567f
C9772 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t0 VSS 0.044954f
C9773 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t8 VSS 0.025429f
C9774 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t12 VSS 0.025112f
C9775 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t11 VSS 0.025112f
C9776 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t16 VSS 0.025112f
C9777 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n4 VSS 0.099955f
C9778 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t18 VSS 0.005219f
C9779 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t10 VSS 0.005219f
C9780 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t17 VSS 0.005219f
C9781 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t7 VSS 0.005219f
C9782 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n5 VSS 0.094428f
C9783 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n6 VSS 0.14768f
C9784 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t9 VSS 0.023483f
C9785 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t15 VSS 0.009014f
C9786 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t13 VSS 0.012448f
C9787 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n7 VSS 0.014328f
C9788 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.t14 VSS 0.009475f
C9789 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n8 VSS 0.01453f
C9790 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n9 VSS 0.049352f
C9791 8bit_ADDER_0.FULL_ADDER_XORED_5.COUT.n10 VSS 0.328192f
C9792 mux8_0.NAND4F_2.Y.n0 VSS 0.530078f
C9793 mux8_0.NAND4F_2.Y.t5 VSS 0.026135f
C9794 mux8_0.NAND4F_2.Y.t6 VSS 0.026135f
C9795 mux8_0.NAND4F_2.Y.n1 VSS 0.060687f
C9796 mux8_0.NAND4F_2.Y.t4 VSS 0.026135f
C9797 mux8_0.NAND4F_2.Y.t3 VSS 0.026135f
C9798 mux8_0.NAND4F_2.Y.n2 VSS 0.060505f
C9799 mux8_0.NAND4F_2.Y.t8 VSS 0.026135f
C9800 mux8_0.NAND4F_2.Y.t7 VSS 0.026135f
C9801 mux8_0.NAND4F_2.Y.n3 VSS 0.060505f
C9802 mux8_0.NAND4F_2.Y.t1 VSS 0.026135f
C9803 mux8_0.NAND4F_2.Y.t2 VSS 0.026135f
C9804 mux8_0.NAND4F_2.Y.n4 VSS 0.060505f
C9805 mux8_0.NAND4F_2.Y.n5 VSS 0.263447f
C9806 mux8_0.NAND4F_2.Y.t0 VSS 0.213114f
C9807 mux8_0.NAND4F_2.Y.t9 VSS 0.034088f
C9808 mux8_0.NAND4F_2.Y.t10 VSS 0.105185f
C9809 mux8_0.NAND4F_2.Y.t11 VSS 0.039267f
C9810 mux8_0.NAND4F_2.Y.n6 VSS 0.131989f
C9811 mux8_0.NAND4F_2.Y.n7 VSS 0.028742f
C9812 mux8_0.NAND4F_2.Y.n8 VSS 1.53344f
C9813 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n0 VSS 0.887305f
C9814 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t1 VSS 0.007677f
C9815 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t2 VSS 0.007677f
C9816 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n1 VSS 0.017083f
C9817 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t6 VSS 0.007677f
C9818 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t4 VSS 0.007677f
C9819 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n2 VSS 0.01713f
C9820 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t3 VSS 0.007677f
C9821 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t5 VSS 0.007677f
C9822 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n3 VSS 0.017083f
C9823 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t0 VSS 0.046356f
C9824 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t8 VSS 0.026222f
C9825 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t15 VSS 0.025896f
C9826 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t14 VSS 0.025896f
C9827 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t7 VSS 0.025896f
C9828 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n4 VSS 0.103072f
C9829 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t12 VSS 0.005381f
C9830 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t16 VSS 0.005381f
C9831 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t18 VSS 0.005381f
C9832 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t13 VSS 0.005381f
C9833 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n5 VSS 0.097373f
C9834 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n6 VSS 0.152286f
C9835 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t10 VSS 0.024216f
C9836 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t9 VSS 0.009295f
C9837 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t11 VSS 0.012836f
C9838 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n7 VSS 0.014774f
C9839 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.t17 VSS 0.00977f
C9840 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n8 VSS 0.014983f
C9841 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n9 VSS 0.050891f
C9842 MULT_0.4bit_ADDER_2.FULL_ADDER_2.COUT.n10 VSS 0.338427f
C9843 mux8_5.NAND4F_0.Y.n0 VSS 0.350455f
C9844 mux8_5.NAND4F_0.Y.t9 VSS 0.022537f
C9845 mux8_5.NAND4F_0.Y.t11 VSS 0.079785f
C9846 mux8_5.NAND4F_0.Y.t10 VSS 0.024808f
C9847 mux8_5.NAND4F_0.Y.n1 VSS 0.070768f
C9848 mux8_5.NAND4F_0.Y.n2 VSS 0.020978f
C9849 mux8_5.NAND4F_0.Y.t5 VSS 0.017278f
C9850 mux8_5.NAND4F_0.Y.t6 VSS 0.017278f
C9851 mux8_5.NAND4F_0.Y.n3 VSS 0.040122f
C9852 mux8_5.NAND4F_0.Y.t1 VSS 0.017278f
C9853 mux8_5.NAND4F_0.Y.t0 VSS 0.017278f
C9854 mux8_5.NAND4F_0.Y.n4 VSS 0.040002f
C9855 mux8_5.NAND4F_0.Y.t8 VSS 0.017278f
C9856 mux8_5.NAND4F_0.Y.t7 VSS 0.017278f
C9857 mux8_5.NAND4F_0.Y.n5 VSS 0.040002f
C9858 mux8_5.NAND4F_0.Y.t2 VSS 0.017278f
C9859 mux8_5.NAND4F_0.Y.t3 VSS 0.017278f
C9860 mux8_5.NAND4F_0.Y.n6 VSS 0.040002f
C9861 mux8_5.NAND4F_0.Y.t4 VSS 0.166327f
C9862 mux8_5.A1.t14 VSS 0.057075f
C9863 mux8_5.A1.t12 VSS 0.05553f
C9864 mux8_5.A1.t13 VSS 0.168161f
C9865 mux8_5.A1.n0 VSS 0.286299f
C9866 mux8_5.A1.t3 VSS 0.016621f
C9867 mux8_5.A1.t4 VSS 0.016621f
C9868 mux8_5.A1.n1 VSS 0.040199f
C9869 mux8_5.A1.t10 VSS 0.016621f
C9870 mux8_5.A1.t6 VSS 0.016621f
C9871 mux8_5.A1.n2 VSS 0.040195f
C9872 mux8_5.A1.n3 VSS 0.288232f
C9873 mux8_5.A1.t5 VSS 0.016621f
C9874 mux8_5.A1.t7 VSS 0.016621f
C9875 mux8_5.A1.n4 VSS 0.033241f
C9876 mux8_5.A1.n5 VSS 0.026112f
C9877 mux8_5.A1.t2 VSS 0.070318f
C9878 mux8_5.A1.t9 VSS 0.070318f
C9879 mux8_5.A1.n6 VSS 0.140637f
C9880 mux8_5.A1.n7 VSS 0.05592f
C9881 mux8_5.A1.t0 VSS 0.070318f
C9882 mux8_5.A1.t1 VSS 0.070318f
C9883 mux8_5.A1.n8 VSS 0.140637f
C9884 mux8_5.A1.n9 VSS 0.061855f
C9885 mux8_5.A1.n10 VSS 0.636828f
C9886 mux8_5.A1.t11 VSS 0.070318f
C9887 mux8_5.A1.t8 VSS 0.070318f
C9888 mux8_5.A1.n11 VSS 0.140637f
C9889 mux8_5.A1.n12 VSS 0.061948f
C9890 mux8_5.A1.n13 VSS 0.408434f
C9891 mux8_5.A1.n14 VSS 0.092045f
C9892 mux8_5.A1.n15 VSS 0.404005f
C9893 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_0.B VSS 0.906354f
C9894 MULT_0.4bit_ADDER_0.FULL_ADDER_2.A VSS 5.06024f
C9895 MULT_0.4bit_ADDER_0.A1.n0 VSS 4.0034f
C9896 MULT_0.4bit_ADDER_0.A1.t12 VSS 0.069048f
C9897 MULT_0.4bit_ADDER_0.A1.t4 VSS 0.026504f
C9898 MULT_0.4bit_ADDER_0.A1.t14 VSS 0.036601f
C9899 MULT_0.4bit_ADDER_0.A1.n1 VSS 0.042128f
C9900 MULT_0.4bit_ADDER_0.A1.t5 VSS 0.027859f
C9901 MULT_0.4bit_ADDER_0.A1.n2 VSS 0.042723f
C9902 MULT_0.4bit_ADDER_0.A1.n3 VSS 0.176842f
C9903 MULT_0.4bit_ADDER_0.FULL_ADDER_2.NAND2_0.B VSS 0.683271f
C9904 MULT_0.4bit_ADDER_0.A1.t6 VSS 0.074769f
C9905 MULT_0.4bit_ADDER_0.A1.t10 VSS 0.073839f
C9906 MULT_0.4bit_ADDER_0.A1.t13 VSS 0.073839f
C9907 MULT_0.4bit_ADDER_0.A1.t11 VSS 0.073839f
C9908 MULT_0.4bit_ADDER_0.A1.n4 VSS 0.2939f
C9909 MULT_0.4bit_ADDER_0.A1.t9 VSS 0.015344f
C9910 MULT_0.4bit_ADDER_0.A1.t8 VSS 0.015344f
C9911 MULT_0.4bit_ADDER_0.A1.t15 VSS 0.015344f
C9912 MULT_0.4bit_ADDER_0.A1.t7 VSS 0.015344f
C9913 MULT_0.4bit_ADDER_0.A1.n5 VSS 0.27765f
C9914 MULT_0.4bit_ADDER_0.A1.n6 VSS 0.4343f
C9915 MULT_0.4bit_ADDER_0.A1.n7 VSS 1.02626f
C9916 MULT_0.4bit_ADDER_0.A1.t1 VSS 0.021891f
C9917 MULT_0.4bit_ADDER_0.A1.t3 VSS 0.021891f
C9918 MULT_0.4bit_ADDER_0.A1.n8 VSS 0.048649f
C9919 MULT_0.4bit_ADDER_0.A1.t0 VSS 0.063431f
C9920 MULT_0.4bit_ADDER_0.A1.t2 VSS 0.0794f
C9921 MULT_0.NAND2_5.Y.n0 VSS 1.19039f
C9922 MULT_0.NAND2_5.Y.n1 VSS 0.18698f
C9923 MULT_0.NAND2_5.Y.t6 VSS 0.023031f
C9924 MULT_0.NAND2_5.Y.t4 VSS 0.023031f
C9925 MULT_0.NAND2_5.Y.n2 VSS 0.051248f
C9926 MULT_0.NAND2_5.Y.t1 VSS 0.023031f
C9927 MULT_0.NAND2_5.Y.t0 VSS 0.023031f
C9928 MULT_0.NAND2_5.Y.n3 VSS 0.051387f
C9929 MULT_0.NAND2_5.Y.t5 VSS 0.023031f
C9930 MULT_0.NAND2_5.Y.t2 VSS 0.023031f
C9931 MULT_0.NAND2_5.Y.n4 VSS 0.051248f
C9932 MULT_0.NAND2_5.Y.t3 VSS 0.138745f
C9933 MULT_0.NAND2_5.Y.t7 VSS 0.029352f
C9934 MULT_0.NAND2_5.Y.t10 VSS 0.040972f
C9935 MULT_0.NAND2_5.Y.t8 VSS 0.040972f
C9936 MULT_0.NAND2_5.Y.n5 VSS 0.133738f
C9937 MULT_0.NAND2_5.Y.t9 VSS 0.046781f
C9938 mux8_0.NAND4F_0.Y.n0 VSS 0.350455f
C9939 mux8_0.NAND4F_0.Y.t10 VSS 0.022537f
C9940 mux8_0.NAND4F_0.Y.t11 VSS 0.079785f
C9941 mux8_0.NAND4F_0.Y.t9 VSS 0.024808f
C9942 mux8_0.NAND4F_0.Y.n1 VSS 0.070768f
C9943 mux8_0.NAND4F_0.Y.n2 VSS 0.020978f
C9944 mux8_0.NAND4F_0.Y.t5 VSS 0.017278f
C9945 mux8_0.NAND4F_0.Y.t6 VSS 0.017278f
C9946 mux8_0.NAND4F_0.Y.n3 VSS 0.040122f
C9947 mux8_0.NAND4F_0.Y.t1 VSS 0.017278f
C9948 mux8_0.NAND4F_0.Y.t0 VSS 0.017278f
C9949 mux8_0.NAND4F_0.Y.n4 VSS 0.040002f
C9950 mux8_0.NAND4F_0.Y.t8 VSS 0.017278f
C9951 mux8_0.NAND4F_0.Y.t7 VSS 0.017278f
C9952 mux8_0.NAND4F_0.Y.n5 VSS 0.040002f
C9953 mux8_0.NAND4F_0.Y.t4 VSS 0.017278f
C9954 mux8_0.NAND4F_0.Y.t3 VSS 0.017278f
C9955 mux8_0.NAND4F_0.Y.n6 VSS 0.040002f
C9956 mux8_0.NAND4F_0.Y.t2 VSS 0.166327f
C9957 left_shifter_0.S1.n0 VSS 16.8575f
C9958 mux8_2.NAND4F_5.A VSS 1.98966f
C9959 left_shifter_0.S1.t4 VSS 0.163797f
C9960 left_shifter_0.S1.t5 VSS 0.482595f
C9961 left_shifter_0.S1.t6 VSS 0.159364f
C9962 left_shifter_0.S1.n1 VSS 0.821633f
C9963 left_shifter_0.S1.t1 VSS 0.07852f
C9964 left_shifter_0.S1.t2 VSS 0.07852f
C9965 left_shifter_0.S1.n2 VSS 0.175162f
C9966 left_shifter_0.S1.t3 VSS 0.284995f
C9967 left_shifter_0.S1.t0 VSS 0.226477f
C9968 mux8_2.A6 VSS 17.6817f
C9969 8bit_ADDER_0.S0.t14 VSS 0.064306f
C9970 8bit_ADDER_0.S0.t12 VSS 0.062566f
C9971 8bit_ADDER_0.S0.t13 VSS 0.189465f
C9972 8bit_ADDER_0.S0.n0 VSS 0.322571f
C9973 8bit_ADDER_0.S0.t9 VSS 0.018726f
C9974 8bit_ADDER_0.S0.t8 VSS 0.018726f
C9975 8bit_ADDER_0.S0.n1 VSS 0.045292f
C9976 8bit_ADDER_0.S0.t0 VSS 0.018726f
C9977 8bit_ADDER_0.S0.t2 VSS 0.018726f
C9978 8bit_ADDER_0.S0.n2 VSS 0.045287f
C9979 8bit_ADDER_0.S0.n3 VSS 0.324749f
C9980 8bit_ADDER_0.S0.t10 VSS 0.018726f
C9981 8bit_ADDER_0.S0.t1 VSS 0.018726f
C9982 8bit_ADDER_0.S0.n4 VSS 0.037453f
C9983 8bit_ADDER_0.S0.n5 VSS 0.02942f
C9984 8bit_ADDER_0.S0.t11 VSS 0.079227f
C9985 8bit_ADDER_0.S0.t3 VSS 0.079227f
C9986 8bit_ADDER_0.S0.n6 VSS 0.158455f
C9987 8bit_ADDER_0.S0.n7 VSS 0.063004f
C9988 8bit_ADDER_0.S0.t7 VSS 0.079227f
C9989 8bit_ADDER_0.S0.t6 VSS 0.079227f
C9990 8bit_ADDER_0.S0.n8 VSS 0.158455f
C9991 8bit_ADDER_0.S0.n9 VSS 0.069691f
C9992 8bit_ADDER_0.S0.n10 VSS 0.717509f
C9993 8bit_ADDER_0.S0.t5 VSS 0.079227f
C9994 8bit_ADDER_0.S0.t4 VSS 0.079227f
C9995 8bit_ADDER_0.S0.n11 VSS 0.158455f
C9996 8bit_ADDER_0.S0.n12 VSS 0.069797f
C9997 8bit_ADDER_0.S0.n13 VSS 0.460179f
C9998 8bit_ADDER_0.S0.n14 VSS 0.103707f
C9999 8bit_ADDER_0.S0.n15 VSS 0.455189f
C10000 AND8_0.S0.n0 VSS 3.31679f
C10001 AND8_0.S0.t5 VSS 0.160494f
C10002 AND8_0.S0.t4 VSS 0.15615f
C10003 AND8_0.S0.t6 VSS 0.472861f
C10004 AND8_0.S0.n1 VSS 0.804994f
C10005 AND8_0.S0.t1 VSS 0.076936f
C10006 AND8_0.S0.t2 VSS 0.076936f
C10007 AND8_0.S0.n2 VSS 0.171447f
C10008 AND8_0.S0.t3 VSS 0.279046f
C10009 AND8_0.S0.t0 VSS 0.221909f
C10010 AND8_0.NOT8_0.A0.n0 VSS 0.588132f
C10011 AND8_0.NOT8_0.A0.t10 VSS 0.014437f
C10012 AND8_0.NOT8_0.A0.t7 VSS 0.020153f
C10013 AND8_0.NOT8_0.A0.t9 VSS 0.020153f
C10014 AND8_0.NOT8_0.A0.n1 VSS 0.065603f
C10015 AND8_0.NOT8_0.A0.t8 VSS 0.023127f
C10016 AND8_0.NOT8_0.A0.n2 VSS 0.20195f
C10017 AND8_0.NOT8_0.A0.t4 VSS 0.068416f
C10018 AND8_0.NOT8_0.A0.t5 VSS 0.011328f
C10019 AND8_0.NOT8_0.A0.t6 VSS 0.011328f
C10020 AND8_0.NOT8_0.A0.n3 VSS 0.025207f
C10021 AND8_0.NOT8_0.A0.t1 VSS 0.011328f
C10022 AND8_0.NOT8_0.A0.t0 VSS 0.011328f
C10023 AND8_0.NOT8_0.A0.n4 VSS 0.025276f
C10024 AND8_0.NOT8_0.A0.t3 VSS 0.011328f
C10025 AND8_0.NOT8_0.A0.t2 VSS 0.011328f
C10026 AND8_0.NOT8_0.A0.n5 VSS 0.025207f
C10027 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n0 VSS 0.860417f
C10028 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t6 VSS 0.007445f
C10029 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t4 VSS 0.007445f
C10030 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n1 VSS 0.016611f
C10031 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t1 VSS 0.007445f
C10032 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t5 VSS 0.007445f
C10033 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n2 VSS 0.016566f
C10034 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t2 VSS 0.007445f
C10035 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t3 VSS 0.007445f
C10036 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n3 VSS 0.016566f
C10037 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t0 VSS 0.044951f
C10038 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t15 VSS 0.025427f
C10039 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t17 VSS 0.025111f
C10040 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t16 VSS 0.025111f
C10041 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t13 VSS 0.025111f
C10042 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n4 VSS 0.099949f
C10043 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t10 VSS 0.005218f
C10044 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t18 VSS 0.005218f
C10045 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t9 VSS 0.005218f
C10046 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t14 VSS 0.005218f
C10047 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n5 VSS 0.094423f
C10048 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n6 VSS 0.147672f
C10049 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t11 VSS 0.023482f
C10050 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t8 VSS 0.009013f
C10051 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t12 VSS 0.012447f
C10052 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n7 VSS 0.014327f
C10053 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.t7 VSS 0.009474f
C10054 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n8 VSS 0.014529f
C10055 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n9 VSS 0.049349f
C10056 8bit_ADDER_0.FULL_ADDER_XORED_7.COUT.n10 VSS 0.328172f
C10057 a_n12314_n26419.n0 VSS 1.48365f
C10058 a_n12314_n26419.n1 VSS 1.48326f
C10059 a_n12314_n26419.t3 VSS 0.093341f
C10060 a_n12314_n26419.t10 VSS 0.093341f
C10061 a_n12314_n26419.t11 VSS 0.093341f
C10062 a_n12314_n26419.n2 VSS 0.202296f
C10063 a_n12314_n26419.t9 VSS 0.093341f
C10064 a_n12314_n26419.t0 VSS 0.093341f
C10065 a_n12314_n26419.n3 VSS 0.202001f
C10066 a_n12314_n26419.t1 VSS 0.093341f
C10067 a_n12314_n26419.t2 VSS 0.093341f
C10068 a_n12314_n26419.n4 VSS 0.202001f
C10069 a_n12314_n26419.t6 VSS 0.093341f
C10070 a_n12314_n26419.t8 VSS 0.093341f
C10071 a_n12314_n26419.n5 VSS 0.202001f
C10072 a_n12314_n26419.t7 VSS 0.093341f
C10073 a_n12314_n26419.t4 VSS 0.093341f
C10074 a_n12314_n26419.n6 VSS 0.202001f
C10075 a_n12314_n26419.n7 VSS 0.20269f
C10076 a_n12314_n26419.t5 VSS 0.093341f
C10077 MULT_0.4bit_ADDER_1.B1.t13 VSS 0.042042f
C10078 MULT_0.4bit_ADDER_1.B1.t18 VSS 0.013691f
C10079 MULT_0.4bit_ADDER_1.B1.t15 VSS 0.018907f
C10080 MULT_0.4bit_ADDER_1.B1.n0 VSS 0.020388f
C10081 MULT_0.4bit_ADDER_1.B1.t22 VSS 0.014075f
C10082 MULT_0.4bit_ADDER_1.B1.n1 VSS 0.035714f
C10083 MULT_0.4bit_ADDER_1.B1.n2 VSS 0.062649f
C10084 MULT_0.4bit_ADDER_1.B1.t17 VSS 0.019196f
C10085 MULT_0.4bit_ADDER_1.B1.t12 VSS 0.038622f
C10086 MULT_0.4bit_ADDER_1.B1.t19 VSS 0.038142f
C10087 MULT_0.4bit_ADDER_1.B1.t20 VSS 0.038142f
C10088 MULT_0.4bit_ADDER_1.B1.t16 VSS 0.038142f
C10089 MULT_0.4bit_ADDER_1.B1.t14 VSS 0.007926f
C10090 MULT_0.4bit_ADDER_1.B1.t21 VSS 0.007926f
C10091 MULT_0.4bit_ADDER_1.B1.t23 VSS 0.007926f
C10092 MULT_0.4bit_ADDER_1.B1.n3 VSS 0.234988f
C10093 MULT_0.4bit_ADDER_1.B1.n4 VSS 0.173079f
C10094 MULT_0.4bit_ADDER_1.B1.n5 VSS 0.094327f
C10095 MULT_0.4bit_ADDER_1.B1.n6 VSS 0.092668f
C10096 MULT_0.4bit_ADDER_1.B1.n7 VSS 0.057001f
C10097 MULT_0.4bit_ADDER_1.B1.n8 VSS 0.074776f
C10098 MULT_0.4bit_ADDER_1.B1.n9 VSS 0.823627f
C10099 MULT_0.4bit_ADDER_1.B1.t0 VSS 0.006869f
C10100 MULT_0.4bit_ADDER_1.B1.t1 VSS 0.006869f
C10101 MULT_0.4bit_ADDER_1.B1.n10 VSS 0.016615f
C10102 MULT_0.4bit_ADDER_1.B1.t7 VSS 0.006869f
C10103 MULT_0.4bit_ADDER_1.B1.t6 VSS 0.006869f
C10104 MULT_0.4bit_ADDER_1.B1.n11 VSS 0.016613f
C10105 MULT_0.4bit_ADDER_1.B1.n12 VSS 0.119127f
C10106 MULT_0.4bit_ADDER_1.B1.t2 VSS 0.006869f
C10107 MULT_0.4bit_ADDER_1.B1.t8 VSS 0.006869f
C10108 MULT_0.4bit_ADDER_1.B1.n13 VSS 0.013739f
C10109 MULT_0.4bit_ADDER_1.B1.n14 VSS 0.010792f
C10110 MULT_0.4bit_ADDER_1.B1.t9 VSS 0.029063f
C10111 MULT_0.4bit_ADDER_1.B1.t4 VSS 0.029063f
C10112 MULT_0.4bit_ADDER_1.B1.n15 VSS 0.058126f
C10113 MULT_0.4bit_ADDER_1.B1.n16 VSS 0.023112f
C10114 MULT_0.4bit_ADDER_1.B1.t10 VSS 0.029063f
C10115 MULT_0.4bit_ADDER_1.B1.t11 VSS 0.029063f
C10116 MULT_0.4bit_ADDER_1.B1.n17 VSS 0.058126f
C10117 MULT_0.4bit_ADDER_1.B1.n18 VSS 0.025565f
C10118 MULT_0.4bit_ADDER_1.B1.n19 VSS 0.263202f
C10119 MULT_0.4bit_ADDER_1.B1.t3 VSS 0.029063f
C10120 MULT_0.4bit_ADDER_1.B1.t5 VSS 0.029063f
C10121 MULT_0.4bit_ADDER_1.B1.n20 VSS 0.058126f
C10122 MULT_0.4bit_ADDER_1.B1.n21 VSS 0.025603f
C10123 MULT_0.4bit_ADDER_1.B1.n22 VSS 0.168806f
C10124 MULT_0.4bit_ADDER_1.B1.n23 VSS 0.038042f
C10125 MULT_0.4bit_ADDER_1.B1.n24 VSS 0.166976f
C10126 mux8_7.NAND4F_9.Y.n0 VSS 0.358256f
C10127 mux8_7.NAND4F_9.Y.t10 VSS 0.017853f
C10128 mux8_7.NAND4F_9.Y.t9 VSS 0.017853f
C10129 mux8_7.NAND4F_9.Y.t14 VSS 0.017853f
C10130 mux8_7.NAND4F_9.Y.t13 VSS 0.017853f
C10131 mux8_7.NAND4F_9.Y.t12 VSS 0.022554f
C10132 mux8_7.NAND4F_9.Y.n1 VSS 0.048188f
C10133 mux8_7.NAND4F_9.Y.n2 VSS 0.030339f
C10134 mux8_7.NAND4F_9.Y.n3 VSS 0.030339f
C10135 mux8_7.NAND4F_9.Y.n4 VSS 0.026149f
C10136 mux8_7.NAND4F_9.Y.t11 VSS 0.014813f
C10137 mux8_7.NAND4F_9.Y.n5 VSS 0.021261f
C10138 mux8_7.NAND4F_9.Y.t4 VSS 0.141821f
C10139 mux8_7.NAND4F_9.Y.t0 VSS 0.017663f
C10140 mux8_7.NAND4F_9.Y.t1 VSS 0.017663f
C10141 mux8_7.NAND4F_9.Y.n6 VSS 0.041015f
C10142 mux8_7.NAND4F_9.Y.t7 VSS 0.017663f
C10143 mux8_7.NAND4F_9.Y.t8 VSS 0.017663f
C10144 mux8_7.NAND4F_9.Y.n7 VSS 0.040893f
C10145 mux8_7.NAND4F_9.Y.t2 VSS 0.017663f
C10146 mux8_7.NAND4F_9.Y.t3 VSS 0.017663f
C10147 mux8_7.NAND4F_9.Y.n8 VSS 0.040893f
C10148 mux8_7.NAND4F_9.Y.t6 VSS 0.017663f
C10149 mux8_7.NAND4F_9.Y.t5 VSS 0.017663f
C10150 mux8_7.NAND4F_9.Y.n9 VSS 0.040893f
C10151 mux8_7.NAND4F_9.Y.n10 VSS 0.168091f
C10152 mux8_8.NAND4F_7.Y.n0 VSS 0.11858f
C10153 mux8_8.NAND4F_7.Y.n1 VSS 0.350455f
C10154 mux8_8.NAND4F_7.Y.t8 VSS 0.168166f
C10155 mux8_8.NAND4F_7.Y.t9 VSS 0.022537f
C10156 mux8_8.NAND4F_7.Y.t11 VSS 0.079785f
C10157 mux8_8.NAND4F_7.Y.t10 VSS 0.024808f
C10158 mux8_8.NAND4F_7.Y.n2 VSS 0.070768f
C10159 mux8_8.NAND4F_7.Y.n3 VSS 0.020978f
C10160 mux8_8.NAND4F_7.Y.t1 VSS 0.017278f
C10161 mux8_8.NAND4F_7.Y.t0 VSS 0.017278f
C10162 mux8_8.NAND4F_7.Y.n4 VSS 0.040122f
C10163 mux8_8.NAND4F_7.Y.t2 VSS 0.017278f
C10164 mux8_8.NAND4F_7.Y.t3 VSS 0.017278f
C10165 mux8_8.NAND4F_7.Y.n5 VSS 0.040002f
C10166 mux8_8.NAND4F_7.Y.t5 VSS 0.017278f
C10167 mux8_8.NAND4F_7.Y.t4 VSS 0.017278f
C10168 mux8_8.NAND4F_7.Y.n6 VSS 0.040002f
C10169 mux8_8.NAND4F_7.Y.t6 VSS 0.017278f
C10170 mux8_8.NAND4F_7.Y.t7 VSS 0.017278f
C10171 mux8_8.NAND4F_7.Y.n7 VSS 0.040002f
C10172 NOT8_0.S6.n0 VSS 1.76051f
C10173 NOT8_0.S6.t6 VSS 0.084969f
C10174 NOT8_0.S6.t5 VSS 0.250343f
C10175 NOT8_0.S6.t4 VSS 0.082669f
C10176 NOT8_0.S6.n1 VSS 0.426218f
C10177 NOT8_0.S6.t1 VSS 0.040732f
C10178 NOT8_0.S6.t2 VSS 0.040732f
C10179 NOT8_0.S6.n2 VSS 0.090768f
C10180 NOT8_0.S6.t3 VSS 0.147733f
C10181 NOT8_0.S6.t0 VSS 0.117484f
C10182 B2.t37 VSS 0.05134f
C10183 B2.t44 VSS 0.071666f
C10184 B2.t42 VSS 0.071666f
C10185 B2.n0 VSS 0.23329f
C10186 B2.t22 VSS 0.08224f
C10187 B2.n1 VSS 0.575854f
C10188 B2.t47 VSS 0.068384f
C10189 B2.t1 VSS 0.137591f
C10190 B2.t25 VSS 0.135879f
C10191 B2.t15 VSS 0.135879f
C10192 B2.t5 VSS 0.135879f
C10193 B2.t12 VSS 0.028237f
C10194 B2.t51 VSS 0.028237f
C10195 B2.t36 VSS 0.028237f
C10196 B2.n2 VSS 0.837136f
C10197 B2.n3 VSS 0.616589f
C10198 B2.n4 VSS 0.336036f
C10199 B2.n5 VSS 0.330126f
C10200 B2.n6 VSS 0.203066f
C10201 B2.n7 VSS 0.230927f
C10202 B2.t46 VSS 0.127063f
C10203 B2.t13 VSS 0.048773f
C10204 B2.t9 VSS 0.067354f
C10205 B2.n8 VSS 0.077524f
C10206 B2.t32 VSS 0.051267f
C10207 B2.n9 VSS 0.07862f
C10208 B2.n10 VSS 0.325046f
C10209 B2.t0 VSS 0.149775f
C10210 B2.t41 VSS 0.048773f
C10211 B2.t34 VSS 0.067354f
C10212 B2.n11 VSS 0.072633f
C10213 B2.t43 VSS 0.050142f
C10214 B2.n12 VSS 0.127229f
C10215 B2.n13 VSS 0.223587f
C10216 B2.n14 VSS 3.26838f
C10217 B2.t3 VSS 0.127063f
C10218 B2.t40 VSS 0.048773f
C10219 B2.t18 VSS 0.067354f
C10220 B2.n15 VSS 0.077524f
C10221 B2.t39 VSS 0.051267f
C10222 B2.n16 VSS 0.07862f
C10223 B2.n17 VSS 0.326238f
C10224 B2.t21 VSS 0.149775f
C10225 B2.t24 VSS 0.048773f
C10226 B2.t8 VSS 0.067354f
C10227 B2.n18 VSS 0.072633f
C10228 B2.t29 VSS 0.050142f
C10229 B2.n19 VSS 0.127229f
C10230 B2.n20 VSS 0.223587f
C10231 B2.n21 VSS 2.93302f
C10232 B2.n22 VSS 22.6259f
C10233 B2.t19 VSS 0.149946f
C10234 B2.t49 VSS 0.064218f
C10235 B2.t52 VSS 0.05134f
C10236 B2.n23 VSS 0.075769f
C10237 B2.t14 VSS 0.050142f
C10238 B2.n24 VSS 0.125081f
C10239 B2.n25 VSS 0.223156f
C10240 B2.n26 VSS 0.318221f
C10241 B2.n27 VSS 3.01592f
C10242 B2.t27 VSS 0.061265f
C10243 B2.t26 VSS 0.065715f
C10244 B2.n28 VSS 0.097922f
C10245 B2.t31 VSS 0.061265f
C10246 B2.t2 VSS 0.061265f
C10247 B2.t4 VSS 0.061265f
C10248 B2.t17 VSS 0.077399f
C10249 B2.n29 VSS 0.165369f
C10250 B2.n30 VSS 0.104117f
C10251 B2.n31 VSS 0.085076f
C10252 B2.n32 VSS 0.04163f
C10253 B2.n33 VSS 6.50337f
C10254 B2.t16 VSS 0.068384f
C10255 B2.t45 VSS 0.137591f
C10256 B2.t50 VSS 0.135879f
C10257 B2.t30 VSS 0.135879f
C10258 B2.t11 VSS 0.135879f
C10259 B2.t28 VSS 0.028237f
C10260 B2.t53 VSS 0.028237f
C10261 B2.t33 VSS 0.028237f
C10262 B2.n34 VSS 0.836925f
C10263 B2.n35 VSS 0.6168f
C10264 B2.n36 VSS 0.336036f
C10265 B2.n37 VSS 0.330126f
C10266 B2.n38 VSS 0.203066f
C10267 B2.n39 VSS 0.261306f
C10268 B2.n40 VSS 1.11027f
C10269 B2.n41 VSS 7.07726f
C10270 B2.t23 VSS 0.05134f
C10271 B2.t7 VSS 0.071666f
C10272 B2.t6 VSS 0.071666f
C10273 B2.n42 VSS 0.23329f
C10274 B2.t48 VSS 0.08224f
C10275 B2.n43 VSS 0.70445f
C10276 B2.n44 VSS 0.457422f
C10277 B2.n45 VSS 5.23113f
C10278 B2.t38 VSS 0.05134f
C10279 B2.t10 VSS 0.071666f
C10280 B2.t35 VSS 0.071666f
C10281 B2.n46 VSS 0.23329f
C10282 B2.t20 VSS 0.08224f
C10283 B2.n47 VSS 0.573448f
C10284 B2.n48 VSS 0.507453f
C10285 B2.n49 VSS 3.84331f
C10286 B2.n50 VSS 0.663052f
C10287 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t12 VSS 0.013766f
C10288 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t17 VSS 0.027698f
C10289 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t19 VSS 0.027354f
C10290 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t18 VSS 0.027354f
C10291 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t16 VSS 0.027354f
C10292 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t13 VSS 0.005684f
C10293 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t23 VSS 0.005684f
C10294 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t22 VSS 0.005684f
C10295 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n0 VSS 0.168523f
C10296 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n1 VSS 0.124125f
C10297 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n2 VSS 0.067647f
C10298 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n3 VSS 0.066457f
C10299 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n4 VSS 0.040879f
C10300 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n5 VSS 0.05311f
C10301 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t14 VSS 0.030151f
C10302 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t21 VSS 0.009818f
C10303 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t20 VSS 0.013559f
C10304 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n6 VSS 0.014622f
C10305 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t15 VSS 0.010094f
C10306 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n7 VSS 0.025612f
C10307 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n8 VSS 0.044927f
C10308 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t10 VSS 0.004926f
C10309 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t11 VSS 0.004926f
C10310 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n9 VSS 0.011915f
C10311 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t4 VSS 0.004926f
C10312 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t7 VSS 0.004926f
C10313 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n10 VSS 0.011914f
C10314 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n11 VSS 0.085433f
C10315 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t9 VSS 0.004926f
C10316 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t3 VSS 0.004926f
C10317 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n12 VSS 0.009853f
C10318 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n13 VSS 0.00774f
C10319 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t0 VSS 0.020843f
C10320 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t5 VSS 0.020843f
C10321 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n14 VSS 0.041685f
C10322 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n15 VSS 0.016575f
C10323 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t1 VSS 0.020843f
C10324 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t2 VSS 0.020843f
C10325 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n16 VSS 0.041685f
C10326 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n17 VSS 0.018334f
C10327 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n18 VSS 0.188757f
C10328 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t6 VSS 0.020843f
C10329 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.t8 VSS 0.020843f
C10330 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n19 VSS 0.041685f
C10331 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n20 VSS 0.018362f
C10332 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n21 VSS 0.12106f
C10333 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n22 VSS 0.027282f
C10334 MULT_0.4bit_ADDER_0.FULL_ADDER_1.XOR2_1.A.n23 VSS 0.119748f
C10335 mux8_8.NAND4F_5.Y.n0 VSS 0.25108f
C10336 mux8_8.NAND4F_5.Y.t10 VSS 0.017162f
C10337 mux8_8.NAND4F_5.Y.t9 VSS 0.050565f
C10338 mux8_8.NAND4F_5.Y.t11 VSS 0.016698f
C10339 mux8_8.NAND4F_5.Y.n1 VSS 0.086077f
C10340 mux8_8.NAND4F_5.Y.t2 VSS 0.099394f
C10341 mux8_8.NAND4F_5.Y.n2 VSS 0.798124f
C10342 mux8_8.NAND4F_5.Y.t0 VSS 0.012379f
C10343 mux8_8.NAND4F_5.Y.t1 VSS 0.012379f
C10344 mux8_8.NAND4F_5.Y.n3 VSS 0.028745f
C10345 mux8_8.NAND4F_5.Y.t6 VSS 0.012379f
C10346 mux8_8.NAND4F_5.Y.t5 VSS 0.012379f
C10347 mux8_8.NAND4F_5.Y.n4 VSS 0.028659f
C10348 mux8_8.NAND4F_5.Y.t7 VSS 0.012379f
C10349 mux8_8.NAND4F_5.Y.t8 VSS 0.012379f
C10350 mux8_8.NAND4F_5.Y.n5 VSS 0.028659f
C10351 mux8_8.NAND4F_5.Y.t3 VSS 0.012379f
C10352 mux8_8.NAND4F_5.Y.t4 VSS 0.012379f
C10353 mux8_8.NAND4F_5.Y.n6 VSS 0.028659f
C10354 mux8_8.NAND4F_5.Y.n7 VSS 0.117805f
C10355 MULT_0.NAND2_11.Y.n0 VSS 1.24545f
C10356 MULT_0.NAND2_11.Y.n1 VSS 0.196221f
C10357 MULT_0.NAND2_11.Y.t6 VSS 0.024169f
C10358 MULT_0.NAND2_11.Y.t5 VSS 0.024169f
C10359 MULT_0.NAND2_11.Y.n2 VSS 0.05378f
C10360 MULT_0.NAND2_11.Y.t1 VSS 0.024169f
C10361 MULT_0.NAND2_11.Y.t0 VSS 0.024169f
C10362 MULT_0.NAND2_11.Y.n3 VSS 0.053926f
C10363 MULT_0.NAND2_11.Y.t4 VSS 0.024169f
C10364 MULT_0.NAND2_11.Y.t2 VSS 0.024169f
C10365 MULT_0.NAND2_11.Y.n4 VSS 0.05378f
C10366 MULT_0.NAND2_11.Y.t3 VSS 0.145599f
C10367 MULT_0.NAND2_11.Y.t10 VSS 0.030802f
C10368 MULT_0.NAND2_11.Y.t9 VSS 0.042997f
C10369 MULT_0.NAND2_11.Y.t7 VSS 0.042997f
C10370 MULT_0.NAND2_11.Y.n5 VSS 0.140346f
C10371 MULT_0.NAND2_11.Y.t8 VSS 0.049092f
C10372 a_n914_3810.n0 VSS 1.45527f
C10373 a_n914_3810.n1 VSS 1.45566f
C10374 a_n914_3810.t3 VSS 0.09158f
C10375 a_n914_3810.t7 VSS 0.09158f
C10376 a_n914_3810.t8 VSS 0.09158f
C10377 a_n914_3810.n2 VSS 0.198865f
C10378 a_n914_3810.t6 VSS 0.09158f
C10379 a_n914_3810.t11 VSS 0.09158f
C10380 a_n914_3810.n3 VSS 0.19819f
C10381 a_n914_3810.t10 VSS 0.09158f
C10382 a_n914_3810.t9 VSS 0.09158f
C10383 a_n914_3810.n4 VSS 0.19819f
C10384 a_n914_3810.t5 VSS 0.09158f
C10385 a_n914_3810.t4 VSS 0.09158f
C10386 a_n914_3810.n5 VSS 0.19819f
C10387 a_n914_3810.t0 VSS 0.09158f
C10388 a_n914_3810.t1 VSS 0.09158f
C10389 a_n914_3810.n6 VSS 0.198479f
C10390 a_n914_3810.n7 VSS 0.19819f
C10391 a_n914_3810.t2 VSS 0.09158f
C10392 mux8_6.NAND4F_5.Y.n0 VSS 0.25108f
C10393 mux8_6.NAND4F_5.Y.t10 VSS 0.017162f
C10394 mux8_6.NAND4F_5.Y.t9 VSS 0.050565f
C10395 mux8_6.NAND4F_5.Y.t11 VSS 0.016698f
C10396 mux8_6.NAND4F_5.Y.n1 VSS 0.086077f
C10397 mux8_6.NAND4F_5.Y.t2 VSS 0.099394f
C10398 mux8_6.NAND4F_5.Y.n2 VSS 0.798124f
C10399 mux8_6.NAND4F_5.Y.t1 VSS 0.012379f
C10400 mux8_6.NAND4F_5.Y.t0 VSS 0.012379f
C10401 mux8_6.NAND4F_5.Y.n3 VSS 0.028745f
C10402 mux8_6.NAND4F_5.Y.t6 VSS 0.012379f
C10403 mux8_6.NAND4F_5.Y.t5 VSS 0.012379f
C10404 mux8_6.NAND4F_5.Y.n4 VSS 0.028659f
C10405 mux8_6.NAND4F_5.Y.t7 VSS 0.012379f
C10406 mux8_6.NAND4F_5.Y.t8 VSS 0.012379f
C10407 mux8_6.NAND4F_5.Y.n5 VSS 0.028659f
C10408 mux8_6.NAND4F_5.Y.t4 VSS 0.012379f
C10409 mux8_6.NAND4F_5.Y.t3 VSS 0.012379f
C10410 mux8_6.NAND4F_5.Y.n6 VSS 0.028659f
C10411 mux8_6.NAND4F_5.Y.n7 VSS 0.117805f
C10412 mux8_6.NAND4F_4.B.n0 VSS 0.921489f
C10413 mux8_6.NAND4F_4.B.t4 VSS 0.03989f
C10414 mux8_6.NAND4F_4.B.t5 VSS 0.123086f
C10415 mux8_6.NAND4F_4.B.t15 VSS 0.04595f
C10416 mux8_6.NAND4F_4.B.n1 VSS 0.154452f
C10417 mux8_6.NAND4F_4.B.n2 VSS 0.033769f
C10418 mux8_6.NAND4F_4.B.t13 VSS 0.03989f
C10419 mux8_6.NAND4F_4.B.t9 VSS 0.123086f
C10420 mux8_6.NAND4F_4.B.t11 VSS 0.04595f
C10421 mux8_6.NAND4F_4.B.n3 VSS 0.154452f
C10422 mux8_6.NAND4F_4.B.n4 VSS 0.032977f
C10423 mux8_6.NAND4F_4.B.t8 VSS 0.03989f
C10424 mux8_6.NAND4F_4.B.t6 VSS 0.123086f
C10425 mux8_6.NAND4F_4.B.t7 VSS 0.04595f
C10426 mux8_6.NAND4F_4.B.n5 VSS 0.154452f
C10427 mux8_6.NAND4F_4.B.n6 VSS 0.033699f
C10428 mux8_6.NAND4F_4.B.n7 VSS 0.612655f
C10429 mux8_6.NAND4F_4.B.t3 VSS 0.020325f
C10430 mux8_6.NAND4F_4.B.t2 VSS 0.020325f
C10431 mux8_6.NAND4F_4.B.n8 VSS 0.045293f
C10432 mux8_6.NAND4F_4.B.t1 VSS 0.073718f
C10433 mux8_6.NAND4F_4.B.t0 VSS 0.058624f
C10434 mux8_6.NAND4F_4.B.n9 VSS 0.607515f
C10435 mux8_6.NAND4F_4.B.t12 VSS 0.03989f
C10436 mux8_6.NAND4F_4.B.t14 VSS 0.123086f
C10437 mux8_6.NAND4F_4.B.t10 VSS 0.04595f
C10438 mux8_6.NAND4F_4.B.n10 VSS 0.154452f
C10439 mux8_6.NAND4F_4.B.n11 VSS 0.033659f
C10440 mux8_6.NAND4F_4.B.n12 VSS 0.776456f
C10441 MULT_0.4bit_ADDER_0.FULL_ADDER_3.NAND2_0.A VSS 0.398199f
C10442 MULT_0.4bit_ADDER_0.B0.n0 VSS 3.4599f
C10443 MULT_0.4bit_ADDER_0.FULL_ADDER_3.B VSS 6.635129f
C10444 MULT_0.4bit_ADDER_0.B0.t0 VSS 0.082848f
C10445 MULT_0.4bit_ADDER_0.B0.t1 VSS 0.104006f
C10446 MULT_0.4bit_ADDER_0.B0.t3 VSS 0.028676f
C10447 MULT_0.4bit_ADDER_0.B0.t2 VSS 0.028676f
C10448 MULT_0.4bit_ADDER_0.B0.n1 VSS 0.063887f
C10449 MULT_0.4bit_ADDER_0.B0.t8 VSS 0.106613f
C10450 MULT_0.4bit_ADDER_0.B0.t15 VSS 0.034718f
C10451 MULT_0.4bit_ADDER_0.B0.t14 VSS 0.047944f
C10452 MULT_0.4bit_ADDER_0.B0.n2 VSS 0.051702f
C10453 MULT_0.4bit_ADDER_0.B0.t4 VSS 0.035692f
C10454 MULT_0.4bit_ADDER_0.B0.n3 VSS 0.090565f
C10455 MULT_0.4bit_ADDER_0.B0.n4 VSS 0.158867f
C10456 MULT_0.4bit_ADDER_0.B0.t10 VSS 0.048677f
C10457 MULT_0.4bit_ADDER_0.B0.t12 VSS 0.09794f
C10458 MULT_0.4bit_ADDER_0.B0.t7 VSS 0.096722f
C10459 MULT_0.4bit_ADDER_0.B0.t6 VSS 0.096722f
C10460 MULT_0.4bit_ADDER_0.B0.t11 VSS 0.096722f
C10461 MULT_0.4bit_ADDER_0.B0.t13 VSS 0.0201f
C10462 MULT_0.4bit_ADDER_0.B0.t5 VSS 0.0201f
C10463 MULT_0.4bit_ADDER_0.B0.t9 VSS 0.0201f
C10464 MULT_0.4bit_ADDER_0.B0.n5 VSS 0.595893f
C10465 MULT_0.4bit_ADDER_0.B0.n6 VSS 0.438902f
C10466 MULT_0.4bit_ADDER_0.B0.n7 VSS 0.239198f
C10467 MULT_0.4bit_ADDER_0.B0.n8 VSS 0.234991f
C10468 MULT_0.4bit_ADDER_0.B0.n9 VSS 0.144547f
C10469 MULT_0.4bit_ADDER_0.B0.n10 VSS 0.189619f
C10470 MULT_0.4bit_ADDER_0.FULL_ADDER_3.XOR2_0.A VSS 0.337212f
C10471 MULT_0.4bit_ADDER_0.B0.n11 VSS 2.09514f
C10472 MULT_0.NAND2_14.Y.n0 VSS 1.18962f
C10473 MULT_0.NAND2_14.Y.n1 VSS 0.18714f
C10474 MULT_0.NAND2_14.Y.t5 VSS 0.023051f
C10475 MULT_0.NAND2_14.Y.t4 VSS 0.023051f
C10476 MULT_0.NAND2_14.Y.n2 VSS 0.051291f
C10477 MULT_0.NAND2_14.Y.t0 VSS 0.023051f
C10478 MULT_0.NAND2_14.Y.t1 VSS 0.023051f
C10479 MULT_0.NAND2_14.Y.n3 VSS 0.051431f
C10480 MULT_0.NAND2_14.Y.t3 VSS 0.023051f
C10481 MULT_0.NAND2_14.Y.t2 VSS 0.023051f
C10482 MULT_0.NAND2_14.Y.n4 VSS 0.051291f
C10483 MULT_0.NAND2_14.Y.t6 VSS 0.138862f
C10484 MULT_0.NAND2_14.Y.t10 VSS 0.029376f
C10485 MULT_0.NAND2_14.Y.t8 VSS 0.041007f
C10486 MULT_0.NAND2_14.Y.t7 VSS 0.041007f
C10487 MULT_0.NAND2_14.Y.n5 VSS 0.133851f
C10488 MULT_0.NAND2_14.Y.t9 VSS 0.04682f
C10489 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n0 VSS 0.941081f
C10490 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t6 VSS 0.008143f
C10491 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t4 VSS 0.008143f
C10492 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n1 VSS 0.018168f
C10493 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t1 VSS 0.008143f
C10494 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t5 VSS 0.008143f
C10495 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n2 VSS 0.018119f
C10496 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t3 VSS 0.008143f
C10497 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t2 VSS 0.008143f
C10498 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n3 VSS 0.018119f
C10499 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t0 VSS 0.049166f
C10500 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t13 VSS 0.027811f
C10501 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t10 VSS 0.027465f
C10502 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t11 VSS 0.027465f
C10503 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t8 VSS 0.027465f
C10504 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n4 VSS 0.109319f
C10505 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t7 VSS 0.005708f
C10506 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t16 VSS 0.005708f
C10507 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t12 VSS 0.005708f
C10508 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t18 VSS 0.005708f
C10509 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n5 VSS 0.103275f
C10510 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n6 VSS 0.161516f
C10511 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t17 VSS 0.025683f
C10512 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t15 VSS 0.009858f
C10513 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t14 VSS 0.013614f
C10514 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n7 VSS 0.01567f
C10515 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.t9 VSS 0.010363f
C10516 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n8 VSS 0.015891f
C10517 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n9 VSS 0.053976f
C10518 MULT_0.4bit_ADDER_0.FULL_ADDER_3.COUT.n10 VSS 0.358938f
C10519 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t14 VSS 0.013766f
C10520 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t18 VSS 0.027698f
C10521 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t21 VSS 0.027354f
C10522 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t22 VSS 0.027354f
C10523 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t15 VSS 0.027354f
C10524 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t13 VSS 0.005684f
C10525 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t20 VSS 0.005684f
C10526 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t19 VSS 0.005684f
C10527 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n0 VSS 0.168523f
C10528 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n1 VSS 0.124125f
C10529 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n2 VSS 0.067647f
C10530 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n3 VSS 0.066457f
C10531 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n4 VSS 0.040879f
C10532 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n5 VSS 0.05311f
C10533 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t12 VSS 0.030151f
C10534 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t16 VSS 0.009818f
C10535 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t17 VSS 0.013559f
C10536 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n6 VSS 0.014622f
C10537 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t23 VSS 0.010094f
C10538 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n7 VSS 0.025612f
C10539 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n8 VSS 0.044927f
C10540 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t5 VSS 0.004926f
C10541 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t4 VSS 0.004926f
C10542 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n9 VSS 0.011915f
C10543 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t6 VSS 0.004926f
C10544 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t10 VSS 0.004926f
C10545 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n10 VSS 0.011914f
C10546 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n11 VSS 0.085433f
C10547 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t3 VSS 0.004926f
C10548 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t7 VSS 0.004926f
C10549 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n12 VSS 0.009853f
C10550 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n13 VSS 0.00774f
C10551 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t0 VSS 0.020843f
C10552 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t9 VSS 0.020843f
C10553 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n14 VSS 0.041685f
C10554 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n15 VSS 0.016575f
C10555 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t2 VSS 0.020843f
C10556 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t1 VSS 0.020843f
C10557 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n16 VSS 0.041685f
C10558 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n17 VSS 0.018334f
C10559 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n18 VSS 0.188757f
C10560 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t8 VSS 0.020843f
C10561 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.t11 VSS 0.020843f
C10562 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n19 VSS 0.041685f
C10563 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n20 VSS 0.018362f
C10564 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n21 VSS 0.12106f
C10565 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n22 VSS 0.027282f
C10566 MULT_0.4bit_ADDER_2.FULL_ADDER_2.XOR2_1.A.n23 VSS 0.119748f
C10567 mux8_5.NAND4F_9.Y.n0 VSS 0.358256f
C10568 mux8_5.NAND4F_9.Y.t13 VSS 0.017853f
C10569 mux8_5.NAND4F_9.Y.t12 VSS 0.017853f
C10570 mux8_5.NAND4F_9.Y.t10 VSS 0.017853f
C10571 mux8_5.NAND4F_9.Y.t9 VSS 0.017853f
C10572 mux8_5.NAND4F_9.Y.t14 VSS 0.022554f
C10573 mux8_5.NAND4F_9.Y.n1 VSS 0.048188f
C10574 mux8_5.NAND4F_9.Y.n2 VSS 0.030339f
C10575 mux8_5.NAND4F_9.Y.n3 VSS 0.030339f
C10576 mux8_5.NAND4F_9.Y.n4 VSS 0.026149f
C10577 mux8_5.NAND4F_9.Y.t11 VSS 0.014813f
C10578 mux8_5.NAND4F_9.Y.n5 VSS 0.021261f
C10579 mux8_5.NAND4F_9.Y.t0 VSS 0.141821f
C10580 mux8_5.NAND4F_9.Y.t3 VSS 0.017663f
C10581 mux8_5.NAND4F_9.Y.t4 VSS 0.017663f
C10582 mux8_5.NAND4F_9.Y.n6 VSS 0.041015f
C10583 mux8_5.NAND4F_9.Y.t7 VSS 0.017663f
C10584 mux8_5.NAND4F_9.Y.t8 VSS 0.017663f
C10585 mux8_5.NAND4F_9.Y.n7 VSS 0.040893f
C10586 mux8_5.NAND4F_9.Y.t5 VSS 0.017663f
C10587 mux8_5.NAND4F_9.Y.t6 VSS 0.017663f
C10588 mux8_5.NAND4F_9.Y.n8 VSS 0.040893f
C10589 mux8_5.NAND4F_9.Y.t2 VSS 0.017663f
C10590 mux8_5.NAND4F_9.Y.t1 VSS 0.017663f
C10591 mux8_5.NAND4F_9.Y.n9 VSS 0.040893f
C10592 mux8_5.NAND4F_9.Y.n10 VSS 0.168091f
C10593 a_n9125_n4534.n0 VSS 1.48326f
C10594 a_n9125_n4534.n1 VSS 1.48365f
C10595 a_n9125_n4534.t8 VSS 0.093341f
C10596 a_n9125_n4534.t11 VSS 0.093341f
C10597 a_n9125_n4534.t6 VSS 0.093341f
C10598 a_n9125_n4534.n2 VSS 0.20269f
C10599 a_n9125_n4534.t5 VSS 0.093341f
C10600 a_n9125_n4534.t10 VSS 0.093341f
C10601 a_n9125_n4534.n3 VSS 0.202001f
C10602 a_n9125_n4534.t3 VSS 0.093341f
C10603 a_n9125_n4534.t4 VSS 0.093341f
C10604 a_n9125_n4534.n4 VSS 0.202001f
C10605 a_n9125_n4534.t2 VSS 0.093341f
C10606 a_n9125_n4534.t0 VSS 0.093341f
C10607 a_n9125_n4534.n5 VSS 0.202001f
C10608 a_n9125_n4534.t7 VSS 0.093341f
C10609 a_n9125_n4534.t1 VSS 0.093341f
C10610 a_n9125_n4534.n6 VSS 0.202001f
C10611 a_n9125_n4534.n7 VSS 0.202296f
C10612 a_n9125_n4534.t9 VSS 0.093341f
C10613 mux8_6.NAND4F_7.Y.n0 VSS 0.11858f
C10614 mux8_6.NAND4F_7.Y.n1 VSS 0.350455f
C10615 mux8_6.NAND4F_7.Y.t4 VSS 0.168166f
C10616 mux8_6.NAND4F_7.Y.t9 VSS 0.022537f
C10617 mux8_6.NAND4F_7.Y.t11 VSS 0.079785f
C10618 mux8_6.NAND4F_7.Y.t10 VSS 0.024808f
C10619 mux8_6.NAND4F_7.Y.n2 VSS 0.070768f
C10620 mux8_6.NAND4F_7.Y.n3 VSS 0.020978f
C10621 mux8_6.NAND4F_7.Y.t1 VSS 0.017278f
C10622 mux8_6.NAND4F_7.Y.t0 VSS 0.017278f
C10623 mux8_6.NAND4F_7.Y.n4 VSS 0.040122f
C10624 mux8_6.NAND4F_7.Y.t2 VSS 0.017278f
C10625 mux8_6.NAND4F_7.Y.t3 VSS 0.017278f
C10626 mux8_6.NAND4F_7.Y.n5 VSS 0.040002f
C10627 mux8_6.NAND4F_7.Y.t8 VSS 0.017278f
C10628 mux8_6.NAND4F_7.Y.t7 VSS 0.017278f
C10629 mux8_6.NAND4F_7.Y.n6 VSS 0.040002f
C10630 mux8_6.NAND4F_7.Y.t6 VSS 0.017278f
C10631 mux8_6.NAND4F_7.Y.t5 VSS 0.017278f
C10632 mux8_6.NAND4F_7.Y.n7 VSS 0.040002f
C10633 NOT8_0.S7.n0 VSS 1.33192f
C10634 NOT8_0.S7.t5 VSS 0.064314f
C10635 NOT8_0.S7.t4 VSS 0.189488f
C10636 NOT8_0.S7.t6 VSS 0.062573f
C10637 NOT8_0.S7.n1 VSS 0.32261f
C10638 NOT8_0.S7.t2 VSS 0.03083f
C10639 NOT8_0.S7.t0 VSS 0.03083f
C10640 NOT8_0.S7.n2 VSS 0.068703f
C10641 NOT8_0.S7.t1 VSS 0.111821f
C10642 NOT8_0.S7.t3 VSS 0.088925f
C10643 a_3493_5534.n0 VSS 1.45566f
C10644 a_3493_5534.n1 VSS 1.45527f
C10645 a_3493_5534.t6 VSS 0.09158f
C10646 a_3493_5534.t5 VSS 0.09158f
C10647 a_3493_5534.t3 VSS 0.09158f
C10648 a_3493_5534.n2 VSS 0.198479f
C10649 a_3493_5534.t4 VSS 0.09158f
C10650 a_3493_5534.t9 VSS 0.09158f
C10651 a_3493_5534.n3 VSS 0.19819f
C10652 a_3493_5534.t11 VSS 0.09158f
C10653 a_3493_5534.t10 VSS 0.09158f
C10654 a_3493_5534.n4 VSS 0.19819f
C10655 a_3493_5534.t7 VSS 0.09158f
C10656 a_3493_5534.t8 VSS 0.09158f
C10657 a_3493_5534.n5 VSS 0.19819f
C10658 a_3493_5534.t1 VSS 0.09158f
C10659 a_3493_5534.t0 VSS 0.09158f
C10660 a_3493_5534.n6 VSS 0.198865f
C10661 a_3493_5534.n7 VSS 0.19819f
C10662 a_3493_5534.t2 VSS 0.09158f
C10663 left_shifter_0.S7.n0 VSS 0.936727f
C10664 left_shifter_0.S7.t5 VSS 0.044962f
C10665 left_shifter_0.S7.t4 VSS 0.132472f
C10666 left_shifter_0.S7.t6 VSS 0.043745f
C10667 left_shifter_0.S7.n1 VSS 0.225538f
C10668 left_shifter_0.S7.t2 VSS 0.021554f
C10669 left_shifter_0.S7.t3 VSS 0.021554f
C10670 left_shifter_0.S7.n2 VSS 0.048082f
C10671 left_shifter_0.S7.t1 VSS 0.078231f
C10672 left_shifter_0.S7.t0 VSS 0.062168f
C10673 mux8_3.NAND4F_4.Y.n0 VSS 0.480308f
C10674 mux8_3.NAND4F_4.Y.t7 VSS 0.023681f
C10675 mux8_3.NAND4F_4.Y.t8 VSS 0.023681f
C10676 mux8_3.NAND4F_4.Y.n1 VSS 0.054989f
C10677 mux8_3.NAND4F_4.Y.t3 VSS 0.023681f
C10678 mux8_3.NAND4F_4.Y.t4 VSS 0.023681f
C10679 mux8_3.NAND4F_4.Y.n2 VSS 0.054824f
C10680 mux8_3.NAND4F_4.Y.t5 VSS 0.023681f
C10681 mux8_3.NAND4F_4.Y.t6 VSS 0.023681f
C10682 mux8_3.NAND4F_4.Y.n3 VSS 0.054824f
C10683 mux8_3.NAND4F_4.Y.t0 VSS 0.023681f
C10684 mux8_3.NAND4F_4.Y.t1 VSS 0.023681f
C10685 mux8_3.NAND4F_4.Y.n4 VSS 0.054824f
C10686 mux8_3.NAND4F_4.Y.n5 VSS 0.238711f
C10687 mux8_3.NAND4F_4.Y.t11 VSS 0.032831f
C10688 mux8_3.NAND4F_4.Y.t9 VSS 0.031942f
C10689 mux8_3.NAND4F_4.Y.t10 VSS 0.096729f
C10690 mux8_3.NAND4F_4.Y.n6 VSS 0.164667f
C10691 mux8_3.NAND4F_4.Y.t2 VSS 0.190137f
C10692 mux8_3.NAND4F_4.Y.n7 VSS 1.51729f
C10693 MULT_0.4bit_ADDER_2.B2.t16 VSS 0.041736f
C10694 MULT_0.4bit_ADDER_2.B2.t18 VSS 0.013591f
C10695 MULT_0.4bit_ADDER_2.B2.t15 VSS 0.018769f
C10696 MULT_0.4bit_ADDER_2.B2.n0 VSS 0.02024f
C10697 MULT_0.4bit_ADDER_2.B2.t14 VSS 0.013973f
C10698 MULT_0.4bit_ADDER_2.B2.n1 VSS 0.035453f
C10699 MULT_0.4bit_ADDER_2.B2.n2 VSS 0.062192f
C10700 MULT_0.4bit_ADDER_2.B2.t21 VSS 0.019056f
C10701 MULT_0.4bit_ADDER_2.B2.t12 VSS 0.038341f
C10702 MULT_0.4bit_ADDER_2.B2.t17 VSS 0.037864f
C10703 MULT_0.4bit_ADDER_2.B2.t19 VSS 0.037864f
C10704 MULT_0.4bit_ADDER_2.B2.t22 VSS 0.037864f
C10705 MULT_0.4bit_ADDER_2.B2.t20 VSS 0.007868f
C10706 MULT_0.4bit_ADDER_2.B2.t13 VSS 0.007868f
C10707 MULT_0.4bit_ADDER_2.B2.t23 VSS 0.007868f
C10708 MULT_0.4bit_ADDER_2.B2.n3 VSS 0.233274f
C10709 MULT_0.4bit_ADDER_2.B2.n4 VSS 0.171817f
C10710 MULT_0.4bit_ADDER_2.B2.n5 VSS 0.093639f
C10711 MULT_0.4bit_ADDER_2.B2.n6 VSS 0.091992f
C10712 MULT_0.4bit_ADDER_2.B2.n7 VSS 0.056586f
C10713 MULT_0.4bit_ADDER_2.B2.n8 VSS 0.07423f
C10714 MULT_0.4bit_ADDER_2.B2.n9 VSS 0.817398f
C10715 MULT_0.4bit_ADDER_2.B2.t8 VSS 0.006819f
C10716 MULT_0.4bit_ADDER_2.B2.t7 VSS 0.006819f
C10717 MULT_0.4bit_ADDER_2.B2.n10 VSS 0.016493f
C10718 MULT_0.4bit_ADDER_2.B2.t0 VSS 0.006819f
C10719 MULT_0.4bit_ADDER_2.B2.t2 VSS 0.006819f
C10720 MULT_0.4bit_ADDER_2.B2.n11 VSS 0.016491f
C10721 MULT_0.4bit_ADDER_2.B2.n12 VSS 0.118258f
C10722 MULT_0.4bit_ADDER_2.B2.t6 VSS 0.006819f
C10723 MULT_0.4bit_ADDER_2.B2.t5 VSS 0.006819f
C10724 MULT_0.4bit_ADDER_2.B2.n13 VSS 0.013639f
C10725 MULT_0.4bit_ADDER_2.B2.n14 VSS 0.010713f
C10726 MULT_0.4bit_ADDER_2.B2.t9 VSS 0.028851f
C10727 MULT_0.4bit_ADDER_2.B2.t1 VSS 0.028851f
C10728 MULT_0.4bit_ADDER_2.B2.n15 VSS 0.057702f
C10729 MULT_0.4bit_ADDER_2.B2.n16 VSS 0.022943f
C10730 MULT_0.4bit_ADDER_2.B2.t10 VSS 0.028851f
C10731 MULT_0.4bit_ADDER_2.B2.t11 VSS 0.028851f
C10732 MULT_0.4bit_ADDER_2.B2.n17 VSS 0.057702f
C10733 MULT_0.4bit_ADDER_2.B2.n18 VSS 0.025378f
C10734 MULT_0.4bit_ADDER_2.B2.n19 VSS 0.261283f
C10735 MULT_0.4bit_ADDER_2.B2.t3 VSS 0.028851f
C10736 MULT_0.4bit_ADDER_2.B2.t4 VSS 0.028851f
C10737 MULT_0.4bit_ADDER_2.B2.n20 VSS 0.057702f
C10738 MULT_0.4bit_ADDER_2.B2.n21 VSS 0.025417f
C10739 MULT_0.4bit_ADDER_2.B2.n22 VSS 0.167575f
C10740 MULT_0.4bit_ADDER_2.B2.n23 VSS 0.037765f
C10741 MULT_0.4bit_ADDER_2.B2.n24 VSS 0.165758f
C10742 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t17 VSS 0.013766f
C10743 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t22 VSS 0.027698f
C10744 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t15 VSS 0.027354f
C10745 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t14 VSS 0.027354f
C10746 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t23 VSS 0.027354f
C10747 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t20 VSS 0.005684f
C10748 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t16 VSS 0.005684f
C10749 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t18 VSS 0.005684f
C10750 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n0 VSS 0.168523f
C10751 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n1 VSS 0.124125f
C10752 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n2 VSS 0.067647f
C10753 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n3 VSS 0.066457f
C10754 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n4 VSS 0.040879f
C10755 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n5 VSS 0.05311f
C10756 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t13 VSS 0.030151f
C10757 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t21 VSS 0.009818f
C10758 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t19 VSS 0.013559f
C10759 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n6 VSS 0.014622f
C10760 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t12 VSS 0.010094f
C10761 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n7 VSS 0.025612f
C10762 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n8 VSS 0.044927f
C10763 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t0 VSS 0.004926f
C10764 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t1 VSS 0.004926f
C10765 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n9 VSS 0.011915f
C10766 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t3 VSS 0.004926f
C10767 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t4 VSS 0.004926f
C10768 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n10 VSS 0.011914f
C10769 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n11 VSS 0.085433f
C10770 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t2 VSS 0.004926f
C10771 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t8 VSS 0.004926f
C10772 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n12 VSS 0.009853f
C10773 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n13 VSS 0.00774f
C10774 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t9 VSS 0.020843f
C10775 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t5 VSS 0.020843f
C10776 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n14 VSS 0.041685f
C10777 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n15 VSS 0.016575f
C10778 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t10 VSS 0.020843f
C10779 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t11 VSS 0.020843f
C10780 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n16 VSS 0.041685f
C10781 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n17 VSS 0.018334f
C10782 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n18 VSS 0.188757f
C10783 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t6 VSS 0.020843f
C10784 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.t7 VSS 0.020843f
C10785 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n19 VSS 0.041685f
C10786 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n20 VSS 0.018362f
C10787 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n21 VSS 0.12106f
C10788 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n22 VSS 0.027282f
C10789 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_1.A.n23 VSS 0.119748f
C10790 MULT_0.NAND2_2.Y.n0 VSS 1.24951f
C10791 MULT_0.NAND2_2.Y.n1 VSS 0.195379f
C10792 MULT_0.NAND2_2.Y.t6 VSS 0.024066f
C10793 MULT_0.NAND2_2.Y.t5 VSS 0.024066f
C10794 MULT_0.NAND2_2.Y.n2 VSS 0.053551f
C10795 MULT_0.NAND2_2.Y.t2 VSS 0.024066f
C10796 MULT_0.NAND2_2.Y.t1 VSS 0.024066f
C10797 MULT_0.NAND2_2.Y.n3 VSS 0.053697f
C10798 MULT_0.NAND2_2.Y.t4 VSS 0.024066f
C10799 MULT_0.NAND2_2.Y.t0 VSS 0.024066f
C10800 MULT_0.NAND2_2.Y.n4 VSS 0.053551f
C10801 MULT_0.NAND2_2.Y.t3 VSS 0.14498f
C10802 MULT_0.NAND2_2.Y.t9 VSS 0.030671f
C10803 MULT_0.NAND2_2.Y.t8 VSS 0.042814f
C10804 MULT_0.NAND2_2.Y.t10 VSS 0.042814f
C10805 MULT_0.NAND2_2.Y.n5 VSS 0.139748f
C10806 MULT_0.NAND2_2.Y.t7 VSS 0.048883f
C10807 B0.t51 VSS 0.042753f
C10808 B0.t31 VSS 0.059679f
C10809 B0.t30 VSS 0.059679f
C10810 B0.n0 VSS 0.194271f
C10811 B0.t14 VSS 0.068485f
C10812 B0.n1 VSS 0.596485f
C10813 B0.t39 VSS 0.042753f
C10814 B0.t44 VSS 0.059679f
C10815 B0.t43 VSS 0.059679f
C10816 B0.n2 VSS 0.194271f
C10817 B0.t28 VSS 0.068485f
C10818 B0.n3 VSS 0.480215f
C10819 B0.n4 VSS 0.553191f
C10820 B0.t27 VSS 0.042753f
C10821 B0.t49 VSS 0.059679f
C10822 B0.t23 VSS 0.059679f
C10823 B0.n5 VSS 0.194271f
C10824 B0.t7 VSS 0.068485f
C10825 B0.n6 VSS 0.481576f
C10826 B0.n7 VSS 0.428f
C10827 B0.n8 VSS 3.52829f
C10828 B0.t52 VSS 0.056946f
C10829 B0.t1 VSS 0.114578f
C10830 B0.t25 VSS 0.113153f
C10831 B0.t18 VSS 0.113153f
C10832 B0.t47 VSS 0.113153f
C10833 B0.t4 VSS 0.023514f
C10834 B0.t38 VSS 0.023514f
C10835 B0.t15 VSS 0.023514f
C10836 B0.n9 VSS 0.69712f
C10837 B0.n10 VSS 0.513461f
C10838 B0.n11 VSS 0.279832f
C10839 B0.n12 VSS 0.274911f
C10840 B0.n13 VSS 0.169102f
C10841 B0.n14 VSS 0.192303f
C10842 B0.t41 VSS 0.124724f
C10843 B0.t22 VSS 0.040615f
C10844 B0.t17 VSS 0.056088f
C10845 B0.n15 VSS 0.060484f
C10846 B0.t37 VSS 0.041756f
C10847 B0.n16 VSS 0.105949f
C10848 B0.n17 VSS 0.186185f
C10849 B0.t19 VSS 0.124724f
C10850 B0.t0 VSS 0.040615f
C10851 B0.t48 VSS 0.056088f
C10852 B0.n18 VSS 0.060484f
C10853 B0.t16 VSS 0.041756f
C10854 B0.n19 VSS 0.105949f
C10855 B0.n20 VSS 0.186182f
C10856 B0.n21 VSS 4.9132f
C10857 B0.t46 VSS 0.124724f
C10858 B0.t24 VSS 0.040615f
C10859 B0.t20 VSS 0.056088f
C10860 B0.n22 VSS 0.060484f
C10861 B0.t42 VSS 0.041756f
C10862 B0.n23 VSS 0.105949f
C10863 B0.n24 VSS 0.186189f
C10864 B0.n25 VSS 3.67188f
C10865 B0.t2 VSS 0.124724f
C10866 B0.t33 VSS 0.040615f
C10867 B0.t10 VSS 0.056088f
C10868 B0.n26 VSS 0.060484f
C10869 B0.t34 VSS 0.041756f
C10870 B0.n27 VSS 0.105949f
C10871 B0.n28 VSS 0.186176f
C10872 B0.n29 VSS 0.804802f
C10873 B0.n30 VSS 19.910698f
C10874 B0.t53 VSS 0.124867f
C10875 B0.t21 VSS 0.053477f
C10876 B0.t36 VSS 0.042753f
C10877 B0.n31 VSS 0.063096f
C10878 B0.t40 VSS 0.041756f
C10879 B0.n32 VSS 0.104161f
C10880 B0.n33 VSS 0.185832f
C10881 B0.n34 VSS 0.273969f
C10882 B0.n35 VSS 2.4511f
C10883 B0.t5 VSS 0.051018f
C10884 B0.t3 VSS 0.054724f
C10885 B0.n36 VSS 0.081544f
C10886 B0.t6 VSS 0.051018f
C10887 B0.t26 VSS 0.051018f
C10888 B0.t29 VSS 0.051018f
C10889 B0.t45 VSS 0.064454f
C10890 B0.n37 VSS 0.13771f
C10891 B0.n38 VSS 0.086703f
C10892 B0.n39 VSS 0.070846f
C10893 B0.n40 VSS 0.034667f
C10894 B0.n41 VSS 0.241588f
C10895 B0.n42 VSS 4.22548f
C10896 B0.t35 VSS 0.056946f
C10897 B0.t11 VSS 0.114578f
C10898 B0.t13 VSS 0.113153f
C10899 B0.t9 VSS 0.113153f
C10900 B0.t50 VSS 0.113153f
C10901 B0.t8 VSS 0.023514f
C10902 B0.t32 VSS 0.023514f
C10903 B0.t12 VSS 0.023514f
C10904 B0.n43 VSS 0.696945f
C10905 B0.n44 VSS 0.513637f
C10906 B0.n45 VSS 0.279832f
C10907 B0.n46 VSS 0.274911f
C10908 B0.n47 VSS 0.169102f
C10909 B0.n48 VSS 0.217601f
C10910 B0.n49 VSS 3.31197f
C10911 B0.n50 VSS 3.2224f
C10912 OR8_0.S5.n0 VSS 3.30271f
C10913 mux8_7.NAND4F_2.A VSS 2.54837f
C10914 OR8_0.S5.t5 VSS 0.159756f
C10915 OR8_0.S5.t6 VSS 0.155431f
C10916 OR8_0.S5.t4 VSS 0.470686f
C10917 OR8_0.S5.n1 VSS 0.801358f
C10918 mux8_7.A3 VSS 17.1499f
C10919 OR8_0.S5.t2 VSS 0.076582f
C10920 OR8_0.S5.t3 VSS 0.076582f
C10921 OR8_0.S5.n2 VSS 0.170658f
C10922 OR8_0.S5.t1 VSS 0.277763f
C10923 OR8_0.S5.t0 VSS 0.220888f
C10924 OR8_0.NOT8_0.S5 VSS 12.4893f
C10925 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t18 VSS 0.013766f
C10926 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t22 VSS 0.027698f
C10927 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t23 VSS 0.027354f
C10928 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t19 VSS 0.027354f
C10929 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t21 VSS 0.027354f
C10930 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t15 VSS 0.005684f
C10931 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t17 VSS 0.005684f
C10932 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t20 VSS 0.005684f
C10933 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n0 VSS 0.168523f
C10934 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n1 VSS 0.124125f
C10935 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n2 VSS 0.067647f
C10936 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n3 VSS 0.066457f
C10937 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n4 VSS 0.040879f
C10938 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n5 VSS 0.05311f
C10939 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t16 VSS 0.030151f
C10940 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t12 VSS 0.009818f
C10941 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t13 VSS 0.013559f
C10942 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n6 VSS 0.014622f
C10943 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t14 VSS 0.010094f
C10944 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n7 VSS 0.025612f
C10945 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n8 VSS 0.044927f
C10946 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t11 VSS 0.004926f
C10947 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t10 VSS 0.004926f
C10948 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n9 VSS 0.011915f
C10949 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t3 VSS 0.004926f
C10950 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t4 VSS 0.004926f
C10951 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n10 VSS 0.011914f
C10952 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n11 VSS 0.085433f
C10953 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t9 VSS 0.004926f
C10954 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t5 VSS 0.004926f
C10955 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n12 VSS 0.009853f
C10956 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n13 VSS 0.00774f
C10957 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t8 VSS 0.020843f
C10958 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t2 VSS 0.020843f
C10959 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n14 VSS 0.041685f
C10960 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n15 VSS 0.016575f
C10961 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t7 VSS 0.020843f
C10962 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t6 VSS 0.020843f
C10963 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n16 VSS 0.041685f
C10964 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n17 VSS 0.018334f
C10965 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n18 VSS 0.188757f
C10966 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t0 VSS 0.020843f
C10967 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.t1 VSS 0.020843f
C10968 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n19 VSS 0.041685f
C10969 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n20 VSS 0.018362f
C10970 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n21 VSS 0.12106f
C10971 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n22 VSS 0.027282f
C10972 8bit_ADDER_0.FULL_ADDER_XORED_7.XOR2_1.A.n23 VSS 0.119748f
C10973 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t15 VSS 0.013766f
C10974 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t17 VSS 0.027698f
C10975 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t20 VSS 0.027354f
C10976 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t22 VSS 0.027354f
C10977 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t21 VSS 0.027354f
C10978 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t14 VSS 0.005684f
C10979 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t19 VSS 0.005684f
C10980 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t18 VSS 0.005684f
C10981 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n0 VSS 0.168523f
C10982 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n1 VSS 0.124125f
C10983 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n2 VSS 0.067647f
C10984 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n3 VSS 0.066457f
C10985 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n4 VSS 0.040879f
C10986 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n5 VSS 0.05311f
C10987 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t13 VSS 0.030151f
C10988 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t12 VSS 0.009818f
C10989 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t16 VSS 0.013559f
C10990 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n6 VSS 0.014622f
C10991 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t23 VSS 0.010094f
C10992 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n7 VSS 0.025612f
C10993 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n8 VSS 0.044927f
C10994 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t8 VSS 0.004926f
C10995 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t7 VSS 0.004926f
C10996 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n9 VSS 0.011915f
C10997 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t3 VSS 0.004926f
C10998 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t2 VSS 0.004926f
C10999 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n10 VSS 0.011914f
C11000 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n11 VSS 0.085433f
C11001 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t0 VSS 0.004926f
C11002 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t6 VSS 0.004926f
C11003 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n12 VSS 0.009853f
C11004 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n13 VSS 0.00774f
C11005 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t9 VSS 0.020843f
C11006 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t1 VSS 0.020843f
C11007 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n14 VSS 0.041685f
C11008 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n15 VSS 0.016575f
C11009 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t11 VSS 0.020843f
C11010 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t10 VSS 0.020843f
C11011 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n16 VSS 0.041685f
C11012 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n17 VSS 0.018334f
C11013 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n18 VSS 0.188757f
C11014 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t5 VSS 0.020843f
C11015 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.t4 VSS 0.020843f
C11016 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n19 VSS 0.041685f
C11017 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n20 VSS 0.018362f
C11018 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n21 VSS 0.12106f
C11019 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n22 VSS 0.027282f
C11020 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_1.A.n23 VSS 0.119748f
C11021 V_FLAG_0.XOR2_2.Y.t13 VSS 0.027208f
C11022 V_FLAG_0.XOR2_2.Y.t12 VSS 0.010444f
C11023 V_FLAG_0.XOR2_2.Y.t15 VSS 0.014422f
C11024 V_FLAG_0.XOR2_2.Y.n0 VSS 0.0166f
C11025 V_FLAG_0.XOR2_2.Y.t14 VSS 0.010978f
C11026 V_FLAG_0.XOR2_2.Y.n1 VSS 0.016835f
C11027 V_FLAG_0.XOR2_2.Y.n2 VSS 0.062222f
C11028 V_FLAG_0.XOR2_2.Y.t2 VSS 0.00524f
C11029 V_FLAG_0.XOR2_2.Y.t1 VSS 0.00524f
C11030 V_FLAG_0.XOR2_2.Y.n3 VSS 0.012674f
C11031 V_FLAG_0.XOR2_2.Y.t7 VSS 0.00524f
C11032 V_FLAG_0.XOR2_2.Y.t10 VSS 0.00524f
C11033 V_FLAG_0.XOR2_2.Y.n4 VSS 0.012673f
C11034 V_FLAG_0.XOR2_2.Y.n5 VSS 0.090874f
C11035 V_FLAG_0.XOR2_2.Y.t0 VSS 0.00524f
C11036 V_FLAG_0.XOR2_2.Y.t11 VSS 0.00524f
C11037 V_FLAG_0.XOR2_2.Y.n6 VSS 0.01048f
C11038 V_FLAG_0.XOR2_2.Y.n7 VSS 0.008233f
C11039 V_FLAG_0.XOR2_2.Y.t4 VSS 0.02217f
C11040 V_FLAG_0.XOR2_2.Y.t8 VSS 0.02217f
C11041 V_FLAG_0.XOR2_2.Y.n8 VSS 0.04434f
C11042 V_FLAG_0.XOR2_2.Y.n9 VSS 0.01763f
C11043 V_FLAG_0.XOR2_2.Y.t5 VSS 0.02217f
C11044 V_FLAG_0.XOR2_2.Y.t3 VSS 0.02217f
C11045 V_FLAG_0.XOR2_2.Y.n10 VSS 0.04434f
C11046 V_FLAG_0.XOR2_2.Y.n11 VSS 0.019501f
C11047 V_FLAG_0.XOR2_2.Y.n12 VSS 0.200779f
C11048 V_FLAG_0.XOR2_2.Y.t9 VSS 0.02217f
C11049 V_FLAG_0.XOR2_2.Y.t6 VSS 0.02217f
C11050 V_FLAG_0.XOR2_2.Y.n13 VSS 0.04434f
C11051 V_FLAG_0.XOR2_2.Y.n14 VSS 0.019531f
C11052 V_FLAG_0.XOR2_2.Y.n15 VSS 0.128771f
C11053 V_FLAG_0.XOR2_2.Y.n16 VSS 0.02902f
C11054 V_FLAG_0.XOR2_2.Y.n17 VSS 0.127428f
C11055 a_n14077_3810.n0 VSS 1.45527f
C11056 a_n14077_3810.n1 VSS 1.45566f
C11057 a_n14077_3810.t0 VSS 0.09158f
C11058 a_n14077_3810.t4 VSS 0.09158f
C11059 a_n14077_3810.t5 VSS 0.09158f
C11060 a_n14077_3810.n2 VSS 0.198865f
C11061 a_n14077_3810.t3 VSS 0.09158f
C11062 a_n14077_3810.t10 VSS 0.09158f
C11063 a_n14077_3810.n3 VSS 0.19819f
C11064 a_n14077_3810.t11 VSS 0.09158f
C11065 a_n14077_3810.t9 VSS 0.09158f
C11066 a_n14077_3810.n4 VSS 0.19819f
C11067 a_n14077_3810.t7 VSS 0.09158f
C11068 a_n14077_3810.t6 VSS 0.09158f
C11069 a_n14077_3810.n5 VSS 0.19819f
C11070 a_n14077_3810.t8 VSS 0.09158f
C11071 a_n14077_3810.t1 VSS 0.09158f
C11072 a_n14077_3810.n6 VSS 0.19819f
C11073 a_n14077_3810.n7 VSS 0.198479f
C11074 a_n14077_3810.t2 VSS 0.09158f
C11075 mux8_4.NAND4F_4.B.n0 VSS 0.921489f
C11076 mux8_4.NAND4F_4.B.t9 VSS 0.03989f
C11077 mux8_4.NAND4F_4.B.t10 VSS 0.123086f
C11078 mux8_4.NAND4F_4.B.t7 VSS 0.04595f
C11079 mux8_4.NAND4F_4.B.n1 VSS 0.154452f
C11080 mux8_4.NAND4F_4.B.n2 VSS 0.033769f
C11081 mux8_4.NAND4F_4.B.t8 VSS 0.03989f
C11082 mux8_4.NAND4F_4.B.t4 VSS 0.123086f
C11083 mux8_4.NAND4F_4.B.t5 VSS 0.04595f
C11084 mux8_4.NAND4F_4.B.n3 VSS 0.154452f
C11085 mux8_4.NAND4F_4.B.n4 VSS 0.032977f
C11086 mux8_4.NAND4F_4.B.t14 VSS 0.03989f
C11087 mux8_4.NAND4F_4.B.t11 VSS 0.123086f
C11088 mux8_4.NAND4F_4.B.t12 VSS 0.04595f
C11089 mux8_4.NAND4F_4.B.n5 VSS 0.154452f
C11090 mux8_4.NAND4F_4.B.n6 VSS 0.033699f
C11091 mux8_4.NAND4F_4.B.n7 VSS 0.612655f
C11092 mux8_4.NAND4F_4.B.t3 VSS 0.020325f
C11093 mux8_4.NAND4F_4.B.t2 VSS 0.020325f
C11094 mux8_4.NAND4F_4.B.n8 VSS 0.045293f
C11095 mux8_4.NAND4F_4.B.t1 VSS 0.073718f
C11096 mux8_4.NAND4F_4.B.t0 VSS 0.058624f
C11097 mux8_4.NAND4F_4.B.n9 VSS 0.607515f
C11098 mux8_4.NAND4F_4.B.t15 VSS 0.03989f
C11099 mux8_4.NAND4F_4.B.t6 VSS 0.123086f
C11100 mux8_4.NAND4F_4.B.t13 VSS 0.04595f
C11101 mux8_4.NAND4F_4.B.n10 VSS 0.154452f
C11102 mux8_4.NAND4F_4.B.n11 VSS 0.033659f
C11103 mux8_4.NAND4F_4.B.n12 VSS 0.776456f
C11104 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t12 VSS 0.013766f
C11105 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t19 VSS 0.027698f
C11106 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t21 VSS 0.027354f
C11107 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t16 VSS 0.027354f
C11108 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t18 VSS 0.027354f
C11109 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t23 VSS 0.005684f
C11110 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t20 VSS 0.005684f
C11111 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t17 VSS 0.005684f
C11112 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n0 VSS 0.168523f
C11113 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n1 VSS 0.124125f
C11114 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n2 VSS 0.067647f
C11115 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n3 VSS 0.066457f
C11116 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n4 VSS 0.040879f
C11117 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n5 VSS 0.05311f
C11118 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t22 VSS 0.030151f
C11119 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t15 VSS 0.009818f
C11120 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t13 VSS 0.013559f
C11121 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n6 VSS 0.014622f
C11122 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t14 VSS 0.010094f
C11123 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n7 VSS 0.025612f
C11124 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n8 VSS 0.044927f
C11125 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t9 VSS 0.004926f
C11126 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t10 VSS 0.004926f
C11127 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n9 VSS 0.011915f
C11128 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t3 VSS 0.004926f
C11129 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t4 VSS 0.004926f
C11130 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n10 VSS 0.011914f
C11131 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n11 VSS 0.085433f
C11132 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t11 VSS 0.004926f
C11133 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t5 VSS 0.004926f
C11134 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n12 VSS 0.009853f
C11135 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n13 VSS 0.00774f
C11136 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t1 VSS 0.020843f
C11137 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t7 VSS 0.020843f
C11138 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n14 VSS 0.041685f
C11139 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n15 VSS 0.016575f
C11140 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t0 VSS 0.020843f
C11141 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t2 VSS 0.020843f
C11142 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n16 VSS 0.041685f
C11143 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n17 VSS 0.018334f
C11144 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n18 VSS 0.188757f
C11145 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t8 VSS 0.020843f
C11146 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.t6 VSS 0.020843f
C11147 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n19 VSS 0.041685f
C11148 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n20 VSS 0.018362f
C11149 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n21 VSS 0.12106f
C11150 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n22 VSS 0.027282f
C11151 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_1.A.n23 VSS 0.119748f
C11152 mux8_8.NAND4F_6.Y.n0 VSS 0.599344f
C11153 mux8_8.NAND4F_6.Y.t2 VSS 0.244548f
C11154 mux8_8.NAND4F_6.Y.t9 VSS 0.038543f
C11155 mux8_8.NAND4F_6.Y.t10 VSS 0.118929f
C11156 mux8_8.NAND4F_6.Y.t11 VSS 0.044398f
C11157 mux8_8.NAND4F_6.Y.n1 VSS 0.149236f
C11158 mux8_8.NAND4F_6.Y.n2 VSS 0.032396f
C11159 mux8_8.NAND4F_6.Y.n3 VSS 1.72835f
C11160 mux8_8.NAND4F_6.Y.t1 VSS 0.029549f
C11161 mux8_8.NAND4F_6.Y.t0 VSS 0.029549f
C11162 mux8_8.NAND4F_6.Y.n4 VSS 0.068617f
C11163 mux8_8.NAND4F_6.Y.t6 VSS 0.029549f
C11164 mux8_8.NAND4F_6.Y.t5 VSS 0.029549f
C11165 mux8_8.NAND4F_6.Y.n5 VSS 0.068411f
C11166 mux8_8.NAND4F_6.Y.t8 VSS 0.029549f
C11167 mux8_8.NAND4F_6.Y.t7 VSS 0.029549f
C11168 mux8_8.NAND4F_6.Y.n6 VSS 0.068411f
C11169 mux8_8.NAND4F_6.Y.t3 VSS 0.029549f
C11170 mux8_8.NAND4F_6.Y.t4 VSS 0.029549f
C11171 mux8_8.NAND4F_6.Y.n7 VSS 0.068411f
C11172 mux8_8.NAND4F_6.Y.n8 VSS 0.281208f
C11173 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n0 VSS 0.967969f
C11174 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t2 VSS 0.008375f
C11175 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t3 VSS 0.008375f
C11176 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n1 VSS 0.018687f
C11177 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t6 VSS 0.008375f
C11178 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t4 VSS 0.008375f
C11179 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n2 VSS 0.018636f
C11180 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t1 VSS 0.008375f
C11181 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t5 VSS 0.008375f
C11182 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n3 VSS 0.018636f
C11183 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t0 VSS 0.05057f
C11184 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t13 VSS 0.028606f
C11185 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t9 VSS 0.02825f
C11186 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t10 VSS 0.02825f
C11187 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t18 VSS 0.02825f
C11188 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n4 VSS 0.112442f
C11189 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t8 VSS 0.005871f
C11190 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t14 VSS 0.005871f
C11191 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t11 VSS 0.005871f
C11192 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t7 VSS 0.005871f
C11193 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n5 VSS 0.106225f
C11194 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n6 VSS 0.166131f
C11195 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t12 VSS 0.026417f
C11196 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t17 VSS 0.01014f
C11197 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t15 VSS 0.014003f
C11198 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n7 VSS 0.016118f
C11199 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.t16 VSS 0.010659f
C11200 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n8 VSS 0.016345f
C11201 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n9 VSS 0.055518f
C11202 MULT_0.4bit_ADDER_0.FULL_ADDER_1.COUT.n10 VSS 0.369194f
C11203 mux8_1.NAND4F_9.Y.n0 VSS 0.358256f
C11204 mux8_1.NAND4F_9.Y.t9 VSS 0.017853f
C11205 mux8_1.NAND4F_9.Y.t10 VSS 0.017853f
C11206 mux8_1.NAND4F_9.Y.t11 VSS 0.017853f
C11207 mux8_1.NAND4F_9.Y.t12 VSS 0.017853f
C11208 mux8_1.NAND4F_9.Y.t13 VSS 0.022554f
C11209 mux8_1.NAND4F_9.Y.n1 VSS 0.048188f
C11210 mux8_1.NAND4F_9.Y.n2 VSS 0.030339f
C11211 mux8_1.NAND4F_9.Y.n3 VSS 0.030339f
C11212 mux8_1.NAND4F_9.Y.n4 VSS 0.026149f
C11213 mux8_1.NAND4F_9.Y.t14 VSS 0.014813f
C11214 mux8_1.NAND4F_9.Y.n5 VSS 0.021261f
C11215 mux8_1.NAND4F_9.Y.t4 VSS 0.141821f
C11216 mux8_1.NAND4F_9.Y.t7 VSS 0.017663f
C11217 mux8_1.NAND4F_9.Y.t8 VSS 0.017663f
C11218 mux8_1.NAND4F_9.Y.n6 VSS 0.041015f
C11219 mux8_1.NAND4F_9.Y.t5 VSS 0.017663f
C11220 mux8_1.NAND4F_9.Y.t6 VSS 0.017663f
C11221 mux8_1.NAND4F_9.Y.n7 VSS 0.040893f
C11222 mux8_1.NAND4F_9.Y.t0 VSS 0.017663f
C11223 mux8_1.NAND4F_9.Y.t1 VSS 0.017663f
C11224 mux8_1.NAND4F_9.Y.n8 VSS 0.040893f
C11225 mux8_1.NAND4F_9.Y.t3 VSS 0.017663f
C11226 mux8_1.NAND4F_9.Y.t2 VSS 0.017663f
C11227 mux8_1.NAND4F_9.Y.n9 VSS 0.040893f
C11228 mux8_1.NAND4F_9.Y.n10 VSS 0.168091f
C11229 mux8_1.NAND4F_7.Y.n0 VSS 0.11858f
C11230 mux8_1.NAND4F_7.Y.n1 VSS 0.350455f
C11231 mux8_1.NAND4F_7.Y.t5 VSS 0.168166f
C11232 mux8_1.NAND4F_7.Y.t9 VSS 0.022537f
C11233 mux8_1.NAND4F_7.Y.t10 VSS 0.079785f
C11234 mux8_1.NAND4F_7.Y.t11 VSS 0.024808f
C11235 mux8_1.NAND4F_7.Y.n2 VSS 0.070768f
C11236 mux8_1.NAND4F_7.Y.n3 VSS 0.020978f
C11237 mux8_1.NAND4F_7.Y.t0 VSS 0.017278f
C11238 mux8_1.NAND4F_7.Y.t1 VSS 0.017278f
C11239 mux8_1.NAND4F_7.Y.n4 VSS 0.040122f
C11240 mux8_1.NAND4F_7.Y.t3 VSS 0.017278f
C11241 mux8_1.NAND4F_7.Y.t2 VSS 0.017278f
C11242 mux8_1.NAND4F_7.Y.n5 VSS 0.040002f
C11243 mux8_1.NAND4F_7.Y.t8 VSS 0.017278f
C11244 mux8_1.NAND4F_7.Y.t7 VSS 0.017278f
C11245 mux8_1.NAND4F_7.Y.n6 VSS 0.040002f
C11246 mux8_1.NAND4F_7.Y.t6 VSS 0.017278f
C11247 mux8_1.NAND4F_7.Y.t4 VSS 0.017278f
C11248 mux8_1.NAND4F_7.Y.n7 VSS 0.040002f
C11249 mux8_1.NAND4F_1.Y.n0 VSS 0.655599f
C11250 mux8_1.NAND4F_1.Y.t4 VSS 0.306614f
C11251 mux8_1.NAND4F_1.Y.t9 VSS 0.132168f
C11252 mux8_1.NAND4F_1.Y.t10 VSS 0.04216f
C11253 mux8_1.NAND4F_1.Y.t11 VSS 0.04216f
C11254 mux8_1.NAND4F_1.Y.n1 VSS 0.049498f
C11255 mux8_1.NAND4F_1.Y.n2 VSS 0.277534f
C11256 mux8_1.NAND4F_1.Y.t0 VSS 0.032323f
C11257 mux8_1.NAND4F_1.Y.t1 VSS 0.032323f
C11258 mux8_1.NAND4F_1.Y.n3 VSS 0.075057f
C11259 mux8_1.NAND4F_1.Y.t3 VSS 0.032323f
C11260 mux8_1.NAND4F_1.Y.t2 VSS 0.032323f
C11261 mux8_1.NAND4F_1.Y.n4 VSS 0.074832f
C11262 mux8_1.NAND4F_1.Y.t7 VSS 0.032323f
C11263 mux8_1.NAND4F_1.Y.t8 VSS 0.032323f
C11264 mux8_1.NAND4F_1.Y.n5 VSS 0.074832f
C11265 mux8_1.NAND4F_1.Y.t5 VSS 0.032323f
C11266 mux8_1.NAND4F_1.Y.t6 VSS 0.032323f
C11267 mux8_1.NAND4F_1.Y.n6 VSS 0.074832f
C11268 mux8_1.NAND4F_1.Y.n7 VSS 0.307603f
C11269 mux8_1.NAND4F_4.B.n0 VSS 0.921489f
C11270 mux8_1.NAND4F_4.B.t10 VSS 0.03989f
C11271 mux8_1.NAND4F_4.B.t14 VSS 0.123086f
C11272 mux8_1.NAND4F_4.B.t12 VSS 0.04595f
C11273 mux8_1.NAND4F_4.B.n1 VSS 0.154452f
C11274 mux8_1.NAND4F_4.B.n2 VSS 0.033769f
C11275 mux8_1.NAND4F_4.B.t9 VSS 0.03989f
C11276 mux8_1.NAND4F_4.B.t8 VSS 0.123086f
C11277 mux8_1.NAND4F_4.B.t11 VSS 0.04595f
C11278 mux8_1.NAND4F_4.B.n3 VSS 0.154452f
C11279 mux8_1.NAND4F_4.B.n4 VSS 0.032977f
C11280 mux8_1.NAND4F_4.B.t15 VSS 0.03989f
C11281 mux8_1.NAND4F_4.B.t7 VSS 0.123086f
C11282 mux8_1.NAND4F_4.B.t5 VSS 0.04595f
C11283 mux8_1.NAND4F_4.B.n5 VSS 0.154452f
C11284 mux8_1.NAND4F_4.B.n6 VSS 0.033699f
C11285 mux8_1.NAND4F_4.B.n7 VSS 0.612655f
C11286 mux8_1.NAND4F_4.B.t1 VSS 0.020325f
C11287 mux8_1.NAND4F_4.B.t3 VSS 0.020325f
C11288 mux8_1.NAND4F_4.B.n8 VSS 0.045293f
C11289 mux8_1.NAND4F_4.B.t2 VSS 0.073718f
C11290 mux8_1.NAND4F_4.B.t0 VSS 0.058624f
C11291 mux8_1.NAND4F_4.B.n9 VSS 0.607515f
C11292 mux8_1.NAND4F_4.B.t4 VSS 0.03989f
C11293 mux8_1.NAND4F_4.B.t13 VSS 0.123086f
C11294 mux8_1.NAND4F_4.B.t6 VSS 0.04595f
C11295 mux8_1.NAND4F_4.B.n10 VSS 0.154452f
C11296 mux8_1.NAND4F_4.B.n11 VSS 0.033659f
C11297 mux8_1.NAND4F_4.B.n12 VSS 0.776456f
C11298 a_n12314_n18115.n0 VSS 1.48365f
C11299 a_n12314_n18115.n1 VSS 1.48326f
C11300 a_n12314_n18115.t1 VSS 0.093341f
C11301 a_n12314_n18115.t6 VSS 0.093341f
C11302 a_n12314_n18115.t8 VSS 0.093341f
C11303 a_n12314_n18115.n2 VSS 0.202296f
C11304 a_n12314_n18115.t7 VSS 0.093341f
C11305 a_n12314_n18115.t3 VSS 0.093341f
C11306 a_n12314_n18115.n3 VSS 0.202001f
C11307 a_n12314_n18115.t4 VSS 0.093341f
C11308 a_n12314_n18115.t5 VSS 0.093341f
C11309 a_n12314_n18115.n4 VSS 0.202001f
C11310 a_n12314_n18115.t9 VSS 0.093341f
C11311 a_n12314_n18115.t10 VSS 0.093341f
C11312 a_n12314_n18115.n5 VSS 0.202001f
C11313 a_n12314_n18115.t11 VSS 0.093341f
C11314 a_n12314_n18115.t0 VSS 0.093341f
C11315 a_n12314_n18115.n6 VSS 0.202001f
C11316 a_n12314_n18115.n7 VSS 0.20269f
C11317 a_n12314_n18115.t2 VSS 0.093341f
C11318 B1.t7 VSS 0.049884f
C11319 B1.t12 VSS 0.069634f
C11320 B1.t11 VSS 0.069634f
C11321 B1.n0 VSS 0.226676f
C11322 B1.t47 VSS 0.079909f
C11323 B1.n1 VSS 0.551146f
C11324 B1.t48 VSS 0.066445f
C11325 B1.t53 VSS 0.13369f
C11326 B1.t28 VSS 0.132027f
C11327 B1.t18 VSS 0.132027f
C11328 B1.t4 VSS 0.132027f
C11329 B1.t49 VSS 0.027436f
C11330 B1.t31 VSS 0.027436f
C11331 B1.t24 VSS 0.027436f
C11332 B1.n2 VSS 0.813405f
C11333 B1.n3 VSS 0.59911f
C11334 B1.n4 VSS 0.32651f
C11335 B1.n5 VSS 0.320768f
C11336 B1.n6 VSS 0.197309f
C11337 B1.n7 VSS 0.224381f
C11338 B1.t40 VSS 0.123461f
C11339 B1.t42 VSS 0.04739f
C11340 B1.t37 VSS 0.065444f
C11341 B1.n8 VSS 0.075326f
C11342 B1.t6 VSS 0.049813f
C11343 B1.n9 VSS 0.076391f
C11344 B1.n10 VSS 0.31699f
C11345 B1.t43 VSS 0.145529f
C11346 B1.t36 VSS 0.04739f
C11347 B1.t30 VSS 0.065444f
C11348 B1.n11 VSS 0.070574f
C11349 B1.t39 VSS 0.048721f
C11350 B1.n12 VSS 0.123623f
C11351 B1.n13 VSS 0.217247f
C11352 B1.n14 VSS 1.53889f
C11353 B1.t9 VSS 0.123461f
C11354 B1.t33 VSS 0.04739f
C11355 B1.t14 VSS 0.065444f
C11356 B1.n15 VSS 0.075326f
C11357 B1.t32 VSS 0.049813f
C11358 B1.n16 VSS 0.076391f
C11359 B1.n17 VSS 0.31699f
C11360 B1.t15 VSS 0.145529f
C11361 B1.t25 VSS 0.04739f
C11362 B1.t3 VSS 0.065444f
C11363 B1.n18 VSS 0.070574f
C11364 B1.t27 VSS 0.048721f
C11365 B1.n19 VSS 0.123623f
C11366 B1.n20 VSS 0.217231f
C11367 B1.n21 VSS 0.957704f
C11368 B1.n22 VSS 2.21734f
C11369 B1.n23 VSS 23.1583f
C11370 B1.t10 VSS 0.145696f
C11371 B1.t35 VSS 0.062397f
C11372 B1.t38 VSS 0.049884f
C11373 B1.n24 VSS 0.073621f
C11374 B1.t2 VSS 0.048721f
C11375 B1.n25 VSS 0.121535f
C11376 B1.n26 VSS 0.21683f
C11377 B1.n27 VSS 0.317894f
C11378 B1.n28 VSS 2.86066f
C11379 B1.t46 VSS 0.059529f
C11380 B1.t45 VSS 0.063852f
C11381 B1.n29 VSS 0.095146f
C11382 B1.t50 VSS 0.059529f
C11383 B1.t13 VSS 0.059529f
C11384 B1.t16 VSS 0.059529f
C11385 B1.t34 VSS 0.075205f
C11386 B1.n30 VSS 0.160682f
C11387 B1.n31 VSS 0.101166f
C11388 B1.n32 VSS 0.082664f
C11389 B1.n33 VSS 0.04045f
C11390 B1.n34 VSS 5.583f
C11391 B1.t26 VSS 0.066445f
C11392 B1.t1 VSS 0.13369f
C11393 B1.t21 VSS 0.132027f
C11394 B1.t0 VSS 0.132027f
C11395 B1.t51 VSS 0.132027f
C11396 B1.t52 VSS 0.027436f
C11397 B1.t22 VSS 0.027436f
C11398 B1.t19 VSS 0.027436f
C11399 B1.n35 VSS 0.8132f
C11400 B1.n36 VSS 0.599315f
C11401 B1.n37 VSS 0.32651f
C11402 B1.n38 VSS 0.320768f
C11403 B1.n39 VSS 0.197309f
C11404 B1.n40 VSS 0.253899f
C11405 B1.n41 VSS 5.32155f
C11406 B1.t23 VSS 0.049884f
C11407 B1.t20 VSS 0.069634f
C11408 B1.t17 VSS 0.069634f
C11409 B1.n42 VSS 0.226676f
C11410 B1.t41 VSS 0.079909f
C11411 B1.n43 VSS 0.673679f
C11412 B1.n44 VSS 4.39263f
C11413 B1.t8 VSS 0.049884f
C11414 B1.t29 VSS 0.069634f
C11415 B1.t5 VSS 0.069634f
C11416 B1.n45 VSS 0.226676f
C11417 B1.t44 VSS 0.079909f
C11418 B1.n46 VSS 0.546091f
C11419 B1.n47 VSS 0.476566f
C11420 B1.n48 VSS 3.96024f
C11421 B1.n49 VSS 0.631599f
C11422 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n0 VSS 0.887305f
C11423 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t2 VSS 0.007677f
C11424 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t0 VSS 0.007677f
C11425 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n1 VSS 0.01713f
C11426 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t6 VSS 0.007677f
C11427 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t1 VSS 0.007677f
C11428 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n2 VSS 0.017083f
C11429 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t4 VSS 0.007677f
C11430 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t3 VSS 0.007677f
C11431 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n3 VSS 0.017083f
C11432 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t5 VSS 0.046356f
C11433 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t15 VSS 0.026222f
C11434 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t14 VSS 0.025896f
C11435 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t12 VSS 0.025896f
C11436 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t13 VSS 0.025896f
C11437 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n4 VSS 0.103072f
C11438 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t8 VSS 0.005381f
C11439 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t9 VSS 0.005381f
C11440 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t11 VSS 0.005381f
C11441 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t10 VSS 0.005381f
C11442 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n5 VSS 0.097373f
C11443 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n6 VSS 0.152286f
C11444 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t7 VSS 0.024216f
C11445 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t16 VSS 0.009295f
C11446 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t17 VSS 0.012836f
C11447 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n7 VSS 0.014774f
C11448 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.t18 VSS 0.00977f
C11449 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n8 VSS 0.014983f
C11450 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n9 VSS 0.050891f
C11451 MULT_0.4bit_ADDER_2.FULL_ADDER_1.COUT.n10 VSS 0.338427f
C11452 mux8_4.NAND4F_9.Y.n0 VSS 0.358256f
C11453 mux8_4.NAND4F_9.Y.t10 VSS 0.017853f
C11454 mux8_4.NAND4F_9.Y.t9 VSS 0.017853f
C11455 mux8_4.NAND4F_9.Y.t14 VSS 0.017853f
C11456 mux8_4.NAND4F_9.Y.t13 VSS 0.017853f
C11457 mux8_4.NAND4F_9.Y.t11 VSS 0.022554f
C11458 mux8_4.NAND4F_9.Y.n1 VSS 0.048188f
C11459 mux8_4.NAND4F_9.Y.n2 VSS 0.030339f
C11460 mux8_4.NAND4F_9.Y.n3 VSS 0.030339f
C11461 mux8_4.NAND4F_9.Y.n4 VSS 0.026149f
C11462 mux8_4.NAND4F_9.Y.t12 VSS 0.014813f
C11463 mux8_4.NAND4F_9.Y.n5 VSS 0.021261f
C11464 mux8_4.NAND4F_9.Y.t0 VSS 0.141821f
C11465 mux8_4.NAND4F_9.Y.t5 VSS 0.017663f
C11466 mux8_4.NAND4F_9.Y.t6 VSS 0.017663f
C11467 mux8_4.NAND4F_9.Y.n6 VSS 0.041015f
C11468 mux8_4.NAND4F_9.Y.t7 VSS 0.017663f
C11469 mux8_4.NAND4F_9.Y.t8 VSS 0.017663f
C11470 mux8_4.NAND4F_9.Y.n7 VSS 0.040893f
C11471 mux8_4.NAND4F_9.Y.t3 VSS 0.017663f
C11472 mux8_4.NAND4F_9.Y.t4 VSS 0.017663f
C11473 mux8_4.NAND4F_9.Y.n8 VSS 0.040893f
C11474 mux8_4.NAND4F_9.Y.t2 VSS 0.017663f
C11475 mux8_4.NAND4F_9.Y.t1 VSS 0.017663f
C11476 mux8_4.NAND4F_9.Y.n9 VSS 0.040893f
C11477 mux8_4.NAND4F_9.Y.n10 VSS 0.168091f
C11478 mux8_4.NAND4F_6.Y.n0 VSS 0.599344f
C11479 mux8_4.NAND4F_6.Y.t2 VSS 0.244548f
C11480 mux8_4.NAND4F_6.Y.t9 VSS 0.038543f
C11481 mux8_4.NAND4F_6.Y.t10 VSS 0.118929f
C11482 mux8_4.NAND4F_6.Y.t11 VSS 0.044398f
C11483 mux8_4.NAND4F_6.Y.n1 VSS 0.149236f
C11484 mux8_4.NAND4F_6.Y.n2 VSS 0.032396f
C11485 mux8_4.NAND4F_6.Y.n3 VSS 1.72835f
C11486 mux8_4.NAND4F_6.Y.t1 VSS 0.029549f
C11487 mux8_4.NAND4F_6.Y.t0 VSS 0.029549f
C11488 mux8_4.NAND4F_6.Y.n4 VSS 0.068617f
C11489 mux8_4.NAND4F_6.Y.t6 VSS 0.029549f
C11490 mux8_4.NAND4F_6.Y.t5 VSS 0.029549f
C11491 mux8_4.NAND4F_6.Y.n5 VSS 0.068411f
C11492 mux8_4.NAND4F_6.Y.t7 VSS 0.029549f
C11493 mux8_4.NAND4F_6.Y.t8 VSS 0.029549f
C11494 mux8_4.NAND4F_6.Y.n6 VSS 0.068411f
C11495 mux8_4.NAND4F_6.Y.t3 VSS 0.029549f
C11496 mux8_4.NAND4F_6.Y.t4 VSS 0.029549f
C11497 mux8_4.NAND4F_6.Y.n7 VSS 0.068411f
C11498 mux8_4.NAND4F_6.Y.n8 VSS 0.281208f
C11499 mux8_5.NAND4F_7.Y.n0 VSS 0.11858f
C11500 mux8_5.NAND4F_7.Y.n1 VSS 0.350455f
C11501 mux8_5.NAND4F_7.Y.t4 VSS 0.168166f
C11502 mux8_5.NAND4F_7.Y.t9 VSS 0.022537f
C11503 mux8_5.NAND4F_7.Y.t11 VSS 0.079785f
C11504 mux8_5.NAND4F_7.Y.t10 VSS 0.024808f
C11505 mux8_5.NAND4F_7.Y.n2 VSS 0.070768f
C11506 mux8_5.NAND4F_7.Y.n3 VSS 0.020978f
C11507 mux8_5.NAND4F_7.Y.t1 VSS 0.017278f
C11508 mux8_5.NAND4F_7.Y.t0 VSS 0.017278f
C11509 mux8_5.NAND4F_7.Y.n4 VSS 0.040122f
C11510 mux8_5.NAND4F_7.Y.t3 VSS 0.017278f
C11511 mux8_5.NAND4F_7.Y.t2 VSS 0.017278f
C11512 mux8_5.NAND4F_7.Y.n5 VSS 0.040002f
C11513 mux8_5.NAND4F_7.Y.t8 VSS 0.017278f
C11514 mux8_5.NAND4F_7.Y.t7 VSS 0.017278f
C11515 mux8_5.NAND4F_7.Y.n6 VSS 0.040002f
C11516 mux8_5.NAND4F_7.Y.t5 VSS 0.017278f
C11517 mux8_5.NAND4F_7.Y.t6 VSS 0.017278f
C11518 mux8_5.NAND4F_7.Y.n7 VSS 0.040002f
C11519 NOT8_0.S4.n0 VSS 2.18109f
C11520 NOT8_0.S4.t6 VSS 0.105501f
C11521 NOT8_0.S4.t5 VSS 0.310838f
C11522 NOT8_0.S4.t4 VSS 0.102646f
C11523 NOT8_0.S4.n1 VSS 0.529212f
C11524 NOT8_0.S4.t3 VSS 0.050574f
C11525 NOT8_0.S4.t2 VSS 0.050574f
C11526 NOT8_0.S4.n2 VSS 0.112702f
C11527 NOT8_0.S4.t1 VSS 0.183433f
C11528 NOT8_0.S4.t0 VSS 0.145873f
C11529 SEL3.t57 VSS 0.011322f
C11530 SEL3.t29 VSS 0.011181f
C11531 SEL3.t50 VSS 0.011181f
C11532 SEL3.t11 VSS 0.011181f
C11533 SEL3.n0 VSS 0.044504f
C11534 SEL3.t15 VSS 0.002324f
C11535 SEL3.t61 VSS 0.002324f
C11536 SEL3.t18 VSS 0.002324f
C11537 SEL3.t81 VSS 0.002324f
C11538 SEL3.n1 VSS 0.042043f
C11539 SEL3.n2 VSS 0.065754f
C11540 SEL3.n3 VSS 0.134841f
C11541 SEL3.t19 VSS 0.010456f
C11542 SEL3.t31 VSS 0.004013f
C11543 SEL3.t36 VSS 0.005542f
C11544 SEL3.n4 VSS 0.006379f
C11545 SEL3.t23 VSS 0.004219f
C11546 SEL3.n5 VSS 0.006469f
C11547 SEL3.n6 VSS 0.021974f
C11548 SEL3.n7 VSS 0.055646f
C11549 SEL3.n8 VSS 0.146125f
C11550 SEL3.t10 VSS 0.011181f
C11551 SEL3.t37 VSS 0.011181f
C11552 SEL3.t80 VSS 0.011322f
C11553 SEL3.t56 VSS 0.011181f
C11554 SEL3.n9 VSS 0.044504f
C11555 SEL3.t72 VSS 0.002324f
C11556 SEL3.t48 VSS 0.002324f
C11557 SEL3.t2 VSS 0.002324f
C11558 SEL3.t25 VSS 0.002324f
C11559 SEL3.n10 VSS 0.042043f
C11560 SEL3.n11 VSS 0.065798f
C11561 SEL3.t13 VSS 0.011181f
C11562 SEL3.t42 VSS 0.011181f
C11563 SEL3.t0 VSS 0.011322f
C11564 SEL3.t58 VSS 0.011181f
C11565 SEL3.n12 VSS 0.044504f
C11566 SEL3.t73 VSS 0.002324f
C11567 SEL3.t51 VSS 0.002324f
C11568 SEL3.t7 VSS 0.002324f
C11569 SEL3.t30 VSS 0.002324f
C11570 SEL3.n13 VSS 0.042043f
C11571 SEL3.n14 VSS 0.065798f
C11572 SEL3.t43 VSS 0.011181f
C11573 SEL3.t9 VSS 0.011181f
C11574 SEL3.t74 VSS 0.011322f
C11575 SEL3.t52 VSS 0.011181f
C11576 SEL3.n15 VSS 0.044504f
C11577 SEL3.t64 VSS 0.002324f
C11578 SEL3.t44 VSS 0.002324f
C11579 SEL3.t32 VSS 0.002324f
C11580 SEL3.t1 VSS 0.002324f
C11581 SEL3.n16 VSS 0.042043f
C11582 SEL3.n17 VSS 0.065798f
C11583 SEL3.t70 VSS 0.011181f
C11584 SEL3.t35 VSS 0.011181f
C11585 SEL3.t78 VSS 0.011322f
C11586 SEL3.t55 VSS 0.011181f
C11587 SEL3.n18 VSS 0.044504f
C11588 SEL3.t68 VSS 0.002324f
C11589 SEL3.t47 VSS 0.002324f
C11590 SEL3.t62 VSS 0.002324f
C11591 SEL3.t24 VSS 0.002324f
C11592 SEL3.n19 VSS 0.042043f
C11593 SEL3.n20 VSS 0.065798f
C11594 SEL3.t4 VSS 0.011181f
C11595 SEL3.t28 VSS 0.011181f
C11596 SEL3.t12 VSS 0.011322f
C11597 SEL3.t65 VSS 0.011181f
C11598 SEL3.n21 VSS 0.044504f
C11599 SEL3.t5 VSS 0.002324f
C11600 SEL3.t59 VSS 0.002324f
C11601 SEL3.t77 VSS 0.002324f
C11602 SEL3.t17 VSS 0.002324f
C11603 SEL3.n22 VSS 0.042043f
C11604 SEL3.n23 VSS 0.065798f
C11605 SEL3.t8 VSS 0.011181f
C11606 SEL3.t33 VSS 0.011181f
C11607 SEL3.t46 VSS 0.011322f
C11608 SEL3.t71 VSS 0.011181f
C11609 SEL3.n24 VSS 0.044504f
C11610 SEL3.t38 VSS 0.002324f
C11611 SEL3.t63 VSS 0.002324f
C11612 SEL3.t82 VSS 0.002324f
C11613 SEL3.t20 VSS 0.002324f
C11614 SEL3.n25 VSS 0.042043f
C11615 SEL3.n26 VSS 0.065798f
C11616 SEL3.n27 VSS 0.742101f
C11617 SEL3.n28 VSS 0.606931f
C11618 SEL3.n29 VSS 0.588633f
C11619 SEL3.t39 VSS 0.011181f
C11620 SEL3.t60 VSS 0.011181f
C11621 SEL3.t21 VSS 0.011322f
C11622 SEL3.t79 VSS 0.011181f
C11623 SEL3.n30 VSS 0.044504f
C11624 SEL3.t14 VSS 0.002324f
C11625 SEL3.t69 VSS 0.002324f
C11626 SEL3.t27 VSS 0.002324f
C11627 SEL3.t54 VSS 0.002324f
C11628 SEL3.n31 VSS 0.042043f
C11629 SEL3.n32 VSS 0.065798f
C11630 SEL3.n33 VSS 0.113445f
C11631 SEL3.n34 VSS 0.590328f
C11632 SEL3.n35 VSS 0.586918f
C11633 SEL3.n36 VSS 0.590713f
C11634 SEL3.n37 VSS 0.290781f
C11635 SEL3.n38 VSS 0.072628f
C11636 SEL3.t3 VSS 0.011181f
C11637 SEL3.t26 VSS 0.011181f
C11638 SEL3.t76 VSS 0.011322f
C11639 SEL3.t49 VSS 0.011181f
C11640 SEL3.n39 VSS 0.044504f
C11641 SEL3.t66 VSS 0.002324f
C11642 SEL3.t40 VSS 0.002324f
C11643 SEL3.t75 VSS 0.002324f
C11644 SEL3.t16 VSS 0.002324f
C11645 SEL3.n40 VSS 0.042043f
C11646 SEL3.n41 VSS 0.065798f
C11647 SEL3.n42 VSS 0.142393f
C11648 SEL3.n43 VSS 0.779154f
C11649 SEL3.t6 VSS 0.005627f
C11650 SEL3.t41 VSS 0.011322f
C11651 SEL3.t83 VSS 0.011181f
C11652 SEL3.t45 VSS 0.011181f
C11653 SEL3.t22 VSS 0.011181f
C11654 SEL3.t67 VSS 0.002324f
C11655 SEL3.t34 VSS 0.002324f
C11656 SEL3.t53 VSS 0.002324f
C11657 SEL3.n44 VSS 0.068886f
C11658 SEL3.n45 VSS 0.050738f
C11659 SEL3.n46 VSS 0.027652f
C11660 SEL3.n47 VSS 0.027165f
C11661 SEL3.n48 VSS 0.01671f
C11662 SEL3.n49 VSS 0.021502f
C11663 SEL3.n50 VSS 0.114785f
C11664 mux8_5.NAND4F_5.Y.n0 VSS 0.25108f
C11665 mux8_5.NAND4F_5.Y.t10 VSS 0.017162f
C11666 mux8_5.NAND4F_5.Y.t9 VSS 0.050565f
C11667 mux8_5.NAND4F_5.Y.t11 VSS 0.016698f
C11668 mux8_5.NAND4F_5.Y.n1 VSS 0.086077f
C11669 mux8_5.NAND4F_5.Y.t2 VSS 0.099394f
C11670 mux8_5.NAND4F_5.Y.n2 VSS 0.798124f
C11671 mux8_5.NAND4F_5.Y.t0 VSS 0.012379f
C11672 mux8_5.NAND4F_5.Y.t1 VSS 0.012379f
C11673 mux8_5.NAND4F_5.Y.n3 VSS 0.028745f
C11674 mux8_5.NAND4F_5.Y.t8 VSS 0.012379f
C11675 mux8_5.NAND4F_5.Y.t7 VSS 0.012379f
C11676 mux8_5.NAND4F_5.Y.n4 VSS 0.028659f
C11677 mux8_5.NAND4F_5.Y.t5 VSS 0.012379f
C11678 mux8_5.NAND4F_5.Y.t6 VSS 0.012379f
C11679 mux8_5.NAND4F_5.Y.n5 VSS 0.028659f
C11680 mux8_5.NAND4F_5.Y.t3 VSS 0.012379f
C11681 mux8_5.NAND4F_5.Y.t4 VSS 0.012379f
C11682 mux8_5.NAND4F_5.Y.n6 VSS 0.028659f
C11683 mux8_5.NAND4F_5.Y.n7 VSS 0.117805f
C11684 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t17 VSS 0.013766f
C11685 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t21 VSS 0.027698f
C11686 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t22 VSS 0.027354f
C11687 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t18 VSS 0.027354f
C11688 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t20 VSS 0.027354f
C11689 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t16 VSS 0.005684f
C11690 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t23 VSS 0.005684f
C11691 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t19 VSS 0.005684f
C11692 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n0 VSS 0.168523f
C11693 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n1 VSS 0.124125f
C11694 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n2 VSS 0.067647f
C11695 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n3 VSS 0.066457f
C11696 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n4 VSS 0.040879f
C11697 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n5 VSS 0.05311f
C11698 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t15 VSS 0.030151f
C11699 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t13 VSS 0.009818f
C11700 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t14 VSS 0.013559f
C11701 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n6 VSS 0.014622f
C11702 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t12 VSS 0.010094f
C11703 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n7 VSS 0.025612f
C11704 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n8 VSS 0.044927f
C11705 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t10 VSS 0.004926f
C11706 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t8 VSS 0.004926f
C11707 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n9 VSS 0.011915f
C11708 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t4 VSS 0.004926f
C11709 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t5 VSS 0.004926f
C11710 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n10 VSS 0.011914f
C11711 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n11 VSS 0.085433f
C11712 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t9 VSS 0.004926f
C11713 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t0 VSS 0.004926f
C11714 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n12 VSS 0.009853f
C11715 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n13 VSS 0.00774f
C11716 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t11 VSS 0.020843f
C11717 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t1 VSS 0.020843f
C11718 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n14 VSS 0.041685f
C11719 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n15 VSS 0.016575f
C11720 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t7 VSS 0.020843f
C11721 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t6 VSS 0.020843f
C11722 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n16 VSS 0.041685f
C11723 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n17 VSS 0.018334f
C11724 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n18 VSS 0.188757f
C11725 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t2 VSS 0.020843f
C11726 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.t3 VSS 0.020843f
C11727 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n19 VSS 0.041685f
C11728 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n20 VSS 0.018362f
C11729 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n21 VSS 0.12106f
C11730 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n22 VSS 0.027282f
C11731 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_1.A.n23 VSS 0.119748f
C11732 a_n4879_2026.n0 VSS 1.48365f
C11733 a_n4879_2026.n1 VSS 1.48326f
C11734 a_n4879_2026.t5 VSS 0.093341f
C11735 a_n4879_2026.t10 VSS 0.093341f
C11736 a_n4879_2026.t9 VSS 0.093341f
C11737 a_n4879_2026.n2 VSS 0.202296f
C11738 a_n4879_2026.t8 VSS 0.093341f
C11739 a_n4879_2026.t4 VSS 0.093341f
C11740 a_n4879_2026.n3 VSS 0.202001f
C11741 a_n4879_2026.t3 VSS 0.093341f
C11742 a_n4879_2026.t11 VSS 0.093341f
C11743 a_n4879_2026.n4 VSS 0.202001f
C11744 a_n4879_2026.t0 VSS 0.093341f
C11745 a_n4879_2026.t1 VSS 0.093341f
C11746 a_n4879_2026.n5 VSS 0.202001f
C11747 a_n4879_2026.t2 VSS 0.093341f
C11748 a_n4879_2026.t6 VSS 0.093341f
C11749 a_n4879_2026.n6 VSS 0.202001f
C11750 a_n4879_2026.n7 VSS 0.20269f
C11751 a_n4879_2026.t7 VSS 0.093341f
C11752 left_shifter_0.S0.n0 VSS 2.34808f
C11753 left_shifter_0.S0.t5 VSS 0.114021f
C11754 left_shifter_0.S0.t6 VSS 0.335938f
C11755 left_shifter_0.S0.t4 VSS 0.110934f
C11756 left_shifter_0.S0.n1 VSS 0.571945f
C11757 left_shifter_0.S0.t3 VSS 0.054658f
C11758 left_shifter_0.S0.t1 VSS 0.054658f
C11759 left_shifter_0.S0.n2 VSS 0.121931f
C11760 left_shifter_0.S0.t2 VSS 0.198387f
C11761 left_shifter_0.S0.t0 VSS 0.157652f
C11762 AND8_0.NOT8_0.A3.n0 VSS 0.694442f
C11763 AND8_0.NOT8_0.A3.t10 VSS 0.016983f
C11764 AND8_0.NOT8_0.A3.t7 VSS 0.023706f
C11765 AND8_0.NOT8_0.A3.t9 VSS 0.023706f
C11766 AND8_0.NOT8_0.A3.n1 VSS 0.07717f
C11767 AND8_0.NOT8_0.A3.t8 VSS 0.027204f
C11768 AND8_0.NOT8_0.A3.n2 VSS 0.237866f
C11769 AND8_0.NOT8_0.A3.t6 VSS 0.080545f
C11770 AND8_0.NOT8_0.A3.t2 VSS 0.013326f
C11771 AND8_0.NOT8_0.A3.t0 VSS 0.013326f
C11772 AND8_0.NOT8_0.A3.n3 VSS 0.029732f
C11773 AND8_0.NOT8_0.A3.t4 VSS 0.013326f
C11774 AND8_0.NOT8_0.A3.t1 VSS 0.013326f
C11775 AND8_0.NOT8_0.A3.n4 VSS 0.029652f
C11776 AND8_0.NOT8_0.A3.t3 VSS 0.013326f
C11777 AND8_0.NOT8_0.A3.t5 VSS 0.013326f
C11778 AND8_0.NOT8_0.A3.n5 VSS 0.029652f
C11779 A3.t30 VSS 0.019493f
C11780 A3.t31 VSS 0.019493f
C11781 A3.t33 VSS 0.019493f
C11782 A3.t17 VSS 0.019493f
C11783 A3.n0 VSS 0.353963f
C11784 A3.t13 VSS 0.093805f
C11785 A3.t41 VSS 0.093805f
C11786 A3.t5 VSS 0.094987f
C11787 A3.t7 VSS 0.093805f
C11788 A3.n1 VSS 0.372133f
C11789 A3.n2 VSS 0.552152f
C11790 A3.t15 VSS 0.087719f
C11791 A3.t28 VSS 0.033671f
C11792 A3.t26 VSS 0.046498f
C11793 A3.n3 VSS 0.053519f
C11794 A3.t19 VSS 0.035392f
C11795 A3.n4 VSS 0.054276f
C11796 A3.n5 VSS 0.22466f
C11797 A3.t21 VSS 0.094987f
C11798 A3.t22 VSS 0.093805f
C11799 A3.t10 VSS 0.093805f
C11800 A3.t43 VSS 0.093805f
C11801 A3.n6 VSS 0.373369f
C11802 A3.t39 VSS 0.019493f
C11803 A3.t23 VSS 0.019493f
C11804 A3.t44 VSS 0.019493f
C11805 A3.t45 VSS 0.019493f
C11806 A3.n7 VSS 0.352726f
C11807 A3.n8 VSS 0.551734f
C11808 A3.n9 VSS 1.09681f
C11809 A3.n10 VSS 1.40614f
C11810 A3.n11 VSS 0.286403f
C11811 A3.t36 VSS 0.087719f
C11812 A3.t16 VSS 0.033671f
C11813 A3.t9 VSS 0.046498f
C11814 A3.n12 VSS 0.053519f
C11815 A3.t32 VSS 0.035392f
C11816 A3.n13 VSS 0.054276f
C11817 A3.n14 VSS 0.22522f
C11818 A3.t40 VSS 0.087719f
C11819 A3.t11 VSS 0.033671f
C11820 A3.t12 VSS 0.046498f
C11821 A3.n15 VSS 0.053519f
C11822 A3.t14 VSS 0.035392f
C11823 A3.n16 VSS 0.054276f
C11824 A3.n17 VSS 0.193368f
C11825 A3.n18 VSS 1.50671f
C11826 A3.n19 VSS 3.44166f
C11827 A3.t38 VSS 0.087719f
C11828 A3.t6 VSS 0.033671f
C11829 A3.t1 VSS 0.046498f
C11830 A3.n20 VSS 0.053519f
C11831 A3.t24 VSS 0.035392f
C11832 A3.n21 VSS 0.054276f
C11833 A3.n22 VSS 0.22522f
C11834 A3.n23 VSS 5.10341f
C11835 A3.n24 VSS 5.10026f
C11836 A3.n25 VSS 2.14728f
C11837 A3.t42 VSS 0.087719f
C11838 A3.t27 VSS 0.033671f
C11839 A3.t29 VSS 0.046498f
C11840 A3.n26 VSS 0.053519f
C11841 A3.t8 VSS 0.035392f
C11842 A3.n27 VSS 0.054276f
C11843 A3.n28 VSS 0.216341f
C11844 A3.n29 VSS 0.362433f
C11845 A3.n30 VSS 0.087728f
C11846 A3.n31 VSS 0.084067f
C11847 A3.n32 VSS 0.009703f
C11848 A3.n33 VSS 0.66893f
C11849 A3.n34 VSS 4.17692f
C11850 A3.n35 VSS 20.733902f
C11851 A3.t25 VSS 0.087717f
C11852 A3.t35 VSS 0.044333f
C11853 A3.t0 VSS 0.035443f
C11854 A3.n36 VSS 0.056283f
C11855 A3.t3 VSS 0.035392f
C11856 A3.n37 VSS 0.051906f
C11857 A3.n38 VSS 0.225331f
C11858 A3.n39 VSS 0.402741f
C11859 A3.n40 VSS 2.73879f
C11860 A3.t2 VSS 0.035093f
C11861 A3.t4 VSS 0.042295f
C11862 A3.t37 VSS 0.042295f
C11863 A3.t34 VSS 0.042295f
C11864 A3.t20 VSS 0.042295f
C11865 A3.t18 VSS 0.053433f
C11866 A3.n41 VSS 0.114164f
C11867 A3.n42 VSS 0.071878f
C11868 A3.n43 VSS 0.071878f
C11869 A3.n44 VSS 0.061949f
C11870 A3.n45 VSS 0.050631f
C11871 A3.n46 VSS 7.05125f
C11872 mux8_1.NAND4F_2.Y.n0 VSS 0.542699f
C11873 mux8_1.NAND4F_2.Y.t4 VSS 0.026757f
C11874 mux8_1.NAND4F_2.Y.t3 VSS 0.026757f
C11875 mux8_1.NAND4F_2.Y.n1 VSS 0.062132f
C11876 mux8_1.NAND4F_2.Y.t6 VSS 0.026757f
C11877 mux8_1.NAND4F_2.Y.t5 VSS 0.026757f
C11878 mux8_1.NAND4F_2.Y.n2 VSS 0.061945f
C11879 mux8_1.NAND4F_2.Y.t7 VSS 0.026757f
C11880 mux8_1.NAND4F_2.Y.t8 VSS 0.026757f
C11881 mux8_1.NAND4F_2.Y.n3 VSS 0.061945f
C11882 mux8_1.NAND4F_2.Y.t2 VSS 0.026757f
C11883 mux8_1.NAND4F_2.Y.t1 VSS 0.026757f
C11884 mux8_1.NAND4F_2.Y.n4 VSS 0.061945f
C11885 mux8_1.NAND4F_2.Y.n5 VSS 0.269719f
C11886 mux8_1.NAND4F_2.Y.t0 VSS 0.218188f
C11887 mux8_1.NAND4F_2.Y.t9 VSS 0.0349f
C11888 mux8_1.NAND4F_2.Y.t11 VSS 0.107689f
C11889 mux8_1.NAND4F_2.Y.t10 VSS 0.040202f
C11890 mux8_1.NAND4F_2.Y.n6 VSS 0.135132f
C11891 mux8_1.NAND4F_2.Y.n7 VSS 0.029427f
C11892 mux8_1.NAND4F_2.Y.n8 VSS 1.56995f
C11893 OR8_0.S0.n0 VSS 3.59161f
C11894 mux8_1.NAND4F_2.A VSS 2.77656f
C11895 OR8_0.NOT8_0.S0 VSS 19.5403f
C11896 OR8_0.S0.t4 VSS 0.174061f
C11897 OR8_0.S0.t5 VSS 0.16935f
C11898 OR8_0.S0.t6 VSS 0.512834f
C11899 OR8_0.S0.n1 VSS 0.873116f
C11900 mux8_1.A3 VSS 24.966f
C11901 OR8_0.S0.t2 VSS 0.08344f
C11902 OR8_0.S0.t1 VSS 0.08344f
C11903 OR8_0.S0.n2 VSS 0.18594f
C11904 OR8_0.S0.t3 VSS 0.302635f
C11905 OR8_0.S0.t0 VSS 0.240668f
C11906 AND8_0.NOT8_0.A1.n0 VSS 0.627733f
C11907 AND8_0.NOT8_0.A1.t9 VSS 0.015463f
C11908 AND8_0.NOT8_0.A1.t10 VSS 0.021586f
C11909 AND8_0.NOT8_0.A1.t8 VSS 0.021586f
C11910 AND8_0.NOT8_0.A1.n1 VSS 0.070267f
C11911 AND8_0.NOT8_0.A1.t7 VSS 0.024771f
C11912 AND8_0.NOT8_0.A1.n2 VSS 0.216729f
C11913 AND8_0.NOT8_0.A1.t0 VSS 0.073261f
C11914 AND8_0.NOT8_0.A1.t6 VSS 0.012134f
C11915 AND8_0.NOT8_0.A1.t4 VSS 0.012134f
C11916 AND8_0.NOT8_0.A1.n3 VSS 0.027073f
C11917 AND8_0.NOT8_0.A1.t2 VSS 0.012134f
C11918 AND8_0.NOT8_0.A1.t5 VSS 0.012134f
C11919 AND8_0.NOT8_0.A1.n4 VSS 0.026999f
C11920 AND8_0.NOT8_0.A1.t1 VSS 0.012134f
C11921 AND8_0.NOT8_0.A1.t3 VSS 0.012134f
C11922 AND8_0.NOT8_0.A1.n5 VSS 0.026999f
C11923 mux8_7.NAND4F_5.Y.n0 VSS 0.25108f
C11924 mux8_7.NAND4F_5.Y.t10 VSS 0.017162f
C11925 mux8_7.NAND4F_5.Y.t9 VSS 0.050565f
C11926 mux8_7.NAND4F_5.Y.t11 VSS 0.016698f
C11927 mux8_7.NAND4F_5.Y.n1 VSS 0.086077f
C11928 mux8_7.NAND4F_5.Y.t2 VSS 0.099394f
C11929 mux8_7.NAND4F_5.Y.n2 VSS 0.798124f
C11930 mux8_7.NAND4F_5.Y.t1 VSS 0.012379f
C11931 mux8_7.NAND4F_5.Y.t0 VSS 0.012379f
C11932 mux8_7.NAND4F_5.Y.n3 VSS 0.028745f
C11933 mux8_7.NAND4F_5.Y.t5 VSS 0.012379f
C11934 mux8_7.NAND4F_5.Y.t4 VSS 0.012379f
C11935 mux8_7.NAND4F_5.Y.n4 VSS 0.028659f
C11936 mux8_7.NAND4F_5.Y.t6 VSS 0.012379f
C11937 mux8_7.NAND4F_5.Y.t7 VSS 0.012379f
C11938 mux8_7.NAND4F_5.Y.n5 VSS 0.028659f
C11939 mux8_7.NAND4F_5.Y.t3 VSS 0.012379f
C11940 mux8_7.NAND4F_5.Y.t8 VSS 0.012379f
C11941 mux8_7.NAND4F_5.Y.n6 VSS 0.028659f
C11942 mux8_7.NAND4F_5.Y.n7 VSS 0.117805f
C11943 mux8_7.NAND4F_4.B.n0 VSS 0.921489f
C11944 mux8_7.NAND4F_4.B.t4 VSS 0.03989f
C11945 mux8_7.NAND4F_4.B.t6 VSS 0.123086f
C11946 mux8_7.NAND4F_4.B.t15 VSS 0.04595f
C11947 mux8_7.NAND4F_4.B.n1 VSS 0.154452f
C11948 mux8_7.NAND4F_4.B.n2 VSS 0.033769f
C11949 mux8_7.NAND4F_4.B.t7 VSS 0.03989f
C11950 mux8_7.NAND4F_4.B.t11 VSS 0.123086f
C11951 mux8_7.NAND4F_4.B.t5 VSS 0.04595f
C11952 mux8_7.NAND4F_4.B.n3 VSS 0.154452f
C11953 mux8_7.NAND4F_4.B.n4 VSS 0.032977f
C11954 mux8_7.NAND4F_4.B.t13 VSS 0.03989f
C11955 mux8_7.NAND4F_4.B.t8 VSS 0.123086f
C11956 mux8_7.NAND4F_4.B.t12 VSS 0.04595f
C11957 mux8_7.NAND4F_4.B.n5 VSS 0.154452f
C11958 mux8_7.NAND4F_4.B.n6 VSS 0.033699f
C11959 mux8_7.NAND4F_4.B.n7 VSS 0.612655f
C11960 mux8_7.NAND4F_4.B.t3 VSS 0.020325f
C11961 mux8_7.NAND4F_4.B.t2 VSS 0.020325f
C11962 mux8_7.NAND4F_4.B.n8 VSS 0.045293f
C11963 mux8_7.NAND4F_4.B.t1 VSS 0.073718f
C11964 mux8_7.NAND4F_4.B.t0 VSS 0.058624f
C11965 mux8_7.NAND4F_4.B.n9 VSS 0.607515f
C11966 mux8_7.NAND4F_4.B.t10 VSS 0.03989f
C11967 mux8_7.NAND4F_4.B.t14 VSS 0.123086f
C11968 mux8_7.NAND4F_4.B.t9 VSS 0.04595f
C11969 mux8_7.NAND4F_4.B.n10 VSS 0.154452f
C11970 mux8_7.NAND4F_4.B.n11 VSS 0.033659f
C11971 mux8_7.NAND4F_4.B.n12 VSS 0.776456f
C11972 A5.t15 VSS 0.028472f
C11973 A5.t17 VSS 0.028472f
C11974 A5.t18 VSS 0.028472f
C11975 A5.t9 VSS 0.028472f
C11976 A5.n0 VSS 0.517003f
C11977 A5.t7 VSS 0.137013f
C11978 A5.t23 VSS 0.137013f
C11979 A5.t2 VSS 0.138739f
C11980 A5.t6 VSS 0.137013f
C11981 A5.n1 VSS 0.543543f
C11982 A5.n2 VSS 0.806481f
C11983 A5.t25 VSS 0.128123f
C11984 A5.t29 VSS 0.04918f
C11985 A5.t27 VSS 0.067916f
C11986 A5.n3 VSS 0.078171f
C11987 A5.t28 VSS 0.051695f
C11988 A5.n4 VSS 0.079276f
C11989 A5.n5 VSS 0.328142f
C11990 A5.t13 VSS 0.138739f
C11991 A5.t4 VSS 0.137013f
C11992 A5.t16 VSS 0.137013f
C11993 A5.t10 VSS 0.137013f
C11994 A5.n6 VSS 0.545349f
C11995 A5.t8 VSS 0.028472f
C11996 A5.t26 VSS 0.028472f
C11997 A5.t0 VSS 0.028472f
C11998 A5.t19 VSS 0.028472f
C11999 A5.n7 VSS 0.515197f
C12000 A5.n8 VSS 0.805871f
C12001 A5.n9 VSS 1.60202f
C12002 A5.n10 VSS 2.05337f
C12003 A5.t24 VSS 0.12812f
C12004 A5.t20 VSS 0.064754f
C12005 A5.t5 VSS 0.051768f
C12006 A5.n11 VSS 0.082208f
C12007 A5.t14 VSS 0.051695f
C12008 A5.n12 VSS 0.075814f
C12009 A5.n13 VSS 0.329122f
C12010 A5.n14 VSS 0.607275f
C12011 A5.n15 VSS 4.21513f
C12012 A5.t1 VSS 0.051258f
C12013 A5.t3 VSS 0.061777f
C12014 A5.t22 VSS 0.061777f
C12015 A5.t21 VSS 0.061777f
C12016 A5.t12 VSS 0.061777f
C12017 A5.t11 VSS 0.078045f
C12018 A5.n16 VSS 0.166749f
C12019 A5.n17 VSS 0.104986f
C12020 A5.n18 VSS 0.104986f
C12021 A5.n19 VSS 0.090484f
C12022 A5.n20 VSS 0.073952f
C12023 A5.n21 VSS 15.018801f
C12024 mux8_0.NAND4F_3.Y.n0 VSS 0.306333f
C12025 mux8_0.NAND4F_3.Y.t7 VSS 0.015103f
C12026 mux8_0.NAND4F_3.Y.t8 VSS 0.015103f
C12027 mux8_0.NAND4F_3.Y.n1 VSS 0.035071f
C12028 mux8_0.NAND4F_3.Y.t3 VSS 0.015103f
C12029 mux8_0.NAND4F_3.Y.t2 VSS 0.015103f
C12030 mux8_0.NAND4F_3.Y.n2 VSS 0.034966f
C12031 mux8_0.NAND4F_3.Y.t0 VSS 0.015103f
C12032 mux8_0.NAND4F_3.Y.t1 VSS 0.015103f
C12033 mux8_0.NAND4F_3.Y.n3 VSS 0.034966f
C12034 mux8_0.NAND4F_3.Y.t5 VSS 0.015103f
C12035 mux8_0.NAND4F_3.Y.t4 VSS 0.015103f
C12036 mux8_0.NAND4F_3.Y.n4 VSS 0.034966f
C12037 mux8_0.NAND4F_3.Y.n5 VSS 0.152246f
C12038 mux8_0.NAND4F_3.Y.t6 VSS 0.143521f
C12039 mux8_0.NAND4F_3.Y.t10 VSS 0.0197f
C12040 mux8_0.NAND4F_3.Y.t11 VSS 0.0197f
C12041 mux8_0.NAND4F_3.Y.n6 VSS 0.023128f
C12042 mux8_0.NAND4F_3.Y.t9 VSS 0.061756f
C12043 mux8_0.NAND4F_3.Y.n7 VSS 0.129679f
C12044 mux8_0.NAND4F_0.C.n0 VSS 1.66671f
C12045 mux8_0.NAND4F_0.C.t9 VSS 0.230719f
C12046 mux8_0.NAND4F_0.C.t12 VSS 0.073597f
C12047 mux8_0.NAND4F_0.C.t10 VSS 0.073597f
C12048 mux8_0.NAND4F_0.C.n1 VSS 0.086405f
C12049 mux8_0.NAND4F_0.C.n2 VSS 0.484461f
C12050 mux8_0.NAND4F_0.C.t8 VSS 0.073597f
C12051 mux8_0.NAND4F_0.C.t11 VSS 0.073597f
C12052 mux8_0.NAND4F_0.C.n3 VSS 0.086405f
C12053 mux8_0.NAND4F_0.C.t5 VSS 0.230719f
C12054 mux8_0.NAND4F_0.C.n4 VSS 0.484492f
C12055 mux8_0.NAND4F_0.C.t4 VSS 0.073597f
C12056 mux8_0.NAND4F_0.C.t6 VSS 0.073597f
C12057 mux8_0.NAND4F_0.C.n5 VSS 0.086405f
C12058 mux8_0.NAND4F_0.C.t7 VSS 0.230719f
C12059 mux8_0.NAND4F_0.C.n6 VSS 0.484506f
C12060 mux8_0.NAND4F_0.C.n7 VSS 1.76702f
C12061 mux8_0.NAND4F_0.C.t2 VSS 0.0375f
C12062 mux8_0.NAND4F_0.C.t3 VSS 0.0375f
C12063 mux8_0.NAND4F_0.C.n8 VSS 0.083565f
C12064 mux8_0.NAND4F_0.C.t1 VSS 0.136011f
C12065 mux8_0.NAND4F_0.C.t0 VSS 0.108161f
C12066 mux8_0.NAND4F_0.C.n9 VSS 3.09373f
C12067 mux8_0.NAND4F_0.C.t14 VSS 0.230719f
C12068 mux8_0.NAND4F_0.C.t15 VSS 0.073597f
C12069 mux8_0.NAND4F_0.C.t13 VSS 0.073597f
C12070 mux8_0.NAND4F_0.C.n10 VSS 0.086405f
C12071 mux8_0.NAND4F_0.C.n11 VSS 0.484478f
C12072 mux8_0.NAND4F_0.C.n12 VSS 2.47931f
C12073 mux8_2.NAND4F_1.Y.n0 VSS 0.655599f
C12074 mux8_2.NAND4F_1.Y.t4 VSS 0.306614f
C12075 mux8_2.NAND4F_1.Y.t11 VSS 0.132168f
C12076 mux8_2.NAND4F_1.Y.t9 VSS 0.04216f
C12077 mux8_2.NAND4F_1.Y.t10 VSS 0.04216f
C12078 mux8_2.NAND4F_1.Y.n1 VSS 0.049498f
C12079 mux8_2.NAND4F_1.Y.n2 VSS 0.277534f
C12080 mux8_2.NAND4F_1.Y.t0 VSS 0.032323f
C12081 mux8_2.NAND4F_1.Y.t1 VSS 0.032323f
C12082 mux8_2.NAND4F_1.Y.n3 VSS 0.075057f
C12083 mux8_2.NAND4F_1.Y.t6 VSS 0.032323f
C12084 mux8_2.NAND4F_1.Y.t5 VSS 0.032323f
C12085 mux8_2.NAND4F_1.Y.n4 VSS 0.074832f
C12086 mux8_2.NAND4F_1.Y.t8 VSS 0.032323f
C12087 mux8_2.NAND4F_1.Y.t7 VSS 0.032323f
C12088 mux8_2.NAND4F_1.Y.n5 VSS 0.074832f
C12089 mux8_2.NAND4F_1.Y.t2 VSS 0.032323f
C12090 mux8_2.NAND4F_1.Y.t3 VSS 0.032323f
C12091 mux8_2.NAND4F_1.Y.n6 VSS 0.074832f
C12092 mux8_2.NAND4F_1.Y.n7 VSS 0.307603f
C12093 XOR8_0.S1.t14 VSS 0.122143f
C12094 XOR8_0.S1.t13 VSS 0.359868f
C12095 XOR8_0.S1.t12 VSS 0.118837f
C12096 XOR8_0.S1.n0 VSS 0.612649f
C12097 XOR8_0.S1.t4 VSS 0.035569f
C12098 XOR8_0.S1.t5 VSS 0.035569f
C12099 XOR8_0.S1.n1 VSS 0.086028f
C12100 XOR8_0.S1.t0 VSS 0.035569f
C12101 XOR8_0.S1.t7 VSS 0.035569f
C12102 XOR8_0.S1.n2 VSS 0.086018f
C12103 XOR8_0.S1.n3 VSS 0.616825f
C12104 XOR8_0.S1.t6 VSS 0.035569f
C12105 XOR8_0.S1.t11 VSS 0.035569f
C12106 XOR8_0.S1.n4 VSS 0.071138f
C12107 XOR8_0.S1.n5 VSS 0.055881f
C12108 XOR8_0.S1.t3 VSS 0.150484f
C12109 XOR8_0.S1.t8 VSS 0.150484f
C12110 XOR8_0.S1.n6 VSS 0.300967f
C12111 XOR8_0.S1.n7 VSS 0.119387f
C12112 XOR8_0.S1.t1 VSS 0.150484f
C12113 XOR8_0.S1.t2 VSS 0.150484f
C12114 XOR8_0.S1.n8 VSS 0.300967f
C12115 XOR8_0.S1.n9 VSS 0.132371f
C12116 XOR8_0.S1.n10 VSS 1.36283f
C12117 XOR8_0.S1.t9 VSS 0.150484f
C12118 XOR8_0.S1.t10 VSS 0.150484f
C12119 XOR8_0.S1.n11 VSS 0.300967f
C12120 XOR8_0.S1.n12 VSS 0.132571f
C12121 XOR8_0.S1.n13 VSS 0.874059f
C12122 XOR8_0.S1.n14 VSS 0.196738f
C12123 XOR8_0.S1.n15 VSS 0.865105f
C12124 mux8_0.NAND4F_8.Y.n0 VSS 0.539804f
C12125 mux8_0.NAND4F_8.Y.t9 VSS 0.026899f
C12126 mux8_0.NAND4F_8.Y.t11 VSS 0.028853f
C12127 mux8_0.NAND4F_8.Y.n1 VSS 0.042994f
C12128 mux8_0.NAND4F_8.Y.t12 VSS 0.026899f
C12129 mux8_0.NAND4F_8.Y.t13 VSS 0.026899f
C12130 mux8_0.NAND4F_8.Y.t14 VSS 0.026899f
C12131 mux8_0.NAND4F_8.Y.t10 VSS 0.033983f
C12132 mux8_0.NAND4F_8.Y.n2 VSS 0.072608f
C12133 mux8_0.NAND4F_8.Y.n3 VSS 0.045714f
C12134 mux8_0.NAND4F_8.Y.n4 VSS 0.037354f
C12135 mux8_0.NAND4F_8.Y.n5 VSS 0.018278f
C12136 mux8_0.NAND4F_8.Y.t2 VSS 0.026614f
C12137 mux8_0.NAND4F_8.Y.t3 VSS 0.026614f
C12138 mux8_0.NAND4F_8.Y.n6 VSS 0.0618f
C12139 mux8_0.NAND4F_8.Y.t0 VSS 0.026614f
C12140 mux8_0.NAND4F_8.Y.t1 VSS 0.026614f
C12141 mux8_0.NAND4F_8.Y.n7 VSS 0.061615f
C12142 mux8_0.NAND4F_8.Y.t5 VSS 0.026614f
C12143 mux8_0.NAND4F_8.Y.t4 VSS 0.026614f
C12144 mux8_0.NAND4F_8.Y.n8 VSS 0.061615f
C12145 mux8_0.NAND4F_8.Y.t6 VSS 0.026614f
C12146 mux8_0.NAND4F_8.Y.t7 VSS 0.026614f
C12147 mux8_0.NAND4F_8.Y.n9 VSS 0.061615f
C12148 mux8_0.NAND4F_8.Y.n10 VSS 0.268281f
C12149 mux8_0.NAND4F_8.Y.t8 VSS 0.21369f
C12150 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t22 VSS 0.013766f
C12151 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t12 VSS 0.027698f
C12152 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t17 VSS 0.027354f
C12153 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t15 VSS 0.027354f
C12154 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t20 VSS 0.027354f
C12155 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t14 VSS 0.005684f
C12156 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t13 VSS 0.005684f
C12157 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t23 VSS 0.005684f
C12158 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n0 VSS 0.168523f
C12159 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n1 VSS 0.124125f
C12160 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n2 VSS 0.067647f
C12161 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n3 VSS 0.066457f
C12162 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n4 VSS 0.040879f
C12163 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n5 VSS 0.05311f
C12164 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t16 VSS 0.030151f
C12165 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t21 VSS 0.009818f
C12166 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t18 VSS 0.013559f
C12167 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n6 VSS 0.014622f
C12168 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t19 VSS 0.010094f
C12169 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n7 VSS 0.025612f
C12170 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n8 VSS 0.044927f
C12171 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t11 VSS 0.004926f
C12172 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t9 VSS 0.004926f
C12173 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n9 VSS 0.011915f
C12174 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t5 VSS 0.004926f
C12175 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t3 VSS 0.004926f
C12176 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n10 VSS 0.011914f
C12177 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n11 VSS 0.085433f
C12178 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t10 VSS 0.004926f
C12179 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t4 VSS 0.004926f
C12180 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n12 VSS 0.009853f
C12181 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n13 VSS 0.00774f
C12182 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t8 VSS 0.020843f
C12183 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t2 VSS 0.020843f
C12184 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n14 VSS 0.041685f
C12185 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n15 VSS 0.016575f
C12186 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t6 VSS 0.020843f
C12187 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t7 VSS 0.020843f
C12188 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n16 VSS 0.041685f
C12189 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n17 VSS 0.018334f
C12190 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n18 VSS 0.188757f
C12191 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t0 VSS 0.020843f
C12192 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.t1 VSS 0.020843f
C12193 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n19 VSS 0.041685f
C12194 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n20 VSS 0.018362f
C12195 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n21 VSS 0.12106f
C12196 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n22 VSS 0.027282f
C12197 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_1.A.n23 VSS 0.119748f
C12198 a_n24624_2026.n0 VSS 1.48326f
C12199 a_n24624_2026.n1 VSS 1.48365f
C12200 a_n24624_2026.t4 VSS 0.093341f
C12201 a_n24624_2026.t9 VSS 0.093341f
C12202 a_n24624_2026.t10 VSS 0.093341f
C12203 a_n24624_2026.n2 VSS 0.20269f
C12204 a_n24624_2026.t1 VSS 0.093341f
C12205 a_n24624_2026.t11 VSS 0.093341f
C12206 a_n24624_2026.n3 VSS 0.202001f
C12207 a_n24624_2026.t2 VSS 0.093341f
C12208 a_n24624_2026.t0 VSS 0.093341f
C12209 a_n24624_2026.n4 VSS 0.202001f
C12210 a_n24624_2026.t7 VSS 0.093341f
C12211 a_n24624_2026.t8 VSS 0.093341f
C12212 a_n24624_2026.n5 VSS 0.202001f
C12213 a_n24624_2026.t3 VSS 0.093341f
C12214 a_n24624_2026.t6 VSS 0.093341f
C12215 a_n24624_2026.n6 VSS 0.202001f
C12216 a_n24624_2026.n7 VSS 0.202296f
C12217 a_n24624_2026.t5 VSS 0.093341f
C12218 AND8_0.NOT8_0.A2.n0 VSS 0.64763f
C12219 AND8_0.NOT8_0.A2.t8 VSS 0.015948f
C12220 AND8_0.NOT8_0.A2.t9 VSS 0.022262f
C12221 AND8_0.NOT8_0.A2.t7 VSS 0.022262f
C12222 AND8_0.NOT8_0.A2.n1 VSS 0.072469f
C12223 AND8_0.NOT8_0.A2.t10 VSS 0.025547f
C12224 AND8_0.NOT8_0.A2.n2 VSS 0.223522f
C12225 AND8_0.NOT8_0.A2.t2 VSS 0.075549f
C12226 AND8_0.NOT8_0.A2.t1 VSS 0.012514f
C12227 AND8_0.NOT8_0.A2.t6 VSS 0.012514f
C12228 AND8_0.NOT8_0.A2.n3 VSS 0.027921f
C12229 AND8_0.NOT8_0.A2.t3 VSS 0.012514f
C12230 AND8_0.NOT8_0.A2.t0 VSS 0.012514f
C12231 AND8_0.NOT8_0.A2.n4 VSS 0.027846f
C12232 AND8_0.NOT8_0.A2.t5 VSS 0.012514f
C12233 AND8_0.NOT8_0.A2.t4 VSS 0.012514f
C12234 AND8_0.NOT8_0.A2.n5 VSS 0.027846f
C12235 A2.t4 VSS 0.102039f
C12236 A2.t38 VSS 0.039167f
C12237 A2.t5 VSS 0.054089f
C12238 A2.n0 VSS 0.062256f
C12239 A2.t35 VSS 0.04117f
C12240 A2.n1 VSS 0.063136f
C12241 A2.n2 VSS 0.261336f
C12242 A2.t2 VSS 0.110493f
C12243 A2.t6 VSS 0.109119f
C12244 A2.t40 VSS 0.109119f
C12245 A2.t25 VSS 0.109119f
C12246 A2.n3 VSS 0.434323f
C12247 A2.t20 VSS 0.022676f
C12248 A2.t8 VSS 0.022676f
C12249 A2.t27 VSS 0.022676f
C12250 A2.t30 VSS 0.022676f
C12251 A2.n4 VSS 0.410309f
C12252 A2.n5 VSS 0.641806f
C12253 A2.n6 VSS 1.27587f
C12254 A2.n7 VSS 1.63542f
C12255 A2.t36 VSS 0.120278f
C12256 A2.t45 VSS 0.039167f
C12257 A2.t1 VSS 0.054089f
C12258 A2.n8 VSS 0.058328f
C12259 A2.t29 VSS 0.040267f
C12260 A2.n9 VSS 0.102173f
C12261 A2.n10 VSS 0.179554f
C12262 A2.t23 VSS 0.102039f
C12263 A2.t3 VSS 0.039167f
C12264 A2.t44 VSS 0.054089f
C12265 A2.n11 VSS 0.062256f
C12266 A2.t15 VSS 0.04117f
C12267 A2.n12 VSS 0.063136f
C12268 A2.n13 VSS 0.252437f
C12269 A2.t31 VSS 0.120278f
C12270 A2.t17 VSS 0.039167f
C12271 A2.t11 VSS 0.054089f
C12272 A2.n14 VSS 0.058328f
C12273 A2.t18 VSS 0.040267f
C12274 A2.n15 VSS 0.102173f
C12275 A2.n16 VSS 0.179554f
C12276 A2.n17 VSS 2.94996f
C12277 A2.t14 VSS 0.120278f
C12278 A2.t37 VSS 0.039167f
C12279 A2.t32 VSS 0.054089f
C12280 A2.n18 VSS 0.058328f
C12281 A2.t39 VSS 0.040267f
C12282 A2.n19 VSS 0.102173f
C12283 A2.n20 VSS 0.179554f
C12284 A2.n21 VSS 5.24226f
C12285 A2.n22 VSS 5.20658f
C12286 A2.n23 VSS 23.4961f
C12287 A2.t21 VSS 0.102036f
C12288 A2.t0 VSS 0.051571f
C12289 A2.t16 VSS 0.041229f
C12290 A2.n24 VSS 0.065472f
C12291 A2.t26 VSS 0.04117f
C12292 A2.n25 VSS 0.060379f
C12293 A2.n26 VSS 0.262117f
C12294 A2.n27 VSS 0.456295f
C12295 A2.n28 VSS 3.01703f
C12296 A2.t9 VSS 0.040822f
C12297 A2.t12 VSS 0.0492f
C12298 A2.t43 VSS 0.0492f
C12299 A2.t41 VSS 0.0492f
C12300 A2.t24 VSS 0.0492f
C12301 A2.t22 VSS 0.062156f
C12302 A2.n29 VSS 0.132801f
C12303 A2.n30 VSS 0.083612f
C12304 A2.n31 VSS 0.083612f
C12305 A2.n32 VSS 0.072062f
C12306 A2.n33 VSS 0.058896f
C12307 A2.n34 VSS 9.15686f
C12308 A2.t28 VSS 0.022676f
C12309 A2.t10 VSS 0.022676f
C12310 A2.t13 VSS 0.022676f
C12311 A2.t42 VSS 0.022676f
C12312 A2.n35 VSS 0.411748f
C12313 A2.t34 VSS 0.109119f
C12314 A2.t19 VSS 0.109119f
C12315 A2.t7 VSS 0.110493f
C12316 A2.t33 VSS 0.109119f
C12317 A2.n36 VSS 0.432884f
C12318 A2.n37 VSS 0.642292f
C12319 A2.n38 VSS 1.59379f
C12320 MULT_0.4bit_ADDER_0.A2.n0 VSS 2.93502f
C12321 MULT_0.4bit_ADDER_0.A2.t3 VSS 0.069415f
C12322 MULT_0.4bit_ADDER_0.A2.t1 VSS 0.019136f
C12323 MULT_0.4bit_ADDER_0.A2.t2 VSS 0.019136f
C12324 MULT_0.4bit_ADDER_0.A2.n1 VSS 0.042666f
C12325 MULT_0.4bit_ADDER_0.A2.t0 VSS 0.055254f
C12326 MULT_0.4bit_ADDER_0.A2.t9 VSS 0.060358f
C12327 MULT_0.4bit_ADDER_0.A2.t10 VSS 0.023168f
C12328 MULT_0.4bit_ADDER_0.A2.t6 VSS 0.031995f
C12329 MULT_0.4bit_ADDER_0.A2.n2 VSS 0.036826f
C12330 MULT_0.4bit_ADDER_0.A2.t14 VSS 0.024353f
C12331 MULT_0.4bit_ADDER_0.A2.n3 VSS 0.037346f
C12332 MULT_0.4bit_ADDER_0.A2.t15 VSS 0.065359f
C12333 MULT_0.4bit_ADDER_0.A2.t11 VSS 0.064546f
C12334 MULT_0.4bit_ADDER_0.A2.t12 VSS 0.064546f
C12335 MULT_0.4bit_ADDER_0.A2.t8 VSS 0.064546f
C12336 MULT_0.4bit_ADDER_0.A2.n4 VSS 0.256911f
C12337 MULT_0.4bit_ADDER_0.A2.t7 VSS 0.013413f
C12338 MULT_0.4bit_ADDER_0.A2.t4 VSS 0.013413f
C12339 MULT_0.4bit_ADDER_0.A2.t13 VSS 0.013413f
C12340 MULT_0.4bit_ADDER_0.A2.t5 VSS 0.013413f
C12341 MULT_0.4bit_ADDER_0.A2.n5 VSS 0.242706f
C12342 MULT_0.4bit_ADDER_0.A2.n6 VSS 0.379641f
C12343 MULT_0.4bit_ADDER_0.A2.n7 VSS 0.897564f
C12344 mux8_1.NAND4F_6.Y.n0 VSS 0.599344f
C12345 mux8_1.NAND4F_6.Y.t3 VSS 0.244548f
C12346 mux8_1.NAND4F_6.Y.t10 VSS 0.038543f
C12347 mux8_1.NAND4F_6.Y.t9 VSS 0.118929f
C12348 mux8_1.NAND4F_6.Y.t11 VSS 0.044398f
C12349 mux8_1.NAND4F_6.Y.n1 VSS 0.149236f
C12350 mux8_1.NAND4F_6.Y.n2 VSS 0.032396f
C12351 mux8_1.NAND4F_6.Y.n3 VSS 1.72835f
C12352 mux8_1.NAND4F_6.Y.t0 VSS 0.029549f
C12353 mux8_1.NAND4F_6.Y.t1 VSS 0.029549f
C12354 mux8_1.NAND4F_6.Y.n4 VSS 0.068617f
C12355 mux8_1.NAND4F_6.Y.t5 VSS 0.029549f
C12356 mux8_1.NAND4F_6.Y.t6 VSS 0.029549f
C12357 mux8_1.NAND4F_6.Y.n5 VSS 0.068411f
C12358 mux8_1.NAND4F_6.Y.t7 VSS 0.029549f
C12359 mux8_1.NAND4F_6.Y.t8 VSS 0.029549f
C12360 mux8_1.NAND4F_6.Y.n6 VSS 0.068411f
C12361 mux8_1.NAND4F_6.Y.t2 VSS 0.029549f
C12362 mux8_1.NAND4F_6.Y.t4 VSS 0.029549f
C12363 mux8_1.NAND4F_6.Y.n7 VSS 0.068411f
C12364 mux8_1.NAND4F_6.Y.n8 VSS 0.281208f
C12365 AND8_0.NOT8_0.A7.n0 VSS 0.651398f
C12366 AND8_0.NOT8_0.A7.t9 VSS 0.016108f
C12367 AND8_0.NOT8_0.A7.t10 VSS 0.022485f
C12368 AND8_0.NOT8_0.A7.t7 VSS 0.022485f
C12369 AND8_0.NOT8_0.A7.n1 VSS 0.073194f
C12370 AND8_0.NOT8_0.A7.t8 VSS 0.025803f
C12371 AND8_0.NOT8_0.A7.n2 VSS 0.22399f
C12372 AND8_0.NOT8_0.A7.t3 VSS 0.076305f
C12373 AND8_0.NOT8_0.A7.t4 VSS 0.012639f
C12374 AND8_0.NOT8_0.A7.t5 VSS 0.012639f
C12375 AND8_0.NOT8_0.A7.n3 VSS 0.028201f
C12376 AND8_0.NOT8_0.A7.t0 VSS 0.012639f
C12377 AND8_0.NOT8_0.A7.t6 VSS 0.012639f
C12378 AND8_0.NOT8_0.A7.n4 VSS 0.028124f
C12379 AND8_0.NOT8_0.A7.t2 VSS 0.012639f
C12380 AND8_0.NOT8_0.A7.t1 VSS 0.012639f
C12381 AND8_0.NOT8_0.A7.n5 VSS 0.028124f
C12382 A7.t24 VSS 0.012518f
C12383 A7.t26 VSS 0.012518f
C12384 A7.t33 VSS 0.012518f
C12385 A7.t12 VSS 0.012518f
C12386 A7.n0 VSS 0.227294f
C12387 A7.t8 VSS 0.060236f
C12388 A7.t36 VSS 0.060236f
C12389 A7.t1 VSS 0.060995f
C12390 A7.t2 VSS 0.060236f
C12391 A7.n1 VSS 0.238962f
C12392 A7.n2 VSS 0.354559f
C12393 A7.t23 VSS 0.030315f
C12394 A7.t45 VSS 0.060995f
C12395 A7.t19 VSS 0.060236f
C12396 A7.t13 VSS 0.060236f
C12397 A7.t5 VSS 0.060236f
C12398 A7.t28 VSS 0.012518f
C12399 A7.t42 VSS 0.012518f
C12400 A7.t4 VSS 0.012518f
C12401 A7.n3 VSS 0.371108f
C12402 A7.n4 VSS 0.273338f
C12403 A7.n5 VSS 0.148967f
C12404 A7.n6 VSS 0.146347f
C12405 A7.n7 VSS 0.09002f
C12406 A7.n8 VSS 0.115839f
C12407 A7.t43 VSS 0.030315f
C12408 A7.t16 VSS 0.060995f
C12409 A7.t39 VSS 0.060236f
C12410 A7.t34 VSS 0.060236f
C12411 A7.t7 VSS 0.060236f
C12412 A7.t32 VSS 0.012518f
C12413 A7.t44 VSS 0.012518f
C12414 A7.t6 VSS 0.012518f
C12415 A7.n9 VSS 0.371108f
C12416 A7.n10 VSS 0.273338f
C12417 A7.n11 VSS 0.148967f
C12418 A7.n12 VSS 0.146347f
C12419 A7.n13 VSS 0.09002f
C12420 A7.n14 VSS 0.115839f
C12421 A7.n15 VSS 2.93873f
C12422 A7.t21 VSS 0.056328f
C12423 A7.t27 VSS 0.021621f
C12424 A7.t29 VSS 0.029858f
C12425 A7.n16 VSS 0.034367f
C12426 A7.t31 VSS 0.022727f
C12427 A7.n17 VSS 0.034853f
C12428 A7.n18 VSS 0.144263f
C12429 A7.t35 VSS 0.060995f
C12430 A7.t15 VSS 0.060236f
C12431 A7.t37 VSS 0.060236f
C12432 A7.t20 VSS 0.060236f
C12433 A7.n19 VSS 0.239756f
C12434 A7.t18 VSS 0.012518f
C12435 A7.t3 VSS 0.012518f
C12436 A7.t17 VSS 0.012518f
C12437 A7.t41 VSS 0.012518f
C12438 A7.n20 VSS 0.2265f
C12439 A7.n21 VSS 0.354291f
C12440 A7.n22 VSS 0.704306f
C12441 A7.n23 VSS 0.901308f
C12442 A7.n24 VSS 1.13841f
C12443 A7.n25 VSS 11.8232f
C12444 A7.t0 VSS 0.056326f
C12445 A7.t11 VSS 0.028468f
C12446 A7.t14 VSS 0.022759f
C12447 A7.n26 VSS 0.036142f
C12448 A7.t30 VSS 0.022727f
C12449 A7.n27 VSS 0.033331f
C12450 A7.n28 VSS 0.144694f
C12451 A7.n29 VSS 0.278948f
C12452 A7.n30 VSS 1.92625f
C12453 A7.t22 VSS 0.022535f
C12454 A7.t25 VSS 0.027159f
C12455 A7.t10 VSS 0.027159f
C12456 A7.t9 VSS 0.027159f
C12457 A7.t40 VSS 0.027159f
C12458 A7.t38 VSS 0.034312f
C12459 A7.n31 VSS 0.073309f
C12460 A7.n32 VSS 0.046156f
C12461 A7.n33 VSS 0.046156f
C12462 A7.n34 VSS 0.03978f
C12463 A7.n35 VSS 0.032512f
C12464 A7.n36 VSS 7.23396f
C12465 XOR8_0.S6.t13 VSS 0.036538f
C12466 XOR8_0.S6.t12 VSS 0.107652f
C12467 XOR8_0.S6.t14 VSS 0.035549f
C12468 XOR8_0.S6.n0 VSS 0.183269f
C12469 XOR8_0.S6.t0 VSS 0.01064f
C12470 XOR8_0.S6.t2 VSS 0.01064f
C12471 XOR8_0.S6.n1 VSS 0.025735f
C12472 XOR8_0.S6.t8 VSS 0.01064f
C12473 XOR8_0.S6.t3 VSS 0.01064f
C12474 XOR8_0.S6.n2 VSS 0.025732f
C12475 XOR8_0.S6.n3 VSS 0.184518f
C12476 XOR8_0.S6.t1 VSS 0.01064f
C12477 XOR8_0.S6.t7 VSS 0.01064f
C12478 XOR8_0.S6.n4 VSS 0.02128f
C12479 XOR8_0.S6.n5 VSS 0.016716f
C12480 XOR8_0.S6.t11 VSS 0.045016f
C12481 XOR8_0.S6.t4 VSS 0.045016f
C12482 XOR8_0.S6.n6 VSS 0.090032f
C12483 XOR8_0.S6.n7 VSS 0.035714f
C12484 XOR8_0.S6.t9 VSS 0.045016f
C12485 XOR8_0.S6.t10 VSS 0.045016f
C12486 XOR8_0.S6.n8 VSS 0.090032f
C12487 XOR8_0.S6.n9 VSS 0.039598f
C12488 XOR8_0.S6.n10 VSS 0.407679f
C12489 XOR8_0.S6.t5 VSS 0.045016f
C12490 XOR8_0.S6.t6 VSS 0.045016f
C12491 XOR8_0.S6.n11 VSS 0.090032f
C12492 XOR8_0.S6.n12 VSS 0.039657f
C12493 XOR8_0.S6.n13 VSS 0.261467f
C12494 XOR8_0.S6.n14 VSS 0.058853f
C12495 XOR8_0.S6.n15 VSS 0.258789f
C12496 MULT_0.4bit_ADDER_1.Cout VSS 1.09361f
C12497 MULT_0.4bit_ADDER_2.B3.n0 VSS 1.31166f
C12498 MULT_0.4bit_ADDER_2.FULL_ADDER_0.NAND2_0.A VSS 0.157675f
C12499 MULT_0.4bit_ADDER_1.FULL_ADDER_0.COUT VSS 0.925405f
C12500 MULT_0.4bit_ADDER_2.B3.t9 VSS 0.042216f
C12501 MULT_0.4bit_ADDER_2.B3.t13 VSS 0.013747f
C12502 MULT_0.4bit_ADDER_2.B3.t15 VSS 0.018984f
C12503 MULT_0.4bit_ADDER_2.B3.n1 VSS 0.020472f
C12504 MULT_0.4bit_ADDER_2.B3.t8 VSS 0.014133f
C12505 MULT_0.4bit_ADDER_2.B3.n2 VSS 0.035861f
C12506 MULT_0.4bit_ADDER_2.B3.n3 VSS 0.062907f
C12507 MULT_0.4bit_ADDER_2.B3.t16 VSS 0.019275f
C12508 MULT_0.4bit_ADDER_2.B3.t7 VSS 0.038781f
C12509 MULT_0.4bit_ADDER_2.B3.t12 VSS 0.038299f
C12510 MULT_0.4bit_ADDER_2.B3.t17 VSS 0.038299f
C12511 MULT_0.4bit_ADDER_2.B3.t18 VSS 0.038299f
C12512 MULT_0.4bit_ADDER_2.B3.t10 VSS 0.007959f
C12513 MULT_0.4bit_ADDER_2.B3.t14 VSS 0.007959f
C12514 MULT_0.4bit_ADDER_2.B3.t11 VSS 0.007959f
C12515 MULT_0.4bit_ADDER_2.B3.n4 VSS 0.235956f
C12516 MULT_0.4bit_ADDER_2.B3.n5 VSS 0.173792f
C12517 MULT_0.4bit_ADDER_2.B3.n6 VSS 0.094715f
C12518 MULT_0.4bit_ADDER_2.B3.n7 VSS 0.09305f
C12519 MULT_0.4bit_ADDER_2.B3.n8 VSS 0.057236f
C12520 MULT_0.4bit_ADDER_2.B3.n9 VSS 0.075084f
C12521 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_0.A VSS 0.133526f
C12522 MULT_0.4bit_ADDER_2.B3.n10 VSS 0.83059f
C12523 MULT_0.4bit_ADDER_2.B3.t2 VSS 0.011355f
C12524 MULT_0.4bit_ADDER_2.B3.t0 VSS 0.011355f
C12525 MULT_0.4bit_ADDER_2.B3.n11 VSS 0.025334f
C12526 MULT_0.4bit_ADDER_2.B3.t6 VSS 0.011355f
C12527 MULT_0.4bit_ADDER_2.B3.t1 VSS 0.011355f
C12528 MULT_0.4bit_ADDER_2.B3.n12 VSS 0.025266f
C12529 MULT_0.4bit_ADDER_2.B3.t5 VSS 0.011355f
C12530 MULT_0.4bit_ADDER_2.B3.t4 VSS 0.011355f
C12531 MULT_0.4bit_ADDER_2.B3.n13 VSS 0.025266f
C12532 MULT_0.4bit_ADDER_2.B3.t3 VSS 0.068559f
C12533 MULT_0.4bit_ADDER_1.A2.n0 VSS 2.79153f
C12534 MULT_0.4bit_ADDER_1.A2.t3 VSS 0.065961f
C12535 MULT_0.4bit_ADDER_1.A2.t1 VSS 0.018184f
C12536 MULT_0.4bit_ADDER_1.A2.t2 VSS 0.018184f
C12537 MULT_0.4bit_ADDER_1.A2.n1 VSS 0.040543f
C12538 MULT_0.4bit_ADDER_1.A2.t0 VSS 0.052505f
C12539 MULT_0.4bit_ADDER_1.A2.t8 VSS 0.057355f
C12540 MULT_0.4bit_ADDER_1.A2.t11 VSS 0.022015f
C12541 MULT_0.4bit_ADDER_1.A2.t9 VSS 0.030403f
C12542 MULT_0.4bit_ADDER_1.A2.n2 VSS 0.034993f
C12543 MULT_0.4bit_ADDER_1.A2.t15 VSS 0.023141f
C12544 MULT_0.4bit_ADDER_1.A2.n3 VSS 0.035488f
C12545 MULT_0.4bit_ADDER_1.A2.t13 VSS 0.062107f
C12546 MULT_0.4bit_ADDER_1.A2.t10 VSS 0.061334f
C12547 MULT_0.4bit_ADDER_1.A2.t12 VSS 0.061334f
C12548 MULT_0.4bit_ADDER_1.A2.t7 VSS 0.061334f
C12549 MULT_0.4bit_ADDER_1.A2.n4 VSS 0.244128f
C12550 MULT_0.4bit_ADDER_1.A2.t5 VSS 0.012746f
C12551 MULT_0.4bit_ADDER_1.A2.t14 VSS 0.012746f
C12552 MULT_0.4bit_ADDER_1.A2.t6 VSS 0.012746f
C12553 MULT_0.4bit_ADDER_1.A2.t4 VSS 0.012746f
C12554 MULT_0.4bit_ADDER_1.A2.n5 VSS 0.23063f
C12555 MULT_0.4bit_ADDER_1.A2.n6 VSS 0.360752f
C12556 MULT_0.4bit_ADDER_1.A2.n7 VSS 0.852904f
C12557 mux8_2.NAND4F_8.Y.n0 VSS 0.539804f
C12558 mux8_2.NAND4F_8.Y.t13 VSS 0.026899f
C12559 mux8_2.NAND4F_8.Y.t14 VSS 0.028853f
C12560 mux8_2.NAND4F_8.Y.n1 VSS 0.042994f
C12561 mux8_2.NAND4F_8.Y.t12 VSS 0.026899f
C12562 mux8_2.NAND4F_8.Y.t11 VSS 0.026899f
C12563 mux8_2.NAND4F_8.Y.t10 VSS 0.026899f
C12564 mux8_2.NAND4F_8.Y.t9 VSS 0.033983f
C12565 mux8_2.NAND4F_8.Y.n2 VSS 0.072608f
C12566 mux8_2.NAND4F_8.Y.n3 VSS 0.045714f
C12567 mux8_2.NAND4F_8.Y.n4 VSS 0.037354f
C12568 mux8_2.NAND4F_8.Y.n5 VSS 0.018278f
C12569 mux8_2.NAND4F_8.Y.t5 VSS 0.026614f
C12570 mux8_2.NAND4F_8.Y.t4 VSS 0.026614f
C12571 mux8_2.NAND4F_8.Y.n6 VSS 0.0618f
C12572 mux8_2.NAND4F_8.Y.t8 VSS 0.026614f
C12573 mux8_2.NAND4F_8.Y.t0 VSS 0.026614f
C12574 mux8_2.NAND4F_8.Y.n7 VSS 0.061615f
C12575 mux8_2.NAND4F_8.Y.t7 VSS 0.026614f
C12576 mux8_2.NAND4F_8.Y.t6 VSS 0.026614f
C12577 mux8_2.NAND4F_8.Y.n8 VSS 0.061615f
C12578 mux8_2.NAND4F_8.Y.t2 VSS 0.026614f
C12579 mux8_2.NAND4F_8.Y.t1 VSS 0.026614f
C12580 mux8_2.NAND4F_8.Y.n9 VSS 0.061615f
C12581 mux8_2.NAND4F_8.Y.n10 VSS 0.268281f
C12582 mux8_2.NAND4F_8.Y.t3 VSS 0.21369f
C12583 XOR8_0.S3.t13 VSS 0.02459f
C12584 XOR8_0.S3.t12 VSS 0.072448f
C12585 XOR8_0.S3.t14 VSS 0.023924f
C12586 XOR8_0.S3.n0 VSS 0.123338f
C12587 XOR8_0.S3.t6 VSS 0.007161f
C12588 XOR8_0.S3.t7 VSS 0.007161f
C12589 XOR8_0.S3.n1 VSS 0.017319f
C12590 XOR8_0.S3.t4 VSS 0.007161f
C12591 XOR8_0.S3.t5 VSS 0.007161f
C12592 XOR8_0.S3.n2 VSS 0.017317f
C12593 XOR8_0.S3.n3 VSS 0.124178f
C12594 XOR8_0.S3.t8 VSS 0.007161f
C12595 XOR8_0.S3.t0 VSS 0.007161f
C12596 XOR8_0.S3.n4 VSS 0.014321f
C12597 XOR8_0.S3.n5 VSS 0.01125f
C12598 XOR8_0.S3.t9 VSS 0.030295f
C12599 XOR8_0.S3.t3 VSS 0.030295f
C12600 XOR8_0.S3.n6 VSS 0.06059f
C12601 XOR8_0.S3.n7 VSS 0.024035f
C12602 XOR8_0.S3.t10 VSS 0.030295f
C12603 XOR8_0.S3.t11 VSS 0.030295f
C12604 XOR8_0.S3.n8 VSS 0.06059f
C12605 XOR8_0.S3.n9 VSS 0.026649f
C12606 XOR8_0.S3.n10 VSS 0.274363f
C12607 XOR8_0.S3.t2 VSS 0.030295f
C12608 XOR8_0.S3.t1 VSS 0.030295f
C12609 XOR8_0.S3.n11 VSS 0.06059f
C12610 XOR8_0.S3.n12 VSS 0.026689f
C12611 XOR8_0.S3.n13 VSS 0.175964f
C12612 XOR8_0.S3.n14 VSS 0.039607f
C12613 XOR8_0.S3.n15 VSS 0.174162f
C12614 mux8_7.NAND4F_7.Y.n0 VSS 0.11858f
C12615 mux8_7.NAND4F_7.Y.n1 VSS 0.350455f
C12616 mux8_7.NAND4F_7.Y.t4 VSS 0.168166f
C12617 mux8_7.NAND4F_7.Y.t9 VSS 0.022537f
C12618 mux8_7.NAND4F_7.Y.t11 VSS 0.079785f
C12619 mux8_7.NAND4F_7.Y.t10 VSS 0.024808f
C12620 mux8_7.NAND4F_7.Y.n2 VSS 0.070768f
C12621 mux8_7.NAND4F_7.Y.n3 VSS 0.020978f
C12622 mux8_7.NAND4F_7.Y.t1 VSS 0.017278f
C12623 mux8_7.NAND4F_7.Y.t0 VSS 0.017278f
C12624 mux8_7.NAND4F_7.Y.n4 VSS 0.040122f
C12625 mux8_7.NAND4F_7.Y.t2 VSS 0.017278f
C12626 mux8_7.NAND4F_7.Y.t3 VSS 0.017278f
C12627 mux8_7.NAND4F_7.Y.n5 VSS 0.040002f
C12628 mux8_7.NAND4F_7.Y.t8 VSS 0.017278f
C12629 mux8_7.NAND4F_7.Y.t7 VSS 0.017278f
C12630 mux8_7.NAND4F_7.Y.n6 VSS 0.040002f
C12631 mux8_7.NAND4F_7.Y.t6 VSS 0.017278f
C12632 mux8_7.NAND4F_7.Y.t5 VSS 0.017278f
C12633 mux8_7.NAND4F_7.Y.n7 VSS 0.040002f
C12634 NOT8_0.S5.n0 VSS 1.86445f
C12635 NOT8_0.S5.t5 VSS 0.090185f
C12636 NOT8_0.S5.t4 VSS 0.265712f
C12637 NOT8_0.S5.t6 VSS 0.087744f
C12638 NOT8_0.S5.n1 VSS 0.452384f
C12639 NOT8_0.S5.t0 VSS 0.043232f
C12640 NOT8_0.S5.t2 VSS 0.043232f
C12641 NOT8_0.S5.n2 VSS 0.09634f
C12642 NOT8_0.S5.t3 VSS 0.156803f
C12643 NOT8_0.S5.t1 VSS 0.124696f
C12644 a_5197_5532.n0 VSS 1.48326f
C12645 a_5197_5532.n1 VSS 1.48365f
C12646 a_5197_5532.t4 VSS 0.093341f
C12647 a_5197_5532.t8 VSS 0.093341f
C12648 a_5197_5532.t9 VSS 0.093341f
C12649 a_5197_5532.n2 VSS 0.202296f
C12650 a_5197_5532.t7 VSS 0.093341f
C12651 a_5197_5532.t5 VSS 0.093341f
C12652 a_5197_5532.n3 VSS 0.202001f
C12653 a_5197_5532.t10 VSS 0.093341f
C12654 a_5197_5532.t11 VSS 0.093341f
C12655 a_5197_5532.n4 VSS 0.20269f
C12656 a_5197_5532.t1 VSS 0.093341f
C12657 a_5197_5532.t3 VSS 0.093341f
C12658 a_5197_5532.n5 VSS 0.202001f
C12659 a_5197_5532.t2 VSS 0.093341f
C12660 a_5197_5532.t0 VSS 0.093341f
C12661 a_5197_5532.n6 VSS 0.202001f
C12662 a_5197_5532.n7 VSS 0.202001f
C12663 a_5197_5532.t6 VSS 0.093341f
C12664 V_FLAG_0.XOR2_0.Y.t13 VSS 0.053228f
C12665 V_FLAG_0.XOR2_0.Y.t15 VSS 0.017333f
C12666 V_FLAG_0.XOR2_0.Y.t14 VSS 0.023937f
C12667 V_FLAG_0.XOR2_0.Y.n0 VSS 0.025813f
C12668 V_FLAG_0.XOR2_0.Y.t12 VSS 0.01782f
C12669 V_FLAG_0.XOR2_0.Y.n1 VSS 0.045216f
C12670 V_FLAG_0.XOR2_0.Y.n2 VSS 0.07946f
C12671 V_FLAG_0.XOR2_0.Y.t11 VSS 0.008697f
C12672 V_FLAG_0.XOR2_0.Y.t6 VSS 0.008697f
C12673 V_FLAG_0.XOR2_0.Y.n3 VSS 0.021035f
C12674 V_FLAG_0.XOR2_0.Y.t5 VSS 0.008697f
C12675 V_FLAG_0.XOR2_0.Y.t0 VSS 0.008697f
C12676 V_FLAG_0.XOR2_0.Y.n4 VSS 0.021032f
C12677 V_FLAG_0.XOR2_0.Y.n5 VSS 0.150821f
C12678 V_FLAG_0.XOR2_0.Y.t10 VSS 0.008697f
C12679 V_FLAG_0.XOR2_0.Y.t2 VSS 0.008697f
C12680 V_FLAG_0.XOR2_0.Y.n6 VSS 0.017394f
C12681 V_FLAG_0.XOR2_0.Y.n7 VSS 0.013663f
C12682 V_FLAG_0.XOR2_0.Y.t9 VSS 0.036795f
C12683 V_FLAG_0.XOR2_0.Y.t4 VSS 0.036795f
C12684 V_FLAG_0.XOR2_0.Y.n8 VSS 0.07359f
C12685 V_FLAG_0.XOR2_0.Y.n9 VSS 0.029261f
C12686 V_FLAG_0.XOR2_0.Y.t8 VSS 0.036795f
C12687 V_FLAG_0.XOR2_0.Y.t7 VSS 0.036795f
C12688 V_FLAG_0.XOR2_0.Y.n10 VSS 0.07359f
C12689 V_FLAG_0.XOR2_0.Y.n11 VSS 0.032366f
C12690 V_FLAG_0.XOR2_0.Y.n12 VSS 0.333229f
C12691 V_FLAG_0.XOR2_0.Y.t1 VSS 0.036795f
C12692 V_FLAG_0.XOR2_0.Y.t3 VSS 0.036795f
C12693 V_FLAG_0.XOR2_0.Y.n13 VSS 0.07359f
C12694 V_FLAG_0.XOR2_0.Y.n14 VSS 0.032415f
C12695 V_FLAG_0.XOR2_0.Y.n15 VSS 0.213718f
C12696 V_FLAG_0.XOR2_0.Y.n16 VSS 0.048164f
C12697 V_FLAG_0.XOR2_0.Y.n17 VSS 0.211401f
C12698 XOR8_0.S4.t13 VSS 0.048734f
C12699 XOR8_0.S4.t12 VSS 0.143586f
C12700 XOR8_0.S4.t14 VSS 0.047415f
C12701 XOR8_0.S4.n0 VSS 0.244444f
C12702 XOR8_0.S4.t3 VSS 0.014192f
C12703 XOR8_0.S4.t5 VSS 0.014192f
C12704 XOR8_0.S4.n1 VSS 0.034325f
C12705 XOR8_0.S4.t9 VSS 0.014192f
C12706 XOR8_0.S4.t11 VSS 0.014192f
C12707 XOR8_0.S4.n2 VSS 0.034321f
C12708 XOR8_0.S4.n3 VSS 0.24611f
C12709 XOR8_0.S4.t4 VSS 0.014192f
C12710 XOR8_0.S4.t10 VSS 0.014192f
C12711 XOR8_0.S4.n4 VSS 0.028384f
C12712 XOR8_0.S4.n5 VSS 0.022296f
C12713 XOR8_0.S4.t2 VSS 0.060042f
C12714 XOR8_0.S4.t6 VSS 0.060042f
C12715 XOR8_0.S4.n6 VSS 0.120084f
C12716 XOR8_0.S4.n7 VSS 0.047635f
C12717 XOR8_0.S4.t0 VSS 0.060042f
C12718 XOR8_0.S4.t1 VSS 0.060042f
C12719 XOR8_0.S4.n8 VSS 0.120084f
C12720 XOR8_0.S4.n9 VSS 0.052815f
C12721 XOR8_0.S4.n10 VSS 0.543762f
C12722 XOR8_0.S4.t8 VSS 0.060042f
C12723 XOR8_0.S4.t7 VSS 0.060042f
C12724 XOR8_0.S4.n11 VSS 0.120084f
C12725 XOR8_0.S4.n12 VSS 0.052895f
C12726 XOR8_0.S4.n13 VSS 0.348745f
C12727 XOR8_0.S4.n14 VSS 0.078497f
C12728 XOR8_0.S4.n15 VSS 0.345173f
C12729 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t5 VSS 0.007073f
C12730 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t3 VSS 0.007073f
C12731 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n0 VSS 0.017105f
C12732 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t9 VSS 0.007073f
C12733 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t11 VSS 0.007073f
C12734 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n1 VSS 0.017107f
C12735 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n2 VSS 0.122656f
C12736 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t7 VSS 0.007073f
C12737 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t10 VSS 0.007073f
C12738 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n3 VSS 0.014146f
C12739 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n4 VSS 0.011112f
C12740 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t8 VSS 0.029924f
C12741 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t0 VSS 0.029924f
C12742 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n5 VSS 0.059848f
C12743 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n6 VSS 0.023796f
C12744 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t6 VSS 0.029924f
C12745 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t4 VSS 0.029924f
C12746 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n7 VSS 0.059848f
C12747 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n8 VSS 0.026362f
C12748 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n9 VSS 0.271f
C12749 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t1 VSS 0.029924f
C12750 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t2 VSS 0.029924f
C12751 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n10 VSS 0.059848f
C12752 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n11 VSS 0.026322f
C12753 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n12 VSS 0.173808f
C12754 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n13 VSS 0.03917f
C12755 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n14 VSS 0.172104f
C12756 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t16 VSS 0.043288f
C12757 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t12 VSS 0.014096f
C12758 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t13 VSS 0.019467f
C12759 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n15 VSS 0.020992f
C12760 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t14 VSS 0.014492f
C12761 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n16 VSS 0.036772f
C12762 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n17 VSS 0.064505f
C12763 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t20 VSS 0.019764f
C12764 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t23 VSS 0.039767f
C12765 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t22 VSS 0.039272f
C12766 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t17 VSS 0.039272f
C12767 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t18 VSS 0.039272f
C12768 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t19 VSS 0.008161f
C12769 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t15 VSS 0.008161f
C12770 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.t21 VSS 0.008161f
C12771 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n18 VSS 0.24195f
C12772 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n19 VSS 0.178207f
C12773 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n20 VSS 0.097121f
C12774 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n21 VSS 0.095413f
C12775 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n22 VSS 0.05869f
C12776 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n23 VSS 0.076991f
C12777 8bit_ADDER_0.FULL_ADDER_XORED_6.XOR2_2.Y.n24 VSS 1.26966f
C12778 a_n4205_3810.n0 VSS 2.91093f
C12779 a_n4205_3810.t1 VSS 0.09158f
C12780 a_n4205_3810.t11 VSS 0.09158f
C12781 a_n4205_3810.t10 VSS 0.09158f
C12782 a_n4205_3810.n1 VSS 0.198865f
C12783 a_n4205_3810.t9 VSS 0.09158f
C12784 a_n4205_3810.t4 VSS 0.09158f
C12785 a_n4205_3810.n2 VSS 0.19819f
C12786 a_n4205_3810.t3 VSS 0.09158f
C12787 a_n4205_3810.t5 VSS 0.09158f
C12788 a_n4205_3810.n3 VSS 0.19819f
C12789 a_n4205_3810.t8 VSS 0.09158f
C12790 a_n4205_3810.t7 VSS 0.09158f
C12791 a_n4205_3810.n4 VSS 0.198479f
C12792 a_n4205_3810.t2 VSS 0.09158f
C12793 a_n4205_3810.t6 VSS 0.09158f
C12794 a_n4205_3810.n5 VSS 0.19819f
C12795 a_n4205_3810.n6 VSS 0.19819f
C12796 a_n4205_3810.t0 VSS 0.09158f
C12797 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n0 VSS 0.967969f
C12798 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t2 VSS 0.008375f
C12799 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t1 VSS 0.008375f
C12800 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n1 VSS 0.018636f
C12801 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t5 VSS 0.008375f
C12802 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t6 VSS 0.008375f
C12803 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n2 VSS 0.018687f
C12804 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t3 VSS 0.008375f
C12805 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t4 VSS 0.008375f
C12806 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n3 VSS 0.018636f
C12807 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t0 VSS 0.05057f
C12808 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t17 VSS 0.028606f
C12809 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t13 VSS 0.02825f
C12810 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t14 VSS 0.02825f
C12811 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t9 VSS 0.02825f
C12812 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n4 VSS 0.112442f
C12813 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t7 VSS 0.005871f
C12814 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t15 VSS 0.005871f
C12815 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t12 VSS 0.005871f
C12816 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t18 VSS 0.005871f
C12817 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n5 VSS 0.106225f
C12818 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n6 VSS 0.166131f
C12819 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t16 VSS 0.026417f
C12820 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t11 VSS 0.01014f
C12821 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t8 VSS 0.014003f
C12822 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n7 VSS 0.016118f
C12823 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.t10 VSS 0.010659f
C12824 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n8 VSS 0.016345f
C12825 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n9 VSS 0.055518f
C12826 MULT_0.4bit_ADDER_1.FULL_ADDER_1.COUT.n10 VSS 0.369194f
C12827 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t16 VSS 0.013766f
C12828 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t19 VSS 0.027698f
C12829 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t12 VSS 0.027354f
C12830 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t23 VSS 0.027354f
C12831 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t18 VSS 0.027354f
C12832 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t21 VSS 0.005684f
C12833 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t15 VSS 0.005684f
C12834 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t17 VSS 0.005684f
C12835 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n0 VSS 0.168523f
C12836 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n1 VSS 0.124125f
C12837 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n2 VSS 0.067647f
C12838 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n3 VSS 0.066457f
C12839 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n4 VSS 0.040879f
C12840 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n5 VSS 0.05311f
C12841 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t22 VSS 0.030151f
C12842 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t14 VSS 0.009818f
C12843 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t13 VSS 0.013559f
C12844 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n6 VSS 0.014622f
C12845 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t20 VSS 0.010094f
C12846 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n7 VSS 0.025612f
C12847 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n8 VSS 0.044927f
C12848 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t0 VSS 0.004926f
C12849 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t1 VSS 0.004926f
C12850 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n9 VSS 0.011915f
C12851 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t9 VSS 0.004926f
C12852 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t11 VSS 0.004926f
C12853 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n10 VSS 0.011914f
C12854 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n11 VSS 0.085433f
C12855 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t2 VSS 0.004926f
C12856 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t10 VSS 0.004926f
C12857 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n12 VSS 0.009853f
C12858 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n13 VSS 0.00774f
C12859 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t5 VSS 0.020843f
C12860 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t7 VSS 0.020843f
C12861 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n14 VSS 0.041685f
C12862 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n15 VSS 0.016575f
C12863 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t3 VSS 0.020843f
C12864 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t4 VSS 0.020843f
C12865 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n16 VSS 0.041685f
C12866 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n17 VSS 0.018334f
C12867 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n18 VSS 0.188757f
C12868 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t6 VSS 0.020843f
C12869 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.t8 VSS 0.020843f
C12870 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n19 VSS 0.041685f
C12871 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n20 VSS 0.018362f
C12872 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n21 VSS 0.12106f
C12873 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n22 VSS 0.027282f
C12874 MULT_0.4bit_ADDER_0.FULL_ADDER_2.XOR2_1.A.n23 VSS 0.119748f
C12875 B6.t2 VSS 0.054102f
C12876 B6.t6 VSS 0.075522f
C12877 B6.t5 VSS 0.075522f
C12878 B6.n0 VSS 0.245841f
C12879 B6.t30 VSS 0.086665f
C12880 B6.n1 VSS 0.612913f
C12881 B6.t36 VSS 0.072063f
C12882 B6.t4 VSS 0.144993f
C12883 B6.t24 VSS 0.14319f
C12884 B6.t7 VSS 0.14319f
C12885 B6.t32 VSS 0.14319f
C12886 B6.t10 VSS 0.029756f
C12887 B6.t26 VSS 0.029756f
C12888 B6.t18 VSS 0.029756f
C12889 B6.n2 VSS 0.882176f
C12890 B6.n3 VSS 0.649763f
C12891 B6.n4 VSS 0.354115f
C12892 B6.n5 VSS 0.347888f
C12893 B6.n6 VSS 0.213991f
C12894 B6.n7 VSS 0.243351f
C12895 B6.t0 VSS 0.158014f
C12896 B6.t15 VSS 0.067673f
C12897 B6.t25 VSS 0.054102f
C12898 B6.n8 VSS 0.079845f
C12899 B6.t34 VSS 0.05284f
C12900 B6.n9 VSS 0.131811f
C12901 B6.n10 VSS 0.235163f
C12902 B6.n11 VSS 0.372034f
C12903 B6.n12 VSS 3.58477f
C12904 B6.t11 VSS 0.064562f
C12905 B6.t9 VSS 0.069251f
C12906 B6.n13 VSS 0.10319f
C12907 B6.t14 VSS 0.064562f
C12908 B6.t22 VSS 0.064562f
C12909 B6.t23 VSS 0.064562f
C12910 B6.t33 VSS 0.081564f
C12911 B6.n14 VSS 0.174267f
C12912 B6.n15 VSS 0.109719f
C12913 B6.n16 VSS 0.089653f
C12914 B6.n17 VSS 0.04387f
C12915 B6.n18 VSS 9.239889f
C12916 B6.t28 VSS 0.072063f
C12917 B6.t13 VSS 0.144993f
C12918 B6.t21 VSS 0.14319f
C12919 B6.t12 VSS 0.14319f
C12920 B6.t31 VSS 0.14319f
C12921 B6.t35 VSS 0.029756f
C12922 B6.t17 VSS 0.029756f
C12923 B6.t1 VSS 0.029756f
C12924 B6.n19 VSS 0.881954f
C12925 B6.n20 VSS 0.649985f
C12926 B6.n21 VSS 0.354115f
C12927 B6.n22 VSS 0.347888f
C12928 B6.n23 VSS 0.213991f
C12929 B6.n24 VSS 0.275365f
C12930 B6.n25 VSS 13.500099f
C12931 B6.t29 VSS 0.054102f
C12932 B6.t16 VSS 0.075522f
C12933 B6.t27 VSS 0.075522f
C12934 B6.n26 VSS 0.245841f
C12935 B6.t8 VSS 0.086665f
C12936 B6.n27 VSS 0.736827f
C12937 B6.n28 VSS 0.462579f
C12938 B6.n29 VSS 9.588349f
C12939 B6.t3 VSS 0.054102f
C12940 B6.t20 VSS 0.075522f
C12941 B6.t37 VSS 0.075522f
C12942 B6.n30 VSS 0.245841f
C12943 B6.t19 VSS 0.086665f
C12944 B6.n31 VSS 0.612032f
C12945 B6.n32 VSS 0.544986f
C12946 B6.n33 VSS 4.3009f
C12947 B6.n34 VSS 0.707456f
C12948 a_n10684_n11063.n0 VSS 1.48326f
C12949 a_n10684_n11063.n1 VSS 1.48365f
C12950 a_n10684_n11063.t5 VSS 0.093341f
C12951 a_n10684_n11063.t8 VSS 0.093341f
C12952 a_n10684_n11063.t7 VSS 0.093341f
C12953 a_n10684_n11063.n2 VSS 0.20269f
C12954 a_n10684_n11063.t2 VSS 0.093341f
C12955 a_n10684_n11063.t0 VSS 0.093341f
C12956 a_n10684_n11063.n3 VSS 0.202001f
C12957 a_n10684_n11063.t1 VSS 0.093341f
C12958 a_n10684_n11063.t3 VSS 0.093341f
C12959 a_n10684_n11063.n4 VSS 0.202001f
C12960 a_n10684_n11063.t10 VSS 0.093341f
C12961 a_n10684_n11063.t9 VSS 0.093341f
C12962 a_n10684_n11063.n5 VSS 0.202001f
C12963 a_n10684_n11063.t4 VSS 0.093341f
C12964 a_n10684_n11063.t11 VSS 0.093341f
C12965 a_n10684_n11063.n6 VSS 0.202001f
C12966 a_n10684_n11063.n7 VSS 0.202296f
C12967 a_n10684_n11063.t6 VSS 0.093341f
C12968 MULT_0.4bit_ADDER_2.FULL_ADDER_3.NAND2_0.B VSS 0.676675f
C12969 MULT_0.inv_8.Y.n0 VSS 4.05379f
C12970 MULT_0.4bit_ADDER_2.FULL_ADDER_3.XOR2_0.B VSS 0.713054f
C12971 MULT_0.4bit_ADDER_2.FULL_ADDER_3.A VSS 2.89793f
C12972 MULT_0.inv_8.Y.t12 VSS 0.054322f
C12973 MULT_0.inv_8.Y.t10 VSS 0.020851f
C12974 MULT_0.inv_8.Y.t13 VSS 0.028795f
C12975 MULT_0.inv_8.Y.n1 VSS 0.033143f
C12976 MULT_0.inv_8.Y.t7 VSS 0.021918f
C12977 MULT_0.inv_8.Y.n2 VSS 0.033612f
C12978 MULT_0.inv_8.Y.t9 VSS 0.058823f
C12979 MULT_0.inv_8.Y.t4 VSS 0.058091f
C12980 MULT_0.inv_8.Y.t11 VSS 0.058091f
C12981 MULT_0.inv_8.Y.t5 VSS 0.058091f
C12982 MULT_0.inv_8.Y.n3 VSS 0.231219f
C12983 MULT_0.inv_8.Y.t8 VSS 0.012072f
C12984 MULT_0.inv_8.Y.t15 VSS 0.012072f
C12985 MULT_0.inv_8.Y.t6 VSS 0.012072f
C12986 MULT_0.inv_8.Y.t14 VSS 0.012072f
C12987 MULT_0.inv_8.Y.n4 VSS 0.218435f
C12988 MULT_0.inv_8.Y.n5 VSS 0.341676f
C12989 MULT_0.inv_8.Y.n6 VSS 0.808123f
C12990 MULT_0.inv_8.Y.t0 VSS 0.017222f
C12991 MULT_0.inv_8.Y.t2 VSS 0.017222f
C12992 MULT_0.inv_8.Y.n7 VSS 0.038274f
C12993 MULT_0.inv_8.Y.t1 VSS 0.049889f
C12994 MULT_0.inv_8.Y.t3 VSS 0.062466f
C12995 B4.t2 VSS 0.051354f
C12996 B4.t7 VSS 0.071686f
C12997 B4.t6 VSS 0.071686f
C12998 B4.n0 VSS 0.233354f
C12999 B4.t30 VSS 0.082263f
C13000 B4.n1 VSS 0.571631f
C13001 B4.n2 VSS 0.653605f
C13002 B4.t35 VSS 0.051354f
C13003 B4.t13 VSS 0.071686f
C13004 B4.t32 VSS 0.071686f
C13005 B4.n3 VSS 0.233354f
C13006 B4.t12 VSS 0.082263f
C13007 B4.n4 VSS 0.569297f
C13008 B4.n5 VSS 0.501485f
C13009 B4.n6 VSS 3.21737f
C13010 B4.t11 VSS 0.051354f
C13011 B4.t31 VSS 0.071686f
C13012 B4.t29 VSS 0.071686f
C13013 B4.n7 VSS 0.233354f
C13014 B4.t23 VSS 0.082263f
C13015 B4.n8 VSS 0.706076f
C13016 B4.n9 VSS 0.417897f
C13017 B4.n10 VSS 6.02383f
C13018 B4.t21 VSS 0.068403f
C13019 B4.t0 VSS 0.137629f
C13020 B4.t4 VSS 0.135917f
C13021 B4.t37 VSS 0.135917f
C13022 B4.t26 VSS 0.135917f
C13023 B4.t36 VSS 0.028245f
C13024 B4.t17 VSS 0.028245f
C13025 B4.t1 VSS 0.028245f
C13026 B4.n11 VSS 0.837158f
C13027 B4.n12 VSS 0.616971f
C13028 B4.n13 VSS 0.336129f
C13029 B4.n14 VSS 0.330218f
C13030 B4.n15 VSS 0.203122f
C13031 B4.n16 VSS 0.261379f
C13032 B4.n17 VSS 8.539599f
C13033 B4.t27 VSS 0.061283f
C13034 B4.t25 VSS 0.065733f
C13035 B4.n18 VSS 0.097949f
C13036 B4.t28 VSS 0.061283f
C13037 B4.t5 VSS 0.061283f
C13038 B4.t8 VSS 0.061283f
C13039 B4.t19 VSS 0.077421f
C13040 B4.n19 VSS 0.165415f
C13041 B4.n20 VSS 0.104146f
C13042 B4.n21 VSS 0.085099f
C13043 B4.n22 VSS 0.041642f
C13044 B4.n23 VSS 6.85914f
C13045 B4.t15 VSS 0.068403f
C13046 B4.t18 VSS 0.137629f
C13047 B4.t22 VSS 0.135917f
C13048 B4.t3 VSS 0.135917f
C13049 B4.t34 VSS 0.135917f
C13050 B4.t24 VSS 0.028245f
C13051 B4.t16 VSS 0.028245f
C13052 B4.t10 VSS 0.028245f
C13053 B4.n24 VSS 0.837369f
C13054 B4.n25 VSS 0.61676f
C13055 B4.n26 VSS 0.336129f
C13056 B4.n27 VSS 0.330218f
C13057 B4.n28 VSS 0.203122f
C13058 B4.n29 VSS 0.230991f
C13059 B4.t14 VSS 0.149988f
C13060 B4.t20 VSS 0.064236f
C13061 B4.t33 VSS 0.051354f
C13062 B4.n30 VSS 0.07579f
C13063 B4.t9 VSS 0.050156f
C13064 B4.n31 VSS 0.125116f
C13065 B4.n32 VSS 0.223218f
C13066 B4.n33 VSS 0.340222f
C13067 B4.n34 VSS 23.331598f
C13068 B4.n35 VSS 3.23022f
C13069 mux8_4.NAND4F_7.Y.n0 VSS 0.11858f
C13070 mux8_4.NAND4F_7.Y.n1 VSS 0.350455f
C13071 mux8_4.NAND4F_7.Y.t2 VSS 0.168166f
C13072 mux8_4.NAND4F_7.Y.t9 VSS 0.022537f
C13073 mux8_4.NAND4F_7.Y.t11 VSS 0.079785f
C13074 mux8_4.NAND4F_7.Y.t10 VSS 0.024808f
C13075 mux8_4.NAND4F_7.Y.n2 VSS 0.070768f
C13076 mux8_4.NAND4F_7.Y.n3 VSS 0.020978f
C13077 mux8_4.NAND4F_7.Y.t1 VSS 0.017278f
C13078 mux8_4.NAND4F_7.Y.t0 VSS 0.017278f
C13079 mux8_4.NAND4F_7.Y.n4 VSS 0.040122f
C13080 mux8_4.NAND4F_7.Y.t7 VSS 0.017278f
C13081 mux8_4.NAND4F_7.Y.t8 VSS 0.017278f
C13082 mux8_4.NAND4F_7.Y.n5 VSS 0.040002f
C13083 mux8_4.NAND4F_7.Y.t6 VSS 0.017278f
C13084 mux8_4.NAND4F_7.Y.t5 VSS 0.017278f
C13085 mux8_4.NAND4F_7.Y.n6 VSS 0.040002f
C13086 mux8_4.NAND4F_7.Y.t3 VSS 0.017278f
C13087 mux8_4.NAND4F_7.Y.t4 VSS 0.017278f
C13088 mux8_4.NAND4F_7.Y.n7 VSS 0.040002f
C13089 NOT8_0.S3.n0 VSS 1.59359f
C13090 NOT8_0.S3.t6 VSS 0.077083f
C13091 NOT8_0.S3.t5 VSS 0.22711f
C13092 NOT8_0.S3.t4 VSS 0.074997f
C13093 NOT8_0.S3.n1 VSS 0.386662f
C13094 NOT8_0.S3.t2 VSS 0.036952f
C13095 NOT8_0.S3.t0 VSS 0.036952f
C13096 NOT8_0.S3.n2 VSS 0.082344f
C13097 NOT8_0.S3.t1 VSS 0.134023f
C13098 NOT8_0.S3.t3 VSS 0.10658f
C13099 mux8_5.NAND4F_3.Y.n0 VSS 0.306333f
C13100 mux8_5.NAND4F_3.Y.t2 VSS 0.015103f
C13101 mux8_5.NAND4F_3.Y.t3 VSS 0.015103f
C13102 mux8_5.NAND4F_3.Y.n1 VSS 0.035071f
C13103 mux8_5.NAND4F_3.Y.t0 VSS 0.015103f
C13104 mux8_5.NAND4F_3.Y.t1 VSS 0.015103f
C13105 mux8_5.NAND4F_3.Y.n2 VSS 0.034966f
C13106 mux8_5.NAND4F_3.Y.t4 VSS 0.015103f
C13107 mux8_5.NAND4F_3.Y.t5 VSS 0.015103f
C13108 mux8_5.NAND4F_3.Y.n3 VSS 0.034966f
C13109 mux8_5.NAND4F_3.Y.t6 VSS 0.015103f
C13110 mux8_5.NAND4F_3.Y.t7 VSS 0.015103f
C13111 mux8_5.NAND4F_3.Y.n4 VSS 0.034966f
C13112 mux8_5.NAND4F_3.Y.n5 VSS 0.152246f
C13113 mux8_5.NAND4F_3.Y.t8 VSS 0.143521f
C13114 mux8_5.NAND4F_3.Y.t9 VSS 0.0197f
C13115 mux8_5.NAND4F_3.Y.t10 VSS 0.0197f
C13116 mux8_5.NAND4F_3.Y.n6 VSS 0.023128f
C13117 mux8_5.NAND4F_3.Y.t11 VSS 0.061756f
C13118 mux8_5.NAND4F_3.Y.n7 VSS 0.129679f
C13119 mux8_5.NAND4F_0.C.n0 VSS 1.72379f
C13120 mux8_5.NAND4F_0.C.t14 VSS 0.238621f
C13121 mux8_5.NAND4F_0.C.t10 VSS 0.076118f
C13122 mux8_5.NAND4F_0.C.t8 VSS 0.076118f
C13123 mux8_5.NAND4F_0.C.n1 VSS 0.089365f
C13124 mux8_5.NAND4F_0.C.n2 VSS 0.501052f
C13125 mux8_5.NAND4F_0.C.t9 VSS 0.076118f
C13126 mux8_5.NAND4F_0.C.t11 VSS 0.076118f
C13127 mux8_5.NAND4F_0.C.n3 VSS 0.089365f
C13128 mux8_5.NAND4F_0.C.t12 VSS 0.238621f
C13129 mux8_5.NAND4F_0.C.n4 VSS 0.501084f
C13130 mux8_5.NAND4F_0.C.t15 VSS 0.076118f
C13131 mux8_5.NAND4F_0.C.t4 VSS 0.076118f
C13132 mux8_5.NAND4F_0.C.n5 VSS 0.089365f
C13133 mux8_5.NAND4F_0.C.t5 VSS 0.238621f
C13134 mux8_5.NAND4F_0.C.n6 VSS 0.501098f
C13135 mux8_5.NAND4F_0.C.n7 VSS 1.82754f
C13136 mux8_5.NAND4F_0.C.t1 VSS 0.038784f
C13137 mux8_5.NAND4F_0.C.t3 VSS 0.038784f
C13138 mux8_5.NAND4F_0.C.n8 VSS 0.086427f
C13139 mux8_5.NAND4F_0.C.t2 VSS 0.140669f
C13140 mux8_5.NAND4F_0.C.t0 VSS 0.111866f
C13141 mux8_5.NAND4F_0.C.n9 VSS 3.19968f
C13142 mux8_5.NAND4F_0.C.t13 VSS 0.238621f
C13143 mux8_5.NAND4F_0.C.t7 VSS 0.076118f
C13144 mux8_5.NAND4F_0.C.t6 VSS 0.076118f
C13145 mux8_5.NAND4F_0.C.n10 VSS 0.089365f
C13146 mux8_5.NAND4F_0.C.n11 VSS 0.50107f
C13147 mux8_5.NAND4F_0.C.n12 VSS 2.56421f
C13148 MULT_0.inv_9.Y.t5 VSS 0.065569f
C13149 MULT_0.inv_9.Y.t4 VSS 0.025168f
C13150 MULT_0.inv_9.Y.t7 VSS 0.034757f
C13151 MULT_0.inv_9.Y.n0 VSS 0.040005f
C13152 MULT_0.inv_9.Y.t14 VSS 0.026455f
C13153 MULT_0.inv_9.Y.n1 VSS 0.04057f
C13154 MULT_0.inv_9.Y.n2 VSS 0.167931f
C13155 MULT_0.inv_9.Y.t12 VSS 0.071001f
C13156 MULT_0.inv_9.Y.t11 VSS 0.070118f
C13157 MULT_0.inv_9.Y.t10 VSS 0.070118f
C13158 MULT_0.inv_9.Y.t15 VSS 0.070118f
C13159 MULT_0.inv_9.Y.n3 VSS 0.279089f
C13160 MULT_0.inv_9.Y.t6 VSS 0.014571f
C13161 MULT_0.inv_9.Y.t13 VSS 0.014571f
C13162 MULT_0.inv_9.Y.t9 VSS 0.014571f
C13163 MULT_0.inv_9.Y.t8 VSS 0.014571f
C13164 MULT_0.inv_9.Y.n4 VSS 0.263659f
C13165 MULT_0.inv_9.Y.n5 VSS 0.412415f
C13166 MULT_0.inv_9.Y.n6 VSS 0.974543f
C13167 MULT_0.inv_9.Y.t1 VSS 0.075398f
C13168 MULT_0.inv_9.Y.t0 VSS 0.060083f
C13169 MULT_0.inv_9.Y.t3 VSS 0.020788f
C13170 MULT_0.inv_9.Y.t2 VSS 0.020788f
C13171 MULT_0.inv_9.Y.n7 VSS 0.046198f
C13172 mux8_4.NAND4F_5.Y.n0 VSS 0.25108f
C13173 mux8_4.NAND4F_5.Y.t10 VSS 0.017162f
C13174 mux8_4.NAND4F_5.Y.t9 VSS 0.050565f
C13175 mux8_4.NAND4F_5.Y.t11 VSS 0.016698f
C13176 mux8_4.NAND4F_5.Y.n1 VSS 0.086077f
C13177 mux8_4.NAND4F_5.Y.t2 VSS 0.099394f
C13178 mux8_4.NAND4F_5.Y.n2 VSS 0.798124f
C13179 mux8_4.NAND4F_5.Y.t0 VSS 0.012379f
C13180 mux8_4.NAND4F_5.Y.t1 VSS 0.012379f
C13181 mux8_4.NAND4F_5.Y.n3 VSS 0.028745f
C13182 mux8_4.NAND4F_5.Y.t6 VSS 0.012379f
C13183 mux8_4.NAND4F_5.Y.t5 VSS 0.012379f
C13184 mux8_4.NAND4F_5.Y.n4 VSS 0.028659f
C13185 mux8_4.NAND4F_5.Y.t7 VSS 0.012379f
C13186 mux8_4.NAND4F_5.Y.t8 VSS 0.012379f
C13187 mux8_4.NAND4F_5.Y.n5 VSS 0.028659f
C13188 mux8_4.NAND4F_5.Y.t3 VSS 0.012379f
C13189 mux8_4.NAND4F_5.Y.t4 VSS 0.012379f
C13190 mux8_4.NAND4F_5.Y.n6 VSS 0.028659f
C13191 mux8_4.NAND4F_5.Y.n7 VSS 0.117805f
C13192 SEL2.t18 VSS 0.025525f
C13193 SEL2.t9 VSS 0.035631f
C13194 SEL2.t48 VSS 0.035631f
C13195 SEL2.n0 VSS 0.1116f
C13196 SEL2.t75 VSS 0.039019f
C13197 SEL2.t107 VSS 0.039309f
C13198 SEL2.t77 VSS 0.139158f
C13199 SEL2.t59 VSS 0.04327f
C13200 SEL2.n1 VSS 0.123432f
C13201 SEL2.n2 VSS 0.036589f
C13202 SEL2.t39 VSS 0.039309f
C13203 SEL2.t58 VSS 0.139158f
C13204 SEL2.t36 VSS 0.04327f
C13205 SEL2.n3 VSS 0.123432f
C13206 SEL2.n4 VSS 0.036555f
C13207 SEL2.n5 VSS 0.087144f
C13208 SEL2.t65 VSS 0.039309f
C13209 SEL2.t33 VSS 0.139158f
C13210 SEL2.t53 VSS 0.04327f
C13211 SEL2.n6 VSS 0.123432f
C13212 SEL2.n7 VSS 0.036571f
C13213 SEL2.n8 VSS 0.05726f
C13214 SEL2.n9 VSS 0.52738f
C13215 SEL2.t91 VSS 0.039309f
C13216 SEL2.t130 VSS 0.139158f
C13217 SEL2.t83 VSS 0.04327f
C13218 SEL2.n10 VSS 0.123432f
C13219 SEL2.n11 VSS 0.036567f
C13220 SEL2.n12 VSS 0.055954f
C13221 SEL2.n13 VSS 0.56381f
C13222 SEL2.n14 VSS 0.893698f
C13223 SEL2.n15 VSS 0.905768f
C13224 SEL2.n16 VSS 0.079769f
C13225 SEL2.n17 VSS 0.086502f
C13226 SEL2.n18 VSS 0.080015f
C13227 SEL2.n19 VSS 0.534409f
C13228 SEL2.t16 VSS 0.025525f
C13229 SEL2.t110 VSS 0.035631f
C13230 SEL2.t26 VSS 0.035631f
C13231 SEL2.n20 VSS 0.1116f
C13232 SEL2.t85 VSS 0.039019f
C13233 SEL2.t3 VSS 0.039309f
C13234 SEL2.t123 VSS 0.139158f
C13235 SEL2.t101 VSS 0.04327f
C13236 SEL2.n21 VSS 0.123432f
C13237 SEL2.n22 VSS 0.036589f
C13238 SEL2.t129 VSS 0.039309f
C13239 SEL2.t99 VSS 0.139158f
C13240 SEL2.t116 VSS 0.04327f
C13241 SEL2.n23 VSS 0.123432f
C13242 SEL2.n24 VSS 0.036555f
C13243 SEL2.n25 VSS 0.087144f
C13244 SEL2.t105 VSS 0.039309f
C13245 SEL2.t60 VSS 0.139158f
C13246 SEL2.t96 VSS 0.04327f
C13247 SEL2.n26 VSS 0.123432f
C13248 SEL2.n27 VSS 0.036571f
C13249 SEL2.n28 VSS 0.05726f
C13250 SEL2.n29 VSS 0.52738f
C13251 SEL2.t139 VSS 0.039309f
C13252 SEL2.t17 VSS 0.139158f
C13253 SEL2.t128 VSS 0.04327f
C13254 SEL2.n30 VSS 0.123432f
C13255 SEL2.n31 VSS 0.036567f
C13256 SEL2.n32 VSS 0.055954f
C13257 SEL2.n33 VSS 0.56381f
C13258 SEL2.n34 VSS 0.893698f
C13259 SEL2.n35 VSS 0.905768f
C13260 SEL2.n36 VSS 0.079769f
C13261 SEL2.n37 VSS 0.086502f
C13262 SEL2.n38 VSS 0.079683f
C13263 SEL2.n39 VSS 0.094336f
C13264 SEL2.n40 VSS 2.25566f
C13265 SEL2.t43 VSS 0.025525f
C13266 SEL2.t6 VSS 0.035631f
C13267 SEL2.t46 VSS 0.035631f
C13268 SEL2.n41 VSS 0.1116f
C13269 SEL2.t21 VSS 0.039019f
C13270 SEL2.t104 VSS 0.039309f
C13271 SEL2.t74 VSS 0.139158f
C13272 SEL2.t56 VSS 0.04327f
C13273 SEL2.n42 VSS 0.123432f
C13274 SEL2.n43 VSS 0.036589f
C13275 SEL2.t82 VSS 0.039309f
C13276 SEL2.t55 VSS 0.139158f
C13277 SEL2.t70 VSS 0.04327f
C13278 SEL2.n44 VSS 0.123432f
C13279 SEL2.n45 VSS 0.036555f
C13280 SEL2.n46 VSS 0.087144f
C13281 SEL2.t61 VSS 0.039309f
C13282 SEL2.t31 VSS 0.139158f
C13283 SEL2.t51 VSS 0.04327f
C13284 SEL2.n47 VSS 0.123432f
C13285 SEL2.n48 VSS 0.036571f
C13286 SEL2.n49 VSS 0.05726f
C13287 SEL2.n50 VSS 0.52738f
C13288 SEL2.t88 VSS 0.039309f
C13289 SEL2.t126 VSS 0.139158f
C13290 SEL2.t80 VSS 0.04327f
C13291 SEL2.n51 VSS 0.123432f
C13292 SEL2.n52 VSS 0.036567f
C13293 SEL2.n53 VSS 0.055954f
C13294 SEL2.n54 VSS 0.56381f
C13295 SEL2.n55 VSS 0.893698f
C13296 SEL2.n56 VSS 0.905768f
C13297 SEL2.n57 VSS 0.079769f
C13298 SEL2.n58 VSS 0.086502f
C13299 SEL2.n59 VSS 0.07989f
C13300 SEL2.n60 VSS 0.096478f
C13301 SEL2.n61 VSS 1.77768f
C13302 SEL2.t15 VSS 0.025525f
C13303 SEL2.t106 VSS 0.035631f
C13304 SEL2.t57 VSS 0.035631f
C13305 SEL2.n62 VSS 0.1116f
C13306 SEL2.t132 VSS 0.039019f
C13307 SEL2.t1 VSS 0.039309f
C13308 SEL2.t10 VSS 0.139158f
C13309 SEL2.t97 VSS 0.04327f
C13310 SEL2.n63 VSS 0.123432f
C13311 SEL2.n64 VSS 0.036589f
C13312 SEL2.t125 VSS 0.039309f
C13313 SEL2.t140 VSS 0.139158f
C13314 SEL2.t114 VSS 0.04327f
C13315 SEL2.n65 VSS 0.123432f
C13316 SEL2.n66 VSS 0.036555f
C13317 SEL2.n67 VSS 0.087144f
C13318 SEL2.t103 VSS 0.039309f
C13319 SEL2.t98 VSS 0.139158f
C13320 SEL2.t92 VSS 0.04327f
C13321 SEL2.n68 VSS 0.123432f
C13322 SEL2.n69 VSS 0.036571f
C13323 SEL2.n70 VSS 0.05726f
C13324 SEL2.n71 VSS 0.52738f
C13325 SEL2.t136 VSS 0.039309f
C13326 SEL2.t38 VSS 0.139158f
C13327 SEL2.t124 VSS 0.04327f
C13328 SEL2.n72 VSS 0.123432f
C13329 SEL2.n73 VSS 0.036567f
C13330 SEL2.n74 VSS 0.055954f
C13331 SEL2.n75 VSS 0.56381f
C13332 SEL2.n76 VSS 0.893698f
C13333 SEL2.n77 VSS 0.905768f
C13334 SEL2.n78 VSS 0.079769f
C13335 SEL2.n79 VSS 0.086502f
C13336 SEL2.n80 VSS 0.08018f
C13337 SEL2.n81 VSS 0.099319f
C13338 SEL2.n82 VSS 1.77102f
C13339 SEL2.t81 VSS 0.025525f
C13340 SEL2.t72 VSS 0.035631f
C13341 SEL2.t141 VSS 0.035631f
C13342 SEL2.n83 VSS 0.1116f
C13343 SEL2.t19 VSS 0.039019f
C13344 SEL2.t0 VSS 0.039309f
C13345 SEL2.t117 VSS 0.139158f
C13346 SEL2.t95 VSS 0.04327f
C13347 SEL2.n84 VSS 0.123432f
C13348 SEL2.n85 VSS 0.036589f
C13349 SEL2.t120 VSS 0.039309f
C13350 SEL2.t93 VSS 0.139158f
C13351 SEL2.t112 VSS 0.04327f
C13352 SEL2.n86 VSS 0.123432f
C13353 SEL2.n87 VSS 0.036555f
C13354 SEL2.n88 VSS 0.087144f
C13355 SEL2.t102 VSS 0.039309f
C13356 SEL2.t52 VSS 0.139158f
C13357 SEL2.t90 VSS 0.04327f
C13358 SEL2.n89 VSS 0.123432f
C13359 SEL2.n90 VSS 0.036571f
C13360 SEL2.n91 VSS 0.05726f
C13361 SEL2.n92 VSS 0.52738f
C13362 SEL2.t135 VSS 0.039309f
C13363 SEL2.t14 VSS 0.139158f
C13364 SEL2.t119 VSS 0.04327f
C13365 SEL2.n93 VSS 0.123432f
C13366 SEL2.n94 VSS 0.036567f
C13367 SEL2.n95 VSS 0.055954f
C13368 SEL2.n96 VSS 0.56381f
C13369 SEL2.n97 VSS 0.893698f
C13370 SEL2.n98 VSS 0.905768f
C13371 SEL2.n99 VSS 0.079769f
C13372 SEL2.n100 VSS 0.086502f
C13373 SEL2.n101 VSS 0.079785f
C13374 SEL2.n102 VSS 0.095408f
C13375 SEL2.n103 VSS 1.76769f
C13376 SEL2.t79 VSS 0.025525f
C13377 SEL2.t71 VSS 0.035631f
C13378 SEL2.t143 VSS 0.035631f
C13379 SEL2.n104 VSS 0.1116f
C13380 SEL2.t84 VSS 0.039019f
C13381 SEL2.t63 VSS 0.039309f
C13382 SEL2.t40 VSS 0.139158f
C13383 SEL2.t30 VSS 0.04327f
C13384 SEL2.n105 VSS 0.123432f
C13385 SEL2.n106 VSS 0.036589f
C13386 SEL2.t11 VSS 0.039309f
C13387 SEL2.t29 VSS 0.139158f
C13388 SEL2.t5 VSS 0.04327f
C13389 SEL2.n107 VSS 0.123432f
C13390 SEL2.n108 VSS 0.036555f
C13391 SEL2.n109 VSS 0.087144f
C13392 SEL2.t35 VSS 0.039309f
C13393 SEL2.t2 VSS 0.139158f
C13394 SEL2.t27 VSS 0.04327f
C13395 SEL2.n110 VSS 0.123432f
C13396 SEL2.n111 VSS 0.036571f
C13397 SEL2.n112 VSS 0.05726f
C13398 SEL2.n113 VSS 0.52738f
C13399 SEL2.t45 VSS 0.039309f
C13400 SEL2.t78 VSS 0.139158f
C13401 SEL2.t42 VSS 0.04327f
C13402 SEL2.n114 VSS 0.123432f
C13403 SEL2.n115 VSS 0.036567f
C13404 SEL2.n116 VSS 0.055954f
C13405 SEL2.n117 VSS 0.56381f
C13406 SEL2.n118 VSS 0.893698f
C13407 SEL2.n119 VSS 0.905768f
C13408 SEL2.n120 VSS 0.079769f
C13409 SEL2.n121 VSS 0.086502f
C13410 SEL2.n122 VSS 0.079768f
C13411 SEL2.n123 VSS 0.095232f
C13412 SEL2.n124 VSS 1.79842f
C13413 SEL2.t64 VSS 0.025525f
C13414 SEL2.t24 VSS 0.035631f
C13415 SEL2.t67 VSS 0.035631f
C13416 SEL2.n125 VSS 0.1116f
C13417 SEL2.t32 VSS 0.039019f
C13418 SEL2.t122 VSS 0.039309f
C13419 SEL2.t47 VSS 0.139158f
C13420 SEL2.t127 VSS 0.04327f
C13421 SEL2.n126 VSS 0.123432f
C13422 SEL2.n127 VSS 0.036589f
C13423 SEL2.t12 VSS 0.039309f
C13424 SEL2.t89 VSS 0.139158f
C13425 SEL2.t25 VSS 0.04327f
C13426 SEL2.n128 VSS 0.123432f
C13427 SEL2.n129 VSS 0.036555f
C13428 SEL2.n130 VSS 0.087144f
C13429 SEL2.t121 VSS 0.039309f
C13430 SEL2.t109 VSS 0.139158f
C13431 SEL2.t142 VSS 0.04327f
C13432 SEL2.n131 VSS 0.123432f
C13433 SEL2.n132 VSS 0.036571f
C13434 SEL2.n133 VSS 0.05726f
C13435 SEL2.n134 VSS 0.52738f
C13436 SEL2.t68 VSS 0.039309f
C13437 SEL2.t134 VSS 0.139158f
C13438 SEL2.t87 VSS 0.04327f
C13439 SEL2.n135 VSS 0.123432f
C13440 SEL2.n136 VSS 0.036567f
C13441 SEL2.n137 VSS 0.055954f
C13442 SEL2.n138 VSS 0.56381f
C13443 SEL2.n139 VSS 0.893698f
C13444 SEL2.n140 VSS 0.905768f
C13445 SEL2.n141 VSS 0.079769f
C13446 SEL2.n142 VSS 0.086502f
C13447 SEL2.n143 VSS 0.08041f
C13448 SEL2.n144 VSS 0.101438f
C13449 SEL2.n145 VSS 1.77552f
C13450 SEL2.t54 VSS 0.025525f
C13451 SEL2.t22 VSS 0.035631f
C13452 SEL2.t62 VSS 0.035631f
C13453 SEL2.n146 VSS 0.1116f
C13454 SEL2.t28 VSS 0.039019f
C13455 SEL2.t8 VSS 0.039309f
C13456 SEL2.t41 VSS 0.139158f
C13457 SEL2.t13 VSS 0.04327f
C13458 SEL2.n147 VSS 0.123432f
C13459 SEL2.n148 VSS 0.036589f
C13460 SEL2.t37 VSS 0.039309f
C13461 SEL2.t73 VSS 0.139158f
C13462 SEL2.t44 VSS 0.04327f
C13463 SEL2.n149 VSS 0.123432f
C13464 SEL2.n150 VSS 0.036555f
C13465 SEL2.n151 VSS 0.087144f
C13466 SEL2.t7 VSS 0.039309f
C13467 SEL2.t94 VSS 0.139158f
C13468 SEL2.t23 VSS 0.04327f
C13469 SEL2.n152 VSS 0.123432f
C13470 SEL2.n153 VSS 0.036571f
C13471 SEL2.n154 VSS 0.05726f
C13472 SEL2.n155 VSS 0.52738f
C13473 SEL2.t108 VSS 0.039309f
C13474 SEL2.t115 VSS 0.139158f
C13475 SEL2.t131 VSS 0.04327f
C13476 SEL2.n156 VSS 0.123432f
C13477 SEL2.n157 VSS 0.036567f
C13478 SEL2.n158 VSS 0.055954f
C13479 SEL2.n159 VSS 0.56381f
C13480 SEL2.n160 VSS 0.893698f
C13481 SEL2.n161 VSS 0.905768f
C13482 SEL2.n162 VSS 0.079769f
C13483 SEL2.n163 VSS 0.086502f
C13484 SEL2.n164 VSS 0.080069f
C13485 SEL2.n165 VSS 0.098255f
C13486 SEL2.n166 VSS 2.22874f
C13487 SEL2.n167 VSS 0.536679f
C13488 SEL2.n168 VSS 0.080371f
C13489 SEL2.t66 VSS 0.039309f
C13490 SEL2.t118 VSS 0.139158f
C13491 SEL2.t138 VSS 0.04327f
C13492 SEL2.n169 VSS 0.123432f
C13493 SEL2.n170 VSS 0.036589f
C13494 SEL2.t69 VSS 0.039309f
C13495 SEL2.t86 VSS 0.139158f
C13496 SEL2.t49 VSS 0.04327f
C13497 SEL2.n171 VSS 0.123432f
C13498 SEL2.n172 VSS 0.036555f
C13499 SEL2.n173 VSS 0.087144f
C13500 SEL2.t100 VSS 0.039309f
C13501 SEL2.t133 VSS 0.139158f
C13502 SEL2.t76 VSS 0.04327f
C13503 SEL2.n174 VSS 0.123432f
C13504 SEL2.n175 VSS 0.036571f
C13505 SEL2.n176 VSS 0.05726f
C13506 SEL2.n177 VSS 0.52738f
C13507 SEL2.t137 VSS 0.039309f
C13508 SEL2.t34 VSS 0.139158f
C13509 SEL2.t113 VSS 0.04327f
C13510 SEL2.n178 VSS 0.123432f
C13511 SEL2.n179 VSS 0.036567f
C13512 SEL2.n180 VSS 0.055954f
C13513 SEL2.n181 VSS 0.56381f
C13514 SEL2.n182 VSS 0.893698f
C13515 SEL2.t20 VSS 0.025525f
C13516 SEL2.t50 VSS 0.035631f
C13517 SEL2.t111 VSS 0.035631f
C13518 SEL2.n183 VSS 0.1116f
C13519 SEL2.n184 VSS 0.086502f
C13520 SEL2.t4 VSS 0.039019f
C13521 SEL2.n185 VSS 0.079769f
C13522 SEL2.n186 VSS 0.905768f
C13523 MULT_0.4bit_ADDER_1.B2.t20 VSS 0.05786f
C13524 MULT_0.4bit_ADDER_1.B2.t12 VSS 0.018842f
C13525 MULT_0.4bit_ADDER_1.B2.t13 VSS 0.02602f
C13526 MULT_0.4bit_ADDER_1.B2.n0 VSS 0.028059f
C13527 MULT_0.4bit_ADDER_1.B2.t16 VSS 0.019371f
C13528 MULT_0.4bit_ADDER_1.B2.n1 VSS 0.049151f
C13529 MULT_0.4bit_ADDER_1.B2.n2 VSS 0.086219f
C13530 MULT_0.4bit_ADDER_1.B2.t15 VSS 0.026418f
C13531 MULT_0.4bit_ADDER_1.B2.t19 VSS 0.053153f
C13532 MULT_0.4bit_ADDER_1.B2.t14 VSS 0.052492f
C13533 MULT_0.4bit_ADDER_1.B2.t23 VSS 0.052492f
C13534 MULT_0.4bit_ADDER_1.B2.t22 VSS 0.052492f
C13535 MULT_0.4bit_ADDER_1.B2.t21 VSS 0.010908f
C13536 MULT_0.4bit_ADDER_1.B2.t17 VSS 0.010908f
C13537 MULT_0.4bit_ADDER_1.B2.t18 VSS 0.010908f
C13538 MULT_0.4bit_ADDER_1.B2.n3 VSS 0.323398f
C13539 MULT_0.4bit_ADDER_1.B2.n4 VSS 0.238197f
C13540 MULT_0.4bit_ADDER_1.B2.n5 VSS 0.129816f
C13541 MULT_0.4bit_ADDER_1.B2.n6 VSS 0.127533f
C13542 MULT_0.4bit_ADDER_1.B2.n7 VSS 0.078447f
C13543 MULT_0.4bit_ADDER_1.B2.n8 VSS 0.102909f
C13544 MULT_0.4bit_ADDER_1.B2.n9 VSS 1.13401f
C13545 MULT_0.4bit_ADDER_1.B2.t8 VSS 0.009454f
C13546 MULT_0.4bit_ADDER_1.B2.t0 VSS 0.009454f
C13547 MULT_0.4bit_ADDER_1.B2.n10 VSS 0.022865f
C13548 MULT_0.4bit_ADDER_1.B2.t3 VSS 0.009454f
C13549 MULT_0.4bit_ADDER_1.B2.t6 VSS 0.009454f
C13550 MULT_0.4bit_ADDER_1.B2.n11 VSS 0.022863f
C13551 MULT_0.4bit_ADDER_1.B2.n12 VSS 0.163946f
C13552 MULT_0.4bit_ADDER_1.B2.t1 VSS 0.009454f
C13553 MULT_0.4bit_ADDER_1.B2.t2 VSS 0.009454f
C13554 MULT_0.4bit_ADDER_1.B2.n13 VSS 0.018908f
C13555 MULT_0.4bit_ADDER_1.B2.n14 VSS 0.014853f
C13556 MULT_0.4bit_ADDER_1.B2.t11 VSS 0.039997f
C13557 MULT_0.4bit_ADDER_1.B2.t4 VSS 0.039997f
C13558 MULT_0.4bit_ADDER_1.B2.n15 VSS 0.079994f
C13559 MULT_0.4bit_ADDER_1.B2.n16 VSS 0.031807f
C13560 MULT_0.4bit_ADDER_1.B2.t9 VSS 0.039997f
C13561 MULT_0.4bit_ADDER_1.B2.t10 VSS 0.039997f
C13562 MULT_0.4bit_ADDER_1.B2.n17 VSS 0.079994f
C13563 MULT_0.4bit_ADDER_1.B2.n18 VSS 0.035183f
C13564 MULT_0.4bit_ADDER_1.B2.n19 VSS 0.362228f
C13565 MULT_0.4bit_ADDER_1.B2.t5 VSS 0.039997f
C13566 MULT_0.4bit_ADDER_1.B2.t7 VSS 0.039997f
C13567 MULT_0.4bit_ADDER_1.B2.n20 VSS 0.079994f
C13568 MULT_0.4bit_ADDER_1.B2.n21 VSS 0.035236f
C13569 MULT_0.4bit_ADDER_1.B2.n22 VSS 0.232317f
C13570 MULT_0.4bit_ADDER_1.B2.n23 VSS 0.052355f
C13571 MULT_0.4bit_ADDER_1.B2.n24 VSS 0.229798f
C13572 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t10 VSS 0.007073f
C13573 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t8 VSS 0.007073f
C13574 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n0 VSS 0.017105f
C13575 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t3 VSS 0.007073f
C13576 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t2 VSS 0.007073f
C13577 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n1 VSS 0.017107f
C13578 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n2 VSS 0.122656f
C13579 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t0 VSS 0.007073f
C13580 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t1 VSS 0.007073f
C13581 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n3 VSS 0.014146f
C13582 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n4 VSS 0.011112f
C13583 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t7 VSS 0.029924f
C13584 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t6 VSS 0.029924f
C13585 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n5 VSS 0.059848f
C13586 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n6 VSS 0.023796f
C13587 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t11 VSS 0.029924f
C13588 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t9 VSS 0.029924f
C13589 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n7 VSS 0.059848f
C13590 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n8 VSS 0.026362f
C13591 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n9 VSS 0.271f
C13592 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t4 VSS 0.029924f
C13593 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t5 VSS 0.029924f
C13594 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n10 VSS 0.059848f
C13595 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n11 VSS 0.026322f
C13596 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n12 VSS 0.173808f
C13597 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n13 VSS 0.03917f
C13598 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n14 VSS 0.172104f
C13599 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t15 VSS 0.043288f
C13600 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t20 VSS 0.014096f
C13601 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t17 VSS 0.019467f
C13602 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n15 VSS 0.020992f
C13603 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t19 VSS 0.014492f
C13604 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n16 VSS 0.036772f
C13605 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n17 VSS 0.064505f
C13606 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t16 VSS 0.019764f
C13607 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t22 VSS 0.039767f
C13608 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t14 VSS 0.039272f
C13609 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t18 VSS 0.039272f
C13610 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t12 VSS 0.039272f
C13611 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t21 VSS 0.008161f
C13612 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t13 VSS 0.008161f
C13613 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.t23 VSS 0.008161f
C13614 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n18 VSS 0.24195f
C13615 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n19 VSS 0.178207f
C13616 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n20 VSS 0.097121f
C13617 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n21 VSS 0.095413f
C13618 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n22 VSS 0.05869f
C13619 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n23 VSS 0.076991f
C13620 8bit_ADDER_0.FULL_ADDER_XORED_0.XOR2_2.Y.n24 VSS 1.26966f
C13621 a_n23950_3810.n0 VSS 2.96691f
C13622 a_n23950_3810.t11 VSS 0.093341f
C13623 a_n23950_3810.t2 VSS 0.093341f
C13624 a_n23950_3810.t1 VSS 0.093341f
C13625 a_n23950_3810.n1 VSS 0.20269f
C13626 a_n23950_3810.t8 VSS 0.093341f
C13627 a_n23950_3810.t7 VSS 0.093341f
C13628 a_n23950_3810.n2 VSS 0.202296f
C13629 a_n23950_3810.t4 VSS 0.093341f
C13630 a_n23950_3810.t6 VSS 0.093341f
C13631 a_n23950_3810.n3 VSS 0.202001f
C13632 a_n23950_3810.t5 VSS 0.093341f
C13633 a_n23950_3810.t3 VSS 0.093341f
C13634 a_n23950_3810.n4 VSS 0.202001f
C13635 a_n23950_3810.t10 VSS 0.093341f
C13636 a_n23950_3810.t9 VSS 0.093341f
C13637 a_n23950_3810.n5 VSS 0.202001f
C13638 a_n23950_3810.n6 VSS 0.202001f
C13639 a_n23950_3810.t0 VSS 0.093341f
C13640 a_n18998_n11063.n0 VSS 1.48365f
C13641 a_n18998_n11063.n1 VSS 1.48326f
C13642 a_n18998_n11063.t6 VSS 0.093341f
C13643 a_n18998_n11063.t1 VSS 0.093341f
C13644 a_n18998_n11063.t2 VSS 0.093341f
C13645 a_n18998_n11063.n2 VSS 0.202296f
C13646 a_n18998_n11063.t0 VSS 0.093341f
C13647 a_n18998_n11063.t11 VSS 0.093341f
C13648 a_n18998_n11063.n3 VSS 0.202001f
C13649 a_n18998_n11063.t10 VSS 0.093341f
C13650 a_n18998_n11063.t9 VSS 0.093341f
C13651 a_n18998_n11063.n4 VSS 0.202001f
C13652 a_n18998_n11063.t4 VSS 0.093341f
C13653 a_n18998_n11063.t3 VSS 0.093341f
C13654 a_n18998_n11063.n5 VSS 0.202001f
C13655 a_n18998_n11063.t8 VSS 0.093341f
C13656 a_n18998_n11063.t5 VSS 0.093341f
C13657 a_n18998_n11063.n6 VSS 0.202001f
C13658 a_n18998_n11063.n7 VSS 0.20269f
C13659 a_n18998_n11063.t7 VSS 0.093341f
C13660 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t17 VSS 0.013766f
C13661 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t20 VSS 0.027698f
C13662 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t13 VSS 0.027354f
C13663 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t12 VSS 0.027354f
C13664 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t14 VSS 0.027354f
C13665 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t21 VSS 0.005684f
C13666 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t23 VSS 0.005684f
C13667 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t22 VSS 0.005684f
C13668 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n0 VSS 0.168523f
C13669 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n1 VSS 0.124125f
C13670 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n2 VSS 0.067647f
C13671 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n3 VSS 0.066457f
C13672 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n4 VSS 0.040879f
C13673 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n5 VSS 0.05311f
C13674 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t16 VSS 0.030151f
C13675 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t18 VSS 0.009818f
C13676 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t19 VSS 0.013559f
C13677 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n6 VSS 0.014622f
C13678 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t15 VSS 0.010094f
C13679 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n7 VSS 0.025612f
C13680 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n8 VSS 0.044927f
C13681 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t11 VSS 0.004926f
C13682 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t10 VSS 0.004926f
C13683 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n9 VSS 0.011915f
C13684 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t7 VSS 0.004926f
C13685 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t5 VSS 0.004926f
C13686 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n10 VSS 0.011914f
C13687 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n11 VSS 0.085433f
C13688 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t9 VSS 0.004926f
C13689 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t8 VSS 0.004926f
C13690 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n12 VSS 0.009853f
C13691 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n13 VSS 0.00774f
C13692 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t0 VSS 0.020843f
C13693 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t4 VSS 0.020843f
C13694 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n14 VSS 0.041685f
C13695 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n15 VSS 0.016575f
C13696 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t2 VSS 0.020843f
C13697 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t1 VSS 0.020843f
C13698 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n16 VSS 0.041685f
C13699 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n17 VSS 0.018334f
C13700 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n18 VSS 0.188757f
C13701 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t3 VSS 0.020843f
C13702 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.t6 VSS 0.020843f
C13703 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n19 VSS 0.041685f
C13704 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n20 VSS 0.018362f
C13705 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n21 VSS 0.12106f
C13706 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n22 VSS 0.027282f
C13707 MULT_0.4bit_ADDER_2.FULL_ADDER_0.XOR2_1.A.n23 VSS 0.119748f
C13708 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n0 VSS 0.967969f
C13709 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t5 VSS 0.008375f
C13710 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t4 VSS 0.008375f
C13711 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n1 VSS 0.018687f
C13712 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t1 VSS 0.008375f
C13713 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t6 VSS 0.008375f
C13714 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n2 VSS 0.018636f
C13715 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t3 VSS 0.008375f
C13716 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t2 VSS 0.008375f
C13717 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n3 VSS 0.018636f
C13718 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t0 VSS 0.05057f
C13719 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t8 VSS 0.028606f
C13720 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t16 VSS 0.02825f
C13721 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t18 VSS 0.02825f
C13722 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t12 VSS 0.02825f
C13723 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n4 VSS 0.112442f
C13724 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t13 VSS 0.005871f
C13725 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t7 VSS 0.005871f
C13726 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t15 VSS 0.005871f
C13727 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t10 VSS 0.005871f
C13728 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n5 VSS 0.106225f
C13729 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n6 VSS 0.166131f
C13730 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t9 VSS 0.026417f
C13731 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t14 VSS 0.01014f
C13732 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t11 VSS 0.014003f
C13733 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n7 VSS 0.016118f
C13734 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.t17 VSS 0.010659f
C13735 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n8 VSS 0.016345f
C13736 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n9 VSS 0.055518f
C13737 MULT_0.4bit_ADDER_1.FULL_ADDER_2.COUT.n10 VSS 0.369194f
C13738 XOR8_0.S0.t13 VSS 0.118279f
C13739 XOR8_0.S0.t14 VSS 0.348483f
C13740 XOR8_0.S0.t12 VSS 0.115077f
C13741 XOR8_0.S0.n0 VSS 0.593267f
C13742 XOR8_0.S0.t0 VSS 0.034444f
C13743 XOR8_0.S0.t1 VSS 0.034444f
C13744 XOR8_0.S0.n1 VSS 0.083306f
C13745 XOR8_0.S0.t11 VSS 0.034444f
C13746 XOR8_0.S0.t9 VSS 0.034444f
C13747 XOR8_0.S0.n2 VSS 0.083297f
C13748 XOR8_0.S0.n3 VSS 0.597311f
C13749 XOR8_0.S0.t2 VSS 0.034444f
C13750 XOR8_0.S0.t10 VSS 0.034444f
C13751 XOR8_0.S0.n4 VSS 0.068887f
C13752 XOR8_0.S0.n5 VSS 0.054113f
C13753 XOR8_0.S0.t3 VSS 0.145723f
C13754 XOR8_0.S0.t8 VSS 0.145723f
C13755 XOR8_0.S0.n6 VSS 0.291446f
C13756 XOR8_0.S0.n7 VSS 0.11561f
C13757 XOR8_0.S0.t4 VSS 0.145723f
C13758 XOR8_0.S0.t5 VSS 0.145723f
C13759 XOR8_0.S0.n8 VSS 0.291446f
C13760 XOR8_0.S0.n9 VSS 0.128183f
C13761 XOR8_0.S0.n10 VSS 1.31971f
C13762 XOR8_0.S0.t7 VSS 0.145723f
C13763 XOR8_0.S0.t6 VSS 0.145723f
C13764 XOR8_0.S0.n11 VSS 0.291446f
C13765 XOR8_0.S0.n12 VSS 0.128377f
C13766 XOR8_0.S0.n13 VSS 0.846407f
C13767 XOR8_0.S0.n14 VSS 0.190514f
C13768 XOR8_0.S0.n15 VSS 0.837736f
C13769 a_n13975_n7799.n0 VSS 1.48365f
C13770 a_n13975_n7799.n1 VSS 1.48326f
C13771 a_n13975_n7799.t3 VSS 0.093341f
C13772 a_n13975_n7799.t1 VSS 0.093341f
C13773 a_n13975_n7799.t0 VSS 0.093341f
C13774 a_n13975_n7799.n2 VSS 0.202296f
C13775 a_n13975_n7799.t2 VSS 0.093341f
C13776 a_n13975_n7799.t9 VSS 0.093341f
C13777 a_n13975_n7799.n3 VSS 0.202001f
C13778 a_n13975_n7799.t10 VSS 0.093341f
C13779 a_n13975_n7799.t11 VSS 0.093341f
C13780 a_n13975_n7799.n4 VSS 0.202001f
C13781 a_n13975_n7799.t8 VSS 0.093341f
C13782 a_n13975_n7799.t7 VSS 0.093341f
C13783 a_n13975_n7799.n5 VSS 0.20269f
C13784 a_n13975_n7799.t4 VSS 0.093341f
C13785 a_n13975_n7799.t6 VSS 0.093341f
C13786 a_n13975_n7799.n6 VSS 0.202001f
C13787 a_n13975_n7799.n7 VSS 0.202001f
C13788 a_n13975_n7799.t5 VSS 0.093341f
C13789 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t16 VSS 0.013766f
C13790 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t22 VSS 0.027698f
C13791 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t13 VSS 0.027354f
C13792 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t12 VSS 0.027354f
C13793 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t21 VSS 0.027354f
C13794 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t20 VSS 0.005684f
C13795 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t14 VSS 0.005684f
C13796 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t17 VSS 0.005684f
C13797 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n0 VSS 0.168523f
C13798 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n1 VSS 0.124125f
C13799 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n2 VSS 0.067647f
C13800 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n3 VSS 0.066457f
C13801 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n4 VSS 0.040879f
C13802 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n5 VSS 0.05311f
C13803 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t15 VSS 0.030151f
C13804 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t19 VSS 0.009818f
C13805 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t18 VSS 0.013559f
C13806 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n6 VSS 0.014622f
C13807 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t23 VSS 0.010094f
C13808 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n7 VSS 0.025612f
C13809 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n8 VSS 0.044927f
C13810 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t7 VSS 0.004926f
C13811 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t8 VSS 0.004926f
C13812 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n9 VSS 0.011915f
C13813 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t1 VSS 0.004926f
C13814 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t2 VSS 0.004926f
C13815 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n10 VSS 0.011914f
C13816 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n11 VSS 0.085433f
C13817 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t6 VSS 0.004926f
C13818 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t0 VSS 0.004926f
C13819 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n12 VSS 0.009853f
C13820 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n13 VSS 0.00774f
C13821 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t11 VSS 0.020843f
C13822 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t3 VSS 0.020843f
C13823 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n14 VSS 0.041685f
C13824 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n15 VSS 0.016575f
C13825 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t9 VSS 0.020843f
C13826 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t10 VSS 0.020843f
C13827 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n16 VSS 0.041685f
C13828 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n17 VSS 0.018334f
C13829 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n18 VSS 0.188757f
C13830 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t5 VSS 0.020843f
C13831 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.t4 VSS 0.020843f
C13832 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n19 VSS 0.041685f
C13833 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n20 VSS 0.018362f
C13834 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n21 VSS 0.12106f
C13835 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n22 VSS 0.027282f
C13836 MULT_0.4bit_ADDER_1.FULL_ADDER_2.XOR2_1.A.n23 VSS 0.119748f
C13837 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t13 VSS 0.013766f
C13838 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t15 VSS 0.027698f
C13839 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t23 VSS 0.027354f
C13840 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t14 VSS 0.027354f
C13841 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t17 VSS 0.027354f
C13842 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t12 VSS 0.005684f
C13843 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t18 VSS 0.005684f
C13844 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t16 VSS 0.005684f
C13845 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n0 VSS 0.168523f
C13846 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n1 VSS 0.124125f
C13847 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n2 VSS 0.067647f
C13848 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n3 VSS 0.066457f
C13849 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n4 VSS 0.040879f
C13850 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n5 VSS 0.05311f
C13851 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t19 VSS 0.030151f
C13852 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t22 VSS 0.009818f
C13853 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t20 VSS 0.013559f
C13854 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n6 VSS 0.014622f
C13855 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t21 VSS 0.010094f
C13856 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n7 VSS 0.025612f
C13857 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n8 VSS 0.044927f
C13858 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t11 VSS 0.004926f
C13859 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t10 VSS 0.004926f
C13860 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n9 VSS 0.011915f
C13861 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t5 VSS 0.004926f
C13862 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t0 VSS 0.004926f
C13863 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n10 VSS 0.011914f
C13864 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n11 VSS 0.085433f
C13865 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t9 VSS 0.004926f
C13866 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t1 VSS 0.004926f
C13867 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n12 VSS 0.009853f
C13868 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n13 VSS 0.00774f
C13869 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t8 VSS 0.020843f
C13870 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t2 VSS 0.020843f
C13871 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n14 VSS 0.041685f
C13872 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n15 VSS 0.016575f
C13873 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t7 VSS 0.020843f
C13874 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t6 VSS 0.020843f
C13875 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n16 VSS 0.041685f
C13876 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n17 VSS 0.018334f
C13877 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n18 VSS 0.188757f
C13878 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t3 VSS 0.020843f
C13879 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.t4 VSS 0.020843f
C13880 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n19 VSS 0.041685f
C13881 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n20 VSS 0.018362f
C13882 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n21 VSS 0.12106f
C13883 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n22 VSS 0.027282f
C13884 8bit_ADDER_0.FULL_ADDER_XORED_2.XOR2_1.A.n23 VSS 0.119748f
C13885 a_n18042_2026.n0 VSS 2.96691f
C13886 a_n18042_2026.t1 VSS 0.093341f
C13887 a_n18042_2026.t9 VSS 0.093341f
C13888 a_n18042_2026.t10 VSS 0.093341f
C13889 a_n18042_2026.n1 VSS 0.20269f
C13890 a_n18042_2026.t5 VSS 0.093341f
C13891 a_n18042_2026.t11 VSS 0.093341f
C13892 a_n18042_2026.n2 VSS 0.202001f
C13893 a_n18042_2026.t3 VSS 0.093341f
C13894 a_n18042_2026.t4 VSS 0.093341f
C13895 a_n18042_2026.n3 VSS 0.202001f
C13896 a_n18042_2026.t6 VSS 0.093341f
C13897 a_n18042_2026.t8 VSS 0.093341f
C13898 a_n18042_2026.n4 VSS 0.202001f
C13899 a_n18042_2026.t2 VSS 0.093341f
C13900 a_n18042_2026.t7 VSS 0.093341f
C13901 a_n18042_2026.n5 VSS 0.202001f
C13902 a_n18042_2026.n6 VSS 0.202296f
C13903 a_n18042_2026.t0 VSS 0.093341f
C13904 mux8_3.NAND4F_8.Y.n0 VSS 0.539804f
C13905 mux8_3.NAND4F_8.Y.t14 VSS 0.026899f
C13906 mux8_3.NAND4F_8.Y.t9 VSS 0.028853f
C13907 mux8_3.NAND4F_8.Y.n1 VSS 0.042994f
C13908 mux8_3.NAND4F_8.Y.t10 VSS 0.026899f
C13909 mux8_3.NAND4F_8.Y.t12 VSS 0.026899f
C13910 mux8_3.NAND4F_8.Y.t11 VSS 0.026899f
C13911 mux8_3.NAND4F_8.Y.t13 VSS 0.033983f
C13912 mux8_3.NAND4F_8.Y.n2 VSS 0.072608f
C13913 mux8_3.NAND4F_8.Y.n3 VSS 0.045714f
C13914 mux8_3.NAND4F_8.Y.n4 VSS 0.037354f
C13915 mux8_3.NAND4F_8.Y.n5 VSS 0.018278f
C13916 mux8_3.NAND4F_8.Y.t3 VSS 0.026614f
C13917 mux8_3.NAND4F_8.Y.t2 VSS 0.026614f
C13918 mux8_3.NAND4F_8.Y.n6 VSS 0.0618f
C13919 mux8_3.NAND4F_8.Y.t0 VSS 0.026614f
C13920 mux8_3.NAND4F_8.Y.t1 VSS 0.026614f
C13921 mux8_3.NAND4F_8.Y.n7 VSS 0.061615f
C13922 mux8_3.NAND4F_8.Y.t7 VSS 0.026614f
C13923 mux8_3.NAND4F_8.Y.t8 VSS 0.026614f
C13924 mux8_3.NAND4F_8.Y.n8 VSS 0.061615f
C13925 mux8_3.NAND4F_8.Y.t6 VSS 0.026614f
C13926 mux8_3.NAND4F_8.Y.t4 VSS 0.026614f
C13927 mux8_3.NAND4F_8.Y.n9 VSS 0.061615f
C13928 mux8_3.NAND4F_8.Y.n10 VSS 0.268281f
C13929 mux8_3.NAND4F_8.Y.t5 VSS 0.21369f
C13930 MULT_0.NAND2_9.Y.n0 VSS 1.19272f
C13931 MULT_0.NAND2_9.Y.n1 VSS 0.186498f
C13932 MULT_0.NAND2_9.Y.t6 VSS 0.022972f
C13933 MULT_0.NAND2_9.Y.t5 VSS 0.022972f
C13934 MULT_0.NAND2_9.Y.n2 VSS 0.051256f
C13935 MULT_0.NAND2_9.Y.t1 VSS 0.022972f
C13936 MULT_0.NAND2_9.Y.t4 VSS 0.022972f
C13937 MULT_0.NAND2_9.Y.n3 VSS 0.051117f
C13938 MULT_0.NAND2_9.Y.t3 VSS 0.022972f
C13939 MULT_0.NAND2_9.Y.t2 VSS 0.022972f
C13940 MULT_0.NAND2_9.Y.n4 VSS 0.051117f
C13941 MULT_0.NAND2_9.Y.t0 VSS 0.13839f
C13942 MULT_0.NAND2_9.Y.t9 VSS 0.029277f
C13943 MULT_0.NAND2_9.Y.t8 VSS 0.040868f
C13944 MULT_0.NAND2_9.Y.t10 VSS 0.040868f
C13945 MULT_0.NAND2_9.Y.n5 VSS 0.133396f
C13946 MULT_0.NAND2_9.Y.t7 VSS 0.046661f
C13947 A1.t13 VSS 0.096296f
C13948 A1.t16 VSS 0.036963f
C13949 A1.t18 VSS 0.051044f
C13950 A1.n0 VSS 0.058752f
C13951 A1.t15 VSS 0.038853f
C13952 A1.n1 VSS 0.059583f
C13953 A1.n2 VSS 0.246626f
C13954 A1.t31 VSS 0.104274f
C13955 A1.t34 VSS 0.102977f
C13956 A1.t39 VSS 0.102977f
C13957 A1.t10 VSS 0.102977f
C13958 A1.n3 VSS 0.409876f
C13959 A1.t22 VSS 0.021399f
C13960 A1.t37 VSS 0.021399f
C13961 A1.t12 VSS 0.021399f
C13962 A1.t17 VSS 0.021399f
C13963 A1.n4 VSS 0.387214f
C13964 A1.n5 VSS 0.60568f
C13965 A1.n6 VSS 1.20405f
C13966 A1.n7 VSS 1.54336f
C13967 A1.t2 VSS 0.096296f
C13968 A1.t21 VSS 0.036963f
C13969 A1.t20 VSS 0.051044f
C13970 A1.n8 VSS 0.058752f
C13971 A1.t36 VSS 0.038853f
C13972 A1.n9 VSS 0.059583f
C13973 A1.n10 VSS 0.247241f
C13974 A1.t9 VSS 0.096296f
C13975 A1.t42 VSS 0.036963f
C13976 A1.t28 VSS 0.051044f
C13977 A1.n11 VSS 0.058752f
C13978 A1.t41 VSS 0.038853f
C13979 A1.n12 VSS 0.059583f
C13980 A1.n13 VSS 0.247241f
C13981 A1.t32 VSS 0.096296f
C13982 A1.t29 VSS 0.036963f
C13983 A1.t0 VSS 0.051044f
C13984 A1.n14 VSS 0.058752f
C13985 A1.t45 VSS 0.038853f
C13986 A1.n15 VSS 0.059583f
C13987 A1.n16 VSS 0.247241f
C13988 A1.t6 VSS 0.096296f
C13989 A1.t4 VSS 0.036963f
C13990 A1.t33 VSS 0.051044f
C13991 A1.n17 VSS 0.058752f
C13992 A1.t3 VSS 0.038853f
C13993 A1.n18 VSS 0.059583f
C13994 A1.n19 VSS 0.247241f
C13995 A1.n20 VSS 7.384779f
C13996 A1.n21 VSS 3.47789f
C13997 A1.n22 VSS 1.25034f
C13998 A1.n23 VSS 22.2531f
C13999 A1.t27 VSS 0.096293f
C14000 A1.t44 VSS 0.048668f
C14001 A1.t1 VSS 0.038908f
C14002 A1.n24 VSS 0.061786f
C14003 A1.t19 VSS 0.038853f
C14004 A1.n25 VSS 0.056981f
C14005 A1.n26 VSS 0.247363f
C14006 A1.n27 VSS 0.422839f
C14007 A1.n28 VSS 2.72407f
C14008 A1.t24 VSS 0.038525f
C14009 A1.t25 VSS 0.04643f
C14010 A1.t11 VSS 0.04643f
C14011 A1.t8 VSS 0.04643f
C14012 A1.t40 VSS 0.04643f
C14013 A1.t35 VSS 0.058657f
C14014 A1.n29 VSS 0.125326f
C14015 A1.n30 VSS 0.078906f
C14016 A1.n31 VSS 0.078906f
C14017 A1.n32 VSS 0.068006f
C14018 A1.n33 VSS 0.055581f
C14019 A1.n34 VSS 7.60877f
C14020 A1.t26 VSS 0.021399f
C14021 A1.t30 VSS 0.021399f
C14022 A1.t43 VSS 0.021399f
C14023 A1.t14 VSS 0.021399f
C14024 A1.n35 VSS 0.388571f
C14025 A1.t23 VSS 0.102977f
C14026 A1.t38 VSS 0.102977f
C14027 A1.t5 VSS 0.104274f
C14028 A1.t7 VSS 0.102977f
C14029 A1.n36 VSS 0.408518f
C14030 A1.n37 VSS 0.606139f
C14031 A1.n38 VSS 1.21854f
C14032 a_n13192_2026.n0 VSS 1.48326f
C14033 a_n13192_2026.n1 VSS 1.48365f
C14034 a_n13192_2026.t7 VSS 0.093341f
C14035 a_n13192_2026.t0 VSS 0.093341f
C14036 a_n13192_2026.t2 VSS 0.093341f
C14037 a_n13192_2026.n2 VSS 0.20269f
C14038 a_n13192_2026.t11 VSS 0.093341f
C14039 a_n13192_2026.t1 VSS 0.093341f
C14040 a_n13192_2026.n3 VSS 0.202001f
C14041 a_n13192_2026.t6 VSS 0.093341f
C14042 a_n13192_2026.t10 VSS 0.093341f
C14043 a_n13192_2026.n4 VSS 0.202001f
C14044 a_n13192_2026.t5 VSS 0.093341f
C14045 a_n13192_2026.t4 VSS 0.093341f
C14046 a_n13192_2026.n5 VSS 0.202001f
C14047 a_n13192_2026.t8 VSS 0.093341f
C14048 a_n13192_2026.t3 VSS 0.093341f
C14049 a_n13192_2026.n6 VSS 0.202001f
C14050 a_n13192_2026.n7 VSS 0.202296f
C14051 a_n13192_2026.t9 VSS 0.093341f
C14052 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n0 VSS 0.860417f
C14053 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t0 VSS 0.007445f
C14054 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t2 VSS 0.007445f
C14055 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n1 VSS 0.016611f
C14056 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t3 VSS 0.007445f
C14057 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t1 VSS 0.007445f
C14058 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n2 VSS 0.016566f
C14059 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t6 VSS 0.007445f
C14060 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t5 VSS 0.007445f
C14061 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n3 VSS 0.016566f
C14062 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t4 VSS 0.044951f
C14063 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t15 VSS 0.025427f
C14064 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t17 VSS 0.025111f
C14065 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t13 VSS 0.025111f
C14066 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t7 VSS 0.025111f
C14067 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n4 VSS 0.099949f
C14068 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t18 VSS 0.005218f
C14069 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t16 VSS 0.005218f
C14070 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t9 VSS 0.005218f
C14071 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t14 VSS 0.005218f
C14072 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n5 VSS 0.094423f
C14073 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n6 VSS 0.147672f
C14074 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t8 VSS 0.023482f
C14075 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t12 VSS 0.009013f
C14076 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t10 VSS 0.012447f
C14077 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n7 VSS 0.014327f
C14078 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.t11 VSS 0.009474f
C14079 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n8 VSS 0.014529f
C14080 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n9 VSS 0.049349f
C14081 8bit_ADDER_0.FULL_ADDER_XORED_4.COUT.n10 VSS 0.328172f
C14082 mux8_5.NAND4F_6.Y.n0 VSS 0.599344f
C14083 mux8_5.NAND4F_6.Y.t0 VSS 0.244548f
C14084 mux8_5.NAND4F_6.Y.t9 VSS 0.038543f
C14085 mux8_5.NAND4F_6.Y.t10 VSS 0.118929f
C14086 mux8_5.NAND4F_6.Y.t11 VSS 0.044398f
C14087 mux8_5.NAND4F_6.Y.n1 VSS 0.149236f
C14088 mux8_5.NAND4F_6.Y.n2 VSS 0.032396f
C14089 mux8_5.NAND4F_6.Y.n3 VSS 1.72835f
C14090 mux8_5.NAND4F_6.Y.t7 VSS 0.029549f
C14091 mux8_5.NAND4F_6.Y.t8 VSS 0.029549f
C14092 mux8_5.NAND4F_6.Y.n4 VSS 0.068617f
C14093 mux8_5.NAND4F_6.Y.t4 VSS 0.029549f
C14094 mux8_5.NAND4F_6.Y.t3 VSS 0.029549f
C14095 mux8_5.NAND4F_6.Y.n5 VSS 0.068411f
C14096 mux8_5.NAND4F_6.Y.t6 VSS 0.029549f
C14097 mux8_5.NAND4F_6.Y.t5 VSS 0.029549f
C14098 mux8_5.NAND4F_6.Y.n6 VSS 0.068411f
C14099 mux8_5.NAND4F_6.Y.t1 VSS 0.029549f
C14100 mux8_5.NAND4F_6.Y.t2 VSS 0.029549f
C14101 mux8_5.NAND4F_6.Y.n7 VSS 0.068411f
C14102 mux8_5.NAND4F_6.Y.n8 VSS 0.281208f
C14103 mux8_7.NAND4F_8.Y.n0 VSS 0.539804f
C14104 mux8_7.NAND4F_8.Y.t9 VSS 0.026899f
C14105 mux8_7.NAND4F_8.Y.t10 VSS 0.028853f
C14106 mux8_7.NAND4F_8.Y.n1 VSS 0.042994f
C14107 mux8_7.NAND4F_8.Y.t11 VSS 0.026899f
C14108 mux8_7.NAND4F_8.Y.t13 VSS 0.026899f
C14109 mux8_7.NAND4F_8.Y.t12 VSS 0.026899f
C14110 mux8_7.NAND4F_8.Y.t14 VSS 0.033983f
C14111 mux8_7.NAND4F_8.Y.n2 VSS 0.072608f
C14112 mux8_7.NAND4F_8.Y.n3 VSS 0.045714f
C14113 mux8_7.NAND4F_8.Y.n4 VSS 0.037354f
C14114 mux8_7.NAND4F_8.Y.n5 VSS 0.018278f
C14115 mux8_7.NAND4F_8.Y.t4 VSS 0.026614f
C14116 mux8_7.NAND4F_8.Y.t3 VSS 0.026614f
C14117 mux8_7.NAND4F_8.Y.n6 VSS 0.0618f
C14118 mux8_7.NAND4F_8.Y.t5 VSS 0.026614f
C14119 mux8_7.NAND4F_8.Y.t6 VSS 0.026614f
C14120 mux8_7.NAND4F_8.Y.n7 VSS 0.061615f
C14121 mux8_7.NAND4F_8.Y.t7 VSS 0.026614f
C14122 mux8_7.NAND4F_8.Y.t8 VSS 0.026614f
C14123 mux8_7.NAND4F_8.Y.n8 VSS 0.061615f
C14124 mux8_7.NAND4F_8.Y.t0 VSS 0.026614f
C14125 mux8_7.NAND4F_8.Y.t1 VSS 0.026614f
C14126 mux8_7.NAND4F_8.Y.n9 VSS 0.061615f
C14127 mux8_7.NAND4F_8.Y.n10 VSS 0.268281f
C14128 mux8_7.NAND4F_8.Y.t2 VSS 0.21369f
C14129 mux8_7.NAND4F_2.Y.n0 VSS 0.530078f
C14130 mux8_7.NAND4F_2.Y.t7 VSS 0.026135f
C14131 mux8_7.NAND4F_2.Y.t8 VSS 0.026135f
C14132 mux8_7.NAND4F_2.Y.n1 VSS 0.060687f
C14133 mux8_7.NAND4F_2.Y.t3 VSS 0.026135f
C14134 mux8_7.NAND4F_2.Y.t2 VSS 0.026135f
C14135 mux8_7.NAND4F_2.Y.n2 VSS 0.060505f
C14136 mux8_7.NAND4F_2.Y.t5 VSS 0.026135f
C14137 mux8_7.NAND4F_2.Y.t6 VSS 0.026135f
C14138 mux8_7.NAND4F_2.Y.n3 VSS 0.060505f
C14139 mux8_7.NAND4F_2.Y.t0 VSS 0.026135f
C14140 mux8_7.NAND4F_2.Y.t4 VSS 0.026135f
C14141 mux8_7.NAND4F_2.Y.n4 VSS 0.060505f
C14142 mux8_7.NAND4F_2.Y.n5 VSS 0.263447f
C14143 mux8_7.NAND4F_2.Y.t1 VSS 0.213114f
C14144 mux8_7.NAND4F_2.Y.t9 VSS 0.034088f
C14145 mux8_7.NAND4F_2.Y.t10 VSS 0.105185f
C14146 mux8_7.NAND4F_2.Y.t11 VSS 0.039267f
C14147 mux8_7.NAND4F_2.Y.n6 VSS 0.131989f
C14148 mux8_7.NAND4F_2.Y.n7 VSS 0.028742f
C14149 mux8_7.NAND4F_2.Y.n8 VSS 1.53344f
C14150 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n0 VSS 0.941081f
C14151 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t0 VSS 0.008143f
C14152 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t1 VSS 0.008143f
C14153 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n1 VSS 0.018168f
C14154 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t5 VSS 0.008143f
C14155 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t2 VSS 0.008143f
C14156 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n2 VSS 0.018119f
C14157 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t3 VSS 0.008143f
C14158 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t4 VSS 0.008143f
C14159 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n3 VSS 0.018119f
C14160 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t6 VSS 0.049166f
C14161 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t13 VSS 0.027811f
C14162 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t10 VSS 0.027465f
C14163 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t12 VSS 0.027465f
C14164 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t9 VSS 0.027465f
C14165 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n4 VSS 0.109319f
C14166 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t17 VSS 0.005708f
C14167 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t14 VSS 0.005708f
C14168 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t8 VSS 0.005708f
C14169 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t15 VSS 0.005708f
C14170 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n5 VSS 0.103275f
C14171 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n6 VSS 0.161516f
C14172 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t18 VSS 0.025683f
C14173 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t7 VSS 0.009858f
C14174 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t16 VSS 0.013614f
C14175 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n7 VSS 0.01567f
C14176 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.t11 VSS 0.010363f
C14177 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n8 VSS 0.015891f
C14178 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n9 VSS 0.053976f
C14179 MULT_0.4bit_ADDER_1.FULL_ADDER_3.COUT.n10 VSS 0.358938f
C14180 mux8_2.NAND4F_5.Y.n0 VSS 0.25108f
C14181 mux8_2.NAND4F_5.Y.t10 VSS 0.017162f
C14182 mux8_2.NAND4F_5.Y.t11 VSS 0.050565f
C14183 mux8_2.NAND4F_5.Y.t9 VSS 0.016698f
C14184 mux8_2.NAND4F_5.Y.n1 VSS 0.086077f
C14185 mux8_2.NAND4F_5.Y.t1 VSS 0.099394f
C14186 mux8_2.NAND4F_5.Y.n2 VSS 0.798124f
C14187 mux8_2.NAND4F_5.Y.t8 VSS 0.012379f
C14188 mux8_2.NAND4F_5.Y.t7 VSS 0.012379f
C14189 mux8_2.NAND4F_5.Y.n3 VSS 0.028745f
C14190 mux8_2.NAND4F_5.Y.t3 VSS 0.012379f
C14191 mux8_2.NAND4F_5.Y.t4 VSS 0.012379f
C14192 mux8_2.NAND4F_5.Y.n4 VSS 0.028659f
C14193 mux8_2.NAND4F_5.Y.t6 VSS 0.012379f
C14194 mux8_2.NAND4F_5.Y.t5 VSS 0.012379f
C14195 mux8_2.NAND4F_5.Y.n5 VSS 0.028659f
C14196 mux8_2.NAND4F_5.Y.t0 VSS 0.012379f
C14197 mux8_2.NAND4F_5.Y.t2 VSS 0.012379f
C14198 mux8_2.NAND4F_5.Y.n6 VSS 0.028659f
C14199 mux8_2.NAND4F_5.Y.n7 VSS 0.117805f
C14200 SEL1.t52 VSS 0.057826f
C14201 SEL1.t95 VSS 0.08072f
C14202 SEL1.t142 VSS 0.08072f
C14203 SEL1.n0 VSS 0.252826f
C14204 SEL1.t35 VSS 0.088396f
C14205 SEL1.t134 VSS 0.279168f
C14206 SEL1.t126 VSS 0.089052f
C14207 SEL1.t29 VSS 0.089052f
C14208 SEL1.n1 VSS 0.10455f
C14209 SEL1.n2 VSS 0.586373f
C14210 SEL1.t53 VSS 0.279168f
C14211 SEL1.t105 VSS 0.089052f
C14212 SEL1.t4 VSS 0.089052f
C14213 SEL1.n3 VSS 0.10455f
C14214 SEL1.n4 VSS 0.586185f
C14215 SEL1.n5 VSS 1.24067f
C14216 SEL1.n6 VSS 2.32934f
C14217 SEL1.t2 VSS 0.089052f
C14218 SEL1.t78 VSS 0.089052f
C14219 SEL1.n7 VSS 0.10455f
C14220 SEL1.t90 VSS 0.279168f
C14221 SEL1.n8 VSS 0.586277f
C14222 SEL1.n9 VSS 0.44444f
C14223 SEL1.t19 VSS 0.089052f
C14224 SEL1.t87 VSS 0.089052f
C14225 SEL1.n10 VSS 0.10455f
C14226 SEL1.t67 VSS 0.279168f
C14227 SEL1.n11 VSS 0.58626f
C14228 SEL1.n12 VSS 0.373286f
C14229 SEL1.n13 VSS 1.46522f
C14230 SEL1.n14 VSS 1.39969f
C14231 SEL1.n15 VSS 0.387297f
C14232 SEL1.n16 VSS 0.180714f
C14233 SEL1.n17 VSS 0.195966f
C14234 SEL1.n18 VSS 0.182076f
C14235 SEL1.t16 VSS 0.057826f
C14236 SEL1.t9 VSS 0.08072f
C14237 SEL1.t69 VSS 0.08072f
C14238 SEL1.n19 VSS 0.252826f
C14239 SEL1.t91 VSS 0.088396f
C14240 SEL1.t41 VSS 0.279168f
C14241 SEL1.t73 VSS 0.089052f
C14242 SEL1.t10 VSS 0.089052f
C14243 SEL1.n20 VSS 0.10455f
C14244 SEL1.n21 VSS 0.586373f
C14245 SEL1.t79 VSS 0.279168f
C14246 SEL1.t92 VSS 0.089052f
C14247 SEL1.t38 VSS 0.089052f
C14248 SEL1.n22 VSS 0.10455f
C14249 SEL1.n23 VSS 0.586185f
C14250 SEL1.n24 VSS 1.24067f
C14251 SEL1.n25 VSS 2.32934f
C14252 SEL1.t135 VSS 0.089052f
C14253 SEL1.t47 VSS 0.089052f
C14254 SEL1.n26 VSS 0.10455f
C14255 SEL1.t129 VSS 0.279168f
C14256 SEL1.n27 VSS 0.586277f
C14257 SEL1.n28 VSS 0.44444f
C14258 SEL1.t111 VSS 0.089052f
C14259 SEL1.t25 VSS 0.089052f
C14260 SEL1.n29 VSS 0.10455f
C14261 SEL1.t85 VSS 0.279168f
C14262 SEL1.n30 VSS 0.58626f
C14263 SEL1.n31 VSS 0.373286f
C14264 SEL1.n32 VSS 1.46522f
C14265 SEL1.n33 VSS 1.39969f
C14266 SEL1.n34 VSS 0.387297f
C14267 SEL1.n35 VSS 0.180714f
C14268 SEL1.n36 VSS 0.195966f
C14269 SEL1.n37 VSS 0.180672f
C14270 SEL1.n38 VSS 1.18334f
C14271 SEL1.t15 VSS 0.057826f
C14272 SEL1.t115 VSS 0.08072f
C14273 SEL1.t31 VSS 0.08072f
C14274 SEL1.n39 VSS 0.252826f
C14275 SEL1.t97 VSS 0.088396f
C14276 SEL1.t75 VSS 0.279168f
C14277 SEL1.t103 VSS 0.089052f
C14278 SEL1.t51 VSS 0.089052f
C14279 SEL1.n40 VSS 0.10455f
C14280 SEL1.n41 VSS 0.586373f
C14281 SEL1.t109 VSS 0.279168f
C14282 SEL1.t130 VSS 0.089052f
C14283 SEL1.t71 VSS 0.089052f
C14284 SEL1.n42 VSS 0.10455f
C14285 SEL1.n43 VSS 0.586185f
C14286 SEL1.n44 VSS 1.24067f
C14287 SEL1.n45 VSS 2.32934f
C14288 SEL1.t128 VSS 0.089052f
C14289 SEL1.t39 VSS 0.089052f
C14290 SEL1.n46 VSS 0.10455f
C14291 SEL1.t21 VSS 0.279168f
C14292 SEL1.n47 VSS 0.586277f
C14293 SEL1.n48 VSS 0.44444f
C14294 SEL1.t102 VSS 0.089052f
C14295 SEL1.t11 VSS 0.089052f
C14296 SEL1.n49 VSS 0.10455f
C14297 SEL1.t131 VSS 0.279168f
C14298 SEL1.n50 VSS 0.58626f
C14299 SEL1.n51 VSS 0.373286f
C14300 SEL1.n52 VSS 1.46522f
C14301 SEL1.n53 VSS 1.39969f
C14302 SEL1.n54 VSS 0.387297f
C14303 SEL1.n55 VSS 0.180714f
C14304 SEL1.n56 VSS 0.195966f
C14305 SEL1.n57 VSS 0.180711f
C14306 SEL1.n58 VSS 0.215745f
C14307 SEL1.n59 VSS 5.09279f
C14308 SEL1.t62 VSS 0.057826f
C14309 SEL1.t6 VSS 0.08072f
C14310 SEL1.t65 VSS 0.08072f
C14311 SEL1.n60 VSS 0.252826f
C14312 SEL1.t24 VSS 0.088396f
C14313 SEL1.t40 VSS 0.279168f
C14314 SEL1.t70 VSS 0.089052f
C14315 SEL1.t5 VSS 0.089052f
C14316 SEL1.n61 VSS 0.10455f
C14317 SEL1.n62 VSS 0.586373f
C14318 SEL1.t76 VSS 0.279168f
C14319 SEL1.t88 VSS 0.089052f
C14320 SEL1.t34 VSS 0.089052f
C14321 SEL1.n63 VSS 0.10455f
C14322 SEL1.n64 VSS 0.586185f
C14323 SEL1.n65 VSS 1.24067f
C14324 SEL1.n66 VSS 2.32934f
C14325 SEL1.t64 VSS 0.089052f
C14326 SEL1.t120 VSS 0.089052f
C14327 SEL1.n67 VSS 0.10455f
C14328 SEL1.t7 VSS 0.279168f
C14329 SEL1.n68 VSS 0.586277f
C14330 SEL1.n69 VSS 0.44444f
C14331 SEL1.t46 VSS 0.089052f
C14332 SEL1.t98 VSS 0.089052f
C14333 SEL1.n70 VSS 0.10455f
C14334 SEL1.t119 VSS 0.279168f
C14335 SEL1.n71 VSS 0.58626f
C14336 SEL1.n72 VSS 0.373286f
C14337 SEL1.n73 VSS 1.46522f
C14338 SEL1.n74 VSS 1.39969f
C14339 SEL1.n75 VSS 0.387297f
C14340 SEL1.n76 VSS 0.180714f
C14341 SEL1.n77 VSS 0.195966f
C14342 SEL1.n78 VSS 0.181393f
C14343 SEL1.n79 VSS 0.222593f
C14344 SEL1.n80 VSS 4.01704f
C14345 SEL1.t14 VSS 0.057826f
C14346 SEL1.t114 VSS 0.08072f
C14347 SEL1.t74 VSS 0.08072f
C14348 SEL1.n81 VSS 0.252826f
C14349 SEL1.t133 VSS 0.088396f
C14350 SEL1.t106 VSS 0.279168f
C14351 SEL1.t101 VSS 0.089052f
C14352 SEL1.t49 VSS 0.089052f
C14353 SEL1.n82 VSS 0.10455f
C14354 SEL1.n83 VSS 0.586373f
C14355 SEL1.t139 VSS 0.279168f
C14356 SEL1.t127 VSS 0.089052f
C14357 SEL1.t68 VSS 0.089052f
C14358 SEL1.n84 VSS 0.10455f
C14359 SEL1.n85 VSS 0.586185f
C14360 SEL1.n86 VSS 1.24067f
C14361 SEL1.n87 VSS 2.32934f
C14362 SEL1.t20 VSS 0.089052f
C14363 SEL1.t77 VSS 0.089052f
C14364 SEL1.n88 VSS 0.10455f
C14365 SEL1.t50 VSS 0.279168f
C14366 SEL1.n89 VSS 0.586277f
C14367 SEL1.n90 VSS 0.44444f
C14368 SEL1.t140 VSS 0.089052f
C14369 SEL1.t60 VSS 0.089052f
C14370 SEL1.n91 VSS 0.10455f
C14371 SEL1.t3 VSS 0.279168f
C14372 SEL1.n92 VSS 0.58626f
C14373 SEL1.n93 VSS 0.373286f
C14374 SEL1.n94 VSS 1.46522f
C14375 SEL1.n95 VSS 1.39969f
C14376 SEL1.n96 VSS 0.387297f
C14377 SEL1.n97 VSS 0.180714f
C14378 SEL1.n98 VSS 0.195966f
C14379 SEL1.n99 VSS 0.180907f
C14380 SEL1.n100 VSS 0.217759f
C14381 SEL1.n101 VSS 4.01483f
C14382 SEL1.t93 VSS 0.057826f
C14383 SEL1.t86 VSS 0.08072f
C14384 SEL1.t136 VSS 0.08072f
C14385 SEL1.n102 VSS 0.252826f
C14386 SEL1.t18 VSS 0.088396f
C14387 SEL1.t72 VSS 0.279168f
C14388 SEL1.t100 VSS 0.089052f
C14389 SEL1.t48 VSS 0.089052f
C14390 SEL1.n103 VSS 0.10455f
C14391 SEL1.n104 VSS 0.586373f
C14392 SEL1.t107 VSS 0.279168f
C14393 SEL1.t122 VSS 0.089052f
C14394 SEL1.t66 VSS 0.089052f
C14395 SEL1.n105 VSS 0.10455f
C14396 SEL1.n106 VSS 0.586185f
C14397 SEL1.n107 VSS 1.24067f
C14398 SEL1.n108 VSS 2.32934f
C14399 SEL1.t63 VSS 0.089052f
C14400 SEL1.t117 VSS 0.089052f
C14401 SEL1.n109 VSS 0.10455f
C14402 SEL1.t57 VSS 0.279168f
C14403 SEL1.n110 VSS 0.586277f
C14404 SEL1.n111 VSS 0.44444f
C14405 SEL1.t43 VSS 0.089052f
C14406 SEL1.t96 VSS 0.089052f
C14407 SEL1.n112 VSS 0.10455f
C14408 SEL1.t13 VSS 0.279168f
C14409 SEL1.n113 VSS 0.58626f
C14410 SEL1.n114 VSS 0.373286f
C14411 SEL1.n115 VSS 1.46522f
C14412 SEL1.n116 VSS 1.39969f
C14413 SEL1.n117 VSS 0.387297f
C14414 SEL1.n118 VSS 0.180714f
C14415 SEL1.n119 VSS 0.195966f
C14416 SEL1.n120 VSS 0.181393f
C14417 SEL1.n121 VSS 0.222593f
C14418 SEL1.n122 VSS 4.0104f
C14419 SEL1.t32 VSS 0.057826f
C14420 SEL1.t28 VSS 0.08072f
C14421 SEL1.t81 VSS 0.08072f
C14422 SEL1.n123 VSS 0.252826f
C14423 SEL1.t94 VSS 0.088396f
C14424 SEL1.t143 VSS 0.279168f
C14425 SEL1.t36 VSS 0.089052f
C14426 SEL1.t121 VSS 0.089052f
C14427 SEL1.n124 VSS 0.10455f
C14428 SEL1.n125 VSS 0.586373f
C14429 SEL1.t42 VSS 0.279168f
C14430 SEL1.t58 VSS 0.089052f
C14431 SEL1.t137 VSS 0.089052f
C14432 SEL1.n126 VSS 0.10455f
C14433 SEL1.n127 VSS 0.586185f
C14434 SEL1.n128 VSS 1.24067f
C14435 SEL1.n129 VSS 2.32934f
C14436 SEL1.t132 VSS 0.089052f
C14437 SEL1.t44 VSS 0.089052f
C14438 SEL1.n130 VSS 0.10455f
C14439 SEL1.t124 VSS 0.279168f
C14440 SEL1.n131 VSS 0.586277f
C14441 SEL1.n132 VSS 0.44444f
C14442 SEL1.t108 VSS 0.089052f
C14443 SEL1.t23 VSS 0.089052f
C14444 SEL1.n133 VSS 0.10455f
C14445 SEL1.t83 VSS 0.279168f
C14446 SEL1.n134 VSS 0.58626f
C14447 SEL1.n135 VSS 0.373286f
C14448 SEL1.n136 VSS 1.46522f
C14449 SEL1.n137 VSS 1.39969f
C14450 SEL1.n138 VSS 0.387297f
C14451 SEL1.n139 VSS 0.180714f
C14452 SEL1.n140 VSS 0.195966f
C14453 SEL1.n141 VSS 0.180519f
C14454 SEL1.n142 VSS 0.213714f
C14455 SEL1.n143 VSS 4.05828f
C14456 SEL1.t12 VSS 0.057826f
C14457 SEL1.t112 VSS 0.08072f
C14458 SEL1.t22 VSS 0.08072f
C14459 SEL1.n144 VSS 0.252826f
C14460 SEL1.t125 VSS 0.088396f
C14461 SEL1.t123 VSS 0.279168f
C14462 SEL1.t0 VSS 0.089052f
C14463 SEL1.t59 VSS 0.089052f
C14464 SEL1.n145 VSS 0.10455f
C14465 SEL1.n146 VSS 0.586373f
C14466 SEL1.t45 VSS 0.279168f
C14467 SEL1.t116 VSS 0.089052f
C14468 SEL1.t27 VSS 0.089052f
C14469 SEL1.n147 VSS 0.10455f
C14470 SEL1.n148 VSS 0.586185f
C14471 SEL1.n149 VSS 1.24067f
C14472 SEL1.n150 VSS 2.32934f
C14473 SEL1.t17 VSS 0.089052f
C14474 SEL1.t113 VSS 0.089052f
C14475 SEL1.n151 VSS 0.10455f
C14476 SEL1.t89 VSS 0.279168f
C14477 SEL1.n152 VSS 0.586277f
C14478 SEL1.n153 VSS 0.44444f
C14479 SEL1.t54 VSS 0.089052f
C14480 SEL1.t138 VSS 0.089052f
C14481 SEL1.n154 VSS 0.10455f
C14482 SEL1.t26 VSS 0.279168f
C14483 SEL1.n155 VSS 0.58626f
C14484 SEL1.n156 VSS 0.373286f
C14485 SEL1.n157 VSS 1.46522f
C14486 SEL1.n158 VSS 1.39969f
C14487 SEL1.n159 VSS 0.387297f
C14488 SEL1.n160 VSS 0.180714f
C14489 SEL1.n161 VSS 0.195966f
C14490 SEL1.n162 VSS 0.181311f
C14491 SEL1.n163 VSS 0.221789f
C14492 SEL1.n164 VSS 4.03611f
C14493 SEL1.t99 VSS 0.057826f
C14494 SEL1.t55 VSS 0.08072f
C14495 SEL1.t104 VSS 0.08072f
C14496 SEL1.n165 VSS 0.252826f
C14497 SEL1.t118 VSS 0.088396f
C14498 SEL1.t110 VSS 0.279168f
C14499 SEL1.t37 VSS 0.089052f
C14500 SEL1.t84 VSS 0.089052f
C14501 SEL1.n166 VSS 0.10455f
C14502 SEL1.n167 VSS 0.586373f
C14503 SEL1.t33 VSS 0.279168f
C14504 SEL1.t1 VSS 0.089052f
C14505 SEL1.t61 VSS 0.089052f
C14506 SEL1.n168 VSS 0.10455f
C14507 SEL1.n169 VSS 0.586185f
C14508 SEL1.n170 VSS 1.24067f
C14509 SEL1.n171 VSS 2.32934f
C14510 SEL1.t56 VSS 0.089052f
C14511 SEL1.t141 VSS 0.089052f
C14512 SEL1.n172 VSS 0.10455f
C14513 SEL1.t80 VSS 0.279168f
C14514 SEL1.n173 VSS 0.586277f
C14515 SEL1.n174 VSS 0.44444f
C14516 SEL1.t82 VSS 0.089052f
C14517 SEL1.t30 VSS 0.089052f
C14518 SEL1.n175 VSS 0.10455f
C14519 SEL1.t8 VSS 0.279168f
C14520 SEL1.n176 VSS 0.58626f
C14521 SEL1.n177 VSS 0.373286f
C14522 SEL1.n178 VSS 1.46522f
C14523 SEL1.n179 VSS 1.39969f
C14524 SEL1.n180 VSS 0.387297f
C14525 SEL1.n181 VSS 0.180714f
C14526 SEL1.n182 VSS 0.195966f
C14527 SEL1.n183 VSS 0.182432f
C14528 SEL1.n184 VSS 5.05492f
C14529 SEL1.n185 VSS 1.20652f
C14530 MULT_0.4bit_ADDER_1.A3.n0 VSS 0.674688f
C14531 MULT_0.inv_13.Y VSS 0.416771f
C14532 MULT_0.4bit_ADDER_1.FULL_ADDER_0.XOR2_0.B VSS 0.273791f
C14533 MULT_0.4bit_ADDER_1.FULL_ADDER_0.A VSS 0.118003f
C14534 MULT_0.4bit_ADDER_1.A3.t6 VSS 0.020858f
C14535 MULT_0.4bit_ADDER_1.A3.t10 VSS 0.008006f
C14536 MULT_0.4bit_ADDER_1.A3.t4 VSS 0.011057f
C14537 MULT_0.4bit_ADDER_1.A3.n1 VSS 0.012726f
C14538 MULT_0.4bit_ADDER_1.A3.t14 VSS 0.008416f
C14539 MULT_0.4bit_ADDER_1.A3.n2 VSS 0.012906f
C14540 MULT_0.4bit_ADDER_1.A3.n3 VSS 0.053421f
C14541 MULT_0.4bit_ADDER_1.FULL_ADDER_0.NAND2_0.B VSS 0.206403f
C14542 MULT_0.4bit_ADDER_1.A3.t9 VSS 0.022586f
C14543 MULT_0.4bit_ADDER_1.A3.t5 VSS 0.022305f
C14544 MULT_0.4bit_ADDER_1.A3.t7 VSS 0.022305f
C14545 MULT_0.4bit_ADDER_1.A3.t12 VSS 0.022305f
C14546 MULT_0.4bit_ADDER_1.A3.n4 VSS 0.088781f
C14547 MULT_0.4bit_ADDER_1.A3.t13 VSS 0.004635f
C14548 MULT_0.4bit_ADDER_1.A3.t8 VSS 0.004635f
C14549 MULT_0.4bit_ADDER_1.A3.t15 VSS 0.004635f
C14550 MULT_0.4bit_ADDER_1.A3.t11 VSS 0.004635f
C14551 MULT_0.4bit_ADDER_1.A3.n5 VSS 0.083872f
C14552 MULT_0.4bit_ADDER_1.A3.n6 VSS 0.131194f
C14553 MULT_0.4bit_ADDER_1.A3.t2 VSS 0.006613f
C14554 MULT_0.4bit_ADDER_1.A3.t1 VSS 0.006613f
C14555 MULT_0.4bit_ADDER_1.A3.n7 VSS 0.014731f
C14556 MULT_0.4bit_ADDER_1.A3.t0 VSS 0.019122f
C14557 MULT_0.4bit_ADDER_1.A3.t3 VSS 0.023985f
C14558 MULT_0.inv_13.A.n0 VSS 1.37982f
C14559 MULT_0.inv_13.A.t1 VSS 0.022953f
C14560 MULT_0.inv_13.A.t2 VSS 0.022953f
C14561 MULT_0.inv_13.A.n1 VSS 0.051213f
C14562 MULT_0.inv_13.A.t5 VSS 0.022953f
C14563 MULT_0.inv_13.A.t0 VSS 0.022953f
C14564 MULT_0.inv_13.A.n2 VSS 0.051074f
C14565 MULT_0.inv_13.A.t3 VSS 0.022953f
C14566 MULT_0.inv_13.A.t4 VSS 0.022953f
C14567 MULT_0.inv_13.A.n3 VSS 0.051074f
C14568 MULT_0.inv_13.A.t10 VSS 0.029252f
C14569 MULT_0.inv_13.A.t9 VSS 0.040833f
C14570 MULT_0.inv_13.A.t7 VSS 0.040833f
C14571 MULT_0.inv_13.A.n4 VSS 0.133283f
C14572 MULT_0.inv_13.A.t8 VSS 0.046622f
C14573 MULT_0.inv_13.A.t6 VSS 0.138274f
C14574 mux8_1.NAND4F_8.Y.n0 VSS 0.539804f
C14575 mux8_1.NAND4F_8.Y.t9 VSS 0.026899f
C14576 mux8_1.NAND4F_8.Y.t14 VSS 0.028853f
C14577 mux8_1.NAND4F_8.Y.n1 VSS 0.042994f
C14578 mux8_1.NAND4F_8.Y.t13 VSS 0.026899f
C14579 mux8_1.NAND4F_8.Y.t12 VSS 0.026899f
C14580 mux8_1.NAND4F_8.Y.t11 VSS 0.026899f
C14581 mux8_1.NAND4F_8.Y.t10 VSS 0.033983f
C14582 mux8_1.NAND4F_8.Y.n2 VSS 0.072608f
C14583 mux8_1.NAND4F_8.Y.n3 VSS 0.045714f
C14584 mux8_1.NAND4F_8.Y.n4 VSS 0.037354f
C14585 mux8_1.NAND4F_8.Y.n5 VSS 0.018278f
C14586 mux8_1.NAND4F_8.Y.t6 VSS 0.026614f
C14587 mux8_1.NAND4F_8.Y.t7 VSS 0.026614f
C14588 mux8_1.NAND4F_8.Y.n6 VSS 0.0618f
C14589 mux8_1.NAND4F_8.Y.t4 VSS 0.026614f
C14590 mux8_1.NAND4F_8.Y.t3 VSS 0.026614f
C14591 mux8_1.NAND4F_8.Y.n7 VSS 0.061615f
C14592 mux8_1.NAND4F_8.Y.t8 VSS 0.026614f
C14593 mux8_1.NAND4F_8.Y.t2 VSS 0.026614f
C14594 mux8_1.NAND4F_8.Y.n8 VSS 0.061615f
C14595 mux8_1.NAND4F_8.Y.t1 VSS 0.026614f
C14596 mux8_1.NAND4F_8.Y.t0 VSS 0.026614f
C14597 mux8_1.NAND4F_8.Y.n9 VSS 0.061615f
C14598 mux8_1.NAND4F_8.Y.n10 VSS 0.268281f
C14599 mux8_1.NAND4F_8.Y.t5 VSS 0.21369f
C14600 mux8_5.NAND4F_8.Y.n0 VSS 0.539804f
C14601 mux8_5.NAND4F_8.Y.t14 VSS 0.026899f
C14602 mux8_5.NAND4F_8.Y.t13 VSS 0.028853f
C14603 mux8_5.NAND4F_8.Y.n1 VSS 0.042994f
C14604 mux8_5.NAND4F_8.Y.t9 VSS 0.026899f
C14605 mux8_5.NAND4F_8.Y.t11 VSS 0.026899f
C14606 mux8_5.NAND4F_8.Y.t10 VSS 0.026899f
C14607 mux8_5.NAND4F_8.Y.t12 VSS 0.033983f
C14608 mux8_5.NAND4F_8.Y.n2 VSS 0.072608f
C14609 mux8_5.NAND4F_8.Y.n3 VSS 0.045714f
C14610 mux8_5.NAND4F_8.Y.n4 VSS 0.037354f
C14611 mux8_5.NAND4F_8.Y.n5 VSS 0.018278f
C14612 mux8_5.NAND4F_8.Y.t6 VSS 0.026614f
C14613 mux8_5.NAND4F_8.Y.t5 VSS 0.026614f
C14614 mux8_5.NAND4F_8.Y.n6 VSS 0.0618f
C14615 mux8_5.NAND4F_8.Y.t7 VSS 0.026614f
C14616 mux8_5.NAND4F_8.Y.t8 VSS 0.026614f
C14617 mux8_5.NAND4F_8.Y.n7 VSS 0.061615f
C14618 mux8_5.NAND4F_8.Y.t3 VSS 0.026614f
C14619 mux8_5.NAND4F_8.Y.t4 VSS 0.026614f
C14620 mux8_5.NAND4F_8.Y.n8 VSS 0.061615f
C14621 mux8_5.NAND4F_8.Y.t0 VSS 0.026614f
C14622 mux8_5.NAND4F_8.Y.t1 VSS 0.026614f
C14623 mux8_5.NAND4F_8.Y.n9 VSS 0.061615f
C14624 mux8_5.NAND4F_8.Y.n10 VSS 0.268281f
C14625 mux8_5.NAND4F_8.Y.t2 VSS 0.21369f
C14626 mux8_2.NAND4F_0.Y.n0 VSS 0.350455f
C14627 mux8_2.NAND4F_0.Y.t11 VSS 0.022537f
C14628 mux8_2.NAND4F_0.Y.t10 VSS 0.079785f
C14629 mux8_2.NAND4F_0.Y.t9 VSS 0.024808f
C14630 mux8_2.NAND4F_0.Y.n1 VSS 0.070768f
C14631 mux8_2.NAND4F_0.Y.n2 VSS 0.020978f
C14632 mux8_2.NAND4F_0.Y.t6 VSS 0.017278f
C14633 mux8_2.NAND4F_0.Y.t5 VSS 0.017278f
C14634 mux8_2.NAND4F_0.Y.n3 VSS 0.040122f
C14635 mux8_2.NAND4F_0.Y.t8 VSS 0.017278f
C14636 mux8_2.NAND4F_0.Y.t7 VSS 0.017278f
C14637 mux8_2.NAND4F_0.Y.n4 VSS 0.040002f
C14638 mux8_2.NAND4F_0.Y.t3 VSS 0.017278f
C14639 mux8_2.NAND4F_0.Y.t4 VSS 0.017278f
C14640 mux8_2.NAND4F_0.Y.n5 VSS 0.040002f
C14641 mux8_2.NAND4F_0.Y.t1 VSS 0.017278f
C14642 mux8_2.NAND4F_0.Y.t0 VSS 0.017278f
C14643 mux8_2.NAND4F_0.Y.n6 VSS 0.040002f
C14644 mux8_2.NAND4F_0.Y.t2 VSS 0.166327f
C14645 VDD.t1247 VSS 0.027215f
C14646 VDD.t375 VSS 0.007233f
C14647 VDD.t1245 VSS 0.007233f
C14648 VDD.n0 VSS 0.016652f
C14649 VDD.n1 VSS 0.129639f
C14650 VDD.t2205 VSS -0.019301f
C14651 VDD.t2207 VSS 0.075145f
C14652 VDD.t1743 VSS 0.075145f
C14653 VDD.t1741 VSS 0.063403f
C14654 VDD.t1945 VSS 0.027215f
C14655 VDD.t1919 VSS 0.007233f
C14656 VDD.t3073 VSS 0.007233f
C14657 VDD.n2 VSS 0.016652f
C14658 VDD.n3 VSS 0.132428f
C14659 VDD.t3039 VSS 0.007233f
C14660 VDD.t645 VSS 0.007233f
C14661 VDD.n4 VSS 0.016652f
C14662 VDD.n5 VSS 0.047679f
C14663 VDD.t643 VSS 0.007233f
C14664 VDD.t2894 VSS 0.007233f
C14665 VDD.n6 VSS 0.016652f
C14666 VDD.n7 VSS 0.073375f
C14667 VDD.t644 VSS 0.042023f
C14668 VDD.t648 VSS 0.075406f
C14669 VDD.t2889 VSS 0.075406f
C14670 VDD.t2891 VSS 0.139422f
C14671 VDD.t1580 VSS 0.139422f
C14672 VDD.t1578 VSS 0.075406f
C14673 VDD.t852 VSS 0.075406f
C14674 VDD.t854 VSS 0.063624f
C14675 VDD.t2900 VSS 0.027188f
C14676 VDD.n8 VSS 0.074488f
C14677 VDD.t1921 VSS 0.027188f
C14678 VDD.n9 VSS 0.074487f
C14679 VDD.t1977 VSS 0.007233f
C14680 VDD.t3043 VSS 0.007233f
C14681 VDD.n10 VSS 0.016652f
C14682 VDD.n11 VSS 0.07634f
C14683 VDD.t2969 VSS 0.007233f
C14684 VDD.t4340 VSS 0.007233f
C14685 VDD.n12 VSS 0.016652f
C14686 VDD.n13 VSS 0.047679f
C14687 VDD.t2944 VSS 0.004807f
C14688 VDD.t2996 VSS 0.004807f
C14689 VDD.n14 VSS 0.010736f
C14690 VDD.t3054 VSS 0.017466f
C14691 VDD.n15 VSS 0.048701f
C14692 VDD.n16 VSS 0.030676f
C14693 VDD.t4405 VSS 0.145552f
C14694 VDD.t4406 VSS 0.004807f
C14695 VDD.t4514 VSS 0.004807f
C14696 VDD.n17 VSS 0.010736f
C14697 VDD.t4457 VSS 0.017466f
C14698 VDD.n18 VSS 0.048701f
C14699 VDD.t3728 VSS 0.004807f
C14700 VDD.t3837 VSS 0.004807f
C14701 VDD.n19 VSS 0.010736f
C14702 VDD.t3761 VSS 0.017466f
C14703 VDD.n20 VSS 0.059157f
C14704 VDD.t3727 VSS 0.137944f
C14705 VDD.n21 VSS 0.135842f
C14706 VDD.n22 VSS 0.031797f
C14707 VDD.n23 VSS 0.030676f
C14708 VDD.n24 VSS 0.028952f
C14709 VDD.n25 VSS 0.135842f
C14710 VDD.t2943 VSS 0.270495f
C14711 VDD.n26 VSS 0.096866f
C14712 VDD.t2888 VSS 0.027204f
C14713 VDD.n27 VSS 0.169958f
C14714 VDD.t4451 VSS 0.007233f
C14715 VDD.t2898 VSS 0.007233f
C14716 VDD.n28 VSS 0.016652f
C14717 VDD.n29 VSS 0.050644f
C14718 VDD.t4339 VSS 0.042023f
C14719 VDD.t4441 VSS 0.075406f
C14720 VDD.t2895 VSS 0.075406f
C14721 VDD.t2901 VSS 0.144962f
C14722 VDD.t1914 VSS 0.14709f
C14723 VDD.t1968 VSS 0.075145f
C14724 VDD.t856 VSS 0.075145f
C14725 VDD.t858 VSS 0.063403f
C14726 VDD.t2887 VSS 0.126024f
C14727 VDD.t2897 VSS 0.075145f
C14728 VDD.t4450 VSS 0.075145f
C14729 VDD.t4362 VSS 0.041877f
C14730 VDD.n30 VSS 0.064693f
C14731 VDD.n31 VSS 0.076519f
C14732 VDD.t859 VSS 0.007233f
C14733 VDD.t4363 VSS 0.007233f
C14734 VDD.n32 VSS 0.016652f
C14735 VDD.n33 VSS 0.047679f
C14736 VDD.t1969 VSS 0.007233f
C14737 VDD.t857 VSS 0.007233f
C14738 VDD.n34 VSS 0.016652f
C14739 VDD.n35 VSS 0.07634f
C14740 VDD.t1915 VSS 0.027188f
C14741 VDD.n36 VSS 0.076455f
C14742 VDD.t2902 VSS 0.027188f
C14743 VDD.n37 VSS 0.076457f
C14744 VDD.t4442 VSS 0.007233f
C14745 VDD.t2896 VSS 0.007233f
C14746 VDD.n38 VSS 0.016652f
C14747 VDD.n39 VSS 0.073375f
C14748 VDD.n40 VSS 0.076519f
C14749 VDD.n41 VSS 0.064809f
C14750 VDD.t2968 VSS 0.063624f
C14751 VDD.t3042 VSS 0.075406f
C14752 VDD.t1976 VSS 0.075406f
C14753 VDD.t1920 VSS 0.141386f
C14754 VDD.t2899 VSS 0.141386f
C14755 VDD.t2893 VSS 0.075406f
C14756 VDD.t642 VSS 0.075406f
C14757 VDD.t640 VSS 0.042023f
C14758 VDD.n42 VSS 0.064809f
C14759 VDD.n43 VSS 0.076519f
C14760 VDD.t855 VSS 0.007233f
C14761 VDD.t641 VSS 0.007233f
C14762 VDD.n44 VSS 0.016652f
C14763 VDD.n45 VSS 0.047679f
C14764 VDD.t1579 VSS 0.007233f
C14765 VDD.t853 VSS 0.007233f
C14766 VDD.n46 VSS 0.016652f
C14767 VDD.n47 VSS 0.07634f
C14768 VDD.t1581 VSS 0.027188f
C14769 VDD.n48 VSS 0.073667f
C14770 VDD.t2892 VSS 0.027188f
C14771 VDD.n49 VSS 0.073669f
C14772 VDD.t649 VSS 0.007233f
C14773 VDD.t2890 VSS 0.007233f
C14774 VDD.n50 VSS 0.016652f
C14775 VDD.n51 VSS 0.073375f
C14776 VDD.n52 VSS 0.076519f
C14777 VDD.n53 VSS 0.064809f
C14778 VDD.t3038 VSS 0.063624f
C14779 VDD.t3072 VSS 0.075406f
C14780 VDD.t1918 VSS 0.075406f
C14781 VDD.t1944 VSS 0.13786f
C14782 VDD.t1246 VSS 0.137401f
C14783 VDD.t1244 VSS 0.075145f
C14784 VDD.t374 VSS 0.075145f
C14785 VDD.t372 VSS 0.041877f
C14786 VDD.n54 VSS 0.064693f
C14787 VDD.n55 VSS 0.076519f
C14788 VDD.t1742 VSS 0.007233f
C14789 VDD.t373 VSS 0.007233f
C14790 VDD.n56 VSS 0.016652f
C14791 VDD.n57 VSS 0.047679f
C14792 VDD.t2208 VSS 0.007233f
C14793 VDD.t1744 VSS 0.007233f
C14794 VDD.n58 VSS 0.016652f
C14795 VDD.n59 VSS 0.07634f
C14796 VDD.t2206 VSS 0.027188f
C14797 VDD.n60 VSS 0.110894f
C14798 VDD.n61 VSS 1.68467f
C14799 VDD.t3333 VSS 0.027215f
C14800 VDD.t931 VSS 0.007233f
C14801 VDD.t3331 VSS 0.007233f
C14802 VDD.n62 VSS 0.016652f
C14803 VDD.n63 VSS 0.129639f
C14804 VDD.t770 VSS -0.019301f
C14805 VDD.t768 VSS 0.075145f
C14806 VDD.t4064 VSS 0.075145f
C14807 VDD.t925 VSS 0.063403f
C14808 VDD.t99 VSS 0.027215f
C14809 VDD.t97 VSS 0.007233f
C14810 VDD.t3045 VSS 0.007233f
C14811 VDD.n64 VSS 0.016652f
C14812 VDD.n65 VSS 0.132428f
C14813 VDD.t3056 VSS 0.007233f
C14814 VDD.t67 VSS 0.007233f
C14815 VDD.n66 VSS 0.016652f
C14816 VDD.n67 VSS 0.047679f
C14817 VDD.t69 VSS 0.007233f
C14818 VDD.t1712 VSS 0.007233f
C14819 VDD.n68 VSS 0.016652f
C14820 VDD.n69 VSS 0.073375f
C14821 VDD.t66 VSS 0.042023f
C14822 VDD.t1419 VSS 0.075406f
C14823 VDD.t1715 VSS 0.075406f
C14824 VDD.t1713 VSS 0.139422f
C14825 VDD.t3357 VSS 0.139422f
C14826 VDD.t3355 VSS 0.075406f
C14827 VDD.t1261 VSS 0.075406f
C14828 VDD.t1273 VSS 0.063624f
C14829 VDD.t1706 VSS 0.027188f
C14830 VDD.n70 VSS 0.074488f
C14831 VDD.t881 VSS 0.027188f
C14832 VDD.n71 VSS 0.074487f
C14833 VDD.t883 VSS 0.007233f
C14834 VDD.t2973 VSS 0.007233f
C14835 VDD.n72 VSS 0.016652f
C14836 VDD.n73 VSS 0.07634f
C14837 VDD.t3013 VSS 0.007233f
C14838 VDD.t4412 VSS 0.007233f
C14839 VDD.n74 VSS 0.016652f
C14840 VDD.n75 VSS 0.047679f
C14841 VDD.t3053 VSS 0.004807f
C14842 VDD.t3050 VSS 0.004807f
C14843 VDD.n76 VSS 0.010736f
C14844 VDD.t2934 VSS 0.017466f
C14845 VDD.n77 VSS 0.048701f
C14846 VDD.n78 VSS 0.030676f
C14847 VDD.t4409 VSS 0.145552f
C14848 VDD.t4462 VSS 0.004807f
C14849 VDD.t4471 VSS 0.004807f
C14850 VDD.n79 VSS 0.010736f
C14851 VDD.t4410 VSS 0.017466f
C14852 VDD.n80 VSS 0.048701f
C14853 VDD.t3766 VSS 0.004807f
C14854 VDD.t3774 VSS 0.004807f
C14855 VDD.n81 VSS 0.010736f
C14856 VDD.t3730 VSS 0.017466f
C14857 VDD.n82 VSS 0.059157f
C14858 VDD.t3729 VSS 0.137944f
C14859 VDD.n83 VSS 0.135842f
C14860 VDD.n84 VSS 0.031797f
C14861 VDD.n85 VSS 0.030676f
C14862 VDD.n86 VSS 0.028952f
C14863 VDD.n87 VSS 0.135842f
C14864 VDD.t2933 VSS 0.270495f
C14865 VDD.n88 VSS 0.096866f
C14866 VDD.t1708 VSS 0.027204f
C14867 VDD.n89 VSS 0.169958f
C14868 VDD.t4378 VSS 0.007233f
C14869 VDD.t1710 VSS 0.007233f
C14870 VDD.n90 VSS 0.016652f
C14871 VDD.n91 VSS 0.050644f
C14872 VDD.t4411 VSS 0.042023f
C14873 VDD.t4512 VSS 0.075406f
C14874 VDD.t1719 VSS 0.075406f
C14875 VDD.t1717 VSS 0.144962f
C14876 VDD.t579 VSS 0.14709f
C14877 VDD.t577 VSS 0.075145f
C14878 VDD.t1269 VSS 0.075145f
C14879 VDD.t1265 VSS 0.063403f
C14880 VDD.t1707 VSS 0.126024f
C14881 VDD.t1709 VSS 0.075145f
C14882 VDD.t4377 VSS 0.075145f
C14883 VDD.t4444 VSS 0.041877f
C14884 VDD.n92 VSS 0.064693f
C14885 VDD.n93 VSS 0.076519f
C14886 VDD.t1266 VSS 0.007233f
C14887 VDD.t4445 VSS 0.007233f
C14888 VDD.n94 VSS 0.016652f
C14889 VDD.n95 VSS 0.047679f
C14890 VDD.t578 VSS 0.007233f
C14891 VDD.t1270 VSS 0.007233f
C14892 VDD.n96 VSS 0.016652f
C14893 VDD.n97 VSS 0.07634f
C14894 VDD.t580 VSS 0.027188f
C14895 VDD.n98 VSS 0.076455f
C14896 VDD.t1718 VSS 0.027188f
C14897 VDD.n99 VSS 0.076457f
C14898 VDD.t4513 VSS 0.007233f
C14899 VDD.t1720 VSS 0.007233f
C14900 VDD.n100 VSS 0.016652f
C14901 VDD.n101 VSS 0.073375f
C14902 VDD.n102 VSS 0.076519f
C14903 VDD.n103 VSS 0.064809f
C14904 VDD.t3012 VSS 0.063624f
C14905 VDD.t2972 VSS 0.075406f
C14906 VDD.t882 VSS 0.075406f
C14907 VDD.t880 VSS 0.141386f
C14908 VDD.t1705 VSS 0.141386f
C14909 VDD.t1711 VSS 0.075406f
C14910 VDD.t68 VSS 0.075406f
C14911 VDD.t72 VSS 0.042023f
C14912 VDD.n104 VSS 0.064809f
C14913 VDD.n105 VSS 0.076519f
C14914 VDD.t1274 VSS 0.007233f
C14915 VDD.t73 VSS 0.007233f
C14916 VDD.n106 VSS 0.016652f
C14917 VDD.n107 VSS 0.047679f
C14918 VDD.t3356 VSS 0.007233f
C14919 VDD.t1262 VSS 0.007233f
C14920 VDD.n108 VSS 0.016652f
C14921 VDD.n109 VSS 0.07634f
C14922 VDD.t3358 VSS 0.027188f
C14923 VDD.n110 VSS 0.073667f
C14924 VDD.t1714 VSS 0.027188f
C14925 VDD.n111 VSS 0.073669f
C14926 VDD.t1420 VSS 0.007233f
C14927 VDD.t1716 VSS 0.007233f
C14928 VDD.n112 VSS 0.016652f
C14929 VDD.n113 VSS 0.073375f
C14930 VDD.n114 VSS 0.076519f
C14931 VDD.n115 VSS 0.064809f
C14932 VDD.t3055 VSS 0.063624f
C14933 VDD.t3044 VSS 0.075406f
C14934 VDD.t96 VSS 0.075406f
C14935 VDD.t98 VSS 0.13786f
C14936 VDD.t3332 VSS 0.137401f
C14937 VDD.t3330 VSS 0.075145f
C14938 VDD.t930 VSS 0.075145f
C14939 VDD.t932 VSS 0.041877f
C14940 VDD.n116 VSS 0.064693f
C14941 VDD.n117 VSS 0.076519f
C14942 VDD.t926 VSS 0.007233f
C14943 VDD.t933 VSS 0.007233f
C14944 VDD.n118 VSS 0.016652f
C14945 VDD.n119 VSS 0.047679f
C14946 VDD.t769 VSS 0.007233f
C14947 VDD.t4065 VSS 0.007233f
C14948 VDD.n120 VSS 0.016652f
C14949 VDD.n121 VSS 0.07634f
C14950 VDD.t771 VSS 0.027188f
C14951 VDD.n122 VSS 0.110894f
C14952 VDD.t1100 VSS 0.004807f
C14953 VDD.t1102 VSS 0.004807f
C14954 VDD.n123 VSS 0.010736f
C14955 VDD.t1104 VSS 0.017466f
C14956 VDD.n124 VSS 0.056287f
C14957 VDD.n125 VSS 0.020342f
C14958 VDD.n126 VSS 0.030311f
C14959 VDD.t1101 VSS 0.089594f
C14960 VDD.n127 VSS 0.035424f
C14961 VDD.t1099 VSS 0.05332f
C14962 VDD.t1103 VSS 0.027493f
C14963 VDD.n128 VSS 0.067089f
C14964 VDD.n129 VSS 0.044915f
C14965 VDD.t1322 VSS 0.081296f
C14966 VDD.t1321 VSS 0.075406f
C14967 VDD.t1320 VSS 0.075406f
C14968 VDD.t1319 VSS 0.075406f
C14969 VDD.t1318 VSS 0.075406f
C14970 VDD.t4314 VSS 0.075406f
C14971 VDD.t4322 VSS 0.075406f
C14972 VDD.t4320 VSS 0.058518f
C14973 VDD.t4316 VSS 0.126462f
C14974 VDD.t4318 VSS 0.05459f
C14975 VDD.n130 VSS 2.52e-19
C14976 VDD.t4315 VSS 0.00575f
C14977 VDD.t4323 VSS 0.00575f
C14978 VDD.n131 VSS 0.0115f
C14979 VDD.n132 VSS 0.012479f
C14980 VDD.t4321 VSS 0.00575f
C14981 VDD.t4319 VSS 0.00575f
C14982 VDD.n133 VSS 0.0115f
C14983 VDD.n134 VSS 0.007448f
C14984 VDD.n135 VSS 0.076419f
C14985 VDD.t4317 VSS 0.01978f
C14986 VDD.n136 VSS 0.014195f
C14987 VDD.n137 VSS -0.011842f
C14988 VDD.n138 VSS 0.077508f
C14989 VDD.n139 VSS 0.837038f
C14990 VDD.n140 VSS 0.45705f
C14991 VDD.n141 VSS 1.37899f
C14992 VDD.t1091 VSS 0.004807f
C14993 VDD.t1093 VSS 0.004807f
C14994 VDD.n142 VSS 0.010725f
C14995 VDD.t1095 VSS 0.017454f
C14996 VDD.n143 VSS 0.059309f
C14997 VDD.n144 VSS 0.019394f
C14998 VDD.t1135 VSS 0.004807f
C14999 VDD.t1136 VSS 0.004807f
C15000 VDD.n145 VSS 0.010725f
C15001 VDD.t1137 VSS 0.017454f
C15002 VDD.n146 VSS 0.048725f
C15003 VDD.t1092 VSS 0.173365f
C15004 VDD.t1090 VSS 0.103373f
C15005 VDD.t1094 VSS 0.116295f
C15006 VDD.n147 VSS 0.110877f
C15007 VDD.n148 VSS 0.035039f
C15008 VDD.n149 VSS 0.039312f
C15009 VDD.n150 VSS 0.017043f
C15010 VDD.n151 VSS 1.61911f
C15011 VDD.t2065 VSS 0.027215f
C15012 VDD.t2028 VSS 0.007233f
C15013 VDD.t414 VSS 0.007233f
C15014 VDD.n152 VSS 0.016652f
C15015 VDD.n153 VSS 0.129639f
C15016 VDD.t490 VSS -0.019301f
C15017 VDD.t492 VSS 0.075145f
C15018 VDD.t271 VSS 0.075145f
C15019 VDD.t273 VSS 0.063403f
C15020 VDD.t416 VSS 0.027215f
C15021 VDD.t418 VSS 0.007233f
C15022 VDD.t2998 VSS 0.007233f
C15023 VDD.n154 VSS 0.016652f
C15024 VDD.n155 VSS 0.132756f
C15025 VDD.t2993 VSS 0.007233f
C15026 VDD.t568 VSS 0.007233f
C15027 VDD.n156 VSS 0.016652f
C15028 VDD.n157 VSS 0.047679f
C15029 VDD.t326 VSS 0.007233f
C15030 VDD.t3765 VSS 0.007233f
C15031 VDD.n158 VSS 0.016652f
C15032 VDD.n159 VSS 0.073624f
C15033 VDD.t567 VSS 0.04195f
C15034 VDD.t569 VSS 0.075275f
C15035 VDD.t3744 VSS 0.075275f
C15036 VDD.t3748 VSS 0.139181f
C15037 VDD.t3265 VSS 0.139181f
C15038 VDD.t3267 VSS 0.075275f
C15039 VDD.t10 VSS 0.075275f
C15040 VDD.t2451 VSS 0.063514f
C15041 VDD.t3779 VSS 0.027188f
C15042 VDD.n160 VSS 0.07466f
C15043 VDD.t280 VSS 0.027188f
C15044 VDD.n161 VSS 0.074656f
C15045 VDD.t282 VSS 0.007233f
C15046 VDD.t2979 VSS 0.007233f
C15047 VDD.n162 VSS 0.016652f
C15048 VDD.n163 VSS 0.076601f
C15049 VDD.t3063 VSS 0.007233f
C15050 VDD.t4388 VSS 0.007233f
C15051 VDD.n164 VSS 0.016652f
C15052 VDD.n165 VSS 0.047822f
C15053 VDD.t3833 VSS 0.027215f
C15054 VDD.t4437 VSS 0.007233f
C15055 VDD.t3771 VSS 0.007233f
C15056 VDD.n166 VSS 0.016652f
C15057 VDD.n167 VSS 0.130541f
C15058 VDD.t4387 VSS 0.04195f
C15059 VDD.t4454 VSS 0.075275f
C15060 VDD.t3801 VSS 0.075275f
C15061 VDD.t3809 VSS 0.145846f
C15062 VDD.t357 VSS 0.145846f
C15063 VDD.t359 VSS 0.075275f
C15064 VDD.t2455 VSS 0.075275f
C15065 VDD.t4 VSS 0.063514f
C15066 VDD.t3832 VSS 0.126243f
C15067 VDD.t3770 VSS 0.075275f
C15068 VDD.t4436 VSS 0.075275f
C15069 VDD.t4349 VSS 0.04195f
C15070 VDD.n168 VSS 0.064751f
C15071 VDD.n169 VSS 0.07665f
C15072 VDD.t5 VSS 0.007233f
C15073 VDD.t4350 VSS 0.007233f
C15074 VDD.n170 VSS 0.016652f
C15075 VDD.n171 VSS 0.047822f
C15076 VDD.t360 VSS 0.007233f
C15077 VDD.t2456 VSS 0.007233f
C15078 VDD.n172 VSS 0.016652f
C15079 VDD.n173 VSS 0.076601f
C15080 VDD.t358 VSS 0.027188f
C15081 VDD.n174 VSS 0.076624f
C15082 VDD.t3810 VSS 0.027188f
C15083 VDD.n175 VSS 0.076629f
C15084 VDD.t4455 VSS 0.007233f
C15085 VDD.t3802 VSS 0.007233f
C15086 VDD.n176 VSS 0.016652f
C15087 VDD.n177 VSS 0.073624f
C15088 VDD.n178 VSS 0.07665f
C15089 VDD.n179 VSS 0.064751f
C15090 VDD.t3062 VSS 0.063514f
C15091 VDD.t2978 VSS 0.075275f
C15092 VDD.t281 VSS 0.075275f
C15093 VDD.t279 VSS 0.141141f
C15094 VDD.t3778 VSS 0.141141f
C15095 VDD.t3764 VSS 0.075275f
C15096 VDD.t325 VSS 0.075275f
C15097 VDD.t323 VSS 0.04195f
C15098 VDD.n180 VSS 0.064751f
C15099 VDD.n181 VSS 0.07665f
C15100 VDD.t2452 VSS 0.007233f
C15101 VDD.t324 VSS 0.007233f
C15102 VDD.n182 VSS 0.016652f
C15103 VDD.n183 VSS 0.047822f
C15104 VDD.t3268 VSS 0.007233f
C15105 VDD.t11 VSS 0.007233f
C15106 VDD.n184 VSS 0.016652f
C15107 VDD.n185 VSS 0.076601f
C15108 VDD.t3266 VSS 0.027188f
C15109 VDD.n186 VSS 0.073849f
C15110 VDD.t3749 VSS 0.027188f
C15111 VDD.n187 VSS 0.073656f
C15112 VDD.t570 VSS 0.007233f
C15113 VDD.t3745 VSS 0.007233f
C15114 VDD.n188 VSS 0.016652f
C15115 VDD.n189 VSS 0.073375f
C15116 VDD.n190 VSS 0.076519f
C15117 VDD.n191 VSS 0.064751f
C15118 VDD.t2992 VSS 0.063514f
C15119 VDD.t2997 VSS 0.075275f
C15120 VDD.t417 VSS 0.075275f
C15121 VDD.t415 VSS 0.137602f
C15122 VDD.t2064 VSS 0.137365f
C15123 VDD.t413 VSS 0.075145f
C15124 VDD.t2027 VSS 0.075145f
C15125 VDD.t2025 VSS 0.041877f
C15126 VDD.n192 VSS 0.064693f
C15127 VDD.n193 VSS 0.076519f
C15128 VDD.t274 VSS 0.007233f
C15129 VDD.t2026 VSS 0.007233f
C15130 VDD.n194 VSS 0.016652f
C15131 VDD.n195 VSS 0.047679f
C15132 VDD.t493 VSS 0.007233f
C15133 VDD.t272 VSS 0.007233f
C15134 VDD.n196 VSS 0.016652f
C15135 VDD.n197 VSS 0.07634f
C15136 VDD.t491 VSS 0.027188f
C15137 VDD.n198 VSS 0.256185f
C15138 VDD.n199 VSS 1.70334f
C15139 VDD.t863 VSS 0.027215f
C15140 VDD.t1454 VSS 0.007233f
C15141 VDD.t865 VSS 0.007233f
C15142 VDD.n200 VSS 0.016652f
C15143 VDD.n201 VSS 0.129639f
C15144 VDD.t912 VSS -0.019301f
C15145 VDD.t910 VSS 0.075145f
C15146 VDD.t2765 VSS 0.075145f
C15147 VDD.t2767 VSS 0.063403f
C15148 VDD.t3339 VSS 0.027215f
C15149 VDD.t3341 VSS 0.007233f
C15150 VDD.t2954 VSS 0.007233f
C15151 VDD.n202 VSS 0.016652f
C15152 VDD.n203 VSS 0.132428f
C15153 VDD.t2942 VSS 0.007233f
C15154 VDD.t328 VSS 0.007233f
C15155 VDD.n204 VSS 0.016652f
C15156 VDD.n205 VSS 0.047679f
C15157 VDD.t566 VSS 0.007233f
C15158 VDD.t420 VSS 0.007233f
C15159 VDD.n206 VSS 0.016652f
C15160 VDD.n207 VSS 0.073375f
C15161 VDD.t327 VSS 0.042023f
C15162 VDD.t329 VSS 0.075406f
C15163 VDD.t431 VSS 0.075406f
C15164 VDD.t433 VSS 0.139422f
C15165 VDD.t3306 VSS 0.139422f
C15166 VDD.t3298 VSS 0.075406f
C15167 VDD.t6 VSS 0.075406f
C15168 VDD.t8 VSS 0.063624f
C15169 VDD.t424 VSS 0.027188f
C15170 VDD.n208 VSS 0.074488f
C15171 VDD.t1223 VSS 0.027188f
C15172 VDD.n209 VSS 0.074487f
C15173 VDD.t1225 VSS 0.007233f
C15174 VDD.t3011 VSS 0.007233f
C15175 VDD.n210 VSS 0.016652f
C15176 VDD.n211 VSS 0.07634f
C15177 VDD.t2958 VSS 0.007233f
C15178 VDD.t4504 VSS 0.007233f
C15179 VDD.n212 VSS 0.016652f
C15180 VDD.n213 VSS 0.047679f
C15181 VDD.t2999 VSS 0.004807f
C15182 VDD.t2950 VSS 0.004807f
C15183 VDD.n214 VSS 0.010736f
C15184 VDD.t3006 VSS 0.017466f
C15185 VDD.n215 VSS 0.048701f
C15186 VDD.n216 VSS 0.030676f
C15187 VDD.t4347 VSS 0.145552f
C15188 VDD.t4359 VSS 0.004807f
C15189 VDD.t4431 VSS 0.004807f
C15190 VDD.n217 VSS 0.010736f
C15191 VDD.t4348 VSS 0.017466f
C15192 VDD.n218 VSS 0.048701f
C15193 VDD.t3726 VSS 0.004807f
C15194 VDD.t3758 VSS 0.004807f
C15195 VDD.n219 VSS 0.010736f
C15196 VDD.t3715 VSS 0.017466f
C15197 VDD.n220 VSS 0.059157f
C15198 VDD.t3714 VSS 0.137944f
C15199 VDD.n221 VSS 0.135842f
C15200 VDD.n222 VSS 0.031797f
C15201 VDD.n223 VSS 0.030676f
C15202 VDD.n224 VSS 0.028952f
C15203 VDD.n225 VSS 0.135842f
C15204 VDD.t2949 VSS 0.270495f
C15205 VDD.n226 VSS 0.096866f
C15206 VDD.t430 VSS 0.027204f
C15207 VDD.n227 VSS 0.169958f
C15208 VDD.t4370 VSS 0.007233f
C15209 VDD.t422 VSS 0.007233f
C15210 VDD.n228 VSS 0.016652f
C15211 VDD.n229 VSS 0.050644f
C15212 VDD.t4503 VSS 0.042023f
C15213 VDD.t4397 VSS 0.075406f
C15214 VDD.t425 VSS 0.075406f
C15215 VDD.t427 VSS 0.144962f
C15216 VDD.t506 VSS 0.14709f
C15217 VDD.t508 VSS 0.075145f
C15218 VDD.t12 VSS 0.075145f
C15219 VDD.t2453 VSS 0.063403f
C15220 VDD.t429 VSS 0.126024f
C15221 VDD.t421 VSS 0.075145f
C15222 VDD.t4369 VSS 0.075145f
C15223 VDD.t4476 VSS 0.041877f
C15224 VDD.n230 VSS 0.064693f
C15225 VDD.n231 VSS 0.076519f
C15226 VDD.t2454 VSS 0.007233f
C15227 VDD.t4477 VSS 0.007233f
C15228 VDD.n232 VSS 0.016652f
C15229 VDD.n233 VSS 0.047679f
C15230 VDD.t509 VSS 0.007233f
C15231 VDD.t13 VSS 0.007233f
C15232 VDD.n234 VSS 0.016652f
C15233 VDD.n235 VSS 0.07634f
C15234 VDD.t507 VSS 0.027188f
C15235 VDD.n236 VSS 0.076455f
C15236 VDD.t428 VSS 0.027188f
C15237 VDD.n237 VSS 0.076457f
C15238 VDD.t4398 VSS 0.007233f
C15239 VDD.t426 VSS 0.007233f
C15240 VDD.n238 VSS 0.016652f
C15241 VDD.n239 VSS 0.073375f
C15242 VDD.n240 VSS 0.076519f
C15243 VDD.n241 VSS 0.064809f
C15244 VDD.t2957 VSS 0.063624f
C15245 VDD.t3010 VSS 0.075406f
C15246 VDD.t1224 VSS 0.075406f
C15247 VDD.t1222 VSS 0.141386f
C15248 VDD.t423 VSS 0.141386f
C15249 VDD.t419 VSS 0.075406f
C15250 VDD.t565 VSS 0.075406f
C15251 VDD.t331 VSS 0.042023f
C15252 VDD.n242 VSS 0.064809f
C15253 VDD.n243 VSS 0.076519f
C15254 VDD.t9 VSS 0.007233f
C15255 VDD.t332 VSS 0.007233f
C15256 VDD.n244 VSS 0.016652f
C15257 VDD.n245 VSS 0.047679f
C15258 VDD.t3299 VSS 0.007233f
C15259 VDD.t7 VSS 0.007233f
C15260 VDD.n246 VSS 0.016652f
C15261 VDD.n247 VSS 0.07634f
C15262 VDD.t3307 VSS 0.027188f
C15263 VDD.n248 VSS 0.073667f
C15264 VDD.t434 VSS 0.027188f
C15265 VDD.n249 VSS 0.073669f
C15266 VDD.t330 VSS 0.007233f
C15267 VDD.t432 VSS 0.007233f
C15268 VDD.n250 VSS 0.016652f
C15269 VDD.n251 VSS 0.073375f
C15270 VDD.n252 VSS 0.076519f
C15271 VDD.n253 VSS 0.064809f
C15272 VDD.t2941 VSS 0.063624f
C15273 VDD.t2953 VSS 0.075406f
C15274 VDD.t3340 VSS 0.075406f
C15275 VDD.t3338 VSS 0.13786f
C15276 VDD.t862 VSS 0.137401f
C15277 VDD.t864 VSS 0.075145f
C15278 VDD.t1453 VSS 0.075145f
C15279 VDD.t1451 VSS 0.041877f
C15280 VDD.n254 VSS 0.064693f
C15281 VDD.n255 VSS 0.076519f
C15282 VDD.t2768 VSS 0.007233f
C15283 VDD.t1452 VSS 0.007233f
C15284 VDD.n256 VSS 0.016652f
C15285 VDD.n257 VSS 0.047679f
C15286 VDD.t911 VSS 0.007233f
C15287 VDD.t2766 VSS 0.007233f
C15288 VDD.n258 VSS 0.016652f
C15289 VDD.n259 VSS 0.07634f
C15290 VDD.t913 VSS 0.027188f
C15291 VDD.n260 VSS 0.110894f
C15292 VDD.t1690 VSS 0.004807f
C15293 VDD.t1692 VSS 0.004807f
C15294 VDD.n261 VSS 0.010736f
C15295 VDD.t1688 VSS 0.017466f
C15296 VDD.n262 VSS 0.056287f
C15297 VDD.n263 VSS 0.020342f
C15298 VDD.n264 VSS 0.030311f
C15299 VDD.t1691 VSS 0.089594f
C15300 VDD.n265 VSS 0.035424f
C15301 VDD.t1689 VSS 0.05332f
C15302 VDD.t1687 VSS 0.027493f
C15303 VDD.n266 VSS 0.067089f
C15304 VDD.n267 VSS 0.044915f
C15305 VDD.t696 VSS 0.081296f
C15306 VDD.t697 VSS 0.075406f
C15307 VDD.t698 VSS 0.075406f
C15308 VDD.t694 VSS 0.075406f
C15309 VDD.t695 VSS 0.075406f
C15310 VDD.t982 VSS 0.075406f
C15311 VDD.t984 VSS 0.075406f
C15312 VDD.t2905 VSS 0.058518f
C15313 VDD.t2907 VSS 0.126462f
C15314 VDD.t2903 VSS 0.05459f
C15315 VDD.n268 VSS 2.52e-19
C15316 VDD.t983 VSS 0.00575f
C15317 VDD.t985 VSS 0.00575f
C15318 VDD.n269 VSS 0.0115f
C15319 VDD.n270 VSS 0.012479f
C15320 VDD.t2906 VSS 0.00575f
C15321 VDD.t2904 VSS 0.00575f
C15322 VDD.n271 VSS 0.0115f
C15323 VDD.n272 VSS 0.007448f
C15324 VDD.n273 VSS 0.076419f
C15325 VDD.t2908 VSS 0.01978f
C15326 VDD.n274 VSS 0.014195f
C15327 VDD.n275 VSS -0.011842f
C15328 VDD.n276 VSS 0.077508f
C15329 VDD.n277 VSS 0.836811f
C15330 VDD.n278 VSS 1.44523f
C15331 VDD.n279 VSS 1.3074f
C15332 VDD.n280 VSS 1.34966f
C15333 VDD.t2570 VSS 0.027215f
C15334 VDD.t1445 VSS 0.007233f
C15335 VDD.t2572 VSS 0.007233f
C15336 VDD.n281 VSS 0.016652f
C15337 VDD.n282 VSS 0.129639f
C15338 VDD.t2284 VSS -0.019301f
C15339 VDD.t2286 VSS 0.075145f
C15340 VDD.t355 VSS 0.075145f
C15341 VDD.t353 VSS 0.063403f
C15342 VDD.t2283 VSS 0.027215f
C15343 VDD.t2281 VSS 0.007233f
C15344 VDD.t3086 VSS 0.007233f
C15345 VDD.n283 VSS 0.016652f
C15346 VDD.n284 VSS 0.132756f
C15347 VDD.t3070 VSS 0.007233f
C15348 VDD.t2660 VSS 0.007233f
C15349 VDD.n285 VSS 0.016652f
C15350 VDD.n286 VSS 0.047679f
C15351 VDD.t2658 VSS 0.007233f
C15352 VDD.t3816 VSS 0.007233f
C15353 VDD.n287 VSS 0.016652f
C15354 VDD.n288 VSS 0.073624f
C15355 VDD.t2659 VSS 0.04195f
C15356 VDD.t2661 VSS 0.075275f
C15357 VDD.t3844 VSS 0.075275f
C15358 VDD.t3862 VSS 0.139181f
C15359 VDD.t3990 VSS 0.139181f
C15360 VDD.t3992 VSS 0.075275f
C15361 VDD.t3163 VSS 0.075275f
C15362 VDD.t3165 VSS 0.063514f
C15363 VDD.t3830 VSS 0.027188f
C15364 VDD.n289 VSS 0.07466f
C15365 VDD.t1065 VSS 0.027188f
C15366 VDD.n290 VSS 0.074656f
C15367 VDD.t1067 VSS 0.007233f
C15368 VDD.t3098 VSS 0.007233f
C15369 VDD.n291 VSS 0.016652f
C15370 VDD.n292 VSS 0.076601f
C15371 VDD.t3021 VSS 0.007233f
C15372 VDD.t4435 VSS 0.007233f
C15373 VDD.n293 VSS 0.016652f
C15374 VDD.n294 VSS 0.047822f
C15375 VDD.t3705 VSS 0.027215f
C15376 VDD.t4470 VSS 0.007233f
C15377 VDD.t3822 VSS 0.007233f
C15378 VDD.n295 VSS 0.016652f
C15379 VDD.n296 VSS 0.130541f
C15380 VDD.t4434 VSS 0.04195f
C15381 VDD.t4499 VSS 0.075275f
C15382 VDD.t3860 VSS 0.075275f
C15383 VDD.t3874 VSS 0.145846f
C15384 VDD.t1860 VSS 0.145846f
C15385 VDD.t1862 VSS 0.075275f
C15386 VDD.t3151 VSS 0.075275f
C15387 VDD.t3155 VSS 0.063514f
C15388 VDD.t3704 VSS 0.126243f
C15389 VDD.t3821 VSS 0.075275f
C15390 VDD.t4469 VSS 0.075275f
C15391 VDD.t4403 VSS 0.04195f
C15392 VDD.n297 VSS 0.064751f
C15393 VDD.n298 VSS 0.07665f
C15394 VDD.t3156 VSS 0.007233f
C15395 VDD.t4404 VSS 0.007233f
C15396 VDD.n299 VSS 0.016652f
C15397 VDD.n300 VSS 0.047822f
C15398 VDD.t1863 VSS 0.007233f
C15399 VDD.t3152 VSS 0.007233f
C15400 VDD.n301 VSS 0.016652f
C15401 VDD.n302 VSS 0.076601f
C15402 VDD.t1861 VSS 0.027188f
C15403 VDD.n303 VSS 0.076624f
C15404 VDD.t3875 VSS 0.027188f
C15405 VDD.n304 VSS 0.076629f
C15406 VDD.t4500 VSS 0.007233f
C15407 VDD.t3861 VSS 0.007233f
C15408 VDD.n305 VSS 0.016652f
C15409 VDD.n306 VSS 0.073624f
C15410 VDD.n307 VSS 0.07665f
C15411 VDD.n308 VSS 0.064751f
C15412 VDD.t3020 VSS 0.063514f
C15413 VDD.t3097 VSS 0.075275f
C15414 VDD.t1066 VSS 0.075275f
C15415 VDD.t1064 VSS 0.141141f
C15416 VDD.t3829 VSS 0.141141f
C15417 VDD.t3815 VSS 0.075275f
C15418 VDD.t2657 VSS 0.075275f
C15419 VDD.t2655 VSS 0.04195f
C15420 VDD.n309 VSS 0.064751f
C15421 VDD.n310 VSS 0.07665f
C15422 VDD.t3166 VSS 0.007233f
C15423 VDD.t2656 VSS 0.007233f
C15424 VDD.n311 VSS 0.016652f
C15425 VDD.n312 VSS 0.047822f
C15426 VDD.t3993 VSS 0.007233f
C15427 VDD.t3164 VSS 0.007233f
C15428 VDD.n313 VSS 0.016652f
C15429 VDD.n314 VSS 0.076601f
C15430 VDD.t3991 VSS 0.027188f
C15431 VDD.n315 VSS 0.073849f
C15432 VDD.t3863 VSS 0.027188f
C15433 VDD.n316 VSS 0.073656f
C15434 VDD.t2662 VSS 0.007233f
C15435 VDD.t3845 VSS 0.007233f
C15436 VDD.n317 VSS 0.016652f
C15437 VDD.n318 VSS 0.073375f
C15438 VDD.n319 VSS 0.076519f
C15439 VDD.n320 VSS 0.064751f
C15440 VDD.t3069 VSS 0.063514f
C15441 VDD.t3085 VSS 0.075275f
C15442 VDD.t2280 VSS 0.075275f
C15443 VDD.t2282 VSS 0.137602f
C15444 VDD.t2569 VSS 0.137365f
C15445 VDD.t2571 VSS 0.075145f
C15446 VDD.t1444 VSS 0.075145f
C15447 VDD.t1442 VSS 0.041877f
C15448 VDD.n321 VSS 0.064693f
C15449 VDD.n322 VSS 0.076519f
C15450 VDD.t354 VSS 0.007233f
C15451 VDD.t1443 VSS 0.007233f
C15452 VDD.n323 VSS 0.016652f
C15453 VDD.n324 VSS 0.047679f
C15454 VDD.t2287 VSS 0.007233f
C15455 VDD.t356 VSS 0.007233f
C15456 VDD.n325 VSS 0.016652f
C15457 VDD.n326 VSS 0.07634f
C15458 VDD.t2285 VSS 0.027188f
C15459 VDD.n327 VSS 0.256185f
C15460 VDD.n328 VSS 1.55094f
C15461 VDD.t167 VSS 0.027215f
C15462 VDD.t3337 VSS 0.007233f
C15463 VDD.t169 VSS 0.007233f
C15464 VDD.n329 VSS 0.016652f
C15465 VDD.n330 VSS 0.129639f
C15466 VDD.t1470 VSS -0.019301f
C15467 VDD.t1472 VSS 0.075145f
C15468 VDD.t1160 VSS 0.075145f
C15469 VDD.t1162 VSS 0.063403f
C15470 VDD.t2491 VSS 0.027215f
C15471 VDD.t2493 VSS 0.007233f
C15472 VDD.t2975 VSS 0.007233f
C15473 VDD.n331 VSS 0.016652f
C15474 VDD.n332 VSS 0.132428f
C15475 VDD.t2956 VSS 0.007233f
C15476 VDD.t2652 VSS 0.007233f
C15477 VDD.n333 VSS 0.016652f
C15478 VDD.n334 VSS 0.047679f
C15479 VDD.t2666 VSS 0.007233f
C15480 VDD.t1134 VSS 0.007233f
C15481 VDD.n335 VSS 0.016652f
C15482 VDD.n336 VSS 0.073375f
C15483 VDD.t2651 VSS 0.042023f
C15484 VDD.t2653 VSS 0.075406f
C15485 VDD.t1513 VSS 0.075406f
C15486 VDD.t1515 VSS 0.139422f
C15487 VDD.t1497 VSS 0.139422f
C15488 VDD.t1495 VSS 0.075406f
C15489 VDD.t3153 VSS 0.075406f
C15490 VDD.t3157 VSS 0.063624f
C15491 VDD.t1506 VSS 0.027188f
C15492 VDD.n337 VSS 0.074488f
C15493 VDD.t3144 VSS 0.027188f
C15494 VDD.n338 VSS 0.074487f
C15495 VDD.t3146 VSS 0.007233f
C15496 VDD.t3023 VSS 0.007233f
C15497 VDD.n339 VSS 0.016652f
C15498 VDD.n340 VSS 0.07634f
C15499 VDD.t2977 VSS 0.007233f
C15500 VDD.t4498 VSS 0.007233f
C15501 VDD.n341 VSS 0.016652f
C15502 VDD.n342 VSS 0.047679f
C15503 VDD.t3000 VSS 0.004807f
C15504 VDD.t2989 VSS 0.004807f
C15505 VDD.n343 VSS 0.010736f
C15506 VDD.t3059 VSS 0.017466f
C15507 VDD.n344 VSS 0.048701f
C15508 VDD.n345 VSS 0.030676f
C15509 VDD.t4357 VSS 0.145552f
C15510 VDD.t4358 VSS 0.004807f
C15511 VDD.t4379 VSS 0.004807f
C15512 VDD.n346 VSS 0.010736f
C15513 VDD.t4482 VSS 0.017466f
C15514 VDD.n347 VSS 0.048701f
C15515 VDD.t3725 VSS 0.004807f
C15516 VDD.t3737 VSS 0.004807f
C15517 VDD.n348 VSS 0.010736f
C15518 VDD.t3836 VSS 0.017466f
C15519 VDD.n349 VSS 0.059157f
C15520 VDD.t3724 VSS 0.137944f
C15521 VDD.n350 VSS 0.135842f
C15522 VDD.n351 VSS 0.031797f
C15523 VDD.n352 VSS 0.030676f
C15524 VDD.n353 VSS 0.028952f
C15525 VDD.n354 VSS 0.135842f
C15526 VDD.t2988 VSS 0.270495f
C15527 VDD.n355 VSS 0.096866f
C15528 VDD.t1512 VSS 0.027204f
C15529 VDD.n356 VSS 0.169958f
C15530 VDD.t4352 VSS 0.007233f
C15531 VDD.t1504 VSS 0.007233f
C15532 VDD.n357 VSS 0.016652f
C15533 VDD.n358 VSS 0.050644f
C15534 VDD.t4497 VSS 0.042023f
C15535 VDD.t4389 VSS 0.075406f
C15536 VDD.t1507 VSS 0.075406f
C15537 VDD.t1509 VSS 0.144962f
C15538 VDD.t1232 VSS 0.14709f
C15539 VDD.t1234 VSS 0.075145f
C15540 VDD.t3159 VSS 0.075145f
C15541 VDD.t3161 VSS 0.063403f
C15542 VDD.t1511 VSS 0.126024f
C15543 VDD.t1503 VSS 0.075145f
C15544 VDD.t4351 VSS 0.075145f
C15545 VDD.t4467 VSS 0.041877f
C15546 VDD.n359 VSS 0.064693f
C15547 VDD.n360 VSS 0.076519f
C15548 VDD.t3162 VSS 0.007233f
C15549 VDD.t4468 VSS 0.007233f
C15550 VDD.n361 VSS 0.016652f
C15551 VDD.n362 VSS 0.047679f
C15552 VDD.t1235 VSS 0.007233f
C15553 VDD.t3160 VSS 0.007233f
C15554 VDD.n363 VSS 0.016652f
C15555 VDD.n364 VSS 0.07634f
C15556 VDD.t1233 VSS 0.027188f
C15557 VDD.n365 VSS 0.076455f
C15558 VDD.t1510 VSS 0.027188f
C15559 VDD.n366 VSS 0.076457f
C15560 VDD.t4390 VSS 0.007233f
C15561 VDD.t1508 VSS 0.007233f
C15562 VDD.n367 VSS 0.016652f
C15563 VDD.n368 VSS 0.073375f
C15564 VDD.n369 VSS 0.076519f
C15565 VDD.n370 VSS 0.064809f
C15566 VDD.t2976 VSS 0.063624f
C15567 VDD.t3022 VSS 0.075406f
C15568 VDD.t3145 VSS 0.075406f
C15569 VDD.t3143 VSS 0.141386f
C15570 VDD.t1505 VSS 0.141386f
C15571 VDD.t1133 VSS 0.075406f
C15572 VDD.t2665 VSS 0.075406f
C15573 VDD.t2663 VSS 0.042023f
C15574 VDD.n371 VSS 0.064809f
C15575 VDD.n372 VSS 0.076519f
C15576 VDD.t3158 VSS 0.007233f
C15577 VDD.t2664 VSS 0.007233f
C15578 VDD.n373 VSS 0.016652f
C15579 VDD.n374 VSS 0.047679f
C15580 VDD.t1496 VSS 0.007233f
C15581 VDD.t3154 VSS 0.007233f
C15582 VDD.n375 VSS 0.016652f
C15583 VDD.n376 VSS 0.07634f
C15584 VDD.t1498 VSS 0.027188f
C15585 VDD.n377 VSS 0.073667f
C15586 VDD.t1516 VSS 0.027188f
C15587 VDD.n378 VSS 0.073669f
C15588 VDD.t2654 VSS 0.007233f
C15589 VDD.t1514 VSS 0.007233f
C15590 VDD.n379 VSS 0.016652f
C15591 VDD.n380 VSS 0.073375f
C15592 VDD.n381 VSS 0.076519f
C15593 VDD.n382 VSS 0.064809f
C15594 VDD.t2955 VSS 0.063624f
C15595 VDD.t2974 VSS 0.075406f
C15596 VDD.t2492 VSS 0.075406f
C15597 VDD.t2490 VSS 0.13786f
C15598 VDD.t166 VSS 0.137401f
C15599 VDD.t168 VSS 0.075145f
C15600 VDD.t3336 VSS 0.075145f
C15601 VDD.t3334 VSS 0.041877f
C15602 VDD.n383 VSS 0.064693f
C15603 VDD.n384 VSS 0.076519f
C15604 VDD.t1163 VSS 0.007233f
C15605 VDD.t3335 VSS 0.007233f
C15606 VDD.n385 VSS 0.016652f
C15607 VDD.n386 VSS 0.047679f
C15608 VDD.t1473 VSS 0.007233f
C15609 VDD.t1161 VSS 0.007233f
C15610 VDD.n387 VSS 0.016652f
C15611 VDD.n388 VSS 0.07634f
C15612 VDD.t1471 VSS 0.027188f
C15613 VDD.n389 VSS 0.110894f
C15614 VDD.t2711 VSS 0.004807f
C15615 VDD.t2707 VSS 0.004807f
C15616 VDD.n390 VSS 0.010736f
C15617 VDD.t2709 VSS 0.017466f
C15618 VDD.n391 VSS 0.056287f
C15619 VDD.n392 VSS 0.020342f
C15620 VDD.n393 VSS 0.030311f
C15621 VDD.t2706 VSS 0.089594f
C15622 VDD.n394 VSS 0.035424f
C15623 VDD.t2710 VSS 0.05332f
C15624 VDD.t2708 VSS 0.027493f
C15625 VDD.n395 VSS 0.067089f
C15626 VDD.n396 VSS 0.044915f
C15627 VDD.t1110 VSS 0.081296f
C15628 VDD.t1111 VSS 0.075406f
C15629 VDD.t1112 VSS 0.075406f
C15630 VDD.t1113 VSS 0.075406f
C15631 VDD.t1114 VSS 0.075406f
C15632 VDD.t742 VSS 0.075406f
C15633 VDD.t734 VSS 0.075406f
C15634 VDD.t738 VSS 0.058518f
C15635 VDD.t740 VSS 0.126462f
C15636 VDD.t736 VSS 0.05459f
C15637 VDD.n397 VSS 2.52e-19
C15638 VDD.t743 VSS 0.00575f
C15639 VDD.t735 VSS 0.00575f
C15640 VDD.n398 VSS 0.0115f
C15641 VDD.n399 VSS 0.012479f
C15642 VDD.t739 VSS 0.00575f
C15643 VDD.t737 VSS 0.00575f
C15644 VDD.n400 VSS 0.0115f
C15645 VDD.n401 VSS 0.007448f
C15646 VDD.n402 VSS 0.076419f
C15647 VDD.t741 VSS 0.01978f
C15648 VDD.n403 VSS 0.014195f
C15649 VDD.n404 VSS -0.011842f
C15650 VDD.n405 VSS 0.077508f
C15651 VDD.n406 VSS 0.836811f
C15652 VDD.n407 VSS 1.27315f
C15653 VDD.n408 VSS 1.3177f
C15654 VDD.n409 VSS 1.33436f
C15655 VDD.t48 VSS 0.027215f
C15656 VDD.t2867 VSS 0.007233f
C15657 VDD.t50 VSS 0.007233f
C15658 VDD.n410 VSS 0.016652f
C15659 VDD.n411 VSS 0.129639f
C15660 VDD.t2037 VSS -0.019301f
C15661 VDD.t2039 VSS 0.075145f
C15662 VDD.t2096 VSS 0.075145f
C15663 VDD.t2098 VSS 0.063403f
C15664 VDD.t52 VSS 0.027215f
C15665 VDD.t54 VSS 0.007233f
C15666 VDD.t2962 VSS 0.007233f
C15667 VDD.n412 VSS 0.016652f
C15668 VDD.n413 VSS 0.132756f
C15669 VDD.t2948 VSS 0.007233f
C15670 VDD.t184 VSS 0.007233f
C15671 VDD.n414 VSS 0.016652f
C15672 VDD.n415 VSS 0.047679f
C15673 VDD.t182 VSS 0.007233f
C15674 VDD.t3763 VSS 0.007233f
C15675 VDD.n416 VSS 0.016652f
C15676 VDD.n417 VSS 0.073624f
C15677 VDD.t183 VSS 0.04195f
C15678 VDD.t185 VSS 0.075275f
C15679 VDD.t3787 VSS 0.075275f
C15680 VDD.t3799 VSS 0.139181f
C15681 VDD.t1201 VSS 0.139181f
C15682 VDD.t1203 VSS 0.075275f
C15683 VDD.t199 VSS 0.075275f
C15684 VDD.t201 VSS 0.063514f
C15685 VDD.t3773 VSS 0.027188f
C15686 VDD.n418 VSS 0.07466f
C15687 VDD.t2112 VSS 0.027188f
C15688 VDD.n419 VSS 0.074656f
C15689 VDD.t845 VSS 0.007233f
C15690 VDD.t2981 VSS 0.007233f
C15691 VDD.n420 VSS 0.016652f
C15692 VDD.n421 VSS 0.076601f
C15693 VDD.t3066 VSS 0.007233f
C15694 VDD.t4382 VSS 0.007233f
C15695 VDD.n422 VSS 0.016652f
C15696 VDD.n423 VSS 0.047822f
C15697 VDD.t3828 VSS 0.027215f
C15698 VDD.t4433 VSS 0.007233f
C15699 VDD.t3768 VSS 0.007233f
C15700 VDD.n424 VSS 0.016652f
C15701 VDD.n425 VSS 0.130541f
C15702 VDD.t4381 VSS 0.04195f
C15703 VDD.t4452 VSS 0.075275f
C15704 VDD.t3796 VSS 0.075275f
C15705 VDD.t3805 VSS 0.145846f
C15706 VDD.t1567 VSS 0.145846f
C15707 VDD.t2790 VSS 0.075275f
C15708 VDD.t207 VSS 0.075275f
C15709 VDD.t2048 VSS 0.063514f
C15710 VDD.t3827 VSS 0.126243f
C15711 VDD.t3767 VSS 0.075275f
C15712 VDD.t4432 VSS 0.075275f
C15713 VDD.t4343 VSS 0.04195f
C15714 VDD.n426 VSS 0.064751f
C15715 VDD.n427 VSS 0.07665f
C15716 VDD.t2049 VSS 0.007233f
C15717 VDD.t4344 VSS 0.007233f
C15718 VDD.n428 VSS 0.016652f
C15719 VDD.n429 VSS 0.047822f
C15720 VDD.t2791 VSS 0.007233f
C15721 VDD.t208 VSS 0.007233f
C15722 VDD.n430 VSS 0.016652f
C15723 VDD.n431 VSS 0.076601f
C15724 VDD.t1568 VSS 0.027188f
C15725 VDD.n432 VSS 0.076624f
C15726 VDD.t3806 VSS 0.027188f
C15727 VDD.n433 VSS 0.076629f
C15728 VDD.t4453 VSS 0.007233f
C15729 VDD.t3797 VSS 0.007233f
C15730 VDD.n434 VSS 0.016652f
C15731 VDD.n435 VSS 0.073624f
C15732 VDD.n436 VSS 0.07665f
C15733 VDD.n437 VSS 0.064751f
C15734 VDD.t3065 VSS 0.063514f
C15735 VDD.t2980 VSS 0.075275f
C15736 VDD.t844 VSS 0.075275f
C15737 VDD.t2111 VSS 0.141141f
C15738 VDD.t3772 VSS 0.141141f
C15739 VDD.t3762 VSS 0.075275f
C15740 VDD.t181 VSS 0.075275f
C15741 VDD.t179 VSS 0.04195f
C15742 VDD.n438 VSS 0.064751f
C15743 VDD.n439 VSS 0.07665f
C15744 VDD.t202 VSS 0.007233f
C15745 VDD.t180 VSS 0.007233f
C15746 VDD.n440 VSS 0.016652f
C15747 VDD.n441 VSS 0.047822f
C15748 VDD.t1204 VSS 0.007233f
C15749 VDD.t200 VSS 0.007233f
C15750 VDD.n442 VSS 0.016652f
C15751 VDD.n443 VSS 0.076601f
C15752 VDD.t1202 VSS 0.027188f
C15753 VDD.n444 VSS 0.073849f
C15754 VDD.t3800 VSS 0.027188f
C15755 VDD.n445 VSS 0.073656f
C15756 VDD.t186 VSS 0.007233f
C15757 VDD.t3788 VSS 0.007233f
C15758 VDD.n446 VSS 0.016652f
C15759 VDD.n447 VSS 0.073375f
C15760 VDD.n448 VSS 0.076519f
C15761 VDD.n449 VSS 0.064751f
C15762 VDD.t2947 VSS 0.063514f
C15763 VDD.t2961 VSS 0.075275f
C15764 VDD.t53 VSS 0.075275f
C15765 VDD.t51 VSS 0.137602f
C15766 VDD.t47 VSS 0.137365f
C15767 VDD.t49 VSS 0.075145f
C15768 VDD.t2866 VSS 0.075145f
C15769 VDD.t2864 VSS 0.041877f
C15770 VDD.n450 VSS 0.064693f
C15771 VDD.n451 VSS 0.076519f
C15772 VDD.t2099 VSS 0.007233f
C15773 VDD.t2865 VSS 0.007233f
C15774 VDD.n452 VSS 0.016652f
C15775 VDD.n453 VSS 0.047679f
C15776 VDD.t2040 VSS 0.007233f
C15777 VDD.t2097 VSS 0.007233f
C15778 VDD.n454 VSS 0.016652f
C15779 VDD.n455 VSS 0.07634f
C15780 VDD.t2038 VSS 0.027188f
C15781 VDD.n456 VSS 0.256185f
C15782 VDD.n457 VSS 1.57623f
C15783 VDD.t957 VSS 0.027215f
C15784 VDD.t2550 VSS 0.007233f
C15785 VDD.t959 VSS 0.007233f
C15786 VDD.n458 VSS 0.016652f
C15787 VDD.n459 VSS 0.129639f
C15788 VDD.t510 VSS -0.019301f
C15789 VDD.t512 VSS 0.075145f
C15790 VDD.t4263 VSS 0.075145f
C15791 VDD.t4261 VSS 0.063403f
C15792 VDD.t1108 VSS 0.027215f
C15793 VDD.t1106 VSS 0.007233f
C15794 VDD.t3029 VSS 0.007233f
C15795 VDD.n460 VSS 0.016652f
C15796 VDD.n461 VSS 0.132428f
C15797 VDD.t3017 VSS 0.007233f
C15798 VDD.t192 VSS 0.007233f
C15799 VDD.n462 VSS 0.016652f
C15800 VDD.n463 VSS 0.047679f
C15801 VDD.t190 VSS 0.007233f
C15802 VDD.t3132 VSS 0.007233f
C15803 VDD.n464 VSS 0.016652f
C15804 VDD.n465 VSS 0.073375f
C15805 VDD.t191 VSS 0.042023f
C15806 VDD.t193 VSS 0.075406f
C15807 VDD.t3127 VSS 0.075406f
C15808 VDD.t3129 VSS 0.139422f
C15809 VDD.t605 VSS 0.139422f
C15810 VDD.t607 VSS 0.075406f
C15811 VDD.t203 VSS 0.075406f
C15812 VDD.t205 VSS 0.063624f
C15813 VDD.t3136 VSS 0.027188f
C15814 VDD.n466 VSS 0.074488f
C15815 VDD.t149 VSS 0.027188f
C15816 VDD.n467 VSS 0.074487f
C15817 VDD.t2647 VSS 0.007233f
C15818 VDD.t2928 VSS 0.007233f
C15819 VDD.n468 VSS 0.016652f
C15820 VDD.n469 VSS 0.07634f
C15821 VDD.t3033 VSS 0.007233f
C15822 VDD.t4425 VSS 0.007233f
C15823 VDD.n470 VSS 0.016652f
C15824 VDD.n471 VSS 0.047679f
C15825 VDD.t2965 VSS 0.004807f
C15826 VDD.t2952 VSS 0.004807f
C15827 VDD.n472 VSS 0.010736f
C15828 VDD.t3007 VSS 0.017466f
C15829 VDD.n473 VSS 0.048701f
C15830 VDD.n474 VSS 0.030676f
C15831 VDD.t4345 VSS 0.145552f
C15832 VDD.t4421 VSS 0.004807f
C15833 VDD.t4426 VSS 0.004807f
C15834 VDD.n475 VSS 0.010736f
C15835 VDD.t4346 VSS 0.017466f
C15836 VDD.n476 VSS 0.048701f
C15837 VDD.t3752 VSS 0.004807f
C15838 VDD.t3757 VSS 0.004807f
C15839 VDD.n477 VSS 0.010736f
C15840 VDD.t3709 VSS 0.017466f
C15841 VDD.n478 VSS 0.059157f
C15842 VDD.t3708 VSS 0.137944f
C15843 VDD.n479 VSS 0.135842f
C15844 VDD.n480 VSS 0.031797f
C15845 VDD.n481 VSS 0.030676f
C15846 VDD.n482 VSS 0.028952f
C15847 VDD.n483 VSS 0.135842f
C15848 VDD.t2951 VSS 0.270495f
C15849 VDD.n484 VSS 0.096866f
C15850 VDD.t3142 VSS 0.027204f
C15851 VDD.n485 VSS 0.169958f
C15852 VDD.t4461 VSS 0.007233f
C15853 VDD.t3134 VSS 0.007233f
C15854 VDD.n486 VSS 0.016652f
C15855 VDD.n487 VSS 0.050644f
C15856 VDD.t4424 VSS 0.042023f
C15857 VDD.t4487 VSS 0.075406f
C15858 VDD.t3137 VSS 0.075406f
C15859 VDD.t3139 VSS 0.144962f
C15860 VDD.t502 VSS 0.14709f
C15861 VDD.t504 VSS 0.075145f
C15862 VDD.t2050 VSS 0.075145f
C15863 VDD.t197 VSS 0.063403f
C15864 VDD.t3141 VSS 0.126024f
C15865 VDD.t3133 VSS 0.075145f
C15866 VDD.t4460 VSS 0.075145f
C15867 VDD.t4395 VSS 0.041877f
C15868 VDD.n488 VSS 0.064693f
C15869 VDD.n489 VSS 0.076519f
C15870 VDD.t198 VSS 0.007233f
C15871 VDD.t4396 VSS 0.007233f
C15872 VDD.n490 VSS 0.016652f
C15873 VDD.n491 VSS 0.047679f
C15874 VDD.t505 VSS 0.007233f
C15875 VDD.t2051 VSS 0.007233f
C15876 VDD.n492 VSS 0.016652f
C15877 VDD.n493 VSS 0.07634f
C15878 VDD.t503 VSS 0.027188f
C15879 VDD.n494 VSS 0.076455f
C15880 VDD.t3140 VSS 0.027188f
C15881 VDD.n495 VSS 0.076457f
C15882 VDD.t4488 VSS 0.007233f
C15883 VDD.t3138 VSS 0.007233f
C15884 VDD.n496 VSS 0.016652f
C15885 VDD.n497 VSS 0.073375f
C15886 VDD.n498 VSS 0.076519f
C15887 VDD.n499 VSS 0.064809f
C15888 VDD.t3032 VSS 0.063624f
C15889 VDD.t2927 VSS 0.075406f
C15890 VDD.t2646 VSS 0.075406f
C15891 VDD.t148 VSS 0.141386f
C15892 VDD.t3135 VSS 0.141386f
C15893 VDD.t3131 VSS 0.075406f
C15894 VDD.t189 VSS 0.075406f
C15895 VDD.t187 VSS 0.042023f
C15896 VDD.n500 VSS 0.064809f
C15897 VDD.n501 VSS 0.076519f
C15898 VDD.t206 VSS 0.007233f
C15899 VDD.t188 VSS 0.007233f
C15900 VDD.n502 VSS 0.016652f
C15901 VDD.n503 VSS 0.047679f
C15902 VDD.t608 VSS 0.007233f
C15903 VDD.t204 VSS 0.007233f
C15904 VDD.n504 VSS 0.016652f
C15905 VDD.n505 VSS 0.07634f
C15906 VDD.t606 VSS 0.027188f
C15907 VDD.n506 VSS 0.073667f
C15908 VDD.t3130 VSS 0.027188f
C15909 VDD.n507 VSS 0.073669f
C15910 VDD.t194 VSS 0.007233f
C15911 VDD.t3128 VSS 0.007233f
C15912 VDD.n508 VSS 0.016652f
C15913 VDD.n509 VSS 0.073375f
C15914 VDD.n510 VSS 0.076519f
C15915 VDD.n511 VSS 0.064809f
C15916 VDD.t3016 VSS 0.063624f
C15917 VDD.t3028 VSS 0.075406f
C15918 VDD.t1105 VSS 0.075406f
C15919 VDD.t1107 VSS 0.13786f
C15920 VDD.t956 VSS 0.137401f
C15921 VDD.t958 VSS 0.075145f
C15922 VDD.t2549 VSS 0.075145f
C15923 VDD.t2547 VSS 0.041877f
C15924 VDD.n512 VSS 0.064693f
C15925 VDD.n513 VSS 0.076519f
C15926 VDD.t4262 VSS 0.007233f
C15927 VDD.t2548 VSS 0.007233f
C15928 VDD.n514 VSS 0.016652f
C15929 VDD.n515 VSS 0.047679f
C15930 VDD.t513 VSS 0.007233f
C15931 VDD.t4264 VSS 0.007233f
C15932 VDD.n516 VSS 0.016652f
C15933 VDD.n517 VSS 0.07634f
C15934 VDD.t511 VSS 0.027188f
C15935 VDD.n518 VSS 0.110894f
C15936 VDD.t2544 VSS 0.004807f
C15937 VDD.t2546 VSS 0.004807f
C15938 VDD.n519 VSS 0.010736f
C15939 VDD.t2542 VSS 0.017466f
C15940 VDD.n520 VSS 0.056287f
C15941 VDD.n521 VSS 0.020342f
C15942 VDD.n522 VSS 0.030311f
C15943 VDD.t2545 VSS 0.089594f
C15944 VDD.n523 VSS 0.035424f
C15945 VDD.t2543 VSS 0.05332f
C15946 VDD.t2541 VSS 0.027493f
C15947 VDD.n524 VSS 0.067089f
C15948 VDD.n525 VSS 0.044915f
C15949 VDD.t3283 VSS 0.081296f
C15950 VDD.t3284 VSS 0.075406f
C15951 VDD.t3285 VSS 0.075406f
C15952 VDD.t3281 VSS 0.075406f
C15953 VDD.t3282 VSS 0.075406f
C15954 VDD.t4251 VSS 0.075406f
C15955 VDD.t4253 VSS 0.075406f
C15956 VDD.t4257 VSS 0.058518f
C15957 VDD.t4259 VSS 0.126462f
C15958 VDD.t4255 VSS 0.05459f
C15959 VDD.n526 VSS 2.52e-19
C15960 VDD.t4252 VSS 0.00575f
C15961 VDD.t4254 VSS 0.00575f
C15962 VDD.n527 VSS 0.0115f
C15963 VDD.n528 VSS 0.012479f
C15964 VDD.t4258 VSS 0.00575f
C15965 VDD.t4256 VSS 0.00575f
C15966 VDD.n529 VSS 0.0115f
C15967 VDD.n530 VSS 0.007448f
C15968 VDD.n531 VSS 0.076419f
C15969 VDD.t4260 VSS 0.01978f
C15970 VDD.n532 VSS 0.014195f
C15971 VDD.n533 VSS -0.011842f
C15972 VDD.n534 VSS 0.077508f
C15973 VDD.n535 VSS 0.836811f
C15974 VDD.n536 VSS 1.33083f
C15975 VDD.n537 VSS 1.22885f
C15976 VDD.n538 VSS 1.34428f
C15977 VDD.t233 VSS 0.027215f
C15978 VDD.t2699 VSS 0.007233f
C15979 VDD.t235 VSS 0.007233f
C15980 VDD.n539 VSS 0.016652f
C15981 VDD.n540 VSS 0.129639f
C15982 VDD.t1153 VSS -0.019301f
C15983 VDD.t1155 VSS 0.075145f
C15984 VDD.t4247 VSS 0.075145f
C15985 VDD.t4245 VSS 0.063403f
C15986 VDD.t3957 VSS 0.027215f
C15987 VDD.t3955 VSS 0.007233f
C15988 VDD.t3090 VSS 0.007233f
C15989 VDD.n541 VSS 0.016652f
C15990 VDD.n542 VSS 0.132756f
C15991 VDD.t3075 VSS 0.007233f
C15992 VDD.t3630 VSS 0.007233f
C15993 VDD.n543 VSS 0.016652f
C15994 VDD.n544 VSS 0.047679f
C15995 VDD.t3628 VSS 0.007233f
C15996 VDD.t3812 VSS 0.007233f
C15997 VDD.n545 VSS 0.016652f
C15998 VDD.n546 VSS 0.073624f
C15999 VDD.t3629 VSS 0.04195f
C16000 VDD.t3633 VSS 0.075275f
C16001 VDD.t3842 VSS 0.075275f
C16002 VDD.t3856 VSS 0.139181f
C16003 VDD.t4130 VSS 0.139181f
C16004 VDD.t4132 VSS 0.075275f
C16005 VDD.t1992 VSS 0.075275f
C16006 VDD.t1996 VSS 0.063514f
C16007 VDD.t3826 VSS 0.027188f
C16008 VDD.n547 VSS 0.07466f
C16009 VDD.t175 VSS 0.027188f
C16010 VDD.n548 VSS 0.074656f
C16011 VDD.t177 VSS 0.007233f
C16012 VDD.t3100 VSS 0.007233f
C16013 VDD.n549 VSS 0.016652f
C16014 VDD.n550 VSS 0.076601f
C16015 VDD.t3025 VSS 0.007233f
C16016 VDD.t4430 VSS 0.007233f
C16017 VDD.n551 VSS 0.016652f
C16018 VDD.n552 VSS 0.047822f
C16019 VDD.t3703 VSS 0.027215f
C16020 VDD.t4466 VSS 0.007233f
C16021 VDD.t3818 VSS 0.007233f
C16022 VDD.n553 VSS 0.016652f
C16023 VDD.n554 VSS 0.130541f
C16024 VDD.t4429 VSS 0.04195f
C16025 VDD.t4495 VSS 0.075275f
C16026 VDD.t3854 VSS 0.075275f
C16027 VDD.t3868 VSS 0.145846f
C16028 VDD.t1486 VSS 0.145846f
C16029 VDD.t1488 VSS 0.075275f
C16030 VDD.t1984 VSS 0.075275f
C16031 VDD.t1986 VSS 0.063514f
C16032 VDD.t3702 VSS 0.126243f
C16033 VDD.t3817 VSS 0.075275f
C16034 VDD.t4465 VSS 0.075275f
C16035 VDD.t4401 VSS 0.04195f
C16036 VDD.n555 VSS 0.064751f
C16037 VDD.n556 VSS 0.07665f
C16038 VDD.t1987 VSS 0.007233f
C16039 VDD.t4402 VSS 0.007233f
C16040 VDD.n557 VSS 0.016652f
C16041 VDD.n558 VSS 0.047822f
C16042 VDD.t1489 VSS 0.007233f
C16043 VDD.t1985 VSS 0.007233f
C16044 VDD.n559 VSS 0.016652f
C16045 VDD.n560 VSS 0.076601f
C16046 VDD.t1487 VSS 0.027188f
C16047 VDD.n561 VSS 0.076624f
C16048 VDD.t3869 VSS 0.027188f
C16049 VDD.n562 VSS 0.076629f
C16050 VDD.t4496 VSS 0.007233f
C16051 VDD.t3855 VSS 0.007233f
C16052 VDD.n563 VSS 0.016652f
C16053 VDD.n564 VSS 0.073624f
C16054 VDD.n565 VSS 0.07665f
C16055 VDD.n566 VSS 0.064751f
C16056 VDD.t3024 VSS 0.063514f
C16057 VDD.t3099 VSS 0.075275f
C16058 VDD.t176 VSS 0.075275f
C16059 VDD.t174 VSS 0.141141f
C16060 VDD.t3825 VSS 0.141141f
C16061 VDD.t3811 VSS 0.075275f
C16062 VDD.t3627 VSS 0.075275f
C16063 VDD.t3625 VSS 0.04195f
C16064 VDD.n567 VSS 0.064751f
C16065 VDD.n568 VSS 0.07665f
C16066 VDD.t1997 VSS 0.007233f
C16067 VDD.t3626 VSS 0.007233f
C16068 VDD.n569 VSS 0.016652f
C16069 VDD.n570 VSS 0.047822f
C16070 VDD.t4133 VSS 0.007233f
C16071 VDD.t1993 VSS 0.007233f
C16072 VDD.n571 VSS 0.016652f
C16073 VDD.n572 VSS 0.076601f
C16074 VDD.t4131 VSS 0.027188f
C16075 VDD.n573 VSS 0.073849f
C16076 VDD.t3857 VSS 0.027188f
C16077 VDD.n574 VSS 0.073656f
C16078 VDD.t3634 VSS 0.007233f
C16079 VDD.t3843 VSS 0.007233f
C16080 VDD.n575 VSS 0.016652f
C16081 VDD.n576 VSS 0.073375f
C16082 VDD.n577 VSS 0.076519f
C16083 VDD.n578 VSS 0.064751f
C16084 VDD.t3074 VSS 0.063514f
C16085 VDD.t3089 VSS 0.075275f
C16086 VDD.t3954 VSS 0.075275f
C16087 VDD.t3956 VSS 0.137602f
C16088 VDD.t232 VSS 0.137365f
C16089 VDD.t234 VSS 0.075145f
C16090 VDD.t2698 VSS 0.075145f
C16091 VDD.t2696 VSS 0.041877f
C16092 VDD.n579 VSS 0.064693f
C16093 VDD.n580 VSS 0.076519f
C16094 VDD.t4246 VSS 0.007233f
C16095 VDD.t2697 VSS 0.007233f
C16096 VDD.n581 VSS 0.016652f
C16097 VDD.n582 VSS 0.047679f
C16098 VDD.t1156 VSS 0.007233f
C16099 VDD.t4248 VSS 0.007233f
C16100 VDD.n583 VSS 0.016652f
C16101 VDD.n584 VSS 0.07634f
C16102 VDD.t1154 VSS 0.027188f
C16103 VDD.n585 VSS 0.256185f
C16104 VDD.n586 VSS 1.58047f
C16105 VDD.t3414 VSS 0.027215f
C16106 VDD.t3578 VSS 0.007233f
C16107 VDD.t3416 VSS 0.007233f
C16108 VDD.n587 VSS 0.016652f
C16109 VDD.n588 VSS 0.129639f
C16110 VDD.t1211 VSS -0.019301f
C16111 VDD.t1213 VSS 0.075145f
C16112 VDD.t1421 VSS 0.075145f
C16113 VDD.t1423 VSS 0.063403f
C16114 VDD.t1367 VSS 0.027215f
C16115 VDD.t1365 VSS 0.007233f
C16116 VDD.t3084 VSS 0.007233f
C16117 VDD.n589 VSS 0.016652f
C16118 VDD.n590 VSS 0.132428f
C16119 VDD.t3068 VSS 0.007233f
C16120 VDD.t3632 VSS 0.007233f
C16121 VDD.n591 VSS 0.016652f
C16122 VDD.n592 VSS 0.047679f
C16123 VDD.t3624 VSS 0.007233f
C16124 VDD.t1369 VSS 0.007233f
C16125 VDD.n593 VSS 0.016652f
C16126 VDD.n594 VSS 0.073375f
C16127 VDD.t3631 VSS 0.041877f
C16128 VDD.t3635 VSS 0.075145f
C16129 VDD.t1380 VSS 0.075145f
C16130 VDD.t1382 VSS 0.138939f
C16131 VDD.t3347 VSS 0.138939f
C16132 VDD.t3349 VSS 0.075145f
C16133 VDD.t1988 VSS 0.075145f
C16134 VDD.t1990 VSS 0.063403f
C16135 VDD.t1373 VSS 0.027188f
C16136 VDD.n595 VSS 0.074488f
C16137 VDD.t2042 VSS 0.027188f
C16138 VDD.n596 VSS 0.074487f
C16139 VDD.t2044 VSS 0.007233f
C16140 VDD.t2987 VSS 0.007233f
C16141 VDD.n597 VSS 0.016652f
C16142 VDD.n598 VSS 0.07634f
C16143 VDD.t3088 VSS 0.007233f
C16144 VDD.t4365 VSS 0.007233f
C16145 VDD.n599 VSS 0.016652f
C16146 VDD.n600 VSS 0.047679f
C16147 VDD.t3003 VSS 0.004807f
C16148 VDD.t2938 VSS 0.004807f
C16149 VDD.n601 VSS 0.010736f
C16150 VDD.t3061 VSS 0.017466f
C16151 VDD.n602 VSS 0.048701f
C16152 VDD.n603 VSS 0.030676f
C16153 VDD.t4355 VSS 0.145552f
C16154 VDD.t4356 VSS 0.004807f
C16155 VDD.t4438 VSS 0.004807f
C16156 VDD.n604 VSS 0.010736f
C16157 VDD.t4481 VSS 0.017466f
C16158 VDD.n605 VSS 0.048701f
C16159 VDD.t3723 VSS 0.004807f
C16160 VDD.t3769 VSS 0.004807f
C16161 VDD.n606 VSS 0.010736f
C16162 VDD.t3831 VSS 0.017466f
C16163 VDD.n607 VSS 0.059157f
C16164 VDD.t3722 VSS 0.137944f
C16165 VDD.n608 VSS 0.135842f
C16166 VDD.n609 VSS 0.031797f
C16167 VDD.n610 VSS 0.030676f
C16168 VDD.n611 VSS 0.028952f
C16169 VDD.n612 VSS 0.135842f
C16170 VDD.t2937 VSS 0.270495f
C16171 VDD.n613 VSS 0.096866f
C16172 VDD.t1379 VSS 0.027204f
C16173 VDD.n614 VSS 0.169958f
C16174 VDD.t4418 VSS 0.007233f
C16175 VDD.t1371 VSS 0.007233f
C16176 VDD.n615 VSS 0.016652f
C16177 VDD.n616 VSS 0.050644f
C16178 VDD.t4364 VSS 0.041877f
C16179 VDD.t4439 VSS 0.075145f
C16180 VDD.t1374 VSS 0.075145f
C16181 VDD.t1376 VSS 0.145593f
C16182 VDD.t872 VSS 0.145593f
C16183 VDD.t874 VSS 0.075145f
C16184 VDD.t1994 VSS 0.075145f
C16185 VDD.t1721 VSS 0.063403f
C16186 VDD.t1378 VSS 0.126024f
C16187 VDD.t1370 VSS 0.075145f
C16188 VDD.t4417 VSS 0.075145f
C16189 VDD.t4510 VSS 0.041877f
C16190 VDD.n617 VSS 0.064693f
C16191 VDD.n618 VSS 0.076519f
C16192 VDD.t1722 VSS 0.007233f
C16193 VDD.t4511 VSS 0.007233f
C16194 VDD.n619 VSS 0.016652f
C16195 VDD.n620 VSS 0.047679f
C16196 VDD.t875 VSS 0.007233f
C16197 VDD.t1995 VSS 0.007233f
C16198 VDD.n621 VSS 0.016652f
C16199 VDD.n622 VSS 0.07634f
C16200 VDD.t873 VSS 0.027188f
C16201 VDD.n623 VSS 0.076455f
C16202 VDD.t1377 VSS 0.027188f
C16203 VDD.n624 VSS 0.076457f
C16204 VDD.t4440 VSS 0.007233f
C16205 VDD.t1375 VSS 0.007233f
C16206 VDD.n625 VSS 0.016652f
C16207 VDD.n626 VSS 0.073375f
C16208 VDD.n627 VSS 0.076519f
C16209 VDD.n628 VSS 0.064693f
C16210 VDD.t3087 VSS 0.063403f
C16211 VDD.t2986 VSS 0.075145f
C16212 VDD.t2043 VSS 0.075145f
C16213 VDD.t2041 VSS 0.140896f
C16214 VDD.t1372 VSS 0.140896f
C16215 VDD.t1368 VSS 0.075145f
C16216 VDD.t3623 VSS 0.075149f
C16217 VDD.t3637 VSS 0.041944f
C16218 VDD.n629 VSS 0.064693f
C16219 VDD.n630 VSS 0.076519f
C16220 VDD.t1991 VSS 0.007233f
C16221 VDD.t3638 VSS 0.007233f
C16222 VDD.n631 VSS 0.016652f
C16223 VDD.n632 VSS 0.047679f
C16224 VDD.t3350 VSS 0.007233f
C16225 VDD.t1989 VSS 0.007233f
C16226 VDD.n633 VSS 0.016652f
C16227 VDD.n634 VSS 0.07634f
C16228 VDD.t3348 VSS 0.027188f
C16229 VDD.n635 VSS 0.073667f
C16230 VDD.t1383 VSS 0.027188f
C16231 VDD.n636 VSS 0.073669f
C16232 VDD.t3636 VSS 0.007233f
C16233 VDD.t1381 VSS 0.007233f
C16234 VDD.n637 VSS 0.016652f
C16235 VDD.n638 VSS 0.073375f
C16236 VDD.n639 VSS 0.076519f
C16237 VDD.n640 VSS 0.064693f
C16238 VDD.t3067 VSS 0.063403f
C16239 VDD.t3083 VSS 0.075145f
C16240 VDD.t1364 VSS 0.075145f
C16241 VDD.t1366 VSS 0.137373f
C16242 VDD.t3413 VSS 0.137373f
C16243 VDD.t3415 VSS 0.075145f
C16244 VDD.t3577 VSS 0.075145f
C16245 VDD.t3575 VSS 0.041877f
C16246 VDD.n641 VSS 0.064693f
C16247 VDD.n642 VSS 0.076519f
C16248 VDD.t1424 VSS 0.007233f
C16249 VDD.t3576 VSS 0.007233f
C16250 VDD.n643 VSS 0.016652f
C16251 VDD.n644 VSS 0.047679f
C16252 VDD.t1214 VSS 0.007233f
C16253 VDD.t1422 VSS 0.007233f
C16254 VDD.n645 VSS 0.016652f
C16255 VDD.n646 VSS 0.07634f
C16256 VDD.t1212 VSS 0.027188f
C16257 VDD.n647 VSS 0.110894f
C16258 VDD.t3346 VSS 0.004807f
C16259 VDD.t1317 VSS 0.004807f
C16260 VDD.n648 VSS 0.010736f
C16261 VDD.t3344 VSS 0.017466f
C16262 VDD.n649 VSS 0.056287f
C16263 VDD.n650 VSS 0.020342f
C16264 VDD.n651 VSS 0.030311f
C16265 VDD.t1316 VSS 0.089594f
C16266 VDD.n652 VSS 0.035424f
C16267 VDD.t3345 VSS 0.05332f
C16268 VDD.t3343 VSS 0.027493f
C16269 VDD.n653 VSS 0.067089f
C16270 VDD.n654 VSS 0.044915f
C16271 VDD.t690 VSS 0.081296f
C16272 VDD.t686 VSS 0.075406f
C16273 VDD.t687 VSS 0.075406f
C16274 VDD.t688 VSS 0.075406f
C16275 VDD.t689 VSS 0.075406f
C16276 VDD.t4305 VSS 0.075406f
C16277 VDD.t4297 VSS 0.075406f
C16278 VDD.t4301 VSS 0.058518f
C16279 VDD.t4303 VSS 0.126462f
C16280 VDD.t4299 VSS 0.05459f
C16281 VDD.n655 VSS 2.52e-19
C16282 VDD.t4306 VSS 0.00575f
C16283 VDD.t4298 VSS 0.00575f
C16284 VDD.n656 VSS 0.0115f
C16285 VDD.n657 VSS 0.012479f
C16286 VDD.t4302 VSS 0.00575f
C16287 VDD.t4300 VSS 0.00575f
C16288 VDD.n658 VSS 0.0115f
C16289 VDD.n659 VSS 0.007448f
C16290 VDD.n660 VSS 0.076419f
C16291 VDD.t4304 VSS 0.01978f
C16292 VDD.n661 VSS 0.014195f
C16293 VDD.n662 VSS -0.011842f
C16294 VDD.n663 VSS 0.077508f
C16295 VDD.n664 VSS 0.836811f
C16296 VDD.n665 VSS 1.3558f
C16297 VDD.n666 VSS 1.17167f
C16298 VDD.n667 VSS 0.059843f
C16299 VDD.t2732 VSS 0.085532f
C16300 VDD.t2004 VSS 0.019227f
C16301 VDD.t2002 VSS 0.019227f
C16302 VDD.n668 VSS 0.05532f
C16303 VDD.t2420 VSS 0.019227f
C16304 VDD.t2419 VSS 0.019227f
C16305 VDD.n669 VSS 0.055358f
C16306 VDD.t2422 VSS 0.085532f
C16307 VDD.n670 VSS 0.178951f
C16308 VDD.n671 VSS 0.108238f
C16309 VDD.t2391 VSS 0.043813f
C16310 VDD.t1461 VSS 0.004807f
C16311 VDD.t1463 VSS 0.004807f
C16312 VDD.n672 VSS 0.010736f
C16313 VDD.t1476 VSS 0.017466f
C16314 VDD.n673 VSS 0.048701f
C16315 VDD.t2389 VSS 0.056456f
C16316 VDD.t2387 VSS 0.061455f
C16317 VDD.t1462 VSS 0.00642f
C16318 VDD.t1460 VSS 0.054398f
C16319 VDD.n674 VSS 0.062239f
C16320 VDD.t1475 VSS 0.086009f
C16321 VDD.n675 VSS 0.063841f
C16322 VDD.t2388 VSS 0.017454f
C16323 VDD.n676 VSS 0.060949f
C16324 VDD.t2390 VSS 0.004807f
C16325 VDD.t2392 VSS 0.004807f
C16326 VDD.n677 VSS 0.010696f
C16327 VDD.n678 VSS 0.052319f
C16328 VDD.t2424 VSS 0.017474f
C16329 VDD.t196 VSS 0.004807f
C16330 VDD.t1821 VSS 0.004807f
C16331 VDD.n679 VSS 0.010696f
C16332 VDD.n680 VSS 0.096107f
C16333 VDD.n681 VSS 0.095147f
C16334 VDD.n682 VSS 0.013667f
C16335 VDD.n683 VSS 7.86e-19
C16336 VDD.t195 VSS 0.040872f
C16337 VDD.t1820 VSS 0.056456f
C16338 VDD.t2423 VSS 0.151258f
C16339 VDD.t560 VSS 0.517243f
C16340 VDD.t561 VSS 0.254838f
C16341 VDD.t562 VSS 0.254838f
C16342 VDD.t3167 VSS 0.254838f
C16343 VDD.t3168 VSS 0.254838f
C16344 VDD.t3169 VSS 0.254838f
C16345 VDD.t1529 VSS 0.254838f
C16346 VDD.t1530 VSS 0.254838f
C16347 VDD.t1528 VSS 0.254838f
C16348 VDD.t2003 VSS 0.254838f
C16349 VDD.t2001 VSS 0.254838f
C16350 VDD.t2421 VSS 0.292552f
C16351 VDD.n684 VSS 0.569521f
C16352 VDD.n685 VSS 0.271667f
C16353 VDD.n686 VSS 0.167926f
C16354 VDD.n687 VSS 0.486632f
C16355 VDD.n688 VSS 0.72887f
C16356 VDD.n689 VSS 1.11637f
C16357 VDD.t4168 VSS 0.027215f
C16358 VDD.t1871 VSS 0.007233f
C16359 VDD.t4170 VSS 0.007233f
C16360 VDD.n690 VSS 0.016652f
C16361 VDD.n691 VSS 0.129639f
C16362 VDD.t4020 VSS -0.019301f
C16363 VDD.t4022 VSS 0.075145f
C16364 VDD.t230 VSS 0.075145f
C16365 VDD.t228 VSS 0.063403f
C16366 VDD.t3574 VSS 0.027215f
C16367 VDD.t3572 VSS 0.007233f
C16368 VDD.t3092 VSS 0.007233f
C16369 VDD.n692 VSS 0.016652f
C16370 VDD.n693 VSS 0.132756f
C16371 VDD.t3081 VSS 0.007233f
C16372 VDD.t3255 VSS 0.007233f
C16373 VDD.n694 VSS 0.016652f
C16374 VDD.n695 VSS 0.047679f
C16375 VDD.t3253 VSS 0.007233f
C16376 VDD.t3808 VSS 0.007233f
C16377 VDD.n696 VSS 0.016652f
C16378 VDD.n697 VSS 0.073624f
C16379 VDD.t3254 VSS 0.04195f
C16380 VDD.t3256 VSS 0.075275f
C16381 VDD.t3838 VSS 0.075275f
C16382 VDD.t3848 VSS 0.139181f
C16383 VDD.t43 VSS 0.139181f
C16384 VDD.t45 VSS 0.075275f
C16385 VDD.t3369 VSS 0.075275f
C16386 VDD.t3373 VSS 0.063514f
C16387 VDD.t3824 VSS 0.027188f
C16388 VDD.n698 VSS 0.07466f
C16389 VDD.t1621 VSS 0.027188f
C16390 VDD.n699 VSS 0.074656f
C16391 VDD.t1623 VSS 0.007233f
C16392 VDD.t2926 VSS 0.007233f
C16393 VDD.n700 VSS 0.016652f
C16394 VDD.n701 VSS 0.076601f
C16395 VDD.t3031 VSS 0.007233f
C16396 VDD.t4428 VSS 0.007233f
C16397 VDD.n702 VSS 0.016652f
C16398 VDD.n703 VSS 0.047822f
C16399 VDD.t3701 VSS 0.027215f
C16400 VDD.t4464 VSS 0.007233f
C16401 VDD.t3814 VSS 0.007233f
C16402 VDD.n704 VSS 0.016652f
C16403 VDD.n705 VSS 0.130541f
C16404 VDD.t4427 VSS 0.04195f
C16405 VDD.t4491 VSS 0.075275f
C16406 VDD.t3846 VSS 0.075275f
C16407 VDD.t3866 VSS 0.145846f
C16408 VDD.t1864 VSS 0.145846f
C16409 VDD.t1866 VSS 0.075275f
C16410 VDD.t3361 VSS 0.075275f
C16411 VDD.t3365 VSS 0.063514f
C16412 VDD.t3700 VSS 0.126243f
C16413 VDD.t3813 VSS 0.075275f
C16414 VDD.t4463 VSS 0.075275f
C16415 VDD.t4399 VSS 0.04195f
C16416 VDD.n706 VSS 0.064751f
C16417 VDD.n707 VSS 0.07665f
C16418 VDD.t3366 VSS 0.007233f
C16419 VDD.t4400 VSS 0.007233f
C16420 VDD.n708 VSS 0.016652f
C16421 VDD.n709 VSS 0.047822f
C16422 VDD.t1867 VSS 0.007233f
C16423 VDD.t3362 VSS 0.007233f
C16424 VDD.n710 VSS 0.016652f
C16425 VDD.n711 VSS 0.076601f
C16426 VDD.t1865 VSS 0.027188f
C16427 VDD.n712 VSS 0.076624f
C16428 VDD.t3867 VSS 0.027188f
C16429 VDD.n713 VSS 0.076629f
C16430 VDD.t4492 VSS 0.007233f
C16431 VDD.t3847 VSS 0.007233f
C16432 VDD.n714 VSS 0.016652f
C16433 VDD.n715 VSS 0.073624f
C16434 VDD.n716 VSS 0.07665f
C16435 VDD.n717 VSS 0.064751f
C16436 VDD.t3030 VSS 0.063514f
C16437 VDD.t2925 VSS 0.075275f
C16438 VDD.t1622 VSS 0.075275f
C16439 VDD.t1620 VSS 0.141141f
C16440 VDD.t3823 VSS 0.141141f
C16441 VDD.t3807 VSS 0.075275f
C16442 VDD.t3252 VSS 0.075275f
C16443 VDD.t3248 VSS 0.04195f
C16444 VDD.n718 VSS 0.064751f
C16445 VDD.n719 VSS 0.07665f
C16446 VDD.t3374 VSS 0.007233f
C16447 VDD.t3249 VSS 0.007233f
C16448 VDD.n720 VSS 0.016652f
C16449 VDD.n721 VSS 0.047822f
C16450 VDD.t46 VSS 0.007233f
C16451 VDD.t3370 VSS 0.007233f
C16452 VDD.n722 VSS 0.016652f
C16453 VDD.n723 VSS 0.076601f
C16454 VDD.t44 VSS 0.027188f
C16455 VDD.n724 VSS 0.073849f
C16456 VDD.t3849 VSS 0.027188f
C16457 VDD.n725 VSS 0.073656f
C16458 VDD.t3257 VSS 0.007233f
C16459 VDD.t3839 VSS 0.007233f
C16460 VDD.n726 VSS 0.016652f
C16461 VDD.n727 VSS 0.073375f
C16462 VDD.n728 VSS 0.076519f
C16463 VDD.n729 VSS 0.064751f
C16464 VDD.t3080 VSS 0.063514f
C16465 VDD.t3091 VSS 0.075275f
C16466 VDD.t3571 VSS 0.075275f
C16467 VDD.t3573 VSS 0.137602f
C16468 VDD.t4167 VSS 0.137365f
C16469 VDD.t4169 VSS 0.075145f
C16470 VDD.t1870 VSS 0.075145f
C16471 VDD.t1868 VSS 0.041877f
C16472 VDD.n730 VSS 0.064693f
C16473 VDD.n731 VSS 0.076519f
C16474 VDD.t229 VSS 0.007233f
C16475 VDD.t1869 VSS 0.007233f
C16476 VDD.n732 VSS 0.016652f
C16477 VDD.n733 VSS 0.047679f
C16478 VDD.t4023 VSS 0.007233f
C16479 VDD.t231 VSS 0.007233f
C16480 VDD.n734 VSS 0.016652f
C16481 VDD.n735 VSS 0.07634f
C16482 VDD.t4021 VSS 0.027188f
C16483 VDD.n736 VSS 0.256185f
C16484 VDD.n737 VSS 1.58763f
C16485 VDD.t796 VSS 0.027215f
C16486 VDD.t1891 VSS 0.007233f
C16487 VDD.t2486 VSS 0.007233f
C16488 VDD.n738 VSS 0.016652f
C16489 VDD.n739 VSS 0.129639f
C16490 VDD.t2786 VSS -0.019301f
C16491 VDD.t2788 VSS 0.075145f
C16492 VDD.t818 VSS 0.075145f
C16493 VDD.t820 VSS 0.063403f
C16494 VDD.t17 VSS 0.027215f
C16495 VDD.t15 VSS 0.007233f
C16496 VDD.t3035 VSS 0.007233f
C16497 VDD.n740 VSS 0.016652f
C16498 VDD.n741 VSS 0.132428f
C16499 VDD.t3019 VSS 0.007233f
C16500 VDD.t3259 VSS 0.007233f
C16501 VDD.n742 VSS 0.016652f
C16502 VDD.n743 VSS 0.047679f
C16503 VDD.t3251 VSS 0.007233f
C16504 VDD.t124 VSS 0.007233f
C16505 VDD.n744 VSS 0.016652f
C16506 VDD.n745 VSS 0.073375f
C16507 VDD.t3258 VSS 0.042023f
C16508 VDD.t3260 VSS 0.075406f
C16509 VDD.t119 VSS 0.075406f
C16510 VDD.t121 VSS 0.139422f
C16511 VDD.t239 VSS 0.139422f
C16512 VDD.t241 VSS 0.075406f
C16513 VDD.t3367 VSS 0.075406f
C16514 VDD.t3371 VSS 0.063624f
C16515 VDD.t128 VSS 0.027188f
C16516 VDD.n746 VSS 0.074488f
C16517 VDD.t410 VSS 0.027188f
C16518 VDD.n747 VSS 0.074487f
C16519 VDD.t412 VSS 0.007233f
C16520 VDD.t2930 VSS 0.007233f
C16521 VDD.n748 VSS 0.016652f
C16522 VDD.n749 VSS 0.07634f
C16523 VDD.t3037 VSS 0.007233f
C16524 VDD.t4423 VSS 0.007233f
C16525 VDD.n750 VSS 0.016652f
C16526 VDD.n751 VSS 0.047679f
C16527 VDD.t3093 VSS 0.004807f
C16528 VDD.t3027 VSS 0.004807f
C16529 VDD.n752 VSS 0.010736f
C16530 VDD.t3094 VSS 0.017466f
C16531 VDD.n753 VSS 0.048701f
C16532 VDD.n754 VSS 0.030676f
C16533 VDD.t4448 VSS 0.145552f
C16534 VDD.t4456 VSS 0.004807f
C16535 VDD.t4505 VSS 0.004807f
C16536 VDD.n755 VSS 0.010736f
C16537 VDD.t4449 VSS 0.017466f
C16538 VDD.n756 VSS 0.048701f
C16539 VDD.t3798 VSS 0.004807f
C16540 VDD.t3876 VSS 0.004807f
C16541 VDD.n757 VSS 0.010736f
C16542 VDD.t3792 VSS 0.017466f
C16543 VDD.n758 VSS 0.059157f
C16544 VDD.t3791 VSS 0.137944f
C16545 VDD.n759 VSS 0.135842f
C16546 VDD.n760 VSS 0.031797f
C16547 VDD.n761 VSS 0.030676f
C16548 VDD.n762 VSS 0.028952f
C16549 VDD.n763 VSS 0.135842f
C16550 VDD.t3026 VSS 0.270495f
C16551 VDD.n764 VSS 0.096866f
C16552 VDD.t134 VSS 0.027204f
C16553 VDD.n765 VSS 0.169958f
C16554 VDD.t4459 VSS 0.007233f
C16555 VDD.t126 VSS 0.007233f
C16556 VDD.n766 VSS 0.016652f
C16557 VDD.n767 VSS 0.050644f
C16558 VDD.t4422 VSS 0.042023f
C16559 VDD.t4485 VSS 0.075406f
C16560 VDD.t129 VSS 0.075406f
C16561 VDD.t131 VSS 0.144962f
C16562 VDD.t2792 VSS 0.14709f
C16563 VDD.t2794 VSS 0.075145f
C16564 VDD.t3359 VSS 0.075145f
C16565 VDD.t3363 VSS 0.063403f
C16566 VDD.t133 VSS 0.126024f
C16567 VDD.t125 VSS 0.075145f
C16568 VDD.t4458 VSS 0.075145f
C16569 VDD.t4391 VSS 0.041877f
C16570 VDD.n768 VSS 0.064693f
C16571 VDD.n769 VSS 0.076519f
C16572 VDD.t3364 VSS 0.007233f
C16573 VDD.t4392 VSS 0.007233f
C16574 VDD.n770 VSS 0.016652f
C16575 VDD.n771 VSS 0.047679f
C16576 VDD.t2795 VSS 0.007233f
C16577 VDD.t3360 VSS 0.007233f
C16578 VDD.n772 VSS 0.016652f
C16579 VDD.n773 VSS 0.07634f
C16580 VDD.t2793 VSS 0.027188f
C16581 VDD.n774 VSS 0.076455f
C16582 VDD.t132 VSS 0.027188f
C16583 VDD.n775 VSS 0.076457f
C16584 VDD.t4486 VSS 0.007233f
C16585 VDD.t130 VSS 0.007233f
C16586 VDD.n776 VSS 0.016652f
C16587 VDD.n777 VSS 0.073375f
C16588 VDD.n778 VSS 0.076519f
C16589 VDD.n779 VSS 0.064809f
C16590 VDD.t3036 VSS 0.063624f
C16591 VDD.t2929 VSS 0.075406f
C16592 VDD.t411 VSS 0.075406f
C16593 VDD.t409 VSS 0.141386f
C16594 VDD.t127 VSS 0.141386f
C16595 VDD.t123 VSS 0.075406f
C16596 VDD.t3250 VSS 0.075406f
C16597 VDD.t3246 VSS 0.042023f
C16598 VDD.n780 VSS 0.064809f
C16599 VDD.n781 VSS 0.076519f
C16600 VDD.t3372 VSS 0.007233f
C16601 VDD.t3247 VSS 0.007233f
C16602 VDD.n782 VSS 0.016652f
C16603 VDD.n783 VSS 0.047679f
C16604 VDD.t242 VSS 0.007233f
C16605 VDD.t3368 VSS 0.007233f
C16606 VDD.n784 VSS 0.016652f
C16607 VDD.n785 VSS 0.07634f
C16608 VDD.t240 VSS 0.027188f
C16609 VDD.n786 VSS 0.073667f
C16610 VDD.t122 VSS 0.027188f
C16611 VDD.n787 VSS 0.073669f
C16612 VDD.t3261 VSS 0.007233f
C16613 VDD.t120 VSS 0.007233f
C16614 VDD.n788 VSS 0.016652f
C16615 VDD.n789 VSS 0.073375f
C16616 VDD.n790 VSS 0.076519f
C16617 VDD.n791 VSS 0.064809f
C16618 VDD.t3018 VSS 0.063624f
C16619 VDD.t3034 VSS 0.075406f
C16620 VDD.t14 VSS 0.075406f
C16621 VDD.t16 VSS 0.13786f
C16622 VDD.t795 VSS 0.137401f
C16623 VDD.t2485 VSS 0.075145f
C16624 VDD.t1890 VSS 0.075145f
C16625 VDD.t1888 VSS 0.041877f
C16626 VDD.n792 VSS 0.064693f
C16627 VDD.n793 VSS 0.076519f
C16628 VDD.t821 VSS 0.007233f
C16629 VDD.t1889 VSS 0.007233f
C16630 VDD.n794 VSS 0.016652f
C16631 VDD.n795 VSS 0.047679f
C16632 VDD.t2789 VSS 0.007233f
C16633 VDD.t819 VSS 0.007233f
C16634 VDD.n796 VSS 0.016652f
C16635 VDD.n797 VSS 0.07634f
C16636 VDD.t2787 VSS 0.027188f
C16637 VDD.n798 VSS 0.110894f
C16638 VDD.t3461 VSS 0.004807f
C16639 VDD.t3457 VSS 0.004807f
C16640 VDD.n799 VSS 0.010736f
C16641 VDD.t3459 VSS 0.017466f
C16642 VDD.n800 VSS 0.056287f
C16643 VDD.n801 VSS 0.020342f
C16644 VDD.n802 VSS 0.030311f
C16645 VDD.t3456 VSS 0.089594f
C16646 VDD.n803 VSS 0.035424f
C16647 VDD.t3460 VSS 0.05332f
C16648 VDD.t3458 VSS 0.027493f
C16649 VDD.n804 VSS 0.067089f
C16650 VDD.n805 VSS 0.044915f
C16651 VDD.t962 VSS 0.081296f
C16652 VDD.t963 VSS 0.075406f
C16653 VDD.t964 VSS 0.075406f
C16654 VDD.t960 VSS 0.075406f
C16655 VDD.t961 VSS 0.075406f
C16656 VDD.t1477 VSS 0.075406f
C16657 VDD.t1479 VSS 0.075406f
C16658 VDD.t1226 VSS 0.058518f
C16659 VDD.t1228 VSS 0.126462f
C16660 VDD.t1481 VSS 0.05459f
C16661 VDD.n806 VSS 2.52e-19
C16662 VDD.t1478 VSS 0.00575f
C16663 VDD.t1480 VSS 0.00575f
C16664 VDD.n807 VSS 0.0115f
C16665 VDD.n808 VSS 0.012479f
C16666 VDD.t1227 VSS 0.00575f
C16667 VDD.t1482 VSS 0.00575f
C16668 VDD.n809 VSS 0.0115f
C16669 VDD.n810 VSS 0.007448f
C16670 VDD.n811 VSS 0.076419f
C16671 VDD.t1229 VSS 0.01978f
C16672 VDD.n812 VSS 0.014195f
C16673 VDD.n813 VSS -0.011842f
C16674 VDD.n814 VSS 0.077508f
C16675 VDD.n815 VSS 0.836811f
C16676 VDD.n816 VSS 1.35111f
C16677 VDD.n817 VSS 1.3368f
C16678 VDD.n818 VSS 1.35832f
C16679 VDD.t3354 VSS 0.027215f
C16680 VDD.t2853 VSS 0.007233f
C16681 VDD.t3352 VSS 0.007233f
C16682 VDD.n819 VSS 0.016652f
C16683 VDD.n820 VSS 0.129639f
C16684 VDD.t921 VSS -0.019301f
C16685 VDD.t923 VSS 0.075145f
C16686 VDD.t1218 VSS 0.075145f
C16687 VDD.t1220 VSS 0.063403f
C16688 VDD.t1726 VSS 0.027215f
C16689 VDD.t1724 VSS 0.007233f
C16690 VDD.t3049 VSS 0.007233f
C16691 VDD.n821 VSS 0.016652f
C16692 VDD.n822 VSS 0.132756f
C16693 VDD.t3041 VSS 0.007233f
C16694 VDD.t2672 VSS 0.007233f
C16695 VDD.n823 VSS 0.016652f
C16696 VDD.n824 VSS 0.047679f
C16697 VDD.t2682 VSS 0.007233f
C16698 VDD.t3739 VSS 0.007233f
C16699 VDD.n825 VSS 0.016652f
C16700 VDD.n826 VSS 0.073624f
C16701 VDD.t2671 VSS 0.04195f
C16702 VDD.t2673 VSS 0.075275f
C16703 VDD.t3706 VSS 0.075275f
C16704 VDD.t3716 VSS 0.139181f
C16705 VDD.t1209 VSS 0.139181f
C16706 VDD.t1207 VSS 0.075275f
C16707 VDD.t2525 VSS 0.075275f
C16708 VDD.t2527 VSS 0.063514f
C16709 VDD.t3743 VSS 0.027188f
C16710 VDD.n827 VSS 0.07466f
C16711 VDD.t1139 VSS 0.027188f
C16712 VDD.n828 VSS 0.074656f
C16713 VDD.t1141 VSS 0.007233f
C16714 VDD.t3005 VSS 0.007233f
C16715 VDD.n829 VSS 0.016652f
C16716 VDD.n830 VSS 0.076601f
C16717 VDD.t2936 VSS 0.007233f
C16718 VDD.t4507 VSS 0.007233f
C16719 VDD.n831 VSS 0.016652f
C16720 VDD.n832 VSS 0.047822f
C16721 VDD.t3776 VSS 0.027215f
C16722 VDD.t4384 VSS 0.007233f
C16723 VDD.t3741 VSS 0.007233f
C16724 VDD.n833 VSS 0.016652f
C16725 VDD.n834 VSS 0.130541f
C16726 VDD.t4506 VSS 0.04195f
C16727 VDD.t4413 VSS 0.075275f
C16728 VDD.t3750 VSS 0.075275f
C16729 VDD.t3755 VSS 0.145846f
C16730 VDD.t3397 VSS 0.145846f
C16731 VDD.t3399 VSS 0.075275f
C16732 VDD.t2533 VSS 0.075275f
C16733 VDD.t2535 VSS 0.063514f
C16734 VDD.t3775 VSS 0.126243f
C16735 VDD.t3740 VSS 0.075275f
C16736 VDD.t4383 VSS 0.075275f
C16737 VDD.t4489 VSS 0.04195f
C16738 VDD.n835 VSS 0.064751f
C16739 VDD.n836 VSS 0.07665f
C16740 VDD.t2536 VSS 0.007233f
C16741 VDD.t4490 VSS 0.007233f
C16742 VDD.n837 VSS 0.016652f
C16743 VDD.n838 VSS 0.047822f
C16744 VDD.t3400 VSS 0.007233f
C16745 VDD.t2534 VSS 0.007233f
C16746 VDD.n839 VSS 0.016652f
C16747 VDD.n840 VSS 0.076601f
C16748 VDD.t3398 VSS 0.027188f
C16749 VDD.n841 VSS 0.076624f
C16750 VDD.t3756 VSS 0.027188f
C16751 VDD.n842 VSS 0.076629f
C16752 VDD.t4414 VSS 0.007233f
C16753 VDD.t3751 VSS 0.007233f
C16754 VDD.n843 VSS 0.016652f
C16755 VDD.n844 VSS 0.073624f
C16756 VDD.n845 VSS 0.07665f
C16757 VDD.n846 VSS 0.064751f
C16758 VDD.t2935 VSS 0.063514f
C16759 VDD.t3004 VSS 0.075275f
C16760 VDD.t1140 VSS 0.075275f
C16761 VDD.t1138 VSS 0.141141f
C16762 VDD.t3742 VSS 0.141141f
C16763 VDD.t3738 VSS 0.075275f
C16764 VDD.t2681 VSS 0.075275f
C16765 VDD.t2679 VSS 0.04195f
C16766 VDD.n847 VSS 0.064751f
C16767 VDD.n848 VSS 0.07665f
C16768 VDD.t2528 VSS 0.007233f
C16769 VDD.t2680 VSS 0.007233f
C16770 VDD.n849 VSS 0.016652f
C16771 VDD.n850 VSS 0.047822f
C16772 VDD.t1208 VSS 0.007233f
C16773 VDD.t2526 VSS 0.007233f
C16774 VDD.n851 VSS 0.016652f
C16775 VDD.n852 VSS 0.076601f
C16776 VDD.t1210 VSS 0.027188f
C16777 VDD.n853 VSS 0.073849f
C16778 VDD.t3717 VSS 0.027188f
C16779 VDD.n854 VSS 0.073656f
C16780 VDD.t2674 VSS 0.007233f
C16781 VDD.t3707 VSS 0.007233f
C16782 VDD.n855 VSS 0.016652f
C16783 VDD.n856 VSS 0.073375f
C16784 VDD.n857 VSS 0.076519f
C16785 VDD.n858 VSS 0.064751f
C16786 VDD.t3040 VSS 0.063514f
C16787 VDD.t3048 VSS 0.075275f
C16788 VDD.t1723 VSS 0.075275f
C16789 VDD.t1725 VSS 0.137602f
C16790 VDD.t3353 VSS 0.137365f
C16791 VDD.t3351 VSS 0.075145f
C16792 VDD.t2852 VSS 0.075145f
C16793 VDD.t2850 VSS 0.041877f
C16794 VDD.n859 VSS 0.064693f
C16795 VDD.n860 VSS 0.076519f
C16796 VDD.t1221 VSS 0.007233f
C16797 VDD.t2851 VSS 0.007233f
C16798 VDD.n861 VSS 0.016652f
C16799 VDD.n862 VSS 0.047679f
C16800 VDD.t924 VSS 0.007233f
C16801 VDD.t1219 VSS 0.007233f
C16802 VDD.n863 VSS 0.016652f
C16803 VDD.n864 VSS 0.07634f
C16804 VDD.t922 VSS 0.027188f
C16805 VDD.n865 VSS 0.256185f
C16806 VDD.n866 VSS 1.52869f
C16807 VDD.t1456 VSS 0.027215f
C16808 VDD.t1194 VSS 0.007233f
C16809 VDD.t1458 VSS 0.007233f
C16810 VDD.n867 VSS 0.016652f
C16811 VDD.n868 VSS 0.129639f
C16812 VDD.t2644 VSS -0.019301f
C16813 VDD.t2642 VSS 0.075145f
C16814 VDD.t3115 VSS 0.075145f
C16815 VDD.t3117 VSS 0.063403f
C16816 VDD.t1647 VSS 0.027215f
C16817 VDD.t1649 VSS 0.007233f
C16818 VDD.t2960 VSS 0.007233f
C16819 VDD.n869 VSS 0.016652f
C16820 VDD.n870 VSS 0.132428f
C16821 VDD.t2946 VSS 0.007233f
C16822 VDD.t2668 VSS 0.007233f
C16823 VDD.n871 VSS 0.016652f
C16824 VDD.n872 VSS 0.047679f
C16825 VDD.t2678 VSS 0.007233f
C16826 VDD.t2797 VSS 0.007233f
C16827 VDD.n873 VSS 0.016652f
C16828 VDD.n874 VSS 0.073375f
C16829 VDD.t2667 VSS 0.042023f
C16830 VDD.t2669 VSS 0.075406f
C16831 VDD.t2808 VSS 0.075406f
C16832 VDD.t2810 VSS 0.139422f
C16833 VDD.t2 VSS 0.139422f
C16834 VDD.t0 VSS 0.075406f
C16835 VDD.t2521 VSS 0.075406f
C16836 VDD.t2523 VSS 0.063624f
C16837 VDD.t2801 VSS 0.027188f
C16838 VDD.n875 VSS 0.074488f
C16839 VDD.t1491 VSS 0.027188f
C16840 VDD.n876 VSS 0.074487f
C16841 VDD.t1493 VSS 0.007233f
C16842 VDD.t3015 VSS 0.007233f
C16843 VDD.n877 VSS 0.016652f
C16844 VDD.n878 VSS 0.07634f
C16845 VDD.t2964 VSS 0.007233f
C16846 VDD.t4502 VSS 0.007233f
C16847 VDD.n879 VSS 0.016652f
C16848 VDD.n880 VSS 0.047679f
C16849 VDD.t3060 VSS 0.004807f
C16850 VDD.t3002 VSS 0.004807f
C16851 VDD.n881 VSS 0.010736f
C16852 VDD.t3064 VSS 0.017466f
C16853 VDD.n882 VSS 0.048701f
C16854 VDD.n883 VSS 0.030676f
C16855 VDD.t4373 VSS 0.145552f
C16856 VDD.t4380 VSS 0.004807f
C16857 VDD.t4443 VSS 0.004807f
C16858 VDD.n884 VSS 0.010736f
C16859 VDD.t4374 VSS 0.017466f
C16860 VDD.n885 VSS 0.048701f
C16861 VDD.t3795 VSS 0.004807f
C16862 VDD.t3879 VSS 0.004807f
C16863 VDD.n886 VSS 0.010736f
C16864 VDD.t3790 VSS 0.017466f
C16865 VDD.n887 VSS 0.059157f
C16866 VDD.t3789 VSS 0.137944f
C16867 VDD.n888 VSS 0.135842f
C16868 VDD.n889 VSS 0.031797f
C16869 VDD.n890 VSS 0.030676f
C16870 VDD.n891 VSS 0.028952f
C16871 VDD.n892 VSS 0.135842f
C16872 VDD.t3001 VSS 0.270495f
C16873 VDD.n893 VSS 0.096866f
C16874 VDD.t2807 VSS 0.027204f
C16875 VDD.n894 VSS 0.169958f
C16876 VDD.t4368 VSS 0.007233f
C16877 VDD.t2799 VSS 0.007233f
C16878 VDD.n895 VSS 0.016652f
C16879 VDD.n896 VSS 0.050644f
C16880 VDD.t4501 VSS 0.042023f
C16881 VDD.t4393 VSS 0.075406f
C16882 VDD.t2802 VSS 0.075406f
C16883 VDD.t2804 VSS 0.144962f
C16884 VDD.t435 VSS 0.14709f
C16885 VDD.t437 VSS 0.075145f
C16886 VDD.t2529 VSS 0.075145f
C16887 VDD.t2531 VSS 0.063403f
C16888 VDD.t2806 VSS 0.126024f
C16889 VDD.t2798 VSS 0.075145f
C16890 VDD.t4367 VSS 0.075145f
C16891 VDD.t4474 VSS 0.041877f
C16892 VDD.n897 VSS 0.064693f
C16893 VDD.n898 VSS 0.076519f
C16894 VDD.t2532 VSS 0.007233f
C16895 VDD.t4475 VSS 0.007233f
C16896 VDD.n899 VSS 0.016652f
C16897 VDD.n900 VSS 0.047679f
C16898 VDD.t438 VSS 0.007233f
C16899 VDD.t2530 VSS 0.007233f
C16900 VDD.n901 VSS 0.016652f
C16901 VDD.n902 VSS 0.07634f
C16902 VDD.t436 VSS 0.027188f
C16903 VDD.n903 VSS 0.076455f
C16904 VDD.t2805 VSS 0.027188f
C16905 VDD.n904 VSS 0.076457f
C16906 VDD.t4394 VSS 0.007233f
C16907 VDD.t2803 VSS 0.007233f
C16908 VDD.n905 VSS 0.016652f
C16909 VDD.n906 VSS 0.073375f
C16910 VDD.n907 VSS 0.076519f
C16911 VDD.n908 VSS 0.064809f
C16912 VDD.t2963 VSS 0.063624f
C16913 VDD.t3014 VSS 0.075406f
C16914 VDD.t1492 VSS 0.075406f
C16915 VDD.t1490 VSS 0.141386f
C16916 VDD.t2800 VSS 0.141386f
C16917 VDD.t2796 VSS 0.075406f
C16918 VDD.t2677 VSS 0.075406f
C16919 VDD.t2675 VSS 0.042023f
C16920 VDD.n909 VSS 0.064809f
C16921 VDD.n910 VSS 0.076519f
C16922 VDD.t2524 VSS 0.007233f
C16923 VDD.t2676 VSS 0.007233f
C16924 VDD.n911 VSS 0.016652f
C16925 VDD.n912 VSS 0.047679f
C16926 VDD.t1 VSS 0.007233f
C16927 VDD.t2522 VSS 0.007233f
C16928 VDD.n913 VSS 0.016652f
C16929 VDD.n914 VSS 0.07634f
C16930 VDD.t3 VSS 0.027188f
C16931 VDD.n915 VSS 0.073667f
C16932 VDD.t2811 VSS 0.027188f
C16933 VDD.n916 VSS 0.073669f
C16934 VDD.t2670 VSS 0.007233f
C16935 VDD.t2809 VSS 0.007233f
C16936 VDD.n917 VSS 0.016652f
C16937 VDD.n918 VSS 0.073375f
C16938 VDD.n919 VSS 0.076519f
C16939 VDD.n920 VSS 0.064809f
C16940 VDD.t2945 VSS 0.063624f
C16941 VDD.t2959 VSS 0.075406f
C16942 VDD.t1648 VSS 0.075406f
C16943 VDD.t1646 VSS 0.13786f
C16944 VDD.t1455 VSS 0.137401f
C16945 VDD.t1457 VSS 0.075145f
C16946 VDD.t1193 VSS 0.075145f
C16947 VDD.t1191 VSS 0.041877f
C16948 VDD.n921 VSS 0.064693f
C16949 VDD.n922 VSS 0.076519f
C16950 VDD.t3118 VSS 0.007233f
C16951 VDD.t1192 VSS 0.007233f
C16952 VDD.n923 VSS 0.016652f
C16953 VDD.n924 VSS 0.047679f
C16954 VDD.t2643 VSS 0.007233f
C16955 VDD.t3116 VSS 0.007233f
C16956 VDD.n925 VSS 0.016652f
C16957 VDD.n926 VSS 0.07634f
C16958 VDD.t2645 VSS 0.027188f
C16959 VDD.n927 VSS 0.110894f
C16960 VDD.t3917 VSS 0.004807f
C16961 VDD.t3919 VSS 0.004807f
C16962 VDD.n928 VSS 0.010736f
C16963 VDD.t3915 VSS 0.017466f
C16964 VDD.n929 VSS 0.056287f
C16965 VDD.n930 VSS 0.020342f
C16966 VDD.n931 VSS 0.030311f
C16967 VDD.t3918 VSS 0.089594f
C16968 VDD.n932 VSS 0.035424f
C16969 VDD.t3916 VSS 0.05332f
C16970 VDD.t3914 VSS 0.027493f
C16971 VDD.n933 VSS 0.067089f
C16972 VDD.n934 VSS 0.044915f
C16973 VDD.t2615 VSS 0.081296f
C16974 VDD.t2616 VSS 0.075406f
C16975 VDD.t2617 VSS 0.075406f
C16976 VDD.t2618 VSS 0.075406f
C16977 VDD.t2619 VSS 0.075406f
C16978 VDD.t3928 VSS 0.075406f
C16979 VDD.t3920 VSS 0.075406f
C16980 VDD.t3924 VSS 0.058518f
C16981 VDD.t3926 VSS 0.126462f
C16982 VDD.t3922 VSS 0.05459f
C16983 VDD.n935 VSS 2.52e-19
C16984 VDD.t3929 VSS 0.00575f
C16985 VDD.t3921 VSS 0.00575f
C16986 VDD.n936 VSS 0.0115f
C16987 VDD.n937 VSS 0.012479f
C16988 VDD.t3925 VSS 0.00575f
C16989 VDD.t3923 VSS 0.00575f
C16990 VDD.n938 VSS 0.0115f
C16991 VDD.n939 VSS 0.007448f
C16992 VDD.n940 VSS 0.076419f
C16993 VDD.t3927 VSS 0.01978f
C16994 VDD.n941 VSS 0.014195f
C16995 VDD.n942 VSS -0.011842f
C16996 VDD.n943 VSS 0.077508f
C16997 VDD.n944 VSS 0.836811f
C16998 VDD.n945 VSS 1.34367f
C16999 VDD.n946 VSS 1.29015f
C17000 VDD.n947 VSS 1.36434f
C17001 VDD.t1351 VSS 0.027215f
C17002 VDD.t657 VSS 0.007233f
C17003 VDD.t1349 VSS 0.007233f
C17004 VDD.n948 VSS 0.016652f
C17005 VDD.n949 VSS 0.129639f
C17006 VDD.t4295 VSS -0.019301f
C17007 VDD.t4293 VSS 0.075145f
C17008 VDD.t1540 VSS 0.075145f
C17009 VDD.t2848 VSS 0.063403f
C17010 VDD.t2210 VSS 0.027215f
C17011 VDD.t2212 VSS 0.007233f
C17012 VDD.t2971 VSS 0.007233f
C17013 VDD.n950 VSS 0.016652f
C17014 VDD.n951 VSS 0.132756f
C17015 VDD.t2985 VSS 0.007233f
C17016 VDD.t3211 VSS 0.007233f
C17017 VDD.n952 VSS 0.016652f
C17018 VDD.n953 VSS 0.047679f
C17019 VDD.t3203 VSS 0.007233f
C17020 VDD.t3878 VSS 0.007233f
C17021 VDD.n954 VSS 0.016652f
C17022 VDD.n955 VSS 0.073624f
C17023 VDD.t3210 VSS 0.04195f
C17024 VDD.t3208 VSS 0.075275f
C17025 VDD.t3735 VSS 0.075275f
C17026 VDD.t3718 VSS 0.139181f
C17027 VDD.t64 VSS 0.139181f
C17028 VDD.t62 VSS 0.075275f
C17029 VDD.t3230 VSS 0.075275f
C17030 VDD.t3226 VSS 0.063514f
C17031 VDD.t3851 VSS 0.027188f
C17032 VDD.n956 VSS 0.07466f
C17033 VDD.t626 VSS 0.027188f
C17034 VDD.n957 VSS 0.074656f
C17035 VDD.t624 VSS 0.007233f
C17036 VDD.t2991 VSS 0.007233f
C17037 VDD.n958 VSS 0.016652f
C17038 VDD.n959 VSS 0.076601f
C17039 VDD.t3052 VSS 0.007233f
C17040 VDD.t4372 VSS 0.007233f
C17041 VDD.n960 VSS 0.016652f
C17042 VDD.n961 VSS 0.047822f
C17043 VDD.t3853 VSS 0.027215f
C17044 VDD.t4336 VSS 0.007233f
C17045 VDD.t3859 VSS 0.007233f
C17046 VDD.n962 VSS 0.016652f
C17047 VDD.n963 VSS 0.130541f
C17048 VDD.t4371 VSS 0.04195f
C17049 VDD.t4483 VSS 0.075275f
C17050 VDD.t3803 VSS 0.075275f
C17051 VDD.t3783 VSS 0.145846f
C17052 VDD.t1248 VSS 0.145846f
C17053 VDD.t1250 VSS 0.075275f
C17054 VDD.t3222 VSS 0.075275f
C17055 VDD.t3218 VSS 0.063514f
C17056 VDD.t3852 VSS 0.126243f
C17057 VDD.t3858 VSS 0.075275f
C17058 VDD.t4335 VSS 0.075275f
C17059 VDD.t4415 VSS 0.04195f
C17060 VDD.n964 VSS 0.064751f
C17061 VDD.n965 VSS 0.07665f
C17062 VDD.t3219 VSS 0.007233f
C17063 VDD.t4416 VSS 0.007233f
C17064 VDD.n966 VSS 0.016652f
C17065 VDD.n967 VSS 0.047822f
C17066 VDD.t1251 VSS 0.007233f
C17067 VDD.t3223 VSS 0.007233f
C17068 VDD.n968 VSS 0.016652f
C17069 VDD.n969 VSS 0.076601f
C17070 VDD.t1249 VSS 0.027188f
C17071 VDD.n970 VSS 0.076624f
C17072 VDD.t3784 VSS 0.027188f
C17073 VDD.n971 VSS 0.076629f
C17074 VDD.t4484 VSS 0.007233f
C17075 VDD.t3804 VSS 0.007233f
C17076 VDD.n972 VSS 0.016652f
C17077 VDD.n973 VSS 0.073624f
C17078 VDD.n974 VSS 0.07665f
C17079 VDD.n975 VSS 0.064751f
C17080 VDD.t3051 VSS 0.063514f
C17081 VDD.t2990 VSS 0.075275f
C17082 VDD.t623 VSS 0.075275f
C17083 VDD.t625 VSS 0.141141f
C17084 VDD.t3850 VSS 0.141141f
C17085 VDD.t3877 VSS 0.075275f
C17086 VDD.t3202 VSS 0.075275f
C17087 VDD.t3206 VSS 0.04195f
C17088 VDD.n976 VSS 0.064751f
C17089 VDD.n977 VSS 0.07665f
C17090 VDD.t3227 VSS 0.007233f
C17091 VDD.t3207 VSS 0.007233f
C17092 VDD.n978 VSS 0.016652f
C17093 VDD.n979 VSS 0.047822f
C17094 VDD.t63 VSS 0.007233f
C17095 VDD.t3231 VSS 0.007233f
C17096 VDD.n980 VSS 0.016652f
C17097 VDD.n981 VSS 0.076601f
C17098 VDD.t65 VSS 0.027188f
C17099 VDD.n982 VSS 0.073849f
C17100 VDD.t3719 VSS 0.027188f
C17101 VDD.n983 VSS 0.073656f
C17102 VDD.t3209 VSS 0.007233f
C17103 VDD.t3736 VSS 0.007233f
C17104 VDD.n984 VSS 0.016652f
C17105 VDD.n985 VSS 0.073375f
C17106 VDD.n986 VSS 0.076519f
C17107 VDD.n987 VSS 0.064751f
C17108 VDD.t2984 VSS 0.063514f
C17109 VDD.t2970 VSS 0.075275f
C17110 VDD.t2211 VSS 0.075275f
C17111 VDD.t2209 VSS 0.137602f
C17112 VDD.t1350 VSS 0.137365f
C17113 VDD.t1348 VSS 0.075145f
C17114 VDD.t656 VSS 0.075145f
C17115 VDD.t658 VSS 0.041877f
C17116 VDD.n988 VSS 0.064693f
C17117 VDD.n989 VSS 0.076519f
C17118 VDD.t2849 VSS 0.007233f
C17119 VDD.t659 VSS 0.007233f
C17120 VDD.n990 VSS 0.016652f
C17121 VDD.n991 VSS 0.047679f
C17122 VDD.t4294 VSS 0.007233f
C17123 VDD.t1541 VSS 0.007233f
C17124 VDD.n992 VSS 0.016652f
C17125 VDD.n993 VSS 0.07634f
C17126 VDD.t4296 VSS 0.027188f
C17127 VDD.n994 VSS 0.256185f
C17128 VDD.n995 VSS 1.50812f
C17129 VDD.t4334 VSS 0.027215f
C17130 VDD.t81 VSS 0.007233f
C17131 VDD.t4332 VSS 0.007233f
C17132 VDD.n996 VSS 0.016652f
C17133 VDD.n997 VSS 0.129639f
C17134 VDD.t916 VSS -0.019301f
C17135 VDD.t914 VSS 0.075145f
C17136 VDD.t2109 VSS 0.075145f
C17137 VDD.t2107 VSS 0.063403f
C17138 VDD.t2032 VSS 0.027215f
C17139 VDD.t2030 VSS 0.007233f
C17140 VDD.t3079 VSS 0.007233f
C17141 VDD.n998 VSS 0.016652f
C17142 VDD.n999 VSS 0.132428f
C17143 VDD.t3102 VSS 0.007233f
C17144 VDD.t3215 VSS 0.007233f
C17145 VDD.n1000 VSS 0.016652f
C17146 VDD.n1001 VSS 0.047679f
C17147 VDD.t3201 VSS 0.007233f
C17148 VDD.t3185 VSS 0.007233f
C17149 VDD.n1002 VSS 0.016652f
C17150 VDD.n1003 VSS 0.073375f
C17151 VDD.t3214 VSS 0.042023f
C17152 VDD.t3212 VSS 0.075406f
C17153 VDD.t3172 VSS 0.075406f
C17154 VDD.t3170 VSS 0.139422f
C17155 VDD.t1532 VSS 0.139422f
C17156 VDD.t1534 VSS 0.075406f
C17157 VDD.t3228 VSS 0.075406f
C17158 VDD.t3224 VSS 0.063624f
C17159 VDD.t3179 VSS 0.027188f
C17160 VDD.n1004 VSS 0.074488f
C17161 VDD.t951 VSS 0.027188f
C17162 VDD.n1005 VSS 0.074487f
C17163 VDD.t949 VSS 0.007233f
C17164 VDD.t2995 VSS 0.007233f
C17165 VDD.n1006 VSS 0.016652f
C17166 VDD.n1007 VSS 0.07634f
C17167 VDD.t3058 VSS 0.007233f
C17168 VDD.t4361 VSS 0.007233f
C17169 VDD.n1008 VSS 0.016652f
C17170 VDD.n1009 VSS 0.047679f
C17171 VDD.t3082 VSS 0.004807f
C17172 VDD.t3071 VSS 0.004807f
C17173 VDD.n1010 VSS 0.010736f
C17174 VDD.t2983 VSS 0.017466f
C17175 VDD.n1011 VSS 0.048701f
C17176 VDD.n1012 VSS 0.030676f
C17177 VDD.t4353 VSS 0.145552f
C17178 VDD.t4354 VSS 0.004807f
C17179 VDD.t4366 VSS 0.004807f
C17180 VDD.n1013 VSS 0.010736f
C17181 VDD.t4478 VSS 0.017466f
C17182 VDD.n1014 VSS 0.048701f
C17183 VDD.t3777 VSS 0.004807f
C17184 VDD.t3782 VSS 0.004807f
C17185 VDD.n1015 VSS 0.010736f
C17186 VDD.t3734 VSS 0.017466f
C17187 VDD.n1016 VSS 0.059157f
C17188 VDD.t3733 VSS 0.137944f
C17189 VDD.n1017 VSS 0.135842f
C17190 VDD.n1018 VSS 0.031797f
C17191 VDD.n1019 VSS 0.030676f
C17192 VDD.n1020 VSS 0.028952f
C17193 VDD.n1021 VSS 0.135842f
C17194 VDD.t2982 VSS 0.270495f
C17195 VDD.n1022 VSS 0.096866f
C17196 VDD.t3181 VSS 0.027204f
C17197 VDD.n1023 VSS 0.169958f
C17198 VDD.t4509 VSS 0.007233f
C17199 VDD.t3183 VSS 0.007233f
C17200 VDD.n1024 VSS 0.016652f
C17201 VDD.n1025 VSS 0.050644f
C17202 VDD.t4360 VSS 0.042023f
C17203 VDD.t4479 VSS 0.075406f
C17204 VDD.t3176 VSS 0.075406f
C17205 VDD.t3174 VSS 0.144962f
C17206 VDD.t793 VSS 0.14709f
C17207 VDD.t791 VSS 0.075145f
C17208 VDD.t3220 VSS 0.075145f
C17209 VDD.t3216 VSS 0.063403f
C17210 VDD.t3180 VSS 0.126024f
C17211 VDD.t3182 VSS 0.075145f
C17212 VDD.t4508 VSS 0.075145f
C17213 VDD.t4407 VSS 0.041877f
C17214 VDD.n1026 VSS 0.064693f
C17215 VDD.n1027 VSS 0.076519f
C17216 VDD.t3217 VSS 0.007233f
C17217 VDD.t4408 VSS 0.007233f
C17218 VDD.n1028 VSS 0.016652f
C17219 VDD.n1029 VSS 0.047679f
C17220 VDD.t792 VSS 0.007233f
C17221 VDD.t3221 VSS 0.007233f
C17222 VDD.n1030 VSS 0.016652f
C17223 VDD.n1031 VSS 0.07634f
C17224 VDD.t794 VSS 0.027188f
C17225 VDD.n1032 VSS 0.076455f
C17226 VDD.t3175 VSS 0.027188f
C17227 VDD.n1033 VSS 0.076457f
C17228 VDD.t4480 VSS 0.007233f
C17229 VDD.t3177 VSS 0.007233f
C17230 VDD.n1034 VSS 0.016652f
C17231 VDD.n1035 VSS 0.073375f
C17232 VDD.n1036 VSS 0.076519f
C17233 VDD.n1037 VSS 0.064809f
C17234 VDD.t3057 VSS 0.063624f
C17235 VDD.t2994 VSS 0.075406f
C17236 VDD.t948 VSS 0.075406f
C17237 VDD.t950 VSS 0.141386f
C17238 VDD.t3178 VSS 0.141386f
C17239 VDD.t3184 VSS 0.075406f
C17240 VDD.t3200 VSS 0.075406f
C17241 VDD.t3204 VSS 0.042023f
C17242 VDD.n1038 VSS 0.064809f
C17243 VDD.n1039 VSS 0.076519f
C17244 VDD.t3225 VSS 0.007233f
C17245 VDD.t3205 VSS 0.007233f
C17246 VDD.n1040 VSS 0.016652f
C17247 VDD.n1041 VSS 0.047679f
C17248 VDD.t1535 VSS 0.007233f
C17249 VDD.t3229 VSS 0.007233f
C17250 VDD.n1042 VSS 0.016652f
C17251 VDD.n1043 VSS 0.07634f
C17252 VDD.t1533 VSS 0.027188f
C17253 VDD.n1044 VSS 0.073667f
C17254 VDD.t3171 VSS 0.027188f
C17255 VDD.n1045 VSS 0.073669f
C17256 VDD.t3213 VSS 0.007233f
C17257 VDD.t3173 VSS 0.007233f
C17258 VDD.n1046 VSS 0.016652f
C17259 VDD.n1047 VSS 0.073375f
C17260 VDD.n1048 VSS 0.076519f
C17261 VDD.n1049 VSS 0.064809f
C17262 VDD.t3101 VSS 0.063624f
C17263 VDD.t3078 VSS 0.075406f
C17264 VDD.t2029 VSS 0.075406f
C17265 VDD.t2031 VSS 0.13786f
C17266 VDD.t4333 VSS 0.137401f
C17267 VDD.t4331 VSS 0.075145f
C17268 VDD.t80 VSS 0.075145f
C17269 VDD.t2397 VSS 0.041877f
C17270 VDD.n1050 VSS 0.064693f
C17271 VDD.n1051 VSS 0.076519f
C17272 VDD.t2108 VSS 0.007233f
C17273 VDD.t2398 VSS 0.007233f
C17274 VDD.n1052 VSS 0.016652f
C17275 VDD.n1053 VSS 0.047679f
C17276 VDD.t915 VSS 0.007233f
C17277 VDD.t2110 VSS 0.007233f
C17278 VDD.n1054 VSS 0.016652f
C17279 VDD.n1055 VSS 0.07634f
C17280 VDD.t917 VSS 0.027188f
C17281 VDD.n1056 VSS 0.110894f
C17282 VDD.t1524 VSS 0.004807f
C17283 VDD.t1520 VSS 0.004807f
C17284 VDD.n1057 VSS 0.010736f
C17285 VDD.t1522 VSS 0.017466f
C17286 VDD.n1058 VSS 0.056287f
C17287 VDD.n1059 VSS 0.020342f
C17288 VDD.n1060 VSS 0.030311f
C17289 VDD.t1519 VSS 0.089594f
C17290 VDD.n1061 VSS 0.035424f
C17291 VDD.t1523 VSS 0.05332f
C17292 VDD.t1521 VSS 0.027493f
C17293 VDD.n1062 VSS 0.067089f
C17294 VDD.n1063 VSS 0.044915f
C17295 VDD.t2116 VSS 0.081296f
C17296 VDD.t2115 VSS 0.075406f
C17297 VDD.t2114 VSS 0.075406f
C17298 VDD.t2113 VSS 0.075406f
C17299 VDD.t2117 VSS 0.075406f
C17300 VDD.t40 VSS 0.075406f
C17301 VDD.t38 VSS 0.075406f
C17302 VDD.t36 VSS 0.058518f
C17303 VDD.t32 VSS 0.126462f
C17304 VDD.t34 VSS 0.05459f
C17305 VDD.n1064 VSS 2.52e-19
C17306 VDD.t41 VSS 0.00575f
C17307 VDD.t39 VSS 0.00575f
C17308 VDD.n1065 VSS 0.0115f
C17309 VDD.n1066 VSS 0.012479f
C17310 VDD.t37 VSS 0.00575f
C17311 VDD.t35 VSS 0.00575f
C17312 VDD.n1067 VSS 0.0115f
C17313 VDD.n1068 VSS 0.007448f
C17314 VDD.n1069 VSS 0.076419f
C17315 VDD.t33 VSS 0.01978f
C17316 VDD.n1070 VSS 0.014195f
C17317 VDD.n1071 VSS -0.011842f
C17318 VDD.n1072 VSS 0.077508f
C17319 VDD.n1073 VSS 0.836811f
C17320 VDD.n1074 VSS 1.3081f
C17321 VDD.n1075 VSS 1.25692f
C17322 VDD.n1076 VSS 1.29212f
C17323 VDD.t1324 VSS 0.027215f
C17324 VDD.t1307 VSS 0.007233f
C17325 VDD.t1326 VSS 0.007233f
C17326 VDD.n1077 VSS 0.016652f
C17327 VDD.n1078 VSS 0.129639f
C17328 VDD.t1599 VSS -0.019301f
C17329 VDD.t1597 VSS 0.075145f
C17330 VDD.t632 VSS 0.075145f
C17331 VDD.t630 VSS 0.063403f
C17332 VDD.t810 VSS 0.027215f
C17333 VDD.t808 VSS 0.007233f
C17334 VDD.t3096 VSS 0.007233f
C17335 VDD.n1079 VSS 0.016652f
C17336 VDD.n1080 VSS 0.132756f
C17337 VDD.t2940 VSS 0.007233f
C17338 VDD.t79 VSS 0.007233f
C17339 VDD.n1081 VSS 0.016652f
C17340 VDD.n1082 VSS 0.047679f
C17341 VDD.t71 VSS 0.007233f
C17342 VDD.t3732 VSS 0.007233f
C17343 VDD.n1083 VSS 0.016652f
C17344 VDD.n1084 VSS 0.073624f
C17345 VDD.t78 VSS 0.04195f
C17346 VDD.t76 VSS 0.075275f
C17347 VDD.t3753 VSS 0.075275f
C17348 VDD.t3746 VSS 0.139181f
C17349 VDD.t3695 VSS 0.139181f
C17350 VDD.t3693 VSS 0.075275f
C17351 VDD.t1263 VSS 0.075275f
C17352 VDD.t1259 VSS 0.063514f
C17353 VDD.t3711 VSS 0.027188f
C17354 VDD.n1085 VSS 0.07466f
C17355 VDD.t1061 VSS 0.027188f
C17356 VDD.n1086 VSS 0.074656f
C17357 VDD.t1063 VSS 0.007233f
C17358 VDD.t2967 VSS 0.007233f
C17359 VDD.n1087 VSS 0.016652f
C17360 VDD.n1088 VSS 0.076601f
C17361 VDD.t3009 VSS 0.007233f
C17362 VDD.t4420 VSS 0.007233f
C17363 VDD.n1089 VSS 0.016652f
C17364 VDD.n1090 VSS 0.047822f
C17365 VDD.t3713 VSS 0.027215f
C17366 VDD.t4386 VSS 0.007233f
C17367 VDD.t3721 VSS 0.007233f
C17368 VDD.n1091 VSS 0.016652f
C17369 VDD.n1092 VSS 0.130541f
C17370 VDD.t4419 VSS 0.04195f
C17371 VDD.t4337 VSS 0.075275f
C17372 VDD.t3864 VSS 0.075275f
C17373 VDD.t3834 VSS 0.145846f
C17374 VDD.t2382 VSS 0.145846f
C17375 VDD.t2380 VSS 0.075275f
C17376 VDD.t1271 VSS 0.075275f
C17377 VDD.t1267 VSS 0.063514f
C17378 VDD.t3712 VSS 0.126243f
C17379 VDD.t3720 VSS 0.075275f
C17380 VDD.t4385 VSS 0.075275f
C17381 VDD.t4446 VSS 0.04195f
C17382 VDD.n1093 VSS 0.064751f
C17383 VDD.n1094 VSS 0.07665f
C17384 VDD.t1268 VSS 0.007233f
C17385 VDD.t4447 VSS 0.007233f
C17386 VDD.n1095 VSS 0.016652f
C17387 VDD.n1096 VSS 0.047822f
C17388 VDD.t2381 VSS 0.007233f
C17389 VDD.t1272 VSS 0.007233f
C17390 VDD.n1097 VSS 0.016652f
C17391 VDD.n1098 VSS 0.076601f
C17392 VDD.t2383 VSS 0.027188f
C17393 VDD.n1099 VSS 0.076624f
C17394 VDD.t3835 VSS 0.027188f
C17395 VDD.n1100 VSS 0.076629f
C17396 VDD.t4338 VSS 0.007233f
C17397 VDD.t3865 VSS 0.007233f
C17398 VDD.n1101 VSS 0.016652f
C17399 VDD.n1102 VSS 0.073624f
C17400 VDD.n1103 VSS 0.07665f
C17401 VDD.n1104 VSS 0.064751f
C17402 VDD.t3008 VSS 0.063514f
C17403 VDD.t2966 VSS 0.075275f
C17404 VDD.t1062 VSS 0.075275f
C17405 VDD.t1060 VSS 0.141141f
C17406 VDD.t3710 VSS 0.141141f
C17407 VDD.t3731 VSS 0.075275f
C17408 VDD.t70 VSS 0.075275f
C17409 VDD.t74 VSS 0.04195f
C17410 VDD.n1105 VSS 0.064751f
C17411 VDD.n1106 VSS 0.07665f
C17412 VDD.t1260 VSS 0.007233f
C17413 VDD.t75 VSS 0.007233f
C17414 VDD.n1107 VSS 0.016652f
C17415 VDD.n1108 VSS 0.047822f
C17416 VDD.t3694 VSS 0.007233f
C17417 VDD.t1264 VSS 0.007233f
C17418 VDD.n1109 VSS 0.016652f
C17419 VDD.n1110 VSS 0.076601f
C17420 VDD.t3696 VSS 0.027188f
C17421 VDD.n1111 VSS 0.073849f
C17422 VDD.t3747 VSS 0.027188f
C17423 VDD.n1112 VSS 0.073656f
C17424 VDD.t77 VSS 0.007233f
C17425 VDD.t3754 VSS 0.007233f
C17426 VDD.n1113 VSS 0.016652f
C17427 VDD.n1114 VSS 0.073375f
C17428 VDD.n1115 VSS 0.076519f
C17429 VDD.n1116 VSS 0.064751f
C17430 VDD.t2939 VSS 0.063514f
C17431 VDD.t3095 VSS 0.075275f
C17432 VDD.t807 VSS 0.075275f
C17433 VDD.t809 VSS 0.137602f
C17434 VDD.t1323 VSS 0.137365f
C17435 VDD.t1325 VSS 0.075145f
C17436 VDD.t1306 VSS 0.075145f
C17437 VDD.t1308 VSS 0.041877f
C17438 VDD.n1117 VSS 0.064693f
C17439 VDD.n1118 VSS 0.076519f
C17440 VDD.t631 VSS 0.007233f
C17441 VDD.t1309 VSS 0.007233f
C17442 VDD.n1119 VSS 0.016652f
C17443 VDD.n1120 VSS 0.047679f
C17444 VDD.t1598 VSS 0.007233f
C17445 VDD.t633 VSS 0.007233f
C17446 VDD.n1121 VSS 0.016652f
C17447 VDD.n1122 VSS 0.07634f
C17448 VDD.t1600 VSS 0.027188f
C17449 VDD.n1123 VSS 0.256185f
C17450 VDD.n1124 VSS 1.31086f
C17451 VDD.n1125 VSS 0.667178f
C17452 VDD.t4125 VSS 0.017458f
C17453 VDD.n1126 VSS 0.052184f
C17454 VDD.t2276 VSS 0.017475f
C17455 VDD.t2272 VSS 0.004807f
C17456 VDD.t2274 VSS 0.004807f
C17457 VDD.n1127 VSS 0.010696f
C17458 VDD.n1128 VSS 0.080765f
C17459 VDD.t3501 VSS 0.004807f
C17460 VDD.t3499 VSS 0.004807f
C17461 VDD.n1129 VSS 0.010736f
C17462 VDD.t3497 VSS 0.017466f
C17463 VDD.n1130 VSS 0.052058f
C17464 VDD.t4124 VSS 0.094682f
C17465 VDD.t4128 VSS 0.056456f
C17466 VDD.t4126 VSS 0.040872f
C17467 VDD.t4127 VSS 0.004807f
C17468 VDD.t4129 VSS 0.004807f
C17469 VDD.n1131 VSS 0.010696f
C17470 VDD.n1132 VSS 0.029338f
C17471 VDD.n1133 VSS 0.023779f
C17472 VDD.n1134 VSS 7.86e-19
C17473 VDD.t2273 VSS 0.043813f
C17474 VDD.t2271 VSS 0.056456f
C17475 VDD.t2275 VSS 0.072023f
C17476 VDD.t3498 VSS 0.09826f
C17477 VDD.t3500 VSS 0.058723f
C17478 VDD.n1135 VSS 0.071067f
C17479 VDD.t3496 VSS 0.099183f
C17480 VDD.n1136 VSS 0.039448f
C17481 VDD.n1137 VSS 0.290581f
C17482 VDD.n1138 VSS 0.41179f
C17483 VDD.n1139 VSS 0.307252f
C17484 VDD.n1140 VSS 0.228067f
C17485 VDD.t3301 VSS 0.010856f
C17486 VDD.t3305 VSS 0.012354f
C17487 VDD.n1141 VSS 0.02321f
C17488 VDD.n1142 VSS 0.043917f
C17489 VDD.t3309 VSS 0.012354f
C17490 VDD.t3303 VSS 0.012354f
C17491 VDD.n1143 VSS 0.024708f
C17492 VDD.n1144 VSS 0.043917f
C17493 VDD.n1145 VSS 0.09494f
C17494 VDD.t3300 VSS 0.190115f
C17495 VDD.t3304 VSS 0.115295f
C17496 VDD.t3308 VSS 0.117748f
C17497 VDD.t3302 VSS 0.117748f
C17498 VDD.t56 VSS 0.117748f
C17499 VDD.t4123 VSS 0.117748f
C17500 VDD.t55 VSS 0.087085f
C17501 VDD.t3450 VSS 0.190115f
C17502 VDD.t3425 VSS 0.115295f
C17503 VDD.t3417 VSS 0.117748f
C17504 VDD.t2292 VSS 0.117748f
C17505 VDD.t278 VSS 0.117748f
C17506 VDD.t1846 VSS 0.117748f
C17507 VDD.t1474 VSS 0.089538f
C17508 VDD.t1392 VSS 0.010856f
C17509 VDD.t1407 VSS 0.012354f
C17510 VDD.n1146 VSS 0.038675f
C17511 VDD.t1411 VSS 0.012354f
C17512 VDD.t1385 VSS 0.012354f
C17513 VDD.n1147 VSS 0.040145f
C17514 VDD.n1148 VSS 0.059265f
C17515 VDD.n1149 VSS 0.244114f
C17516 VDD.n1150 VSS 0.244114f
C17517 VDD.n1151 VSS 0.244114f
C17518 VDD.n1152 VSS 0.244114f
C17519 VDD.n1153 VSS 0.244114f
C17520 VDD.n1154 VSS 0.244114f
C17521 VDD.n1155 VSS 0.244114f
C17522 VDD.n1156 VSS 0.538951f
C17523 VDD.t3441 VSS 0.010856f
C17524 VDD.t3428 VSS 0.012354f
C17525 VDD.n1157 VSS 0.038675f
C17526 VDD.t3422 VSS 0.012354f
C17527 VDD.t3445 VSS 0.012354f
C17528 VDD.n1158 VSS 0.040145f
C17529 VDD.n1159 VSS 0.059265f
C17530 VDD.t1450 VSS 0.088051f
C17531 VDD.t1116 VSS 0.010856f
C17532 VDD.t1145 VSS 0.012354f
C17533 VDD.n1160 VSS 0.038675f
C17534 VDD.t1124 VSS 0.012354f
C17535 VDD.t1147 VSS 0.012354f
C17536 VDD.n1161 VSS 0.040145f
C17537 VDD.n1162 VSS 0.059265f
C17538 VDD.n1163 VSS 0.532668f
C17539 VDD.n1164 VSS 0.597315f
C17540 VDD.t4211 VSS 0.017474f
C17541 VDD.t4213 VSS 0.004807f
C17542 VDD.t4229 VSS 0.004807f
C17543 VDD.n1165 VSS 0.010696f
C17544 VDD.n1166 VSS 0.09764f
C17545 VDD.t990 VSS 0.017474f
C17546 VDD.t1035 VSS 0.004807f
C17547 VDD.t584 VSS 0.004807f
C17548 VDD.n1167 VSS 0.010696f
C17549 VDD.n1168 VSS 0.097619f
C17550 VDD.t1665 VSS 0.053549f
C17551 VDD.t2235 VSS 0.017474f
C17552 VDD.t2241 VSS 0.004807f
C17553 VDD.t1666 VSS 0.004807f
C17554 VDD.n1169 VSS 0.010696f
C17555 VDD.n1170 VSS 0.09764f
C17556 VDD.n1171 VSS 0.336014f
C17557 VDD.n1172 VSS 0.848376f
C17558 VDD.t256 VSS 0.010856f
C17559 VDD.t246 VSS 0.012354f
C17560 VDD.n1173 VSS 0.038675f
C17561 VDD.t250 VSS 0.012354f
C17562 VDD.t252 VSS 0.012354f
C17563 VDD.n1174 VSS 0.040145f
C17564 VDD.n1175 VSS 0.059265f
C17565 VDD.t2918 VSS 0.012354f
C17566 VDD.t2920 VSS 0.012354f
C17567 VDD.n1176 VSS 0.040938f
C17568 VDD.t2922 VSS 0.012354f
C17569 VDD.t2912 VSS 0.010856f
C17570 VDD.n1177 VSS 0.038523f
C17571 VDD.n1178 VSS 0.058757f
C17572 VDD.t1853 VSS 0.088051f
C17573 VDD.t1938 VSS 0.532028f
C17574 VDD.t1912 VSS 0.116575f
C17575 VDD.t1936 VSS 0.119055f
C17576 VDD.t1940 VSS 0.119055f
C17577 VDD.t746 VSS 0.119055f
C17578 VDD.t745 VSS 0.119055f
C17579 VDD.t744 VSS 0.090532f
C17580 VDD.t639 VSS 0.010856f
C17581 VDD.t1608 VSS 0.012354f
C17582 VDD.n1179 VSS 0.038675f
C17583 VDD.t1612 VSS 0.012354f
C17584 VDD.t635 VSS 0.012354f
C17585 VDD.n1180 VSS 0.040145f
C17586 VDD.n1181 VSS 0.059265f
C17587 VDD.n1182 VSS 0.301692f
C17588 VDD.t441 VSS 0.004807f
C17589 VDD.t442 VSS 0.004807f
C17590 VDD.n1183 VSS 0.010736f
C17591 VDD.t440 VSS 0.017466f
C17592 VDD.n1184 VSS 0.059057f
C17593 VDD.n1185 VSS 0.047231f
C17594 VDD.t2369 VSS 0.017474f
C17595 VDD.t2375 VSS 0.004807f
C17596 VDD.t2328 VSS 0.004807f
C17597 VDD.n1186 VSS 0.010696f
C17598 VDD.n1187 VSS 0.09764f
C17599 VDD.t524 VSS 0.017474f
C17600 VDD.t515 VSS 0.004807f
C17601 VDD.t522 VSS 0.004807f
C17602 VDD.n1188 VSS 0.010696f
C17603 VDD.n1189 VSS 0.097619f
C17604 VDD.t439 VSS 0.227821f
C17605 VDD.t2368 VSS 0.169702f
C17606 VDD.t2374 VSS 0.070832f
C17607 VDD.t2327 VSS 0.054969f
C17608 VDD.t523 VSS 0.118791f
C17609 VDD.t521 VSS 0.070832f
C17610 VDD.t514 VSS 0.051279f
C17611 VDD.n1190 VSS 0.007974f
C17612 VDD.n1191 VSS 0.024454f
C17613 VDD.n1192 VSS 0.173847f
C17614 VDD.n1193 VSS 0.815703f
C17615 VDD.t2336 VSS 0.017474f
C17616 VDD.t2361 VSS 0.004807f
C17617 VDD.t2359 VSS 0.004807f
C17618 VDD.n1194 VSS 0.010696f
C17619 VDD.n1195 VSS 0.09764f
C17620 VDD.n1196 VSS 0.201715f
C17621 VDD.t1663 VSS 0.122298f
C17622 VDD.t1655 VSS 0.072923f
C17623 VDD.t2229 VSS 0.052793f
C17624 VDD.t1664 VSS 0.017474f
C17625 VDD.t2230 VSS 0.004807f
C17626 VDD.t1656 VSS 0.004807f
C17627 VDD.n1197 VSS 0.010696f
C17628 VDD.n1198 VSS 0.097619f
C17629 VDD.n1199 VSS 0.024454f
C17630 VDD.n1200 VSS 0.009019f
C17631 VDD.t2358 VSS 0.056591f
C17632 VDD.t2360 VSS 0.072923f
C17633 VDD.t2335 VSS 0.173952f
C17634 VDD.t1125 VSS 0.299488f
C17635 VDD.t1127 VSS 0.004807f
C17636 VDD.t1128 VSS 0.004807f
C17637 VDD.n1201 VSS 0.010736f
C17638 VDD.t1126 VSS 0.017466f
C17639 VDD.n1202 VSS 0.059057f
C17640 VDD.n1203 VSS 0.044914f
C17641 VDD.n1204 VSS 0.835655f
C17642 VDD.n1205 VSS 0.8887f
C17643 VDD.n1206 VSS 0.26475f
C17644 VDD.t4218 VSS 0.017474f
C17645 VDD.t4238 VSS 0.004807f
C17646 VDD.t4236 VSS 0.004807f
C17647 VDD.n1207 VSS 0.010696f
C17648 VDD.n1208 VSS 0.09764f
C17649 VDD.n1209 VSS 0.201748f
C17650 VDD.t2351 VSS 0.118791f
C17651 VDD.t2349 VSS 0.070832f
C17652 VDD.t2322 VSS 0.051279f
C17653 VDD.t2352 VSS 0.017474f
C17654 VDD.t2323 VSS 0.004807f
C17655 VDD.t2350 VSS 0.004807f
C17656 VDD.n1210 VSS 0.010696f
C17657 VDD.n1211 VSS 0.097619f
C17658 VDD.n1212 VSS 0.024454f
C17659 VDD.n1213 VSS 0.007974f
C17660 VDD.t4235 VSS 0.054969f
C17661 VDD.t4237 VSS 0.070832f
C17662 VDD.t4217 VSS 0.168226f
C17663 VDD.t3147 VSS 0.231917f
C17664 VDD.t3148 VSS 0.004807f
C17665 VDD.t3149 VSS 0.004807f
C17666 VDD.n1214 VSS 0.010736f
C17667 VDD.t3150 VSS 0.017466f
C17668 VDD.n1215 VSS 0.059057f
C17669 VDD.n1216 VSS 0.044645f
C17670 VDD.n1217 VSS 1.00467f
C17671 VDD.n1218 VSS 0.654849f
C17672 VDD.t2372 VSS 0.118791f
C17673 VDD.t2366 VSS 0.070832f
C17674 VDD.t2356 VSS 0.051279f
C17675 VDD.t4069 VSS 0.017474f
C17676 VDD.t4076 VSS 0.004807f
C17677 VDD.t4104 VSS 0.004807f
C17678 VDD.n1219 VSS 0.010696f
C17679 VDD.n1220 VSS 0.09764f
C17680 VDD.n1221 VSS 0.173847f
C17681 VDD.t2373 VSS 0.017474f
C17682 VDD.t2357 VSS 0.004807f
C17683 VDD.t2367 VSS 0.004807f
C17684 VDD.n1222 VSS 0.010696f
C17685 VDD.n1223 VSS 0.097619f
C17686 VDD.n1224 VSS 0.024454f
C17687 VDD.n1225 VSS 0.007974f
C17688 VDD.t4103 VSS 0.054969f
C17689 VDD.t4075 VSS 0.070832f
C17690 VDD.t4068 VSS 0.167488f
C17691 VDD.t2620 VSS 0.233965f
C17692 VDD.t2623 VSS 0.004807f
C17693 VDD.t2621 VSS 0.004807f
C17694 VDD.n1226 VSS 0.010736f
C17695 VDD.t2622 VSS 0.017466f
C17696 VDD.n1227 VSS 0.059057f
C17697 VDD.n1228 VSS 0.044658f
C17698 VDD.n1229 VSS 0.313597f
C17699 VDD.n1230 VSS 0.186353f
C17700 VDD.t2599 VSS 0.017474f
C17701 VDD.t472 VSS 0.004807f
C17702 VDD.t470 VSS 0.004807f
C17703 VDD.n1231 VSS 0.010696f
C17704 VDD.n1232 VSS 0.09764f
C17705 VDD.n1233 VSS 0.198901f
C17706 VDD.t1669 VSS 0.118791f
C17707 VDD.t1667 VSS 0.070832f
C17708 VDD.t2242 VSS 0.051279f
C17709 VDD.t1670 VSS 0.017474f
C17710 VDD.t2243 VSS 0.004807f
C17711 VDD.t1668 VSS 0.004807f
C17712 VDD.n1234 VSS 0.010696f
C17713 VDD.n1235 VSS 0.097619f
C17714 VDD.n1236 VSS 0.024454f
C17715 VDD.n1237 VSS 0.007974f
C17716 VDD.t469 VSS 0.054969f
C17717 VDD.t471 VSS 0.070832f
C17718 VDD.t2598 VSS 0.168964f
C17719 VDD.t1086 VSS 0.229869f
C17720 VDD.t1088 VSS 0.004807f
C17721 VDD.t1089 VSS 0.004807f
C17722 VDD.n1238 VSS 0.010736f
C17723 VDD.t1087 VSS 0.017466f
C17724 VDD.n1239 VSS 0.059084f
C17725 VDD.n1240 VSS 0.044768f
C17726 VDD.n1241 VSS 1.39038f
C17727 VDD.n1242 VSS 0.877131f
C17728 VDD.t547 VSS 0.118791f
C17729 VDD.t543 VSS 0.070832f
C17730 VDD.t535 VSS 0.051279f
C17731 VDD.t2586 VSS 0.017474f
C17732 VDD.t2591 VSS 0.004807f
C17733 VDD.t2614 VSS 0.004807f
C17734 VDD.n1243 VSS 0.010696f
C17735 VDD.n1244 VSS 0.09764f
C17736 VDD.n1245 VSS 0.173847f
C17737 VDD.t548 VSS 0.017474f
C17738 VDD.t536 VSS 0.004807f
C17739 VDD.t544 VSS 0.004807f
C17740 VDD.n1246 VSS 0.010696f
C17741 VDD.n1247 VSS 0.097619f
C17742 VDD.n1248 VSS 0.024454f
C17743 VDD.n1249 VSS 0.007974f
C17744 VDD.t2613 VSS 0.054969f
C17745 VDD.t2590 VSS 0.070832f
C17746 VDD.t2585 VSS 0.167857f
C17747 VDD.t811 VSS 0.232941f
C17748 VDD.t813 VSS 0.004807f
C17749 VDD.t814 VSS 0.004807f
C17750 VDD.n1250 VSS 0.010736f
C17751 VDD.t812 VSS 0.017466f
C17752 VDD.n1251 VSS 0.059057f
C17753 VDD.n1252 VSS 0.044651f
C17754 VDD.n1253 VSS 0.453843f
C17755 VDD.n1254 VSS 0.342027f
C17756 VDD.t4224 VSS 0.017474f
C17757 VDD.t4193 VSS 0.004807f
C17758 VDD.t4191 VSS 0.004807f
C17759 VDD.n1255 VSS 0.010696f
C17760 VDD.n1256 VSS 0.09764f
C17761 VDD.n1257 VSS 0.201767f
C17762 VDD.t2607 VSS 0.106518f
C17763 VDD.t2601 VSS 0.063514f
C17764 VDD.t2583 VSS 0.045981f
C17765 VDD.t2608 VSS 0.017474f
C17766 VDD.t2584 VSS 0.004807f
C17767 VDD.t2602 VSS 0.004807f
C17768 VDD.n1258 VSS 0.010696f
C17769 VDD.n1259 VSS 0.097619f
C17770 VDD.n1260 VSS 0.024454f
C17771 VDD.n1261 VSS 0.004315f
C17772 VDD.t4190 VSS 0.049289f
C17773 VDD.t4192 VSS 0.037537f
C17774 VDD.t4223 VSS 0.091822f
C17775 VDD.t2077 VSS 0.245355f
C17776 VDD.t2078 VSS 0.004807f
C17777 VDD.t2079 VSS 0.004807f
C17778 VDD.n1262 VSS 0.010736f
C17779 VDD.t2080 VSS 0.017466f
C17780 VDD.n1263 VSS 0.059057f
C17781 VDD.n1264 VSS 0.044832f
C17782 VDD.n1265 VSS 1.00745f
C17783 VDD.n1266 VSS 0.65801f
C17784 VDD.t476 VSS 0.106518f
C17785 VDD.t473 VSS 0.063514f
C17786 VDD.t463 VSS 0.045981f
C17787 VDD.t4082 VSS 0.017474f
C17788 VDD.t4094 VSS 0.004807f
C17789 VDD.t4114 VSS 0.004807f
C17790 VDD.n1267 VSS 0.010696f
C17791 VDD.n1268 VSS 0.09764f
C17792 VDD.n1269 VSS 0.173847f
C17793 VDD.t477 VSS 0.017474f
C17794 VDD.t464 VSS 0.004807f
C17795 VDD.t474 VSS 0.004807f
C17796 VDD.n1270 VSS 0.010696f
C17797 VDD.n1271 VSS 0.097619f
C17798 VDD.n1272 VSS 0.024454f
C17799 VDD.n1273 VSS 0.004315f
C17800 VDD.t4113 VSS 0.049289f
C17801 VDD.t4093 VSS 0.037537f
C17802 VDD.t4081 VSS 0.092153f
C17803 VDD.t4273 VSS 0.245685f
C17804 VDD.t4324 VSS 0.004807f
C17805 VDD.t4274 VSS 0.004807f
C17806 VDD.n1274 VSS 0.010736f
C17807 VDD.t4275 VSS 0.017466f
C17808 VDD.n1275 VSS 0.059057f
C17809 VDD.n1276 VSS 0.044832f
C17810 VDD.n1277 VSS 0.315345f
C17811 VDD.n1278 VSS 0.186353f
C17812 VDD.t2137 VSS 0.017474f
C17813 VDD.t2177 VSS 0.004807f
C17814 VDD.t2135 VSS 0.004807f
C17815 VDD.n1279 VSS 0.010696f
C17816 VDD.n1280 VSS 0.09764f
C17817 VDD.n1281 VSS 0.198923f
C17818 VDD.t1674 VSS 0.118791f
C17819 VDD.t1681 VSS 0.070832f
C17820 VDD.t2236 VSS 0.051279f
C17821 VDD.t1675 VSS 0.017474f
C17822 VDD.t2237 VSS 0.004807f
C17823 VDD.t1682 VSS 0.004807f
C17824 VDD.n1282 VSS 0.010696f
C17825 VDD.n1283 VSS 0.097619f
C17826 VDD.n1284 VSS 0.024454f
C17827 VDD.n1285 VSS 0.007974f
C17828 VDD.t2134 VSS 0.054969f
C17829 VDD.t2176 VSS 0.070832f
C17830 VDD.t2136 VSS 0.169333f
C17831 VDD.t725 VSS 0.228845f
C17832 VDD.t727 VSS 0.004807f
C17833 VDD.t728 VSS 0.004807f
C17834 VDD.n1286 VSS 0.010736f
C17835 VDD.t726 VSS 0.017466f
C17836 VDD.n1287 VSS 0.059057f
C17837 VDD.n1288 VSS 0.044625f
C17838 VDD.n1289 VSS 1.38878f
C17839 VDD.n1290 VSS 0.876344f
C17840 VDD.t533 VSS 0.118791f
C17841 VDD.t555 VSS 0.070832f
C17842 VDD.t259 VSS 0.051279f
C17843 VDD.t2175 VSS 0.017474f
C17844 VDD.t2171 VSS 0.004807f
C17845 VDD.t2144 VSS 0.004807f
C17846 VDD.n1291 VSS 0.010696f
C17847 VDD.n1292 VSS 0.09764f
C17848 VDD.n1293 VSS 0.173847f
C17849 VDD.t534 VSS 0.017474f
C17850 VDD.t260 VSS 0.004807f
C17851 VDD.t556 VSS 0.004807f
C17852 VDD.n1294 VSS 0.010696f
C17853 VDD.n1295 VSS 0.097619f
C17854 VDD.n1296 VSS 0.024454f
C17855 VDD.n1297 VSS 0.007974f
C17856 VDD.t2143 VSS 0.054969f
C17857 VDD.t2170 VSS 0.070832f
C17858 VDD.t2174 VSS 0.167857f
C17859 VDD.t2632 VSS 0.232941f
C17860 VDD.t2635 VSS 0.004807f
C17861 VDD.t2633 VSS 0.004807f
C17862 VDD.n1298 VSS 0.010736f
C17863 VDD.t2634 VSS 0.017466f
C17864 VDD.n1299 VSS 0.059057f
C17865 VDD.n1300 VSS 0.044651f
C17866 VDD.n1301 VSS 0.455276f
C17867 VDD.n1302 VSS 0.342027f
C17868 VDD.t4187 VSS 0.017474f
C17869 VDD.t4220 VSS 0.004807f
C17870 VDD.t4242 VSS 0.004807f
C17871 VDD.n1303 VSS 0.010696f
C17872 VDD.n1304 VSS 0.09764f
C17873 VDD.n1305 VSS 0.20174f
C17874 VDD.t2172 VSS 0.118791f
C17875 VDD.t2178 VSS 0.070832f
C17876 VDD.t2138 VSS 0.051279f
C17877 VDD.t2173 VSS 0.017474f
C17878 VDD.t2139 VSS 0.004807f
C17879 VDD.t2179 VSS 0.004807f
C17880 VDD.n1306 VSS 0.010696f
C17881 VDD.n1307 VSS 0.097619f
C17882 VDD.n1308 VSS 0.024454f
C17883 VDD.n1309 VSS 0.007974f
C17884 VDD.t4241 VSS 0.054969f
C17885 VDD.t4219 VSS 0.070832f
C17886 VDD.t4186 VSS 0.169333f
C17887 VDD.t3930 VSS 0.228845f
C17888 VDD.t3932 VSS 0.004807f
C17889 VDD.t3933 VSS 0.004807f
C17890 VDD.n1310 VSS 0.010736f
C17891 VDD.t3931 VSS 0.017466f
C17892 VDD.n1311 VSS 0.059057f
C17893 VDD.n1312 VSS 0.044625f
C17894 VDD.n1313 VSS 1.00478f
C17895 VDD.n1314 VSS 0.654698f
C17896 VDD.t2124 VSS 0.118791f
C17897 VDD.t2141 VSS 0.070832f
C17898 VDD.t2145 VSS 0.051279f
C17899 VDD.t4112 VSS 0.017474f
C17900 VDD.t4108 VSS 0.004807f
C17901 VDD.t4080 VSS 0.004807f
C17902 VDD.n1315 VSS 0.010696f
C17903 VDD.n1316 VSS 0.09764f
C17904 VDD.n1317 VSS 0.173847f
C17905 VDD.t2125 VSS 0.017474f
C17906 VDD.t2146 VSS 0.004807f
C17907 VDD.t2142 VSS 0.004807f
C17908 VDD.n1318 VSS 0.010696f
C17909 VDD.n1319 VSS 0.097619f
C17910 VDD.n1320 VSS 0.024454f
C17911 VDD.n1321 VSS 0.007974f
C17912 VDD.t4079 VSS 0.054969f
C17913 VDD.t4107 VSS 0.070832f
C17914 VDD.t4111 VSS 0.166381f
C17915 VDD.t2683 VSS 0.237037f
C17916 VDD.t2685 VSS 0.004807f
C17917 VDD.t2686 VSS 0.004807f
C17918 VDD.n1322 VSS 0.010736f
C17919 VDD.t2684 VSS 0.017466f
C17920 VDD.n1323 VSS 0.059057f
C17921 VDD.n1324 VSS 0.044677f
C17922 VDD.n1325 VSS 0.316425f
C17923 VDD.n1326 VSS 0.326881f
C17924 VDD.t3323 VSS 0.017476f
C17925 VDD.t3321 VSS 0.004807f
C17926 VDD.t3315 VSS 0.004807f
C17927 VDD.n1327 VSS 0.010696f
C17928 VDD.n1328 VSS 0.099623f
C17929 VDD.t4053 VSS 0.017474f
C17930 VDD.t4059 VSS 0.004807f
C17931 VDD.t4057 VSS 0.004807f
C17932 VDD.n1329 VSS 0.010696f
C17933 VDD.n1330 VSS 0.099467f
C17934 VDD.t946 VSS 0.052737f
C17935 VDD.t945 VSS 0.017462f
C17936 VDD.n1331 VSS 0.526294f
C17937 VDD.t2075 VSS 0.017476f
C17938 VDD.t2071 VSS 0.004807f
C17939 VDD.t2073 VSS 0.004807f
C17940 VDD.n1332 VSS 0.010696f
C17941 VDD.n1333 VSS 0.098224f
C17942 VDD.t966 VSS 0.017474f
C17943 VDD.t970 VSS 0.004807f
C17944 VDD.t968 VSS 0.004807f
C17945 VDD.n1334 VSS 0.010696f
C17946 VDD.n1335 VSS 0.099162f
C17947 VDD.t2437 VSS 0.052737f
C17948 VDD.t2444 VSS 0.017476f
C17949 VDD.t2442 VSS 0.004807f
C17950 VDD.t2438 VSS 0.004807f
C17951 VDD.n1336 VSS 0.010696f
C17952 VDD.n1337 VSS 0.099623f
C17953 VDD.n1338 VSS 0.322573f
C17954 VDD.n1339 VSS 0.165156f
C17955 VDD.t837 VSS 0.017462f
C17956 VDD.t1284 VSS 0.017474f
C17957 VDD.t1286 VSS 0.004807f
C17958 VDD.t1282 VSS 0.004807f
C17959 VDD.n1340 VSS 0.010696f
C17960 VDD.n1341 VSS 0.097619f
C17961 VDD.t4016 VSS 0.052737f
C17962 VDD.t4009 VSS 0.017476f
C17963 VDD.t4007 VSS 0.004807f
C17964 VDD.t4017 VSS 0.004807f
C17965 VDD.n1342 VSS 0.010696f
C17966 VDD.n1343 VSS 0.099623f
C17967 VDD.n1344 VSS 0.326881f
C17968 VDD.n1345 VSS 0.325933f
C17969 VDD.n1346 VSS 0.272753f
C17970 VDD.n1347 VSS 0.165156f
C17971 VDD.n1348 VSS 0.177022f
C17972 VDD.n1349 VSS 0.325933f
C17973 VDD.n1350 VSS 0.272753f
C17974 VDD.n1351 VSS 0.165156f
C17975 VDD.n1352 VSS 0.177022f
C17976 VDD.n1353 VSS 0.247768f
C17977 VDD.t2307 VSS 0.010856f
C17978 VDD.t2311 VSS 0.012354f
C17979 VDD.n1354 VSS 0.038675f
C17980 VDD.t2309 VSS 0.012354f
C17981 VDD.t2313 VSS 0.012354f
C17982 VDD.n1355 VSS 0.040145f
C17983 VDD.n1356 VSS 0.059265f
C17984 VDD.t1333 VSS 0.012354f
C17985 VDD.t1341 VSS 0.012354f
C17986 VDD.n1357 VSS 0.040938f
C17987 VDD.t1339 VSS 0.012354f
C17988 VDD.t1343 VSS 0.010856f
C17989 VDD.n1358 VSS 0.038523f
C17990 VDD.n1359 VSS 0.058757f
C17991 VDD.t3342 VSS 0.088051f
C17992 VDD.t216 VSS 0.010856f
C17993 VDD.t2418 VSS 0.012354f
C17994 VDD.n1360 VSS 0.038675f
C17995 VDD.t212 VSS 0.012354f
C17996 VDD.t214 VSS 0.012354f
C17997 VDD.n1361 VSS 0.040145f
C17998 VDD.n1362 VSS 0.059265f
C17999 VDD.n1363 VSS 0.667524f
C18000 VDD.n1364 VSS 0.166576f
C18001 VDD.t218 VSS 0.017462f
C18002 VDD.t4182 VSS 0.017474f
C18003 VDD.t4174 VSS 0.004807f
C18004 VDD.t4176 VSS 0.004807f
C18005 VDD.n1365 VSS 0.010696f
C18006 VDD.n1366 VSS 0.097619f
C18007 VDD.t1299 VSS 0.052737f
C18008 VDD.t1294 VSS 0.017476f
C18009 VDD.t1296 VSS 0.004807f
C18010 VDD.t1300 VSS 0.004807f
C18011 VDD.n1367 VSS 0.010696f
C18012 VDD.n1368 VSS 0.099623f
C18013 VDD.n1369 VSS 0.327492f
C18014 VDD.t1290 VSS 0.010856f
C18015 VDD.t1298 VSS 0.012354f
C18016 VDD.n1370 VSS 0.038675f
C18017 VDD.t1302 VSS 0.012354f
C18018 VDD.t1292 VSS 0.012354f
C18019 VDD.n1371 VSS 0.040145f
C18020 VDD.n1372 VSS 0.059265f
C18021 VDD.t290 VSS 0.012354f
C18022 VDD.t286 VSS 0.012354f
C18023 VDD.n1373 VSS 0.040938f
C18024 VDD.t288 VSS 0.012354f
C18025 VDD.t292 VSS 0.010856f
C18026 VDD.n1374 VSS 0.038523f
C18027 VDD.n1375 VSS 0.058757f
C18028 VDD.t1924 VSS 0.192225f
C18029 VDD.t1982 VSS 0.116575f
C18030 VDD.t1974 VSS 0.119055f
C18031 VDD.t1962 VSS 0.119055f
C18032 VDD.t309 VSS 0.119055f
C18033 VDD.t310 VSS 0.119055f
C18034 VDD.t308 VSS 0.088051f
C18035 VDD.t1925 VSS 0.010856f
C18036 VDD.t1983 VSS 0.012354f
C18037 VDD.n1376 VSS 0.038675f
C18038 VDD.t1975 VSS 0.012354f
C18039 VDD.t1963 VSS 0.012354f
C18040 VDD.n1377 VSS 0.040145f
C18041 VDD.n1378 VSS 0.059265f
C18042 VDD.t2059 VSS 0.012354f
C18043 VDD.t2061 VSS 0.012354f
C18044 VDD.n1379 VSS 0.040938f
C18045 VDD.t1602 VSS 0.012354f
C18046 VDD.t2055 VSS 0.010856f
C18047 VDD.n1380 VSS 0.038523f
C18048 VDD.n1381 VSS 0.058757f
C18049 VDD.n1382 VSS 0.479072f
C18050 VDD.n1383 VSS -0.041546f
C18051 VDD.t367 VSS 0.090532f
C18052 VDD.t368 VSS 0.119055f
C18053 VDD.t1539 VSS 0.119055f
C18054 VDD.t2058 VSS 0.119055f
C18055 VDD.t2060 VSS 0.119055f
C18056 VDD.t1601 VSS 0.116575f
C18057 VDD.t2054 VSS 0.254852f
C18058 VDD.t1289 VSS 0.254852f
C18059 VDD.t1297 VSS 0.116575f
C18060 VDD.t1301 VSS 0.119055f
C18061 VDD.t1291 VSS 0.119055f
C18062 VDD.t306 VSS 0.119055f
C18063 VDD.t307 VSS 0.119055f
C18064 VDD.t305 VSS 0.088051f
C18065 VDD.t3287 VSS 0.119055f
C18066 VDD.t3286 VSS 0.119055f
C18067 VDD.t213 VSS 0.119055f
C18068 VDD.t211 VSS 0.119055f
C18069 VDD.t2417 VSS 0.116575f
C18070 VDD.t215 VSS 0.362126f
C18071 VDD.t291 VSS 0.362126f
C18072 VDD.t287 VSS 0.116575f
C18073 VDD.t285 VSS 0.119055f
C18074 VDD.t289 VSS 0.119055f
C18075 VDD.t2863 VSS 0.119055f
C18076 VDD.t2862 VSS 0.119055f
C18077 VDD.t2650 VSS 0.090532f
C18078 VDD.n1384 VSS -0.041546f
C18079 VDD.n1385 VSS 0.479072f
C18080 VDD.n1386 VSS 0.22487f
C18081 VDD.n1387 VSS 0.290998f
C18082 VDD.n1388 VSS 0.646669f
C18083 VDD.t222 VSS 0.017474f
C18084 VDD.t224 VSS 0.004807f
C18085 VDD.t226 VSS 0.004807f
C18086 VDD.n1389 VSS 0.010696f
C18087 VDD.n1390 VSS 0.097975f
C18088 VDD.n1391 VSS 0.046984f
C18089 VDD.t1911 VSS 0.017462f
C18090 VDD.t2057 VSS 0.017474f
C18091 VDD.t1604 VSS 0.004807f
C18092 VDD.t2053 VSS 0.004807f
C18093 VDD.n1392 VSS 0.010696f
C18094 VDD.n1393 VSS 0.097619f
C18095 VDD.t221 VSS 0.19396f
C18096 VDD.t223 VSS 0.067957f
C18097 VDD.t225 VSS 0.052737f
C18098 VDD.t2247 VSS 0.017474f
C18099 VDD.t2249 VSS 0.004807f
C18100 VDD.t2426 VSS 0.004807f
C18101 VDD.n1394 VSS 0.010696f
C18102 VDD.n1395 VSS 0.099162f
C18103 VDD.n1396 VSS 0.02587f
C18104 VDD.n1397 VSS 0.006536f
C18105 VDD.t2248 VSS 0.049198f
C18106 VDD.t2425 VSS 0.067957f
C18107 VDD.t2246 VSS 0.176263f
C18108 VDD.t1910 VSS 0.176263f
C18109 VDD.t1980 VSS 0.067957f
C18110 VDD.t1978 VSS 0.052737f
C18111 VDD.t1295 VSS 0.067957f
C18112 VDD.t1293 VSS 0.256608f
C18113 VDD.t2056 VSS 0.256608f
C18114 VDD.t2052 VSS 0.067957f
C18115 VDD.t1603 VSS 0.049198f
C18116 VDD.n1398 VSS 0.006536f
C18117 VDD.n1399 VSS 0.024888f
C18118 VDD.t1981 VSS 0.004807f
C18119 VDD.t1979 VSS 0.004807f
C18120 VDD.n1400 VSS 0.010696f
C18121 VDD.n1401 VSS 0.036584f
C18122 VDD.n1402 VSS 0.092113f
C18123 VDD.n1403 VSS 0.273535f
C18124 VDD.n1404 VSS 0.336089f
C18125 VDD.n1405 VSS 0.374912f
C18126 VDD.n1406 VSS 0.323484f
C18127 VDD.n1407 VSS 0.175602f
C18128 VDD.n1408 VSS 0.166576f
C18129 VDD.n1409 VSS 0.356684f
C18130 VDD.n1410 VSS 0.374912f
C18131 VDD.n1411 VSS 0.323484f
C18132 VDD.n1412 VSS 0.175602f
C18133 VDD.n1413 VSS 0.137976f
C18134 VDD.t4005 VSS 0.017476f
C18135 VDD.t4003 VSS 0.004807f
C18136 VDD.t4001 VSS 0.004807f
C18137 VDD.n1414 VSS 0.010696f
C18138 VDD.n1415 VSS 0.098224f
C18139 VDD.t3410 VSS 0.017474f
C18140 VDD.t3408 VSS 0.004807f
C18141 VDD.t3412 VSS 0.004807f
C18142 VDD.n1416 VSS 0.010696f
C18143 VDD.n1417 VSS 0.099162f
C18144 VDD.t1942 VSS 0.052737f
C18145 VDD.t1929 VSS 0.017462f
C18146 VDD.t2105 VSS 0.017474f
C18147 VDD.t2103 VSS 0.004807f
C18148 VDD.t2101 VSS 0.004807f
C18149 VDD.n1418 VSS 0.010696f
C18150 VDD.n1419 VSS 0.097975f
C18151 VDD.t869 VSS 0.017474f
C18152 VDD.t867 VSS 0.004807f
C18153 VDD.t871 VSS 0.004807f
C18154 VDD.n1420 VSS 0.010696f
C18155 VDD.n1421 VSS 0.099162f
C18156 VDD.t2104 VSS 0.19396f
C18157 VDD.t2102 VSS 0.067957f
C18158 VDD.t2100 VSS 0.052737f
C18159 VDD.t1930 VSS 0.067957f
C18160 VDD.t1928 VSS 0.176263f
C18161 VDD.t868 VSS 0.176263f
C18162 VDD.t870 VSS 0.067957f
C18163 VDD.t866 VSS 0.049198f
C18164 VDD.n1422 VSS 0.006536f
C18165 VDD.n1423 VSS 0.02587f
C18166 VDD.n1424 VSS 0.047051f
C18167 VDD.t1935 VSS 0.010856f
C18168 VDD.t1947 VSS 0.012354f
C18169 VDD.n1425 VSS 0.038675f
C18170 VDD.t1955 VSS 0.012354f
C18171 VDD.t1959 VSS 0.012354f
C18172 VDD.n1426 VSS 0.040145f
C18173 VDD.n1427 VSS 0.059265f
C18174 VDD.t1934 VSS 0.192225f
C18175 VDD.t1946 VSS 0.116575f
C18176 VDD.t1954 VSS 0.119055f
C18177 VDD.t1958 VSS 0.119055f
C18178 VDD.t907 VSS 0.119055f
C18179 VDD.t906 VSS 0.119055f
C18180 VDD.t905 VSS 0.088051f
C18181 VDD.t1313 VSS 0.090532f
C18182 VDD.t2440 VSS 0.010856f
C18183 VDD.t2450 VSS 0.012354f
C18184 VDD.n1428 VSS 0.038675f
C18185 VDD.t2448 VSS 0.012354f
C18186 VDD.t2446 VSS 0.012354f
C18187 VDD.n1429 VSS 0.040145f
C18188 VDD.n1430 VSS 0.059265f
C18189 VDD.n1431 VSS 0.356684f
C18190 VDD.t941 VSS 0.010856f
C18191 VDD.t937 VSS 0.012354f
C18192 VDD.n1432 VSS 0.038675f
C18193 VDD.t939 VSS 0.012354f
C18194 VDD.t935 VSS 0.012354f
C18195 VDD.n1433 VSS 0.040145f
C18196 VDD.n1434 VSS 0.059265f
C18197 VDD.t3658 VSS 0.012354f
C18198 VDD.t3654 VSS 0.012354f
C18199 VDD.n1435 VSS 0.040938f
C18200 VDD.t3656 VSS 0.012354f
C18201 VDD.t3666 VSS 0.010856f
C18202 VDD.n1436 VSS 0.038523f
C18203 VDD.n1437 VSS 0.058757f
C18204 VDD.t1314 VSS 0.119055f
C18205 VDD.t1315 VSS 0.119055f
C18206 VDD.t1815 VSS 0.119055f
C18207 VDD.t160 VSS 0.119055f
C18208 VDD.t156 VSS 0.116575f
C18209 VDD.t150 VSS 0.362126f
C18210 VDD.t940 VSS 0.362126f
C18211 VDD.t936 VSS 0.116575f
C18212 VDD.t938 VSS 0.119055f
C18213 VDD.t934 VSS 0.119055f
C18214 VDD.t2728 VSS 0.119055f
C18215 VDD.t2727 VSS 0.119055f
C18216 VDD.t2726 VSS 0.088051f
C18217 VDD.t4050 VSS 0.532028f
C18218 VDD.t4054 VSS 0.116575f
C18219 VDD.t4060 VSS 0.119055f
C18220 VDD.t4062 VSS 0.119055f
C18221 VDD.t3455 VSS 0.119055f
C18222 VDD.t3453 VSS 0.119055f
C18223 VDD.t3454 VSS 0.090532f
C18224 VDD.t3319 VSS 0.010856f
C18225 VDD.t3317 VSS 0.012354f
C18226 VDD.n1438 VSS 0.038675f
C18227 VDD.t3313 VSS 0.012354f
C18228 VDD.t3311 VSS 0.012354f
C18229 VDD.n1439 VSS 0.040145f
C18230 VDD.n1440 VSS 0.059265f
C18231 VDD.n1441 VSS 0.22487f
C18232 VDD.t4063 VSS 0.012354f
C18233 VDD.t4061 VSS 0.012354f
C18234 VDD.n1442 VSS 0.040938f
C18235 VDD.t4055 VSS 0.012354f
C18236 VDD.t4051 VSS 0.010856f
C18237 VDD.n1443 VSS 0.038523f
C18238 VDD.n1444 VSS 0.058757f
C18239 VDD.n1445 VSS 0.479072f
C18240 VDD.n1446 VSS -0.041546f
C18241 VDD.t2430 VSS 0.088051f
C18242 VDD.t2431 VSS 0.119055f
C18243 VDD.t2432 VSS 0.119055f
C18244 VDD.t3310 VSS 0.119055f
C18245 VDD.t3312 VSS 0.119055f
C18246 VDD.t3316 VSS 0.116575f
C18247 VDD.t3318 VSS 0.254852f
C18248 VDD.t3665 VSS 0.254852f
C18249 VDD.t3655 VSS 0.116575f
C18250 VDD.t3653 VSS 0.119055f
C18251 VDD.t3657 VSS 0.119055f
C18252 VDD.t2484 VSS 0.119055f
C18253 VDD.t1548 VSS 0.119055f
C18254 VDD.t1549 VSS 0.090532f
C18255 VDD.n1447 VSS -0.041546f
C18256 VDD.n1448 VSS 0.479072f
C18257 VDD.n1449 VSS 0.22487f
C18258 VDD.n1450 VSS 0.376311f
C18259 VDD.n1451 VSS 0.174791f
C18260 VDD.n1452 VSS 0.167387f
C18261 VDD.n1453 VSS 0.376311f
C18262 VDD.t29 VSS 0.010856f
C18263 VDD.t19 VSS 0.012354f
C18264 VDD.n1454 VSS 0.038675f
C18265 VDD.t23 VSS 0.012354f
C18266 VDD.t27 VSS 0.012354f
C18267 VDD.n1455 VSS 0.040145f
C18268 VDD.n1456 VSS 0.059265f
C18269 VDD.t4035 VSS 0.012354f
C18270 VDD.t4037 VSS 0.012354f
C18271 VDD.n1457 VSS 0.040938f
C18272 VDD.t4029 VSS 0.012354f
C18273 VDD.t4033 VSS 0.010856f
C18274 VDD.n1458 VSS 0.038523f
C18275 VDD.n1459 VSS 0.058757f
C18276 VDD.t1916 VSS 0.192225f
C18277 VDD.t1970 VSS 0.116575f
C18278 VDD.t1960 VSS 0.119055f
C18279 VDD.t1948 VSS 0.119055f
C18280 VDD.t1701 VSS 0.119055f
C18281 VDD.t1836 VSS 0.119055f
C18282 VDD.t1190 VSS 0.088051f
C18283 VDD.t1917 VSS 0.010856f
C18284 VDD.t1971 VSS 0.012354f
C18285 VDD.n1460 VSS 0.038675f
C18286 VDD.t1961 VSS 0.012354f
C18287 VDD.t1949 VSS 0.012354f
C18288 VDD.n1461 VSS 0.040145f
C18289 VDD.n1462 VSS 0.059265f
C18290 VDD.t1591 VSS 0.012354f
C18291 VDD.t598 VSS 0.012354f
C18292 VDD.n1463 VSS 0.040938f
C18293 VDD.t600 VSS 0.012354f
C18294 VDD.t604 VSS 0.010856f
C18295 VDD.n1464 VSS 0.038523f
C18296 VDD.n1465 VSS 0.058757f
C18297 VDD.t2742 VSS 0.017474f
C18298 VDD.t2744 VSS 0.004807f
C18299 VDD.t2746 VSS 0.004807f
C18300 VDD.n1466 VSS 0.010696f
C18301 VDD.n1467 VSS 0.097975f
C18302 VDD.n1468 VSS 0.047061f
C18303 VDD.t1967 VSS 0.017462f
C18304 VDD.t1593 VSS 0.017474f
C18305 VDD.t602 VSS 0.004807f
C18306 VDD.t1589 VSS 0.004807f
C18307 VDD.n1469 VSS 0.010696f
C18308 VDD.n1470 VSS 0.097619f
C18309 VDD.t2741 VSS 0.19396f
C18310 VDD.t2743 VSS 0.067957f
C18311 VDD.t2745 VSS 0.052737f
C18312 VDD.t2216 VSS 0.017474f
C18313 VDD.t2218 VSS 0.004807f
C18314 VDD.t2214 VSS 0.004807f
C18315 VDD.n1471 VSS 0.010696f
C18316 VDD.n1472 VSS 0.099162f
C18317 VDD.n1473 VSS 0.02587f
C18318 VDD.n1474 VSS 0.006536f
C18319 VDD.t2217 VSS 0.049198f
C18320 VDD.t2213 VSS 0.067957f
C18321 VDD.t2215 VSS 0.176263f
C18322 VDD.t1966 VSS 0.176263f
C18323 VDD.t1956 VSS 0.067957f
C18324 VDD.t1952 VSS 0.052737f
C18325 VDD.t2716 VSS 0.454462f
C18326 VDD.t2712 VSS 0.067957f
C18327 VDD.t2724 VSS 0.049198f
C18328 VDD.t4244 VSS 0.017476f
C18329 VDD.t4250 VSS 0.004807f
C18330 VDD.t3937 VSS 0.004807f
C18331 VDD.n1475 VSS 0.010696f
C18332 VDD.n1476 VSS 0.099623f
C18333 VDD.n1477 VSS 0.026083f
C18334 VDD.t2717 VSS 0.017474f
C18335 VDD.t2725 VSS 0.004807f
C18336 VDD.t2713 VSS 0.004807f
C18337 VDD.n1478 VSS 0.010696f
C18338 VDD.n1479 VSS 0.099467f
C18339 VDD.n1480 VSS 0.025249f
C18340 VDD.n1481 VSS 0.006536f
C18341 VDD.t3936 VSS 0.052737f
C18342 VDD.t4249 VSS 0.067957f
C18343 VDD.t4243 VSS 0.256608f
C18344 VDD.t2250 VSS 0.256608f
C18345 VDD.t1050 VSS 0.067957f
C18346 VDD.t1048 VSS 0.049198f
C18347 VDD.t4149 VSS 0.017462f
C18348 VDD.n1482 VSS 0.357653f
C18349 VDD.n1483 VSS 0.32785f
C18350 VDD.n1484 VSS 0.137976f
C18351 VDD.n1485 VSS 0.092113f
C18352 VDD.t4155 VSS 0.004807f
C18353 VDD.t4153 VSS 0.004807f
C18354 VDD.n1486 VSS 0.010696f
C18355 VDD.n1487 VSS 0.036584f
C18356 VDD.t2251 VSS 0.017474f
C18357 VDD.t1049 VSS 0.004807f
C18358 VDD.t1051 VSS 0.004807f
C18359 VDD.n1488 VSS 0.010696f
C18360 VDD.n1489 VSS 0.097619f
C18361 VDD.n1490 VSS 0.024888f
C18362 VDD.n1491 VSS 0.006536f
C18363 VDD.t4152 VSS 0.052737f
C18364 VDD.t4154 VSS 0.067957f
C18365 VDD.t4148 VSS 0.176263f
C18366 VDD.t142 VSS 0.176263f
C18367 VDD.t146 VSS 0.067957f
C18368 VDD.t144 VSS 0.049198f
C18369 VDD.t574 VSS 0.017476f
C18370 VDD.t572 VSS 0.004807f
C18371 VDD.t576 VSS 0.004807f
C18372 VDD.n1492 VSS 0.010696f
C18373 VDD.n1493 VSS 0.098224f
C18374 VDD.n1494 VSS 0.040206f
C18375 VDD.t143 VSS 0.017474f
C18376 VDD.t145 VSS 0.004807f
C18377 VDD.t147 VSS 0.004807f
C18378 VDD.n1495 VSS 0.010696f
C18379 VDD.n1496 VSS 0.099162f
C18380 VDD.n1497 VSS 0.02587f
C18381 VDD.n1498 VSS 0.006536f
C18382 VDD.t575 VSS 0.052737f
C18383 VDD.t571 VSS 0.067957f
C18384 VDD.t573 VSS 0.324211f
C18385 VDD.t4030 VSS 0.324211f
C18386 VDD.t4024 VSS 0.067957f
C18387 VDD.t4026 VSS 0.049198f
C18388 VDD.t21 VSS 0.017476f
C18389 VDD.t25 VSS 0.004807f
C18390 VDD.t31 VSS 0.004807f
C18391 VDD.n1499 VSS 0.010696f
C18392 VDD.n1500 VSS 0.099623f
C18393 VDD.n1501 VSS 0.026083f
C18394 VDD.t4031 VSS 0.017474f
C18395 VDD.t4027 VSS 0.004807f
C18396 VDD.t4025 VSS 0.004807f
C18397 VDD.n1502 VSS 0.010696f
C18398 VDD.n1503 VSS 0.099467f
C18399 VDD.n1504 VSS 0.025249f
C18400 VDD.n1505 VSS 0.006536f
C18401 VDD.t30 VSS 0.052737f
C18402 VDD.t24 VSS 0.067957f
C18403 VDD.t20 VSS 0.256608f
C18404 VDD.t668 VSS 0.256608f
C18405 VDD.t662 VSS 0.067957f
C18406 VDD.t660 VSS 0.049198f
C18407 VDD.t3670 VSS 0.017462f
C18408 VDD.n1506 VSS 0.323543f
C18409 VDD.n1507 VSS 0.32785f
C18410 VDD.n1508 VSS 0.137976f
C18411 VDD.n1509 VSS 0.092113f
C18412 VDD.t3674 VSS 0.004807f
C18413 VDD.t3678 VSS 0.004807f
C18414 VDD.n1510 VSS 0.010696f
C18415 VDD.n1511 VSS 0.036584f
C18416 VDD.t669 VSS 0.017474f
C18417 VDD.t661 VSS 0.004807f
C18418 VDD.t663 VSS 0.004807f
C18419 VDD.n1512 VSS 0.010696f
C18420 VDD.n1513 VSS 0.097619f
C18421 VDD.n1514 VSS 0.024888f
C18422 VDD.n1515 VSS 0.006536f
C18423 VDD.t3677 VSS 0.052737f
C18424 VDD.t3673 VSS 0.067957f
C18425 VDD.t3669 VSS 0.176263f
C18426 VDD.t4048 VSS 0.176263f
C18427 VDD.t4046 VSS 0.067957f
C18428 VDD.t4044 VSS 0.049198f
C18429 VDD.t4041 VSS 0.017476f
C18430 VDD.t4039 VSS 0.004807f
C18431 VDD.t4043 VSS 0.004807f
C18432 VDD.n1516 VSS 0.010696f
C18433 VDD.n1517 VSS 0.098224f
C18434 VDD.n1518 VSS 0.040206f
C18435 VDD.t4049 VSS 0.017474f
C18436 VDD.t4045 VSS 0.004807f
C18437 VDD.t4047 VSS 0.004807f
C18438 VDD.n1519 VSS 0.010696f
C18439 VDD.n1520 VSS 0.099162f
C18440 VDD.n1521 VSS 0.02587f
C18441 VDD.n1522 VSS 0.006536f
C18442 VDD.t4042 VSS 0.052737f
C18443 VDD.t4038 VSS 0.067957f
C18444 VDD.t4040 VSS 0.324211f
C18445 VDD.t3279 VSS 0.324211f
C18446 VDD.t3273 VSS 0.067957f
C18447 VDD.t3269 VSS 0.049198f
C18448 VDD.t104 VSS 0.017476f
C18449 VDD.t106 VSS 0.004807f
C18450 VDD.t108 VSS 0.004807f
C18451 VDD.n1523 VSS 0.010696f
C18452 VDD.n1524 VSS 0.099623f
C18453 VDD.n1525 VSS 0.026083f
C18454 VDD.t3280 VSS 0.017474f
C18455 VDD.t3270 VSS 0.004807f
C18456 VDD.t3274 VSS 0.004807f
C18457 VDD.n1526 VSS 0.010696f
C18458 VDD.n1527 VSS 0.099467f
C18459 VDD.n1528 VSS 0.025249f
C18460 VDD.n1529 VSS 0.006536f
C18461 VDD.t107 VSS 0.052737f
C18462 VDD.t105 VSS 0.067957f
C18463 VDD.t103 VSS 0.256608f
C18464 VDD.t3895 VSS 0.256608f
C18465 VDD.t3889 VSS 0.067957f
C18466 VDD.t3887 VSS 0.049198f
C18467 VDD.t4292 VSS 0.017462f
C18468 VDD.n1530 VSS 0.357653f
C18469 VDD.n1531 VSS 0.32785f
C18470 VDD.n1532 VSS 0.137976f
C18471 VDD.n1533 VSS 0.092113f
C18472 VDD.t4280 VSS 0.004807f
C18473 VDD.t4286 VSS 0.004807f
C18474 VDD.n1534 VSS 0.010696f
C18475 VDD.n1535 VSS 0.036584f
C18476 VDD.t3896 VSS 0.017474f
C18477 VDD.t3888 VSS 0.004807f
C18478 VDD.t3890 VSS 0.004807f
C18479 VDD.n1536 VSS 0.010696f
C18480 VDD.n1537 VSS 0.097619f
C18481 VDD.n1538 VSS 0.024888f
C18482 VDD.n1539 VSS 0.006536f
C18483 VDD.t4285 VSS 0.052737f
C18484 VDD.t4279 VSS 0.067957f
C18485 VDD.t4291 VSS 0.176263f
C18486 VDD.t4269 VSS 0.176263f
C18487 VDD.t4267 VSS 0.067957f
C18488 VDD.t4265 VSS 0.049198f
C18489 VDD.t3682 VSS 0.017476f
C18490 VDD.t3684 VSS 0.004807f
C18491 VDD.t3686 VSS 0.004807f
C18492 VDD.n1540 VSS 0.010696f
C18493 VDD.n1541 VSS 0.098224f
C18494 VDD.n1542 VSS 0.040206f
C18495 VDD.t4270 VSS 0.017474f
C18496 VDD.t4266 VSS 0.004807f
C18497 VDD.t4268 VSS 0.004807f
C18498 VDD.n1543 VSS 0.010696f
C18499 VDD.n1544 VSS 0.099162f
C18500 VDD.n1545 VSS 0.02587f
C18501 VDD.n1546 VSS 0.006536f
C18502 VDD.t3685 VSS 0.052737f
C18503 VDD.t3683 VSS 0.067957f
C18504 VDD.t3681 VSS 0.324211f
C18505 VDD.t2503 VSS 0.324211f
C18506 VDD.t2499 VSS 0.067957f
C18507 VDD.t2497 VSS 0.049198f
C18508 VDD.t3193 VSS 0.017476f
C18509 VDD.t3195 VSS 0.004807f
C18510 VDD.t3187 VSS 0.004807f
C18511 VDD.n1547 VSS 0.010696f
C18512 VDD.n1548 VSS 0.099623f
C18513 VDD.n1549 VSS 0.026083f
C18514 VDD.t2504 VSS 0.017474f
C18515 VDD.t2498 VSS 0.004807f
C18516 VDD.t2500 VSS 0.004807f
C18517 VDD.n1550 VSS 0.010696f
C18518 VDD.n1551 VSS 0.099467f
C18519 VDD.n1552 VSS 0.025249f
C18520 VDD.n1553 VSS 0.006536f
C18521 VDD.t3186 VSS 0.052737f
C18522 VDD.t3194 VSS 0.067957f
C18523 VDD.t3192 VSS 0.256608f
C18524 VDD.t1592 VSS 0.256608f
C18525 VDD.t1588 VSS 0.067957f
C18526 VDD.t601 VSS 0.049198f
C18527 VDD.n1554 VSS 0.006536f
C18528 VDD.n1555 VSS 0.024888f
C18529 VDD.t1957 VSS 0.004807f
C18530 VDD.t1953 VSS 0.004807f
C18531 VDD.n1556 VSS 0.010696f
C18532 VDD.n1557 VSS 0.036584f
C18533 VDD.n1558 VSS 0.092113f
C18534 VDD.n1559 VSS 0.27508f
C18535 VDD.n1560 VSS 0.32785f
C18536 VDD.n1561 VSS 0.709936f
C18537 VDD.n1562 VSS 0.326043f
C18538 VDD.n1563 VSS 0.479072f
C18539 VDD.n1564 VSS -0.041546f
C18540 VDD.t1041 VSS 0.090532f
C18541 VDD.t1042 VSS 0.119055f
C18542 VDD.t1043 VSS 0.119055f
C18543 VDD.t1590 VSS 0.119055f
C18544 VDD.t597 VSS 0.119055f
C18545 VDD.t599 VSS 0.116575f
C18546 VDD.t603 VSS 0.254852f
C18547 VDD.t3188 VSS 0.254852f
C18548 VDD.t3196 VSS 0.116575f
C18549 VDD.t3198 VSS 0.119055f
C18550 VDD.t3190 VSS 0.119055f
C18551 VDD.t1080 VSS 0.119055f
C18552 VDD.t1081 VSS 0.119055f
C18553 VDD.t1347 VSS 0.088051f
C18554 VDD.t3189 VSS 0.010856f
C18555 VDD.t3197 VSS 0.012354f
C18556 VDD.n1565 VSS 0.038675f
C18557 VDD.t3199 VSS 0.012354f
C18558 VDD.t3191 VSS 0.012354f
C18559 VDD.n1566 VSS 0.040145f
C18560 VDD.n1567 VSS 0.059265f
C18561 VDD.n1568 VSS 0.22487f
C18562 VDD.t2508 VSS 0.012354f
C18563 VDD.t2502 VSS 0.012354f
C18564 VDD.n1569 VSS 0.040938f
C18565 VDD.t2506 VSS 0.012354f
C18566 VDD.t2510 VSS 0.010856f
C18567 VDD.n1570 VSS 0.038523f
C18568 VDD.n1571 VSS 0.058757f
C18569 VDD.n1572 VSS 0.479072f
C18570 VDD.n1573 VSS -0.041546f
C18571 VDD.t699 VSS 0.090532f
C18572 VDD.t1699 VSS 0.119055f
C18573 VDD.t1700 VSS 0.119055f
C18574 VDD.t2507 VSS 0.119055f
C18575 VDD.t2501 VSS 0.119055f
C18576 VDD.t2505 VSS 0.116575f
C18577 VDD.t2509 VSS 0.362126f
C18578 VDD.t4289 VSS 0.362126f
C18579 VDD.t4281 VSS 0.116575f
C18580 VDD.t4283 VSS 0.119055f
C18581 VDD.t4287 VSS 0.119055f
C18582 VDD.t2434 VSS 0.119055f
C18583 VDD.t3382 VSS 0.119055f
C18584 VDD.t2433 VSS 0.088051f
C18585 VDD.t4290 VSS 0.010856f
C18586 VDD.t4282 VSS 0.012354f
C18587 VDD.n1574 VSS 0.038675f
C18588 VDD.t4284 VSS 0.012354f
C18589 VDD.t4288 VSS 0.012354f
C18590 VDD.n1575 VSS 0.040145f
C18591 VDD.n1576 VSS 0.059265f
C18592 VDD.n1577 VSS 0.22487f
C18593 VDD.t3892 VSS 0.012354f
C18594 VDD.t3884 VSS 0.012354f
C18595 VDD.n1578 VSS 0.040938f
C18596 VDD.t3886 VSS 0.012354f
C18597 VDD.t3894 VSS 0.010856f
C18598 VDD.n1579 VSS 0.038523f
C18599 VDD.n1580 VSS 0.058757f
C18600 VDD.n1581 VSS 0.479072f
C18601 VDD.n1582 VSS -0.041546f
C18602 VDD.t1838 VSS 0.090532f
C18603 VDD.t1837 VSS 0.119055f
C18604 VDD.t1839 VSS 0.119055f
C18605 VDD.t3891 VSS 0.119055f
C18606 VDD.t3883 VSS 0.119055f
C18607 VDD.t3885 VSS 0.116575f
C18608 VDD.t3893 VSS 0.254852f
C18609 VDD.t109 VSS 0.254852f
C18610 VDD.t113 VSS 0.116575f
C18611 VDD.t111 VSS 0.119055f
C18612 VDD.t115 VSS 0.119055f
C18613 VDD.t3620 VSS 0.119055f
C18614 VDD.t3621 VSS 0.119055f
C18615 VDD.t3622 VSS 0.088051f
C18616 VDD.t110 VSS 0.010856f
C18617 VDD.t114 VSS 0.012354f
C18618 VDD.n1583 VSS 0.038675f
C18619 VDD.t112 VSS 0.012354f
C18620 VDD.t116 VSS 0.012354f
C18621 VDD.n1584 VSS 0.040145f
C18622 VDD.n1585 VSS 0.059265f
C18623 VDD.t3272 VSS 0.012354f
C18624 VDD.t3278 VSS 0.012354f
C18625 VDD.n1586 VSS 0.040938f
C18626 VDD.t3276 VSS 0.012354f
C18627 VDD.t3495 VSS 0.010856f
C18628 VDD.n1587 VSS 0.038523f
C18629 VDD.n1588 VSS 0.058757f
C18630 VDD.n1589 VSS 0.22487f
C18631 VDD.n1590 VSS 0.479072f
C18632 VDD.n1591 VSS -0.041546f
C18633 VDD.t3691 VSS 0.090532f
C18634 VDD.t3689 VSS 0.119055f
C18635 VDD.t3688 VSS 0.119055f
C18636 VDD.t3271 VSS 0.119055f
C18637 VDD.t3277 VSS 0.119055f
C18638 VDD.t3275 VSS 0.116575f
C18639 VDD.t3494 VSS 0.362126f
C18640 VDD.t3667 VSS 0.362126f
C18641 VDD.t3671 VSS 0.116575f
C18642 VDD.t3675 VSS 0.119055f
C18643 VDD.t3679 VSS 0.119055f
C18644 VDD.t60 VSS 0.119055f
C18645 VDD.t59 VSS 0.119055f
C18646 VDD.t61 VSS 0.088051f
C18647 VDD.t3668 VSS 0.010856f
C18648 VDD.t3672 VSS 0.012354f
C18649 VDD.n1592 VSS 0.038675f
C18650 VDD.t3676 VSS 0.012354f
C18651 VDD.t3680 VSS 0.012354f
C18652 VDD.n1593 VSS 0.040145f
C18653 VDD.n1594 VSS 0.059265f
C18654 VDD.n1595 VSS 0.22487f
C18655 VDD.t665 VSS 0.012354f
C18656 VDD.t671 VSS 0.012354f
C18657 VDD.n1596 VSS 0.040938f
C18658 VDD.t673 VSS 0.012354f
C18659 VDD.t667 VSS 0.010856f
C18660 VDD.n1597 VSS 0.038523f
C18661 VDD.n1598 VSS 0.058757f
C18662 VDD.n1599 VSS 0.479072f
C18663 VDD.n1600 VSS -0.041546f
C18664 VDD.t1439 VSS 0.090532f
C18665 VDD.t1440 VSS 0.119055f
C18666 VDD.t2396 VSS 0.119055f
C18667 VDD.t664 VSS 0.119055f
C18668 VDD.t670 VSS 0.119055f
C18669 VDD.t672 VSS 0.116575f
C18670 VDD.t666 VSS 0.254852f
C18671 VDD.t28 VSS 0.254852f
C18672 VDD.t18 VSS 0.116575f
C18673 VDD.t22 VSS 0.119055f
C18674 VDD.t26 VSS 0.119055f
C18675 VDD.t3290 VSS 0.119055f
C18676 VDD.t3288 VSS 0.119055f
C18677 VDD.t3289 VSS 0.088051f
C18678 VDD.t2720 VSS 0.532028f
C18679 VDD.t2714 VSS 0.116575f
C18680 VDD.t2722 VSS 0.119055f
C18681 VDD.t2718 VSS 0.119055f
C18682 VDD.t2861 VSS 0.119055f
C18683 VDD.t2860 VSS 0.119055f
C18684 VDD.t2859 VSS 0.090532f
C18685 VDD.t4311 VSS 0.010856f
C18686 VDD.t4272 VSS 0.012354f
C18687 VDD.n1601 VSS 0.038675f
C18688 VDD.t3935 VSS 0.012354f
C18689 VDD.t4313 VSS 0.012354f
C18690 VDD.n1602 VSS 0.040145f
C18691 VDD.n1603 VSS 0.059265f
C18692 VDD.n1604 VSS 0.22487f
C18693 VDD.t2719 VSS 0.012354f
C18694 VDD.t2723 VSS 0.012354f
C18695 VDD.n1605 VSS 0.040938f
C18696 VDD.t2715 VSS 0.012354f
C18697 VDD.t2721 VSS 0.010856f
C18698 VDD.n1606 VSS 0.038523f
C18699 VDD.n1607 VSS 0.058757f
C18700 VDD.n1608 VSS 0.479072f
C18701 VDD.n1609 VSS -0.041546f
C18702 VDD.t2868 VSS 0.088051f
C18703 VDD.t2870 VSS 0.119055f
C18704 VDD.t2869 VSS 0.119055f
C18705 VDD.t4312 VSS 0.119055f
C18706 VDD.t3934 VSS 0.119055f
C18707 VDD.t4271 VSS 0.116575f
C18708 VDD.t4310 VSS 0.254852f
C18709 VDD.t1052 VSS 0.254852f
C18710 VDD.t1046 VSS 0.116575f
C18711 VDD.t1044 VSS 0.119055f
C18712 VDD.t1054 VSS 0.119055f
C18713 VDD.t277 VSS 0.119055f
C18714 VDD.t276 VSS 0.119055f
C18715 VDD.t275 VSS 0.090532f
C18716 VDD.t4161 VSS 0.010856f
C18717 VDD.t4151 VSS 0.012354f
C18718 VDD.n1610 VSS 0.038675f
C18719 VDD.t4157 VSS 0.012354f
C18720 VDD.t4159 VSS 0.012354f
C18721 VDD.n1611 VSS 0.040145f
C18722 VDD.n1612 VSS 0.059265f
C18723 VDD.n1613 VSS 0.22487f
C18724 VDD.t1055 VSS 0.012354f
C18725 VDD.t1045 VSS 0.012354f
C18726 VDD.n1614 VSS 0.040938f
C18727 VDD.t1047 VSS 0.012354f
C18728 VDD.t1053 VSS 0.010856f
C18729 VDD.n1615 VSS 0.038523f
C18730 VDD.n1616 VSS 0.058757f
C18731 VDD.n1617 VSS 0.479072f
C18732 VDD.n1618 VSS -0.041546f
C18733 VDD.t1344 VSS 0.088051f
C18734 VDD.t1346 VSS 0.119055f
C18735 VDD.t1345 VSS 0.119055f
C18736 VDD.t4158 VSS 0.119055f
C18737 VDD.t4156 VSS 0.119055f
C18738 VDD.t4150 VSS 0.116575f
C18739 VDD.t4160 VSS 0.362126f
C18740 VDD.t4032 VSS 0.362126f
C18741 VDD.t4028 VSS 0.116575f
C18742 VDD.t4036 VSS 0.119055f
C18743 VDD.t4034 VSS 0.119055f
C18744 VDD.t1040 VSS 0.119055f
C18745 VDD.t733 VSS 0.119055f
C18746 VDD.t732 VSS 0.090532f
C18747 VDD.n1619 VSS -0.041546f
C18748 VDD.n1620 VSS 0.479072f
C18749 VDD.n1621 VSS 0.22487f
C18750 VDD.n1622 VSS 0.322085f
C18751 VDD.n1623 VSS 0.985447f
C18752 VDD.n1624 VSS 0.837497f
C18753 VDD.n1625 VSS 0.98386f
C18754 VDD.n1626 VSS 0.322085f
C18755 VDD.n1627 VSS 0.22487f
C18756 VDD.t1816 VSS 0.012354f
C18757 VDD.t161 VSS 0.012354f
C18758 VDD.n1628 VSS 0.040938f
C18759 VDD.t157 VSS 0.012354f
C18760 VDD.t151 VSS 0.010856f
C18761 VDD.n1629 VSS 0.038523f
C18762 VDD.n1630 VSS 0.058757f
C18763 VDD.n1631 VSS 0.479072f
C18764 VDD.n1632 VSS -0.041546f
C18765 VDD.t2858 VSS 0.088051f
C18766 VDD.t2649 VSS 0.119055f
C18767 VDD.t2857 VSS 0.119055f
C18768 VDD.t2445 VSS 0.119055f
C18769 VDD.t2447 VSS 0.119055f
C18770 VDD.t2449 VSS 0.116575f
C18771 VDD.t2439 VSS 0.254852f
C18772 VDD.t1287 VSS 0.254852f
C18773 VDD.t1275 VSS 0.116575f
C18774 VDD.t1277 VSS 0.119055f
C18775 VDD.t1279 VSS 0.119055f
C18776 VDD.t1616 VSS 0.119055f
C18777 VDD.t1109 VSS 0.119055f
C18778 VDD.t1615 VSS 0.090532f
C18779 VDD.t833 VSS 0.010856f
C18780 VDD.t831 VSS 0.012354f
C18781 VDD.n1633 VSS 0.038675f
C18782 VDD.t841 VSS 0.012354f
C18783 VDD.t839 VSS 0.012354f
C18784 VDD.n1634 VSS 0.040145f
C18785 VDD.n1635 VSS 0.059265f
C18786 VDD.n1636 VSS 0.22487f
C18787 VDD.t1280 VSS 0.012354f
C18788 VDD.t1278 VSS 0.012354f
C18789 VDD.n1637 VSS 0.040938f
C18790 VDD.t1276 VSS 0.012354f
C18791 VDD.t1288 VSS 0.010856f
C18792 VDD.n1638 VSS 0.038523f
C18793 VDD.n1639 VSS 0.058757f
C18794 VDD.n1640 VSS 0.479072f
C18795 VDD.n1641 VSS -0.041546f
C18796 VDD.t100 VSS 0.088051f
C18797 VDD.t101 VSS 0.119055f
C18798 VDD.t102 VSS 0.119055f
C18799 VDD.t838 VSS 0.119055f
C18800 VDD.t840 VSS 0.119055f
C18801 VDD.t830 VSS 0.116575f
C18802 VDD.t832 VSS 0.362126f
C18803 VDD.t1898 VSS 0.362126f
C18804 VDD.t1902 VSS 0.116575f
C18805 VDD.t1896 VSS 0.119055f
C18806 VDD.t1904 VSS 0.119055f
C18807 VDD.t2024 VSS 0.119055f
C18808 VDD.t2022 VSS 0.119055f
C18809 VDD.t2023 VSS 0.090532f
C18810 VDD.t4015 VSS 0.010856f
C18811 VDD.t4019 VSS 0.012354f
C18812 VDD.n1642 VSS 0.038675f
C18813 VDD.t4013 VSS 0.012354f
C18814 VDD.t4011 VSS 0.012354f
C18815 VDD.n1643 VSS 0.040145f
C18816 VDD.n1644 VSS 0.059265f
C18817 VDD.t1905 VSS 0.012354f
C18818 VDD.t1897 VSS 0.012354f
C18819 VDD.n1645 VSS 0.040938f
C18820 VDD.t1903 VSS 0.012354f
C18821 VDD.t1899 VSS 0.010856f
C18822 VDD.n1646 VSS 0.038523f
C18823 VDD.n1647 VSS 0.058757f
C18824 VDD.n1648 VSS 0.22487f
C18825 VDD.n1649 VSS 0.479072f
C18826 VDD.n1650 VSS -0.041546f
C18827 VDD.t1650 VSS 0.088051f
C18828 VDD.t1651 VSS 0.119055f
C18829 VDD.t1652 VSS 0.119055f
C18830 VDD.t4010 VSS 0.119055f
C18831 VDD.t4012 VSS 0.119055f
C18832 VDD.t4018 VSS 0.116575f
C18833 VDD.t4014 VSS 0.254852f
C18834 VDD.t2014 VSS 0.254852f
C18835 VDD.t2016 VSS 0.116575f
C18836 VDD.t2018 VSS 0.119055f
C18837 VDD.t2008 VSS 0.119055f
C18838 VDD.t1241 VSS 0.119055f
C18839 VDD.t1243 VSS 0.119055f
C18840 VDD.t1242 VSS 0.090532f
C18841 VDD.t2781 VSS 0.010856f
C18842 VDD.t2777 VSS 0.012354f
C18843 VDD.n1651 VSS 0.038675f
C18844 VDD.t2775 VSS 0.012354f
C18845 VDD.t2773 VSS 0.012354f
C18846 VDD.n1652 VSS 0.040145f
C18847 VDD.n1653 VSS 0.059265f
C18848 VDD.n1654 VSS 0.22487f
C18849 VDD.t2009 VSS 0.012354f
C18850 VDD.t2019 VSS 0.012354f
C18851 VDD.n1655 VSS 0.040938f
C18852 VDD.t2017 VSS 0.012354f
C18853 VDD.t2015 VSS 0.010856f
C18854 VDD.n1656 VSS 0.038523f
C18855 VDD.n1657 VSS 0.058757f
C18856 VDD.n1658 VSS 0.479072f
C18857 VDD.n1659 VSS -0.041546f
C18858 VDD.t4307 VSS 0.088051f
C18859 VDD.t4308 VSS 0.119055f
C18860 VDD.t4309 VSS 0.119055f
C18861 VDD.t2772 VSS 0.119055f
C18862 VDD.t2774 VSS 0.119055f
C18863 VDD.t2776 VSS 0.116575f
C18864 VDD.t2780 VSS 0.362126f
C18865 VDD.t1074 VSS 0.362126f
C18866 VDD.t1882 VSS 0.116575f
C18867 VDD.t1884 VSS 0.119055f
C18868 VDD.t1072 VSS 0.119055f
C18869 VDD.t1537 VSS 0.119055f
C18870 VDD.t1538 VSS 0.119055f
C18871 VDD.t1536 VSS 0.090532f
C18872 VDD.t3519 VSS 0.010856f
C18873 VDD.t3515 VSS 0.012354f
C18874 VDD.n1660 VSS 0.038675f
C18875 VDD.t3513 VSS 0.012354f
C18876 VDD.t3523 VSS 0.012354f
C18877 VDD.n1661 VSS 0.040145f
C18878 VDD.n1662 VSS 0.059265f
C18879 VDD.n1663 VSS 0.22487f
C18880 VDD.t1073 VSS 0.012354f
C18881 VDD.t1885 VSS 0.012354f
C18882 VDD.n1664 VSS 0.040938f
C18883 VDD.t1883 VSS 0.012354f
C18884 VDD.t1075 VSS 0.010856f
C18885 VDD.n1665 VSS 0.038523f
C18886 VDD.n1666 VSS 0.058757f
C18887 VDD.n1667 VSS 0.479072f
C18888 VDD.n1668 VSS -0.041546f
C18889 VDD.t2005 VSS 0.088051f
C18890 VDD.t2006 VSS 0.119055f
C18891 VDD.t2007 VSS 0.119055f
C18892 VDD.t3522 VSS 0.119055f
C18893 VDD.t3512 VSS 0.119055f
C18894 VDD.t3514 VSS 0.116575f
C18895 VDD.t3518 VSS 0.254852f
C18896 VDD.t3387 VSS 0.254852f
C18897 VDD.t3389 VSS 0.116575f
C18898 VDD.t3393 VSS 0.119055f
C18899 VDD.t3391 VSS 0.119055f
C18900 VDD.t2734 VSS 0.119055f
C18901 VDD.t2033 VSS 0.119055f
C18902 VDD.t2733 VSS 0.090532f
C18903 VDD.n1669 VSS -0.041546f
C18904 VDD.t3392 VSS 0.012354f
C18905 VDD.t3394 VSS 0.012354f
C18906 VDD.n1670 VSS 0.040938f
C18907 VDD.t3390 VSS 0.012354f
C18908 VDD.t3388 VSS 0.010856f
C18909 VDD.n1671 VSS 0.038523f
C18910 VDD.n1672 VSS 0.058757f
C18911 VDD.n1673 VSS 0.479072f
C18912 VDD.n1674 VSS 0.325106f
C18913 VDD.n1675 VSS 0.705706f
C18914 VDD.n1676 VSS 0.326881f
C18915 VDD.n1677 VSS 0.274887f
C18916 VDD.n1678 VSS 0.092113f
C18917 VDD.t1931 VSS 0.004807f
C18918 VDD.t1943 VSS 0.004807f
C18919 VDD.n1679 VSS 0.010696f
C18920 VDD.n1680 VSS 0.036584f
C18921 VDD.t3396 VSS 0.017474f
C18922 VDD.t3386 VSS 0.004807f
C18923 VDD.t3384 VSS 0.004807f
C18924 VDD.n1681 VSS 0.010696f
C18925 VDD.n1682 VSS 0.097619f
C18926 VDD.n1683 VSS 0.024888f
C18927 VDD.n1684 VSS 0.006536f
C18928 VDD.t3385 VSS 0.049198f
C18929 VDD.t3383 VSS 0.067957f
C18930 VDD.t3395 VSS 0.256608f
C18931 VDD.t3524 VSS 0.256608f
C18932 VDD.t3520 VSS 0.067957f
C18933 VDD.t3516 VSS 0.052737f
C18934 VDD.t3525 VSS 0.017476f
C18935 VDD.t3521 VSS 0.004807f
C18936 VDD.t3517 VSS 0.004807f
C18937 VDD.n1685 VSS 0.010696f
C18938 VDD.n1686 VSS 0.099623f
C18939 VDD.n1687 VSS 0.026083f
C18940 VDD.t1077 VSS 0.017474f
C18941 VDD.t1887 VSS 0.004807f
C18942 VDD.t1079 VSS 0.004807f
C18943 VDD.n1688 VSS 0.010696f
C18944 VDD.n1689 VSS 0.099467f
C18945 VDD.n1690 VSS 0.025249f
C18946 VDD.n1691 VSS 0.006536f
C18947 VDD.t1886 VSS 0.049198f
C18948 VDD.t1078 VSS 0.067957f
C18949 VDD.t1076 VSS 0.324211f
C18950 VDD.t4004 VSS 0.324211f
C18951 VDD.t4002 VSS 0.067957f
C18952 VDD.t4000 VSS 0.052737f
C18953 VDD.t4006 VSS 0.067957f
C18954 VDD.t4008 VSS 0.256608f
C18955 VDD.t2020 VSS 0.256608f
C18956 VDD.t2010 VSS 0.067957f
C18957 VDD.t2012 VSS 0.049198f
C18958 VDD.t2785 VSS 0.017462f
C18959 VDD.n1692 VSS 0.092113f
C18960 VDD.t2783 VSS 0.004807f
C18961 VDD.t2779 VSS 0.004807f
C18962 VDD.n1693 VSS 0.010696f
C18963 VDD.n1694 VSS 0.036584f
C18964 VDD.t2021 VSS 0.017474f
C18965 VDD.t2013 VSS 0.004807f
C18966 VDD.t2011 VSS 0.004807f
C18967 VDD.n1695 VSS 0.010696f
C18968 VDD.n1696 VSS 0.097619f
C18969 VDD.n1697 VSS 0.024888f
C18970 VDD.n1698 VSS 0.006536f
C18971 VDD.t2778 VSS 0.052737f
C18972 VDD.t2782 VSS 0.067957f
C18973 VDD.t2784 VSS 0.176263f
C18974 VDD.t3409 VSS 0.176263f
C18975 VDD.t3411 VSS 0.067957f
C18976 VDD.t3407 VSS 0.049198f
C18977 VDD.n1699 VSS 0.006536f
C18978 VDD.n1700 VSS 0.02587f
C18979 VDD.n1701 VSS 0.040206f
C18980 VDD.n1702 VSS 0.166576f
C18981 VDD.n1703 VSS 0.526294f
C18982 VDD.n1704 VSS 0.98386f
C18983 VDD.n1705 VSS 0.837497f
C18984 VDD.n1706 VSS 0.985447f
C18985 VDD.n1707 VSS 0.848376f
C18986 VDD.n1708 VSS 0.175602f
C18987 VDD.n1709 VSS 0.026083f
C18988 VDD.t284 VSS 0.017474f
C18989 VDD.t294 VSS 0.004807f
C18990 VDD.t296 VSS 0.004807f
C18991 VDD.n1710 VSS 0.010696f
C18992 VDD.n1711 VSS 0.099467f
C18993 VDD.n1712 VSS 0.025249f
C18994 VDD.n1713 VSS 0.006536f
C18995 VDD.t293 VSS 0.049198f
C18996 VDD.t295 VSS 0.067957f
C18997 VDD.t283 VSS 0.324211f
C18998 VDD.t712 VSS 0.324211f
C18999 VDD.t714 VSS 0.067957f
C19000 VDD.t716 VSS 0.052737f
C19001 VDD.t713 VSS 0.017476f
C19002 VDD.t715 VSS 0.004807f
C19003 VDD.t717 VSS 0.004807f
C19004 VDD.n1714 VSS 0.010696f
C19005 VDD.n1715 VSS 0.098224f
C19006 VDD.n1716 VSS 0.040206f
C19007 VDD.t2520 VSS 0.017474f
C19008 VDD.t2516 VSS 0.004807f
C19009 VDD.t2518 VSS 0.004807f
C19010 VDD.n1717 VSS 0.010696f
C19011 VDD.n1718 VSS 0.099162f
C19012 VDD.n1719 VSS 0.02587f
C19013 VDD.n1720 VSS 0.006536f
C19014 VDD.t2515 VSS 0.049198f
C19015 VDD.t2517 VSS 0.067957f
C19016 VDD.t2519 VSS 0.176263f
C19017 VDD.t217 VSS 0.176263f
C19018 VDD.t219 VSS 0.067957f
C19019 VDD.t209 VSS 0.052737f
C19020 VDD.t459 VSS 0.049198f
C19021 VDD.t701 VSS 0.017462f
C19022 VDD.t244 VSS 0.017476f
C19023 VDD.t248 VSS 0.004807f
C19024 VDD.t254 VSS 0.004807f
C19025 VDD.n1721 VSS 0.010696f
C19026 VDD.n1722 VSS 0.099623f
C19027 VDD.t2910 VSS 0.017474f
C19028 VDD.t2916 VSS 0.004807f
C19029 VDD.t2914 VSS 0.004807f
C19030 VDD.n1723 VSS 0.010696f
C19031 VDD.n1724 VSS 0.099467f
C19032 VDD.t461 VSS 0.067957f
C19033 VDD.t449 VSS 0.256608f
C19034 VDD.t243 VSS 0.256608f
C19035 VDD.t247 VSS 0.067957f
C19036 VDD.t253 VSS 0.052737f
C19037 VDD.t4325 VSS 0.049198f
C19038 VDD.t723 VSS 0.017476f
C19039 VDD.t721 VSS 0.004807f
C19040 VDD.t719 VSS 0.004807f
C19041 VDD.n1725 VSS 0.010696f
C19042 VDD.n1726 VSS 0.098224f
C19043 VDD.n1727 VSS 0.342174f
C19044 VDD.n1728 VSS 0.336089f
C19045 VDD.t2562 VSS 0.017462f
C19046 VDD.t497 VSS 0.017474f
C19047 VDD.t2738 VSS 0.004807f
C19048 VDD.t2740 VSS 0.004807f
C19049 VDD.n1729 VSS 0.010696f
C19050 VDD.n1730 VSS 0.097619f
C19051 VDD.t4327 VSS 0.067957f
C19052 VDD.t4329 VSS 0.176263f
C19053 VDD.t2561 VSS 0.176263f
C19054 VDD.t2565 VSS 0.067957f
C19055 VDD.t2563 VSS 0.052737f
C19056 VDD.t1972 VSS 0.454462f
C19057 VDD.t1926 VSS 0.067957f
C19058 VDD.t1932 VSS 0.049198f
C19059 VDD.t1610 VSS 0.017476f
C19060 VDD.t637 VSS 0.004807f
C19061 VDD.t1606 VSS 0.004807f
C19062 VDD.n1731 VSS 0.010696f
C19063 VDD.n1732 VSS 0.099623f
C19064 VDD.n1733 VSS 0.026083f
C19065 VDD.t1973 VSS 0.017474f
C19066 VDD.t1933 VSS 0.004807f
C19067 VDD.t1927 VSS 0.004807f
C19068 VDD.n1734 VSS 0.010696f
C19069 VDD.n1735 VSS 0.099467f
C19070 VDD.n1736 VSS 0.025249f
C19071 VDD.n1737 VSS 0.006536f
C19072 VDD.t1605 VSS 0.052737f
C19073 VDD.t636 VSS 0.067957f
C19074 VDD.t1609 VSS 0.256608f
C19075 VDD.t496 VSS 0.256608f
C19076 VDD.t2739 VSS 0.067957f
C19077 VDD.t2737 VSS 0.049198f
C19078 VDD.n1738 VSS 0.006536f
C19079 VDD.n1739 VSS 0.024888f
C19080 VDD.t2566 VSS 0.004807f
C19081 VDD.t2564 VSS 0.004807f
C19082 VDD.n1740 VSS 0.010696f
C19083 VDD.n1741 VSS 0.036584f
C19084 VDD.n1742 VSS 0.092113f
C19085 VDD.n1743 VSS 0.137976f
C19086 VDD.n1744 VSS 0.167387f
C19087 VDD.n1745 VSS 0.040206f
C19088 VDD.t4330 VSS 0.017474f
C19089 VDD.t4326 VSS 0.004807f
C19090 VDD.t4328 VSS 0.004807f
C19091 VDD.n1746 VSS 0.010696f
C19092 VDD.n1747 VSS 0.099162f
C19093 VDD.n1748 VSS 0.02587f
C19094 VDD.n1749 VSS 0.006536f
C19095 VDD.t718 VSS 0.052737f
C19096 VDD.t720 VSS 0.067957f
C19097 VDD.t722 VSS 0.324211f
C19098 VDD.t2909 VSS 0.324211f
C19099 VDD.t2913 VSS 0.067957f
C19100 VDD.t2915 VSS 0.049198f
C19101 VDD.n1750 VSS 0.006536f
C19102 VDD.n1751 VSS 0.025249f
C19103 VDD.n1752 VSS 0.026083f
C19104 VDD.n1753 VSS 0.174791f
C19105 VDD.n1754 VSS 0.313107f
C19106 VDD.n1755 VSS 0.336089f
C19107 VDD.n1756 VSS 0.137976f
C19108 VDD.n1757 VSS 0.092113f
C19109 VDD.t703 VSS 0.004807f
C19110 VDD.t707 VSS 0.004807f
C19111 VDD.n1758 VSS 0.010696f
C19112 VDD.n1759 VSS 0.036584f
C19113 VDD.t450 VSS 0.017474f
C19114 VDD.t460 VSS 0.004807f
C19115 VDD.t462 VSS 0.004807f
C19116 VDD.n1760 VSS 0.010696f
C19117 VDD.n1761 VSS 0.097619f
C19118 VDD.n1762 VSS 0.024888f
C19119 VDD.n1763 VSS 0.006536f
C19120 VDD.t706 VSS 0.052737f
C19121 VDD.t702 VSS 0.067957f
C19122 VDD.t700 VSS 0.176263f
C19123 VDD.t1082 VSS 0.176263f
C19124 VDD.t563 VSS 0.067957f
C19125 VDD.t1084 VSS 0.049198f
C19126 VDD.t118 VSS 0.017476f
C19127 VDD.t1130 VSS 0.004807f
C19128 VDD.t1132 VSS 0.004807f
C19129 VDD.n1764 VSS 0.010696f
C19130 VDD.n1765 VSS 0.098224f
C19131 VDD.n1766 VSS 0.040206f
C19132 VDD.t1083 VSS 0.017474f
C19133 VDD.t1085 VSS 0.004807f
C19134 VDD.t564 VSS 0.004807f
C19135 VDD.n1767 VSS 0.010696f
C19136 VDD.n1768 VSS 0.099162f
C19137 VDD.n1769 VSS 0.02587f
C19138 VDD.n1770 VSS 0.006536f
C19139 VDD.t1131 VSS 0.052737f
C19140 VDD.t1129 VSS 0.067957f
C19141 VDD.t117 VSS 0.324211f
C19142 VDD.t1336 VSS 0.324211f
C19143 VDD.t1334 VSS 0.067957f
C19144 VDD.t1330 VSS 0.049198f
C19145 VDD.t2315 VSS 0.017476f
C19146 VDD.t2303 VSS 0.004807f
C19147 VDD.t2305 VSS 0.004807f
C19148 VDD.n1771 VSS 0.010696f
C19149 VDD.n1772 VSS 0.099623f
C19150 VDD.n1773 VSS 0.026083f
C19151 VDD.t1337 VSS 0.017474f
C19152 VDD.t1331 VSS 0.004807f
C19153 VDD.t1335 VSS 0.004807f
C19154 VDD.n1774 VSS 0.010696f
C19155 VDD.n1775 VSS 0.099467f
C19156 VDD.n1776 VSS 0.025249f
C19157 VDD.n1777 VSS 0.006536f
C19158 VDD.t2304 VSS 0.052737f
C19159 VDD.t2302 VSS 0.067957f
C19160 VDD.t2314 VSS 0.256608f
C19161 VDD.t4181 VSS 0.256608f
C19162 VDD.t4175 VSS 0.067957f
C19163 VDD.t4173 VSS 0.049198f
C19164 VDD.n1778 VSS 0.006536f
C19165 VDD.n1779 VSS 0.024888f
C19166 VDD.t220 VSS 0.004807f
C19167 VDD.t210 VSS 0.004807f
C19168 VDD.n1780 VSS 0.010696f
C19169 VDD.n1781 VSS 0.036584f
C19170 VDD.n1782 VSS 0.092113f
C19171 VDD.n1783 VSS 0.137976f
C19172 VDD.n1784 VSS 0.336089f
C19173 VDD.n1785 VSS 0.342174f
C19174 VDD.n1786 VSS 0.334821f
C19175 VDD.n1787 VSS 0.22487f
C19176 VDD.t4178 VSS 0.012354f
C19177 VDD.t4184 VSS 0.012354f
C19178 VDD.n1788 VSS 0.040938f
C19179 VDD.t4172 VSS 0.012354f
C19180 VDD.t4180 VSS 0.010856f
C19181 VDD.n1789 VSS 0.038523f
C19182 VDD.n1790 VSS 0.058757f
C19183 VDD.n1791 VSS 0.479072f
C19184 VDD.n1792 VSS -0.041546f
C19185 VDD.t1152 VSS 0.090532f
C19186 VDD.t1151 VSS 0.119055f
C19187 VDD.t986 VSS 0.119055f
C19188 VDD.t4177 VSS 0.119055f
C19189 VDD.t4183 VSS 0.119055f
C19190 VDD.t4171 VSS 0.116575f
C19191 VDD.t4179 VSS 0.254852f
C19192 VDD.t2306 VSS 0.254852f
C19193 VDD.t2310 VSS 0.116575f
C19194 VDD.t2308 VSS 0.119055f
C19195 VDD.t2312 VSS 0.119055f
C19196 VDD.t1525 VSS 0.119055f
C19197 VDD.t1526 VSS 0.119055f
C19198 VDD.t1527 VSS 0.088051f
C19199 VDD.t2395 VSS 0.119055f
C19200 VDD.t2394 VSS 0.119055f
C19201 VDD.t251 VSS 0.119055f
C19202 VDD.t249 VSS 0.119055f
C19203 VDD.t245 VSS 0.116575f
C19204 VDD.t255 VSS 0.254852f
C19205 VDD.t453 VSS 0.254852f
C19206 VDD.t457 VSS 0.116575f
C19207 VDD.t455 VSS 0.119055f
C19208 VDD.t451 VSS 0.119055f
C19209 VDD.t2268 VSS 0.119055f
C19210 VDD.t2269 VSS 0.119055f
C19211 VDD.t2270 VSS 0.090532f
C19212 VDD.t3989 VSS 0.010856f
C19213 VDD.t705 VSS 0.012354f
C19214 VDD.n1793 VSS 0.038675f
C19215 VDD.t709 VSS 0.012354f
C19216 VDD.t711 VSS 0.012354f
C19217 VDD.n1794 VSS 0.040145f
C19218 VDD.n1795 VSS 0.059265f
C19219 VDD.t452 VSS 0.012354f
C19220 VDD.t456 VSS 0.012354f
C19221 VDD.n1796 VSS 0.040938f
C19222 VDD.t458 VSS 0.012354f
C19223 VDD.t454 VSS 0.010856f
C19224 VDD.n1797 VSS 0.038523f
C19225 VDD.n1798 VSS 0.058757f
C19226 VDD.n1799 VSS 0.22487f
C19227 VDD.n1800 VSS 0.479072f
C19228 VDD.n1801 VSS -0.041546f
C19229 VDD.t929 VSS 0.088051f
C19230 VDD.t927 VSS 0.119055f
C19231 VDD.t928 VSS 0.119055f
C19232 VDD.t710 VSS 0.119055f
C19233 VDD.t708 VSS 0.119055f
C19234 VDD.t704 VSS 0.116575f
C19235 VDD.t3988 VSS 0.362126f
C19236 VDD.t1342 VSS 0.362126f
C19237 VDD.t1338 VSS 0.116575f
C19238 VDD.t1340 VSS 0.119055f
C19239 VDD.t1332 VSS 0.119055f
C19240 VDD.t4162 VSS 0.119055f
C19241 VDD.t4164 VSS 0.119055f
C19242 VDD.t4163 VSS 0.090532f
C19243 VDD.n1802 VSS -0.041546f
C19244 VDD.n1803 VSS 0.479072f
C19245 VDD.n1804 VSS 0.22487f
C19246 VDD.n1805 VSS 0.293085f
C19247 VDD.n1806 VSS 0.278804f
C19248 VDD.n1807 VSS 0.827977f
C19249 VDD.n1808 VSS 0.985447f
C19250 VDD.n1809 VSS 0.837497f
C19251 VDD.n1810 VSS 0.98386f
C19252 VDD.n1811 VSS 0.526294f
C19253 VDD.n1812 VSS 0.177022f
C19254 VDD.n1813 VSS 0.026083f
C19255 VDD.t1893 VSS 0.017474f
C19256 VDD.t1901 VSS 0.004807f
C19257 VDD.t1895 VSS 0.004807f
C19258 VDD.n1814 VSS 0.010696f
C19259 VDD.n1815 VSS 0.099467f
C19260 VDD.n1816 VSS 0.025249f
C19261 VDD.n1817 VSS 0.006536f
C19262 VDD.t1900 VSS 0.049198f
C19263 VDD.t1894 VSS 0.067957f
C19264 VDD.t1892 VSS 0.324211f
C19265 VDD.t1695 VSS 0.324211f
C19266 VDD.t1693 VSS 0.067957f
C19267 VDD.t1697 VSS 0.052737f
C19268 VDD.t1696 VSS 0.017476f
C19269 VDD.t1694 VSS 0.004807f
C19270 VDD.t1698 VSS 0.004807f
C19271 VDD.n1818 VSS 0.010696f
C19272 VDD.n1819 VSS 0.098224f
C19273 VDD.n1820 VSS 0.040206f
C19274 VDD.t1465 VSS 0.017474f
C19275 VDD.t1467 VSS 0.004807f
C19276 VDD.t1469 VSS 0.004807f
C19277 VDD.n1821 VSS 0.010696f
C19278 VDD.n1822 VSS 0.099162f
C19279 VDD.n1823 VSS 0.02587f
C19280 VDD.n1824 VSS 0.006536f
C19281 VDD.t1466 VSS 0.049198f
C19282 VDD.t1468 VSS 0.067957f
C19283 VDD.t1464 VSS 0.176263f
C19284 VDD.t836 VSS 0.176263f
C19285 VDD.t834 VSS 0.067957f
C19286 VDD.t842 VSS 0.052737f
C19287 VDD.t2441 VSS 0.067957f
C19288 VDD.t2443 VSS 0.256608f
C19289 VDD.t1283 VSS 0.256608f
C19290 VDD.t1281 VSS 0.067957f
C19291 VDD.t1285 VSS 0.049198f
C19292 VDD.n1825 VSS 0.006536f
C19293 VDD.n1826 VSS 0.024888f
C19294 VDD.t835 VSS 0.004807f
C19295 VDD.t843 VSS 0.004807f
C19296 VDD.n1827 VSS 0.010696f
C19297 VDD.n1828 VSS 0.036584f
C19298 VDD.n1829 VSS 0.092113f
C19299 VDD.n1830 VSS 0.137976f
C19300 VDD.n1831 VSS 0.326881f
C19301 VDD.n1832 VSS 0.174791f
C19302 VDD.n1833 VSS 0.026083f
C19303 VDD.t153 VSS 0.017474f
C19304 VDD.t155 VSS 0.004807f
C19305 VDD.t159 VSS 0.004807f
C19306 VDD.n1834 VSS 0.010696f
C19307 VDD.n1835 VSS 0.099467f
C19308 VDD.n1836 VSS 0.025249f
C19309 VDD.n1837 VSS 0.006536f
C19310 VDD.t154 VSS 0.049198f
C19311 VDD.t158 VSS 0.067957f
C19312 VDD.t152 VSS 0.324211f
C19313 VDD.t2074 VSS 0.324211f
C19314 VDD.t2070 VSS 0.067957f
C19315 VDD.t2072 VSS 0.052737f
C19316 VDD.t942 VSS 0.067957f
C19317 VDD.t944 VSS 0.176263f
C19318 VDD.t965 VSS 0.176263f
C19319 VDD.t967 VSS 0.067957f
C19320 VDD.t969 VSS 0.049198f
C19321 VDD.n1838 VSS 0.006536f
C19322 VDD.n1839 VSS 0.02587f
C19323 VDD.n1840 VSS 0.040206f
C19324 VDD.n1841 VSS 0.167387f
C19325 VDD.n1842 VSS 0.137976f
C19326 VDD.n1843 VSS 0.092113f
C19327 VDD.t943 VSS 0.004807f
C19328 VDD.t947 VSS 0.004807f
C19329 VDD.n1844 VSS 0.010696f
C19330 VDD.n1845 VSS 0.036584f
C19331 VDD.t3660 VSS 0.017474f
C19332 VDD.t3664 VSS 0.004807f
C19333 VDD.t3662 VSS 0.004807f
C19334 VDD.n1846 VSS 0.010696f
C19335 VDD.n1847 VSS 0.097619f
C19336 VDD.n1848 VSS 0.024888f
C19337 VDD.n1849 VSS 0.006536f
C19338 VDD.t3663 VSS 0.049198f
C19339 VDD.t3661 VSS 0.067957f
C19340 VDD.t3659 VSS 0.256608f
C19341 VDD.t3322 VSS 0.256608f
C19342 VDD.t3320 VSS 0.067957f
C19343 VDD.t3314 VSS 0.052737f
C19344 VDD.t4052 VSS 0.454462f
C19345 VDD.t4056 VSS 0.067957f
C19346 VDD.t4058 VSS 0.049198f
C19347 VDD.n1850 VSS 0.006536f
C19348 VDD.n1851 VSS 0.025249f
C19349 VDD.n1852 VSS 0.026083f
C19350 VDD.n1853 VSS 0.186353f
C19351 VDD.n1854 VSS 0.277926f
C19352 VDD.t1353 VSS 0.004807f
C19353 VDD.t1357 VSS 0.004807f
C19354 VDD.n1855 VSS 0.010736f
C19355 VDD.t1355 VSS 0.017466f
C19356 VDD.n1856 VSS 0.054891f
C19357 VDD.t1352 VSS 0.109586f
C19358 VDD.t1356 VSS 0.053772f
C19359 VDD.t828 VSS 0.090299f
C19360 VDD.t826 VSS 0.044589f
C19361 VDD.t829 VSS 0.004807f
C19362 VDD.t827 VSS 0.004807f
C19363 VDD.n1857 VSS 0.010736f
C19364 VDD.t825 VSS 0.017466f
C19365 VDD.n1858 VSS 0.054891f
C19366 VDD.n1859 VSS 0.054877f
C19367 VDD.t824 VSS 0.095016f
C19368 VDD.t678 VSS 0.42081f
C19369 VDD.t676 VSS 0.206484f
C19370 VDD.t674 VSS 0.192109f
C19371 VDD.t1571 VSS 0.088326f
C19372 VDD.t1569 VSS 0.041419f
C19373 VDD.t1573 VSS 0.089823f
C19374 VDD.t3488 VSS 0.117695f
C19375 VDD.t3486 VSS 0.055923f
C19376 VDD.t3489 VSS 0.004807f
C19377 VDD.t3487 VSS 0.004807f
C19378 VDD.n1860 VSS 0.010736f
C19379 VDD.t3485 VSS 0.017466f
C19380 VDD.n1861 VSS 0.054891f
C19381 VDD.n1862 VSS 0.259532f
C19382 VDD.t2638 VSS 0.004807f
C19383 VDD.t2637 VSS 0.004807f
C19384 VDD.n1863 VSS 0.010736f
C19385 VDD.t2636 VSS 0.017466f
C19386 VDD.n1864 VSS 0.054891f
C19387 VDD.t2384 VSS 0.004807f
C19388 VDD.t2386 VSS 0.004807f
C19389 VDD.n1865 VSS 0.010736f
C19390 VDD.t2385 VSS 0.017466f
C19391 VDD.n1866 VSS 0.054891f
C19392 VDD.n1867 VSS 0.016863f
C19393 VDD.t679 VSS 0.004807f
C19394 VDD.t677 VSS 0.004807f
C19395 VDD.n1868 VSS 0.010736f
C19396 VDD.t675 VSS 0.017466f
C19397 VDD.n1869 VSS 0.054891f
C19398 VDD.n1870 VSS 0.016863f
C19399 VDD.t3483 VSS 0.004807f
C19400 VDD.t3482 VSS 0.004807f
C19401 VDD.n1871 VSS 0.010736f
C19402 VDD.t3481 VSS 0.017466f
C19403 VDD.n1872 VSS 0.054891f
C19404 VDD.n1873 VSS 0.178625f
C19405 VDD.n1874 VSS 0.24945f
C19406 VDD.n1875 VSS 0.016863f
C19407 VDD.n1876 VSS 0.423791f
C19408 VDD.n1877 VSS 0.016863f
C19409 VDD.n1878 VSS 0.252735f
C19410 VDD.t1572 VSS 0.004807f
C19411 VDD.t1570 VSS 0.004807f
C19412 VDD.n1879 VSS 0.010736f
C19413 VDD.t1574 VSS 0.017466f
C19414 VDD.n1880 VSS 0.054891f
C19415 VDD.n1881 VSS 0.050916f
C19416 VDD.n1882 VSS 0.404067f
C19417 VDD.n1883 VSS 0.056662f
C19418 VDD.t3484 VSS 0.129226f
C19419 VDD.n1884 VSS 0.105853f
C19420 VDD.n1885 VSS 0.149767f
C19421 VDD.t1354 VSS 0.121592f
C19422 VDD.n1886 VSS 0.058448f
C19423 VDD.n1887 VSS 0.575022f
C19424 VDD.t1025 VSS 0.017474f
C19425 VDD.t998 VSS 0.004807f
C19426 VDD.t1020 VSS 0.004807f
C19427 VDD.n1888 VSS 0.010696f
C19428 VDD.n1889 VSS 0.097039f
C19429 VDD.n1890 VSS 0.064426f
C19430 VDD.n1891 VSS 0.457559f
C19431 VDD.t4240 VSS 0.017474f
C19432 VDD.t4189 VSS 0.004807f
C19433 VDD.t4209 VSS 0.004807f
C19434 VDD.n1892 VSS 0.010696f
C19435 VDD.n1893 VSS 0.09735f
C19436 VDD.t2321 VSS 0.017474f
C19437 VDD.t2365 VSS 0.004807f
C19438 VDD.t2371 VSS 0.004807f
C19439 VDD.n1894 VSS 0.010696f
C19440 VDD.n1895 VSS 0.097619f
C19441 VDD.t2225 VSS 0.094682f
C19442 VDD.t2238 VSS 0.056456f
C19443 VDD.t1661 VSS 0.043813f
C19444 VDD.t2226 VSS 0.017474f
C19445 VDD.t2239 VSS 0.004807f
C19446 VDD.t1662 VSS 0.004807f
C19447 VDD.n1896 VSS 0.010696f
C19448 VDD.n1897 VSS 0.09764f
C19449 VDD.n1898 VSS 0.012276f
C19450 VDD.n1899 VSS 7.86e-19
C19451 VDD.t997 VSS 0.040872f
C19452 VDD.t1019 VSS 0.057424f
C19453 VDD.t1024 VSS 0.235213f
C19454 VDD.t4239 VSS 0.235803f
C19455 VDD.t4188 VSS 0.056456f
C19456 VDD.t4208 VSS 0.043813f
C19457 VDD.t2157 VSS 0.040872f
C19458 VDD.t4117 VSS 0.017474f
C19459 VDD.t4067 VSS 0.004807f
C19460 VDD.t4071 VSS 0.004807f
C19461 VDD.n1900 VSS 0.010696f
C19462 VDD.n1901 VSS 0.09764f
C19463 VDD.n1902 VSS 0.486739f
C19464 VDD.t1634 VSS 0.017474f
C19465 VDD.t1641 VSS 0.004807f
C19466 VDD.t2198 VSS 0.004807f
C19467 VDD.n1903 VSS 0.010696f
C19468 VDD.n1904 VSS 0.09764f
C19469 VDD.t2162 VSS 0.057482f
C19470 VDD.t2126 VSS 0.23847f
C19471 VDD.t1633 VSS 0.238735f
C19472 VDD.t1640 VSS 0.056456f
C19473 VDD.t2197 VSS 0.043813f
C19474 VDD.t3543 VSS 0.040872f
C19475 VDD.t2831 VSS 0.017474f
C19476 VDD.t2833 VSS 0.004807f
C19477 VDD.t2820 VSS 0.004807f
C19478 VDD.n1905 VSS 0.010696f
C19479 VDD.n1906 VSS 0.09764f
C19480 VDD.t2301 VSS 0.017474f
C19481 VDD.t3420 VSS 0.004807f
C19482 VDD.t3435 VSS 0.004807f
C19483 VDD.n1907 VSS 0.010696f
C19484 VDD.n1908 VSS 0.09764f
C19485 VDD.t3556 VSS 0.056456f
C19486 VDD.t3568 VSS 0.271991f
C19487 VDD.t2300 VSS 0.271991f
C19488 VDD.t3419 VSS 0.056456f
C19489 VDD.t3434 VSS 0.043813f
C19490 VDD.t1402 VSS 0.094682f
C19491 VDD.t1178 VSS 0.056456f
C19492 VDD.t1414 VSS 0.040872f
C19493 VDD.n1909 VSS 7.86e-19
C19494 VDD.n1910 VSS 0.01242f
C19495 VDD.t1403 VSS 0.017474f
C19496 VDD.t1415 VSS 0.004807f
C19497 VDD.t1179 VSS 0.004807f
C19498 VDD.n1911 VSS 0.010696f
C19499 VDD.n1912 VSS 0.096895f
C19500 VDD.n1913 VSS 0.073583f
C19501 VDD.n1914 VSS 0.876375f
C19502 VDD.t3569 VSS 0.017474f
C19503 VDD.t3544 VSS 0.004807f
C19504 VDD.t3557 VSS 0.004807f
C19505 VDD.n1915 VSS 0.010696f
C19506 VDD.n1916 VSS 0.096315f
C19507 VDD.n1917 VSS 0.06611f
C19508 VDD.n1918 VSS 0.013f
C19509 VDD.n1919 VSS 7.86e-19
C19510 VDD.t2819 VSS 0.043813f
C19511 VDD.t2832 VSS 0.056456f
C19512 VDD.t2830 VSS 0.270505f
C19513 VDD.t889 VSS 0.270006f
C19514 VDD.t3974 VSS 0.057424f
C19515 VDD.t903 VSS 0.040872f
C19516 VDD.t398 VSS 0.017474f
C19517 VDD.t382 VSS 0.004807f
C19518 VDD.t394 VSS 0.004807f
C19519 VDD.n1920 VSS 0.010696f
C19520 VDD.n1921 VSS 0.09764f
C19521 VDD.t890 VSS 0.017474f
C19522 VDD.t904 VSS 0.004807f
C19523 VDD.t3975 VSS 0.004807f
C19524 VDD.n1922 VSS 0.010696f
C19525 VDD.n1923 VSS 0.097185f
C19526 VDD.n1924 VSS 0.067245f
C19527 VDD.n1925 VSS 0.01213f
C19528 VDD.n1926 VSS 7.86e-19
C19529 VDD.t393 VSS 0.043813f
C19530 VDD.t381 VSS 0.056456f
C19531 VDD.t397 VSS 0.248629f
C19532 VDD.t3592 VSS 0.257948f
C19533 VDD.t3613 VSS 0.059127f
C19534 VDD.t3600 VSS 0.040872f
C19535 VDD.n1927 VSS 7.86e-19
C19536 VDD.n1928 VSS 0.01271f
C19537 VDD.t3593 VSS 0.017474f
C19538 VDD.t3601 VSS 0.004807f
C19539 VDD.t3614 VSS 0.004807f
C19540 VDD.n1929 VSS 0.010696f
C19541 VDD.n1930 VSS 0.096605f
C19542 VDD.n1931 VSS 0.063324f
C19543 VDD.n1932 VSS 0.465658f
C19544 VDD.n1933 VSS 0.45058f
C19545 VDD.t2127 VSS 0.017474f
C19546 VDD.t2158 VSS 0.004807f
C19547 VDD.t2163 VSS 0.004807f
C19548 VDD.n1934 VSS 0.010696f
C19549 VDD.n1935 VSS 0.096605f
C19550 VDD.n1936 VSS 0.063071f
C19551 VDD.n1937 VSS 0.01271f
C19552 VDD.n1938 VSS 7.86e-19
C19553 VDD.t4070 VSS 0.043813f
C19554 VDD.t4066 VSS 0.056456f
C19555 VDD.t4116 VSS 0.219572f
C19556 VDD.t2592 VSS 0.223466f
C19557 VDD.t485 VSS 0.058219f
C19558 VDD.t481 VSS 0.040872f
C19559 VDD.t258 VSS 0.017474f
C19560 VDD.t520 VSS 0.004807f
C19561 VDD.t532 VSS 0.004807f
C19562 VDD.n1939 VSS 0.010696f
C19563 VDD.n1940 VSS 0.09764f
C19564 VDD.t2593 VSS 0.017474f
C19565 VDD.t482 VSS 0.004807f
C19566 VDD.t486 VSS 0.004807f
C19567 VDD.n1941 VSS 0.010696f
C19568 VDD.n1942 VSS 0.09588f
C19569 VDD.n1943 VSS 0.062944f
C19570 VDD.n1944 VSS 0.013435f
C19571 VDD.n1945 VSS 7.86e-19
C19572 VDD.t531 VSS 0.043813f
C19573 VDD.t519 VSS 0.056456f
C19574 VDD.t257 VSS 0.24522f
C19575 VDD.t2320 VSS 0.245934f
C19576 VDD.t2370 VSS 0.057651f
C19577 VDD.t2364 VSS 0.040872f
C19578 VDD.n1946 VSS 7.86e-19
C19579 VDD.n1947 VSS 0.024888f
C19580 VDD.n1948 VSS 0.063796f
C19581 VDD.n1949 VSS 0.338659f
C19582 VDD.n1950 VSS 0.981836f
C19583 VDD.n1951 VSS 1.08047f
C19584 VDD.n1952 VSS 0.030311f
C19585 VDD.t1653 VSS 0.126462f
C19586 VDD.t1654 VSS 0.075406f
C19587 VDD.t1671 VSS 0.075406f
C19588 VDD.t1676 VSS 0.075406f
C19589 VDD.t2233 VSS 0.075406f
C19590 VDD.t587 VSS 0.075406f
C19591 VDD.t589 VSS 0.075406f
C19592 VDD.t1006 VSS 0.058518f
C19593 VDD.t1030 VSS 0.126462f
C19594 VDD.t1009 VSS 0.05459f
C19595 VDD.n1953 VSS 2.52e-19
C19596 VDD.t588 VSS 0.00575f
C19597 VDD.t590 VSS 0.00575f
C19598 VDD.n1954 VSS 0.0115f
C19599 VDD.n1955 VSS 0.012479f
C19600 VDD.t1007 VSS 0.00575f
C19601 VDD.t1010 VSS 0.00575f
C19602 VDD.n1956 VSS 0.0115f
C19603 VDD.n1957 VSS 0.007448f
C19604 VDD.n1958 VSS 0.076419f
C19605 VDD.t1031 VSS 0.01978f
C19606 VDD.n1959 VSS 0.014195f
C19607 VDD.n1960 VSS -0.012705f
C19608 VDD.n1961 VSS 0.360694f
C19609 VDD.n1962 VSS 0.58185f
C19610 VDD.t4197 VSS 0.012354f
C19611 VDD.t4215 VSS 0.012354f
C19612 VDD.n1963 VSS 0.040118f
C19613 VDD.t4195 VSS 0.010856f
C19614 VDD.t4231 VSS 0.012354f
C19615 VDD.n1964 VSS 0.038648f
C19616 VDD.n1965 VSS 0.059315f
C19617 VDD.t1672 VSS 0.189904f
C19618 VDD.t1657 VSS 0.115167f
C19619 VDD.t1659 VSS 0.117618f
C19620 VDD.t1679 VSS 0.117618f
C19621 VDD.t1149 VSS 0.117618f
C19622 VDD.t1150 VSS 0.117618f
C19623 VDD.t1148 VSS 0.086988f
C19624 VDD.t1660 VSS 0.012354f
C19625 VDD.t1680 VSS 0.012354f
C19626 VDD.n1966 VSS 0.040118f
C19627 VDD.t1673 VSS 0.010856f
C19628 VDD.t1658 VSS 0.012354f
C19629 VDD.n1967 VSS 0.038648f
C19630 VDD.n1968 VSS 0.059315f
C19631 VDD.t988 VSS 0.012354f
C19632 VDD.t596 VSS 0.010856f
C19633 VDD.n1969 VSS 0.038523f
C19634 VDD.t1038 VSS 0.012354f
C19635 VDD.t592 VSS 0.012354f
C19636 VDD.n1970 VSS 0.040938f
C19637 VDD.n1971 VSS 0.058757f
C19638 VDD.n1972 VSS 0.479077f
C19639 VDD.n1973 VSS -0.042265f
C19640 VDD.t3690 VSS 0.089438f
C19641 VDD.t3692 VSS 0.117618f
C19642 VDD.t3687 VSS 0.117618f
C19643 VDD.t1037 VSS 0.117618f
C19644 VDD.t591 VSS 0.117618f
C19645 VDD.t987 VSS 0.115167f
C19646 VDD.t595 VSS 1.02168f
C19647 VDD.t4194 VSS 1.02235f
C19648 VDD.t4230 VSS 0.115423f
C19649 VDD.t4196 VSS 0.117879f
C19650 VDD.t4214 VSS 0.117879f
C19651 VDD.t1303 VSS 0.117879f
C19652 VDD.t1304 VSS 0.117879f
C19653 VDD.t1305 VSS 0.087181f
C19654 VDD.t3452 VSS 0.089637f
C19655 VDD.t4078 VSS 0.012354f
C19656 VDD.t4090 VSS 0.012354f
C19657 VDD.n1974 VSS 0.040118f
C19658 VDD.t4074 VSS 0.010856f
C19659 VDD.t4120 VSS 0.012354f
C19660 VDD.n1975 VSS 0.038648f
C19661 VDD.n1976 VSS 0.059315f
C19662 VDD.t2181 VSS 0.012354f
C19663 VDD.t2154 VSS 0.010856f
C19664 VDD.n1977 VSS 0.038523f
C19665 VDD.t2133 VSS 0.012354f
C19666 VDD.t2152 VSS 0.012354f
C19667 VDD.n1978 VSS 0.040938f
C19668 VDD.n1979 VSS 0.058757f
C19669 VDD.n1980 VSS 0.556637f
C19670 VDD.t2196 VSS 0.012354f
C19671 VDD.t1632 VSS 0.012354f
C19672 VDD.n1981 VSS 0.040118f
C19673 VDD.t2200 VSS 0.010856f
C19674 VDD.t2194 VSS 0.012354f
C19675 VDD.n1982 VSS 0.038648f
C19676 VDD.n1983 VSS 0.059315f
C19677 VDD.t42 VSS 0.117879f
C19678 VDD.t3490 VSS 0.117879f
C19679 VDD.t2132 VSS 0.117879f
C19680 VDD.t2151 VSS 0.117879f
C19681 VDD.t2180 VSS 0.115423f
C19682 VDD.t2153 VSS 0.992821f
C19683 VDD.t2199 VSS 0.992821f
C19684 VDD.t2193 VSS 0.115423f
C19685 VDD.t2195 VSS 0.117879f
C19686 VDD.t1631 VSS 0.117879f
C19687 VDD.t627 VSS 0.117879f
C19688 VDD.t628 VSS 0.117879f
C19689 VDD.t629 VSS 0.087181f
C19690 VDD.t1828 VSS 0.089637f
C19691 VDD.t2813 VSS 0.012354f
C19692 VDD.t2815 VSS 0.012354f
C19693 VDD.n1984 VSS 0.040118f
C19694 VDD.t2844 VSS 0.010856f
C19695 VDD.t2826 VSS 0.012354f
C19696 VDD.n1985 VSS 0.038648f
C19697 VDD.n1986 VSS 0.059315f
C19698 VDD.t3549 VSS 0.012354f
C19699 VDD.t3540 VSS 0.010856f
C19700 VDD.n1987 VSS 0.038523f
C19701 VDD.t3563 VSS 0.012354f
C19702 VDD.t3538 VSS 0.012354f
C19703 VDD.n1988 VSS 0.040938f
C19704 VDD.n1989 VSS 0.058757f
C19705 VDD.t2291 VSS 0.012354f
C19706 VDD.t2297 VSS 0.012354f
C19707 VDD.n1990 VSS 0.040118f
C19708 VDD.t2289 VSS 0.010856f
C19709 VDD.t3443 VSS 0.012354f
C19710 VDD.n1991 VSS 0.038648f
C19711 VDD.n1992 VSS 0.059315f
C19712 VDD.t1397 VSS 0.012354f
C19713 VDD.t1181 VSS 0.010856f
C19714 VDD.n1993 VSS 0.038523f
C19715 VDD.t1413 VSS 0.012354f
C19716 VDD.t1177 VSS 0.012354f
C19717 VDD.n1994 VSS 0.040938f
C19718 VDD.n1995 VSS 0.058757f
C19719 VDD.t1829 VSS 0.117879f
C19720 VDD.t1830 VSS 0.117879f
C19721 VDD.t3562 VSS 0.117879f
C19722 VDD.t3537 VSS 0.117879f
C19723 VDD.t3548 VSS 0.115423f
C19724 VDD.t3539 VSS 0.902282f
C19725 VDD.t2288 VSS 0.901611f
C19726 VDD.t3442 VSS 0.115167f
C19727 VDD.t2290 VSS 0.117618f
C19728 VDD.t2296 VSS 0.117618f
C19729 VDD.t1594 VSS 0.117618f
C19730 VDD.t1595 VSS 0.117618f
C19731 VDD.t1596 VSS 0.086988f
C19732 VDD.t1180 VSS 0.189904f
C19733 VDD.t1396 VSS 0.115167f
C19734 VDD.t1176 VSS 0.117618f
C19735 VDD.t1412 VSS 0.117618f
C19736 VDD.t973 VSS 0.117618f
C19737 VDD.t972 VSS 0.117618f
C19738 VDD.t971 VSS 0.089438f
C19739 VDD.n1996 VSS -0.042265f
C19740 VDD.n1997 VSS 0.479077f
C19741 VDD.n1998 VSS 0.512919f
C19742 VDD.n1999 VSS 0.700061f
C19743 VDD.n2000 VSS 0.22487f
C19744 VDD.n2001 VSS 0.479077f
C19745 VDD.n2002 VSS -0.042134f
C19746 VDD.t2641 VSS 0.087181f
C19747 VDD.t2640 VSS 0.117879f
C19748 VDD.t2639 VSS 0.117879f
C19749 VDD.t2814 VSS 0.117879f
C19750 VDD.t2812 VSS 0.117879f
C19751 VDD.t2825 VSS 0.115423f
C19752 VDD.t2843 VSS 0.895419f
C19753 VDD.t897 VSS 0.895419f
C19754 VDD.t3968 VSS 0.115423f
C19755 VDD.t893 VSS 0.117879f
C19756 VDD.t3979 VSS 0.117879f
C19757 VDD.t1835 VSS 0.117879f
C19758 VDD.t1459 VSS 0.117879f
C19759 VDD.t3291 VSS 0.089637f
C19760 VDD.t384 VSS 0.012354f
C19761 VDD.t386 VSS 0.012354f
C19762 VDD.n2003 VSS 0.040118f
C19763 VDD.t377 VSS 0.010856f
C19764 VDD.t402 VSS 0.012354f
C19765 VDD.n2004 VSS 0.038648f
C19766 VDD.n2005 VSS 0.059315f
C19767 VDD.t3969 VSS 0.012354f
C19768 VDD.t898 VSS 0.010856f
C19769 VDD.n2006 VSS 0.038523f
C19770 VDD.t3980 VSS 0.012354f
C19771 VDD.t894 VSS 0.012354f
C19772 VDD.n2007 VSS 0.040938f
C19773 VDD.n2008 VSS 0.058757f
C19774 VDD.n2009 VSS 0.22487f
C19775 VDD.n2010 VSS 0.479077f
C19776 VDD.n2011 VSS -0.042134f
C19777 VDD.t1819 VSS 0.087181f
C19778 VDD.t1818 VSS 0.117879f
C19779 VDD.t1817 VSS 0.117879f
C19780 VDD.t385 VSS 0.117879f
C19781 VDD.t383 VSS 0.117879f
C19782 VDD.t401 VSS 0.115423f
C19783 VDD.t376 VSS 0.910121f
C19784 VDD.t3579 VSS 0.910121f
C19785 VDD.t3584 VSS 0.115423f
C19786 VDD.t3618 VSS 0.117879f
C19787 VDD.t3604 VSS 0.117879f
C19788 VDD.t3526 VSS 0.117879f
C19789 VDD.t4165 VSS 0.117879f
C19790 VDD.t4166 VSS 0.089637f
C19791 VDD.n2012 VSS -0.042134f
C19792 VDD.t3585 VSS 0.012354f
C19793 VDD.t3580 VSS 0.010856f
C19794 VDD.n2013 VSS 0.038523f
C19795 VDD.t3605 VSS 0.012354f
C19796 VDD.t3619 VSS 0.012354f
C19797 VDD.n2014 VSS 0.040938f
C19798 VDD.n2015 VSS 0.058757f
C19799 VDD.n2016 VSS 0.479077f
C19800 VDD.n2017 VSS 0.22487f
C19801 VDD.n2018 VSS 0.570273f
C19802 VDD.n2019 VSS 0.565642f
C19803 VDD.n2020 VSS 0.22487f
C19804 VDD.n2021 VSS 0.479077f
C19805 VDD.n2022 VSS -0.042134f
C19806 VDD.t2762 VSS 0.087181f
C19807 VDD.t2764 VSS 0.117879f
C19808 VDD.t2763 VSS 0.117879f
C19809 VDD.t4089 VSS 0.117879f
C19810 VDD.t4077 VSS 0.117879f
C19811 VDD.t4119 VSS 0.115423f
C19812 VDD.t4073 VSS 0.877041f
C19813 VDD.t479 VSS 0.877041f
C19814 VDD.t483 VSS 0.115423f
C19815 VDD.t2609 VSS 0.117879f
C19816 VDD.t2588 VSS 0.117879f
C19817 VDD.t2871 VSS 0.117879f
C19818 VDD.t1237 VSS 0.117879f
C19819 VDD.t1236 VSS 0.089637f
C19820 VDD.t538 VSS 0.012354f
C19821 VDD.t540 VSS 0.012354f
C19822 VDD.n2023 VSS 0.040118f
C19823 VDD.t270 VSS 0.010856f
C19824 VDD.t526 VSS 0.012354f
C19825 VDD.n2024 VSS 0.038648f
C19826 VDD.n2025 VSS 0.059315f
C19827 VDD.t484 VSS 0.012354f
C19828 VDD.t480 VSS 0.010856f
C19829 VDD.n2026 VSS 0.038523f
C19830 VDD.t2589 VSS 0.012354f
C19831 VDD.t2610 VSS 0.012354f
C19832 VDD.n2027 VSS 0.040938f
C19833 VDD.n2028 VSS 0.058757f
C19834 VDD.n2029 VSS 0.22487f
C19835 VDD.n2030 VSS 0.479077f
C19836 VDD.n2031 VSS -0.042134f
C19837 VDD.t2416 VSS 0.087181f
C19838 VDD.t2415 VSS 0.117879f
C19839 VDD.t2414 VSS 0.117879f
C19840 VDD.t539 VSS 0.117879f
C19841 VDD.t537 VSS 0.117879f
C19842 VDD.t525 VSS 0.115423f
C19843 VDD.t269 VSS 1.1086f
C19844 VDD.t2318 VSS 1.1086f
C19845 VDD.t2345 VSS 0.115423f
C19846 VDD.t2316 VSS 0.117879f
C19847 VDD.t1831 VSS 0.117879f
C19848 VDD.t2459 VSS 0.117879f
C19849 VDD.t2458 VSS 0.117879f
C19850 VDD.t2457 VSS 0.089637f
C19851 VDD.n2032 VSS -0.042134f
C19852 VDD.t2346 VSS 0.012354f
C19853 VDD.t2319 VSS 0.010856f
C19854 VDD.n2033 VSS 0.038523f
C19855 VDD.t1832 VSS 0.012354f
C19856 VDD.t2317 VSS 0.012354f
C19857 VDD.n2034 VSS 0.040938f
C19858 VDD.n2035 VSS 0.058757f
C19859 VDD.n2036 VSS 0.479077f
C19860 VDD.n2037 VSS 0.22487f
C19861 VDD.n2038 VSS 0.486456f
C19862 VDD.n2039 VSS 0.154688f
C19863 VDD.t1029 VSS 0.004807f
C19864 VDD.t1023 VSS 0.004807f
C19865 VDD.n2040 VSS 0.010736f
C19866 VDD.t1028 VSS 0.017466f
C19867 VDD.n2041 VSS 0.059157f
C19868 VDD.t365 VSS 1.52631f
C19869 VDD.t361 VSS 0.9101f
C19870 VDD.t363 VSS 1.02386f
C19871 VDD.t1704 VSS 0.004807f
C19872 VDD.t1702 VSS 0.004807f
C19873 VDD.n2042 VSS 0.010736f
C19874 VDD.t1703 VSS 0.017466f
C19875 VDD.n2043 VSS 0.048701f
C19876 VDD.n2044 VSS 0.011913f
C19877 VDD.n2045 VSS 0.001485f
C19878 VDD.n2046 VSS 0.001485f
C19879 VDD.t366 VSS 0.004807f
C19880 VDD.t362 VSS 0.004807f
C19881 VDD.n2047 VSS 0.010736f
C19882 VDD.t364 VSS 0.017466f
C19883 VDD.n2048 VSS 0.048701f
C19884 VDD.n2049 VSS 0.011913f
C19885 VDD.n2050 VSS 0.058133f
C19886 VDD.t2332 VSS 0.004807f
C19887 VDD.t2329 VSS 0.004807f
C19888 VDD.n2051 VSS 0.010736f
C19889 VDD.t2331 VSS 0.017466f
C19890 VDD.n2052 VSS 0.059157f
C19891 VDD.n2053 VSS 0.00433f
C19892 VDD.n2054 VSS 0.001485f
C19893 VDD.t478 VSS 0.004807f
C19894 VDD.t466 VSS 0.004807f
C19895 VDD.n2055 VSS 0.010736f
C19896 VDD.t475 VSS 0.017466f
C19897 VDD.n2056 VSS 0.059157f
C19898 VDD.n2057 VSS 0.00433f
C19899 VDD.n2058 VSS 0.001485f
C19900 VDD.t2165 VSS 0.004807f
C19901 VDD.t2159 VSS 0.004807f
C19902 VDD.n2059 VSS 0.010736f
C19903 VDD.t2164 VSS 0.017466f
C19904 VDD.n2060 VSS 0.059157f
C19905 VDD.n2061 VSS 0.00433f
C19906 VDD.n2062 VSS 0.001485f
C19907 VDD.t3589 VSS 0.004807f
C19908 VDD.t3581 VSS 0.004807f
C19909 VDD.n2063 VSS 0.010736f
C19910 VDD.t3588 VSS 0.017466f
C19911 VDD.n2064 VSS 0.059157f
C19912 VDD.n2065 VSS 0.00433f
C19913 VDD.n2066 VSS 0.001485f
C19914 VDD.t3963 VSS 0.004807f
C19915 VDD.t900 VSS 0.004807f
C19916 VDD.n2067 VSS 0.010736f
C19917 VDD.t902 VSS 0.017466f
C19918 VDD.n2068 VSS 0.059157f
C19919 VDD.n2069 VSS 0.00433f
C19920 VDD.n2070 VSS 0.001485f
C19921 VDD.t3532 VSS 0.004807f
C19922 VDD.t3527 VSS 0.004807f
C19923 VDD.n2071 VSS 0.010736f
C19924 VDD.t3531 VSS 0.017466f
C19925 VDD.n2072 VSS 0.059157f
C19926 VDD.n2073 VSS 0.00433f
C19927 VDD.n2074 VSS 0.001485f
C19928 VDD.t1390 VSS 0.004807f
C19929 VDD.t1388 VSS 0.004807f
C19930 VDD.n2075 VSS 0.010736f
C19931 VDD.t1389 VSS 0.017466f
C19932 VDD.n2076 VSS 0.059157f
C19933 VDD.n2077 VSS 0.00433f
C19934 VDD.t3106 VSS 0.004807f
C19935 VDD.t3110 VSS 0.004807f
C19936 VDD.n2078 VSS 0.010736f
C19937 VDD.t3108 VSS 0.017466f
C19938 VDD.n2079 VSS 0.054891f
C19939 VDD.t3109 VSS 0.006126f
C19940 VDD.t3105 VSS 0.008551f
C19941 VDD.t3107 VSS 0.008551f
C19942 VDD.n2080 VSS 0.027836f
C19943 VDD.t4515 VSS 0.009813f
C19944 VDD.n2081 VSS 0.069974f
C19945 VDD.t2000 VSS 0.004807f
C19946 VDD.t1998 VSS 0.004807f
C19947 VDD.n2082 VSS 0.010736f
C19948 VDD.t1999 VSS 0.017466f
C19949 VDD.n2083 VSS 0.048701f
C19950 VDD.n2084 VSS 0.011913f
C19951 VDD.n2085 VSS 0.058133f
C19952 VDD.n2086 VSS 0.154553f
C19953 VDD.t2496 VSS 0.004807f
C19954 VDD.t2494 VSS 0.004807f
C19955 VDD.n2087 VSS 0.010736f
C19956 VDD.t2495 VSS 0.017466f
C19957 VDD.n2088 VSS 0.048701f
C19958 VDD.n2089 VSS 0.011913f
C19959 VDD.n2090 VSS 0.058133f
C19960 VDD.n2091 VSS 0.12226f
C19961 VDD.t747 VSS 0.004807f
C19962 VDD.t800 VSS 0.004807f
C19963 VDD.n2092 VSS 0.010736f
C19964 VDD.t952 VSS 0.017466f
C19965 VDD.n2093 VSS 0.048701f
C19966 VDD.n2094 VSS 0.011913f
C19967 VDD.n2095 VSS 0.058133f
C19968 VDD.n2096 VSS 0.122181f
C19969 VDD.t682 VSS 0.004807f
C19970 VDD.t680 VSS 0.004807f
C19971 VDD.n2097 VSS 0.010736f
C19972 VDD.t681 VSS 0.017466f
C19973 VDD.n2098 VSS 0.048701f
C19974 VDD.n2099 VSS 0.011913f
C19975 VDD.n2100 VSS 0.058133f
C19976 VDD.n2101 VSS 0.154553f
C19977 VDD.t3493 VSS 0.004807f
C19978 VDD.t3491 VSS 0.004807f
C19979 VDD.n2102 VSS 0.010736f
C19980 VDD.t3492 VSS 0.017466f
C19981 VDD.n2103 VSS 0.048701f
C19982 VDD.n2104 VSS 0.011913f
C19983 VDD.n2105 VSS 0.058133f
C19984 VDD.n2106 VSS 0.154553f
C19985 VDD.t1189 VSS 0.004807f
C19986 VDD.t1187 VSS 0.004807f
C19987 VDD.n2107 VSS 0.010736f
C19988 VDD.t1188 VSS 0.017466f
C19989 VDD.n2108 VSS 0.048701f
C19990 VDD.n2109 VSS 0.011913f
C19991 VDD.n2110 VSS 0.058133f
C19992 VDD.n2111 VSS 0.211653f
C19993 VDD.n2112 VSS 0.04206f
C19994 VDD.n2113 VSS 0.012347f
C19995 VDD.n2114 VSS 0.982039f
C19996 VDD.n2115 VSS 0.00433f
C19997 VDD.n2116 VSS 0.058133f
C19998 VDD.n2117 VSS 0.457412f
C19999 VDD.n2118 VSS 0.384103f
C20000 VDD.n2119 VSS 0.154553f
C20001 VDD.t1238 VSS 0.004807f
C20002 VDD.t1240 VSS 0.004807f
C20003 VDD.n2120 VSS 0.010725f
C20004 VDD.t1239 VSS 0.017454f
C20005 VDD.n2121 VSS 0.048725f
C20006 VDD.t135 VSS 1.52631f
C20007 VDD.t467 VSS 0.9101f
C20008 VDD.t137 VSS 1.02386f
C20009 VDD.t1036 VSS 0.004807f
C20010 VDD.t1008 VSS 0.004807f
C20011 VDD.n2122 VSS 0.010725f
C20012 VDD.t1001 VSS 0.017454f
C20013 VDD.n2123 VSS 0.059309f
C20014 VDD.n2124 VSS 0.004283f
C20015 VDD.t2355 VSS 0.004807f
C20016 VDD.t2330 VSS 0.004807f
C20017 VDD.n2125 VSS 0.010725f
C20018 VDD.t2326 VSS 0.017454f
C20019 VDD.n2126 VSS 0.059309f
C20020 VDD.n2127 VSS 0.004283f
C20021 VDD.t2587 VSS 0.004807f
C20022 VDD.t468 VSS 0.004807f
C20023 VDD.n2128 VSS 0.010725f
C20024 VDD.t465 VSS 0.017454f
C20025 VDD.n2129 VSS 0.059309f
C20026 VDD.n2130 VSS 0.004283f
C20027 VDD.t2182 VSS 0.004807f
C20028 VDD.t2150 VSS 0.004807f
C20029 VDD.n2131 VSS 0.010725f
C20030 VDD.t2149 VSS 0.017454f
C20031 VDD.n2132 VSS 0.059309f
C20032 VDD.n2133 VSS 0.004283f
C20033 VDD.t3595 VSS 0.004807f
C20034 VDD.t3617 VSS 0.004807f
C20035 VDD.n2134 VSS 0.010725f
C20036 VDD.t3612 VSS 0.017454f
C20037 VDD.n2135 VSS 0.059309f
C20038 VDD.n2136 VSS 0.004283f
C20039 VDD.t3976 VSS 0.004807f
C20040 VDD.t901 VSS 0.004807f
C20041 VDD.n2137 VSS 0.010725f
C20042 VDD.t899 VSS 0.017454f
C20043 VDD.n2138 VSS 0.059309f
C20044 VDD.n2139 VSS 0.004283f
C20045 VDD.t3547 VSS 0.004807f
C20046 VDD.t3528 VSS 0.004807f
C20047 VDD.n2140 VSS 0.010725f
C20048 VDD.t3570 VSS 0.017454f
C20049 VDD.n2141 VSS 0.059309f
C20050 VDD.n2142 VSS 0.004283f
C20051 VDD.t1395 VSS 0.004807f
C20052 VDD.t1169 VSS 0.004807f
C20053 VDD.n2143 VSS 0.010725f
C20054 VDD.t1418 VSS 0.017454f
C20055 VDD.n2144 VSS 0.059309f
C20056 VDD.n2145 VSS 0.004283f
C20057 VDD.n2146 VSS 0.001403f
C20058 VDD.n2147 VSS 0.001403f
C20059 VDD.n2148 VSS 0.001403f
C20060 VDD.n2149 VSS 0.001403f
C20061 VDD.n2150 VSS 0.001403f
C20062 VDD.t1184 VSS 0.004807f
C20063 VDD.t1186 VSS 0.004807f
C20064 VDD.n2151 VSS 0.010725f
C20065 VDD.t1185 VSS 0.017454f
C20066 VDD.n2152 VSS 0.048725f
C20067 VDD.t136 VSS 0.004807f
C20068 VDD.t1206 VSS 0.004807f
C20069 VDD.n2153 VSS 0.010725f
C20070 VDD.t138 VSS 0.017454f
C20071 VDD.n2154 VSS 0.048725f
C20072 VDD.n2155 VSS 0.011995f
C20073 VDD.n2156 VSS 0.060165f
C20074 VDD.t1312 VSS 0.004807f
C20075 VDD.t1311 VSS 0.004807f
C20076 VDD.n2157 VSS 0.010725f
C20077 VDD.t1310 VSS 0.017454f
C20078 VDD.n2158 VSS 0.048725f
C20079 VDD.n2159 VSS 0.011995f
C20080 VDD.n2160 VSS 0.058133f
C20081 VDD.n2161 VSS 0.251569f
C20082 VDD.t817 VSS 0.004807f
C20083 VDD.t816 VSS 0.004807f
C20084 VDD.n2162 VSS 0.010725f
C20085 VDD.t815 VSS 0.017454f
C20086 VDD.n2163 VSS 0.048725f
C20087 VDD.n2164 VSS 0.011995f
C20088 VDD.n2165 VSS 0.058133f
C20089 VDD.n2166 VSS 0.154553f
C20090 VDD.t1197 VSS 0.004807f
C20091 VDD.t2063 VSS 0.004807f
C20092 VDD.n2167 VSS 0.010725f
C20093 VDD.t2062 VSS 0.017454f
C20094 VDD.n2168 VSS 0.048725f
C20095 VDD.n2169 VSS 0.011995f
C20096 VDD.n2170 VSS 0.058133f
C20097 VDD.n2171 VSS 0.121944f
C20098 VDD.t2553 VSS 0.004807f
C20099 VDD.t2552 VSS 0.004807f
C20100 VDD.n2172 VSS 0.010725f
C20101 VDD.t2551 VSS 0.017454f
C20102 VDD.n2173 VSS 0.048725f
C20103 VDD.n2174 VSS 0.011995f
C20104 VDD.n2175 VSS 0.058133f
C20105 VDD.n2176 VSS 0.122497f
C20106 VDD.n2177 VSS 0.154553f
C20107 VDD.n2178 VSS 0.058133f
C20108 VDD.n2179 VSS 0.011995f
C20109 VDD.n2180 VSS 0.001403f
C20110 VDD.t3264 VSS 0.004807f
C20111 VDD.t3263 VSS 0.004807f
C20112 VDD.n2181 VSS 0.010725f
C20113 VDD.t3262 VSS 0.017454f
C20114 VDD.n2182 VSS 0.048725f
C20115 VDD.n2183 VSS 0.058133f
C20116 VDD.n2184 VSS 0.011995f
C20117 VDD.n2185 VSS 0.001403f
C20118 VDD.t3112 VSS 0.004807f
C20119 VDD.t3114 VSS 0.004807f
C20120 VDD.n2186 VSS 0.010725f
C20121 VDD.t3104 VSS 0.017454f
C20122 VDD.n2187 VSS 0.054915f
C20123 VDD.t3113 VSS 0.006126f
C20124 VDD.t3111 VSS 0.008551f
C20125 VDD.t3103 VSS 0.008551f
C20126 VDD.n2188 VSS 0.027836f
C20127 VDD.t4516 VSS 0.009813f
C20128 VDD.n2189 VSS 0.069974f
C20129 VDD.n2190 VSS 0.04206f
C20130 VDD.n2191 VSS 0.012347f
C20131 VDD.n2192 VSS 0.982039f
C20132 VDD.n2193 VSS 0.001403f
C20133 VDD.n2194 VSS 0.011995f
C20134 VDD.n2195 VSS 0.058133f
C20135 VDD.n2196 VSS 0.095336f
C20136 VDD.n2197 VSS 0.50585f
C20137 VDD.n2198 VSS 0.54253f
C20138 VDD.n2199 VSS 0.106429f
C20139 VDD.t2344 VSS 0.004807f
C20140 VDD.t2348 VSS 0.004807f
C20141 VDD.n2200 VSS 0.010736f
C20142 VDD.t2340 VSS 0.017466f
C20143 VDD.n2201 VSS 0.054891f
C20144 VDD.t1011 VSS 0.231315f
C20145 VDD.t2582 VSS 0.004807f
C20146 VDD.t2600 VSS 0.004807f
C20147 VDD.n2202 VSS 0.010736f
C20148 VDD.t2581 VSS 0.017466f
C20149 VDD.n2203 VSS 0.054891f
C20150 VDD.n2204 VSS 0.016863f
C20151 VDD.t3611 VSS 0.004807f
C20152 VDD.t3594 VSS 0.004807f
C20153 VDD.n2205 VSS 0.010736f
C20154 VDD.t3610 VSS 0.017466f
C20155 VDD.n2206 VSS 0.054891f
C20156 VDD.n2207 VSS 0.016863f
C20157 VDD.t3971 VSS 0.004807f
C20158 VDD.t888 VSS 0.004807f
C20159 VDD.n2208 VSS 0.010736f
C20160 VDD.t3970 VSS 0.017466f
C20161 VDD.n2209 VSS 0.054891f
C20162 VDD.n2210 VSS 0.016863f
C20163 VDD.t2121 VSS 0.004807f
C20164 VDD.t2140 VSS 0.004807f
C20165 VDD.n2211 VSS 0.010736f
C20166 VDD.t2118 VSS 0.017466f
C20167 VDD.n2212 VSS 0.054891f
C20168 VDD.t3546 VSS 0.004807f
C20169 VDD.t3561 VSS 0.004807f
C20170 VDD.n2213 VSS 0.010736f
C20171 VDD.t3559 VSS 0.017466f
C20172 VDD.n2214 VSS 0.054891f
C20173 VDD.t1167 VSS 0.117695f
C20174 VDD.t1393 VSS 0.055923f
C20175 VDD.t1168 VSS 0.004807f
C20176 VDD.t1394 VSS 0.004807f
C20177 VDD.n2215 VSS 0.010736f
C20178 VDD.t1166 VSS 0.017466f
C20179 VDD.n2216 VSS 0.054891f
C20180 VDD.n2217 VSS 0.056662f
C20181 VDD.t1165 VSS 0.129226f
C20182 VDD.t3545 VSS 0.088326f
C20183 VDD.t3560 VSS 0.041419f
C20184 VDD.t2343 VSS 0.433154f
C20185 VDD.t1013 VSS 0.185052f
C20186 VDD.t2347 VSS 0.185052f
C20187 VDD.t887 VSS 0.134934f
C20188 VDD.t2339 VSS 0.052046f
C20189 VDD.n2218 VSS 0.244544f
C20190 VDD.t3558 VSS 0.089823f
C20191 VDD.n2219 VSS 0.050916f
C20192 VDD.n2220 VSS 0.221778f
C20193 VDD.n2221 VSS 0.121572f
C20194 VDD.n2222 VSS 0.1278f
C20195 VDD.n2223 VSS 0.092985f
C20196 VDD.n2224 VSS 0.016863f
C20197 VDD.t1014 VSS 0.004807f
C20198 VDD.t1039 VSS 0.004807f
C20199 VDD.n2225 VSS 0.010736f
C20200 VDD.t1012 VSS 0.017466f
C20201 VDD.n2226 VSS 0.054891f
C20202 VDD.n2227 VSS 0.016863f
C20203 VDD.n2228 VSS 0.404443f
C20204 VDD.n2229 VSS 0.221605f
C20205 VDD.n2230 VSS 0.016863f
C20206 VDD.n2231 VSS 0.865667f
C20207 VDD.n2232 VSS 2.10742f
C20208 VDD.n2233 VSS 0.094628f
C20209 VDD.n2234 VSS 0.221778f
C20210 VDD.t2279 VSS 0.004807f
C20211 VDD.t2278 VSS 0.004807f
C20212 VDD.n2235 VSS 0.010736f
C20213 VDD.t2277 VSS 0.017466f
C20214 VDD.n2236 VSS 0.054891f
C20215 VDD.t789 VSS 0.117695f
C20216 VDD.t787 VSS 0.055923f
C20217 VDD.t790 VSS 0.004807f
C20218 VDD.t788 VSS 0.004807f
C20219 VDD.n2237 VSS 0.010736f
C20220 VDD.t786 VSS 0.017466f
C20221 VDD.n2238 VSS 0.054891f
C20222 VDD.n2239 VSS 0.056662f
C20223 VDD.t785 VSS 0.129226f
C20224 VDD.t319 VSS 0.088326f
C20225 VDD.t317 VSS 0.041419f
C20226 VDD.t320 VSS 0.004807f
C20227 VDD.t318 VSS 0.004807f
C20228 VDD.n2240 VSS 0.010736f
C20229 VDD.t322 VSS 0.017466f
C20230 VDD.n2241 VSS 0.054891f
C20231 VDD.n2242 VSS 0.050916f
C20232 VDD.t321 VSS 0.089823f
C20233 VDD.t2482 VSS 0.433154f
C20234 VDD.t315 VSS 0.185052f
C20235 VDD.t2480 VSS 0.185052f
C20236 VDD.t313 VSS 0.134934f
C20237 VDD.n2243 VSS 0.244544f
C20238 VDD.t2478 VSS 0.052046f
C20239 VDD.t311 VSS 0.231315f
C20240 VDD.n2244 VSS 0.221605f
C20241 VDD.t316 VSS 0.004807f
C20242 VDD.t314 VSS 0.004807f
C20243 VDD.n2245 VSS 0.010736f
C20244 VDD.t312 VSS 0.017466f
C20245 VDD.n2246 VSS 0.054891f
C20246 VDD.n2247 VSS 0.016863f
C20247 VDD.t1547 VSS 0.004807f
C20248 VDD.t1546 VSS 0.004807f
C20249 VDD.n2248 VSS 0.010736f
C20250 VDD.t1545 VSS 0.017466f
C20251 VDD.n2249 VSS 0.054891f
C20252 VDD.n2250 VSS 0.016863f
C20253 VDD.t729 VSS 0.004807f
C20254 VDD.t731 VSS 0.004807f
C20255 VDD.n2251 VSS 0.010736f
C20256 VDD.t730 VSS 0.017466f
C20257 VDD.n2252 VSS 0.054891f
C20258 VDD.t2483 VSS 0.004807f
C20259 VDD.t2481 VSS 0.004807f
C20260 VDD.n2253 VSS 0.010736f
C20261 VDD.t2479 VSS 0.017466f
C20262 VDD.n2254 VSS 0.054891f
C20263 VDD.n2255 VSS 0.016863f
C20264 VDD.n2256 VSS 0.237366f
C20265 VDD.n2257 VSS 0.125401f
C20266 VDD.n2258 VSS 0.092985f
C20267 VDD.n2259 VSS 0.016863f
C20268 VDD.t371 VSS 0.004807f
C20269 VDD.t370 VSS 0.004807f
C20270 VDD.n2260 VSS 0.010736f
C20271 VDD.t369 VSS 0.017466f
C20272 VDD.n2261 VSS 0.054891f
C20273 VDD.n2262 VSS 0.016863f
C20274 VDD.n2263 VSS 0.404443f
C20275 VDD.n2264 VSS 0.016863f
C20276 VDD.n2265 VSS 0.072977f
C20277 VDD.n2266 VSS 0.344202f
C20278 VDD.n2267 VSS 0.030311f
C20279 VDD.t3446 VSS 0.126462f
C20280 VDD.t3449 VSS 0.075406f
C20281 VDD.t2298 VSS 0.075406f
C20282 VDD.t2299 VSS 0.075406f
C20283 VDD.t3429 VSS 0.075406f
C20284 VDD.t1170 VSS 0.075406f
C20285 VDD.t1172 VSS 0.075406f
C20286 VDD.t1398 VSS 0.058518f
C20287 VDD.t1416 VSS 0.126462f
C20288 VDD.t1400 VSS 0.05459f
C20289 VDD.n2268 VSS 2.52e-19
C20290 VDD.t1171 VSS 0.00575f
C20291 VDD.t1173 VSS 0.00575f
C20292 VDD.n2269 VSS 0.0115f
C20293 VDD.n2270 VSS 0.012479f
C20294 VDD.t1399 VSS 0.00575f
C20295 VDD.t1401 VSS 0.00575f
C20296 VDD.n2271 VSS 0.0115f
C20297 VDD.n2272 VSS 0.007448f
C20298 VDD.n2273 VSS 0.076419f
C20299 VDD.t1417 VSS 0.01978f
C20300 VDD.n2274 VSS 0.014195f
C20301 VDD.n2275 VSS -0.012705f
C20302 VDD.n2276 VSS 0.394106f
C20303 VDD.n2277 VSS 0.030311f
C20304 VDD.t2838 VSS 0.126462f
C20305 VDD.t2816 VSS 0.075406f
C20306 VDD.t2821 VSS 0.075406f
C20307 VDD.t2822 VSS 0.075406f
C20308 VDD.t2829 VSS 0.075406f
C20309 VDD.t3535 VSS 0.075406f
C20310 VDD.t3541 VSS 0.075406f
C20311 VDD.t3550 VSS 0.058518f
C20312 VDD.t3566 VSS 0.126462f
C20313 VDD.t3552 VSS 0.05459f
C20314 VDD.n2278 VSS 2.52e-19
C20315 VDD.t3536 VSS 0.00575f
C20316 VDD.t3542 VSS 0.00575f
C20317 VDD.n2279 VSS 0.0115f
C20318 VDD.n2280 VSS 0.012479f
C20319 VDD.t3551 VSS 0.00575f
C20320 VDD.t3553 VSS 0.00575f
C20321 VDD.n2281 VSS 0.0115f
C20322 VDD.n2282 VSS 0.007448f
C20323 VDD.n2283 VSS 0.076419f
C20324 VDD.t3567 VSS 0.01978f
C20325 VDD.n2284 VSS 0.014195f
C20326 VDD.n2285 VSS -0.012705f
C20327 VDD.n2286 VSS 0.753036f
C20328 VDD.n2287 VSS 0.030311f
C20329 VDD.t389 VSS 0.126462f
C20330 VDD.t390 VSS 0.075406f
C20331 VDD.t399 VSS 0.075406f
C20332 VDD.t400 VSS 0.075406f
C20333 VDD.t378 VSS 0.075406f
C20334 VDD.t3961 VSS 0.075406f
C20335 VDD.t3964 VSS 0.075406f
C20336 VDD.t3977 VSS 0.058518f
C20337 VDD.t895 VSS 0.126462f
C20338 VDD.t3983 VSS 0.05459f
C20339 VDD.n2288 VSS 2.52e-19
C20340 VDD.t3962 VSS 0.00575f
C20341 VDD.t3965 VSS 0.00575f
C20342 VDD.n2289 VSS 0.0115f
C20343 VDD.n2290 VSS 0.012479f
C20344 VDD.t3978 VSS 0.00575f
C20345 VDD.t3984 VSS 0.00575f
C20346 VDD.n2291 VSS 0.0115f
C20347 VDD.n2292 VSS 0.007448f
C20348 VDD.n2293 VSS 0.076419f
C20349 VDD.t896 VSS 0.01978f
C20350 VDD.n2294 VSS 0.014195f
C20351 VDD.n2295 VSS -0.012705f
C20352 VDD.n2296 VSS 0.759366f
C20353 VDD.n2297 VSS 0.030311f
C20354 VDD.t1642 VSS 0.126462f
C20355 VDD.t1643 VSS 0.075406f
C20356 VDD.t2203 VSS 0.075406f
C20357 VDD.t2204 VSS 0.075406f
C20358 VDD.t1637 VSS 0.075406f
C20359 VDD.t3606 VSS 0.075406f
C20360 VDD.t3608 VSS 0.075406f
C20361 VDD.t3586 VSS 0.058518f
C20362 VDD.t3598 VSS 0.126462f
C20363 VDD.t3590 VSS 0.05459f
C20364 VDD.n2298 VSS 2.52e-19
C20365 VDD.t3607 VSS 0.00575f
C20366 VDD.t3609 VSS 0.00575f
C20367 VDD.n2299 VSS 0.0115f
C20368 VDD.n2300 VSS 0.012479f
C20369 VDD.t3587 VSS 0.00575f
C20370 VDD.t3591 VSS 0.00575f
C20371 VDD.n2301 VSS 0.0115f
C20372 VDD.n2302 VSS 0.007448f
C20373 VDD.n2303 VSS 0.076419f
C20374 VDD.t3599 VSS 0.01978f
C20375 VDD.n2304 VSS 0.014195f
C20376 VDD.n2305 VSS -0.012705f
C20377 VDD.n2306 VSS 0.550475f
C20378 VDD.n2307 VSS 0.661458f
C20379 VDD.n2308 VSS 0.030311f
C20380 VDD.t4095 VSS 0.126462f
C20381 VDD.t4098 VSS 0.075406f
C20382 VDD.t4115 VSS 0.075406f
C20383 VDD.t4118 VSS 0.075406f
C20384 VDD.t4072 VSS 0.075406f
C20385 VDD.t2160 VSS 0.075406f
C20386 VDD.t2166 VSS 0.075406f
C20387 VDD.t2122 VSS 0.058518f
C20388 VDD.t2147 VSS 0.126462f
C20389 VDD.t2128 VSS 0.05459f
C20390 VDD.n2309 VSS 2.52e-19
C20391 VDD.t2161 VSS 0.00575f
C20392 VDD.t2167 VSS 0.00575f
C20393 VDD.n2310 VSS 0.0115f
C20394 VDD.n2311 VSS 0.012479f
C20395 VDD.t2123 VSS 0.00575f
C20396 VDD.t2129 VSS 0.00575f
C20397 VDD.n2312 VSS 0.0115f
C20398 VDD.n2313 VSS 0.007448f
C20399 VDD.n2314 VSS 0.076419f
C20400 VDD.t2148 VSS 0.01978f
C20401 VDD.n2315 VSS 0.014195f
C20402 VDD.n2316 VSS -0.012705f
C20403 VDD.n2317 VSS 0.596411f
C20404 VDD.n2318 VSS 0.030311f
C20405 VDD.t527 VSS 0.126462f
C20406 VDD.t528 VSS 0.075406f
C20407 VDD.t551 VSS 0.075406f
C20408 VDD.t552 VSS 0.075406f
C20409 VDD.t516 VSS 0.075406f
C20410 VDD.t2605 VSS 0.075406f
C20411 VDD.t2611 VSS 0.075406f
C20412 VDD.t2575 VSS 0.058518f
C20413 VDD.t2596 VSS 0.126462f
C20414 VDD.t2577 VSS 0.05459f
C20415 VDD.n2319 VSS 2.52e-19
C20416 VDD.t2606 VSS 0.00575f
C20417 VDD.t2612 VSS 0.00575f
C20418 VDD.n2320 VSS 0.0115f
C20419 VDD.n2321 VSS 0.012479f
C20420 VDD.t2576 VSS 0.00575f
C20421 VDD.t2578 VSS 0.00575f
C20422 VDD.n2322 VSS 0.0115f
C20423 VDD.n2323 VSS 0.007448f
C20424 VDD.n2324 VSS 0.076419f
C20425 VDD.t2597 VSS 0.01978f
C20426 VDD.n2325 VSS 0.014195f
C20427 VDD.n2326 VSS -0.012705f
C20428 VDD.n2327 VSS 0.755669f
C20429 VDD.n2328 VSS 0.030311f
C20430 VDD.t4227 VSS 0.126462f
C20431 VDD.t4234 VSS 0.075406f
C20432 VDD.t4198 VSS 0.075406f
C20433 VDD.t4201 VSS 0.075406f
C20434 VDD.t4216 VSS 0.075406f
C20435 VDD.t2376 VSS 0.075406f
C20436 VDD.t2378 VSS 0.075406f
C20437 VDD.t2333 VSS 0.058518f
C20438 VDD.t2362 VSS 0.126462f
C20439 VDD.t2337 VSS 0.05459f
C20440 VDD.n2329 VSS 2.52e-19
C20441 VDD.t2377 VSS 0.00575f
C20442 VDD.t2379 VSS 0.00575f
C20443 VDD.n2330 VSS 0.0115f
C20444 VDD.n2331 VSS 0.012479f
C20445 VDD.t2334 VSS 0.00575f
C20446 VDD.t2338 VSS 0.00575f
C20447 VDD.n2332 VSS 0.0115f
C20448 VDD.n2333 VSS 0.007448f
C20449 VDD.n2334 VSS 0.076419f
C20450 VDD.t2363 VSS 0.01978f
C20451 VDD.n2335 VSS 0.014195f
C20452 VDD.n2336 VSS -0.012705f
C20453 VDD.n2337 VSS 0.574483f
C20454 VDD.n2338 VSS 1.23571f
C20455 VDD.n2339 VSS 0.930271f
C20456 VDD.n2340 VSS 1.47494f
C20457 VDD.n2341 VSS 1.34255f
C20458 VDD.n2342 VSS 0.970482f
C20459 VDD.n2343 VSS 0.856497f
C20460 VDD.n2344 VSS 0.97219f
C20461 VDD.n2345 VSS 0.865236f
C20462 VDD.n2346 VSS 0.444376f
C20463 VDD.n2347 VSS 0.132031f
C20464 VDD.n2348 VSS 0.306798f
C20465 VDD.n2349 VSS 0.22487f
C20466 VDD.t1941 VSS 0.012354f
C20467 VDD.t1937 VSS 0.012354f
C20468 VDD.n2350 VSS 0.040938f
C20469 VDD.t1913 VSS 0.012354f
C20470 VDD.t1939 VSS 0.010856f
C20471 VDD.n2351 VSS 0.038523f
C20472 VDD.n2352 VSS 0.058757f
C20473 VDD.n2353 VSS 0.479072f
C20474 VDD.n2354 VSS -0.041546f
C20475 VDD.t2036 VSS 0.088051f
C20476 VDD.t2035 VSS 0.119055f
C20477 VDD.t2034 VSS 0.119055f
C20478 VDD.t634 VSS 0.119055f
C20479 VDD.t1611 VSS 0.119055f
C20480 VDD.t1607 VSS 0.116575f
C20481 VDD.t638 VSS 0.254852f
C20482 VDD.t494 VSS 0.254852f
C20483 VDD.t2735 VSS 0.116575f
C20484 VDD.t500 VSS 0.119055f
C20485 VDD.t498 VSS 0.119055f
C20486 VDD.t693 VSS 0.119055f
C20487 VDD.t692 VSS 0.119055f
C20488 VDD.t691 VSS 0.090532f
C20489 VDD.t2560 VSS 0.010856f
C20490 VDD.t2568 VSS 0.012354f
C20491 VDD.n2355 VSS 0.038675f
C20492 VDD.t2556 VSS 0.012354f
C20493 VDD.t2558 VSS 0.012354f
C20494 VDD.n2356 VSS 0.040145f
C20495 VDD.n2357 VSS 0.059265f
C20496 VDD.n2358 VSS 0.22487f
C20497 VDD.t499 VSS 0.012354f
C20498 VDD.t501 VSS 0.012354f
C20499 VDD.n2359 VSS 0.040938f
C20500 VDD.t2736 VSS 0.012354f
C20501 VDD.t495 VSS 0.010856f
C20502 VDD.n2360 VSS 0.038523f
C20503 VDD.n2361 VSS 0.058757f
C20504 VDD.n2362 VSS 0.479072f
C20505 VDD.n2363 VSS -0.041546f
C20506 VDD.t2847 VSS 0.088051f
C20507 VDD.t2846 VSS 0.119055f
C20508 VDD.t2845 VSS 0.119055f
C20509 VDD.t2557 VSS 0.119055f
C20510 VDD.t2555 VSS 0.119055f
C20511 VDD.t2567 VSS 0.116575f
C20512 VDD.t2559 VSS 0.362126f
C20513 VDD.t2911 VSS 0.362126f
C20514 VDD.t2921 VSS 0.116575f
C20515 VDD.t2919 VSS 0.119055f
C20516 VDD.t2917 VSS 0.119055f
C20517 VDD.t2429 VSS 0.119055f
C20518 VDD.t2428 VSS 0.119055f
C20519 VDD.t2427 VSS 0.090532f
C20520 VDD.n2364 VSS -0.041546f
C20521 VDD.n2365 VSS 0.479072f
C20522 VDD.n2366 VSS 0.22487f
C20523 VDD.n2367 VSS 0.289805f
C20524 VDD.n2368 VSS 1.02856f
C20525 VDD.t2240 VSS 0.069002f
C20526 VDD.t2234 VSS 0.171787f
C20527 VDD.t162 VSS 0.238557f
C20528 VDD.t164 VSS 0.004807f
C20529 VDD.t165 VSS 0.004807f
C20530 VDD.n2369 VSS 0.010736f
C20531 VDD.t163 VSS 0.017466f
C20532 VDD.n2370 VSS 0.059057f
C20533 VDD.n2371 VSS 0.044667f
C20534 VDD.n2372 VSS 0.763609f
C20535 VDD.n2373 VSS 0.699488f
C20536 VDD.n2374 VSS 0.173847f
C20537 VDD.t1022 VSS 0.017474f
C20538 VDD.t992 VSS 0.004807f
C20539 VDD.t1000 VSS 0.004807f
C20540 VDD.n2375 VSS 0.010696f
C20541 VDD.n2376 VSS 0.097619f
C20542 VDD.n2377 VSS 0.024454f
C20543 VDD.n2378 VSS 0.007059f
C20544 VDD.t991 VSS 0.049955f
C20545 VDD.t999 VSS 0.069002f
C20546 VDD.t1021 VSS 0.3637f
C20547 VDD.t1058 VSS 0.004807f
C20548 VDD.t1059 VSS 0.004807f
C20549 VDD.n2379 VSS 0.010736f
C20550 VDD.t1057 VSS 0.017466f
C20551 VDD.n2380 VSS 0.059057f
C20552 VDD.n2381 VSS 0.044188f
C20553 VDD.n2382 VSS 0.319849f
C20554 VDD.t1056 VSS 0.130817f
C20555 VDD.t4210 VSS 0.164959f
C20556 VDD.t4212 VSS 0.069002f
C20557 VDD.t4228 VSS 0.053549f
C20558 VDD.t236 VSS 0.126864f
C20559 VDD.t237 VSS 0.004807f
C20560 VDD.t238 VSS 0.004807f
C20561 VDD.n2383 VSS 0.010736f
C20562 VDD.t1329 VSS 0.017466f
C20563 VDD.n2384 VSS 0.059057f
C20564 VDD.n2385 VSS 1.14539f
C20565 VDD.t554 VSS 0.017474f
C20566 VDD.t264 VSS 0.004807f
C20567 VDD.t518 VSS 0.004807f
C20568 VDD.n2386 VSS 0.010696f
C20569 VDD.n2387 VSS 0.09764f
C20570 VDD.t1027 VSS 0.017474f
C20571 VDD.t996 VSS 0.004807f
C20572 VDD.t1003 VSS 0.004807f
C20573 VDD.n2388 VSS 0.010696f
C20574 VDD.n2389 VSS 0.097619f
C20575 VDD.t553 VSS 0.161006f
C20576 VDD.t263 VSS 0.069002f
C20577 VDD.t517 VSS 0.053549f
C20578 VDD.t1017 VSS 0.115723f
C20579 VDD.t1015 VSS 0.069002f
C20580 VDD.t593 VSS 0.049955f
C20581 VDD.t4088 VSS 0.017474f
C20582 VDD.t4086 VSS 0.004807f
C20583 VDD.t4092 VSS 0.004807f
C20584 VDD.n2390 VSS 0.010696f
C20585 VDD.n2391 VSS 0.09764f
C20586 VDD.n2392 VSS 0.201578f
C20587 VDD.t1018 VSS 0.017474f
C20588 VDD.t594 VSS 0.004807f
C20589 VDD.t1016 VSS 0.004807f
C20590 VDD.n2393 VSS 0.010696f
C20591 VDD.n2394 VSS 0.097619f
C20592 VDD.n2395 VSS 0.024454f
C20593 VDD.n2396 VSS 0.007059f
C20594 VDD.t4091 VSS 0.053549f
C20595 VDD.t4085 VSS 0.069002f
C20596 VDD.t4087 VSS 0.167115f
C20597 VDD.t1157 VSS 0.132973f
C20598 VDD.t1205 VSS 0.004807f
C20599 VDD.t1158 VSS 0.004807f
C20600 VDD.n2397 VSS 0.010736f
C20601 VDD.t1159 VSS 0.017466f
C20602 VDD.n2398 VSS 0.059057f
C20603 VDD.n2399 VSS 0.044188f
C20604 VDD.n2400 VSS 0.417243f
C20605 VDD.t1026 VSS 0.461094f
C20606 VDD.t1002 VSS 0.069002f
C20607 VDD.t995 VSS 0.049955f
C20608 VDD.n2401 VSS 0.007059f
C20609 VDD.n2402 VSS 0.024454f
C20610 VDD.n2403 VSS 0.173847f
C20611 VDD.n2404 VSS 0.767891f
C20612 VDD.n2405 VSS 0.378545f
C20613 VDD.n2406 VSS 0.044188f
C20614 VDD.n2407 VSS 0.31302f
C20615 VDD.t989 VSS 0.356872f
C20616 VDD.t583 VSS 0.069002f
C20617 VDD.t1034 VSS 0.049955f
C20618 VDD.n2408 VSS 0.007059f
C20619 VDD.n2409 VSS 0.024454f
C20620 VDD.n2410 VSS 0.173847f
C20621 VDD.n2411 VSS 0.368537f
C20622 VDD.n2412 VSS 0.356333f
C20623 VDD.n2413 VSS 0.331071f
C20624 VDD.t2473 VSS 0.017476f
C20625 VDD.t2477 VSS 0.004807f
C20626 VDD.t2475 VSS 0.004807f
C20627 VDD.n2414 VSS 0.010696f
C20628 VDD.n2415 VSS 0.098224f
C20629 VDD.n2416 VSS 0.048045f
C20630 VDD.t1120 VSS 0.017462f
C20631 VDD.t2406 VSS 0.017474f
C20632 VDD.t2402 VSS 0.004807f
C20633 VDD.t2408 VSS 0.004807f
C20634 VDD.n2417 VSS 0.010696f
C20635 VDD.n2418 VSS 0.097619f
C20636 VDD.t405 VSS 0.052737f
C20637 VDD.t404 VSS 0.017476f
C20638 VDD.t408 VSS 0.004807f
C20639 VDD.t406 VSS 0.004807f
C20640 VDD.n2419 VSS 0.010696f
C20641 VDD.n2420 VSS 0.099623f
C20642 VDD.n2421 VSS 0.194608f
C20643 VDD.t2753 VSS 0.010856f
C20644 VDD.t2749 VSS 0.012354f
C20645 VDD.n2422 VSS 0.038675f
C20646 VDD.t2755 VSS 0.012354f
C20647 VDD.t2751 VSS 0.012354f
C20648 VDD.n2423 VSS 0.040145f
C20649 VDD.n2424 VSS 0.059265f
C20650 VDD.t3905 VSS 0.012354f
C20651 VDD.t3901 VSS 0.012354f
C20652 VDD.n2425 VSS 0.040938f
C20653 VDD.t3913 VSS 0.012354f
C20654 VDD.t3903 VSS 0.010856f
C20655 VDD.n2426 VSS 0.038523f
C20656 VDD.n2427 VSS 0.058757f
C20657 VDD.t773 VSS 0.088051f
C20658 VDD.t3949 VSS 0.010856f
C20659 VDD.t3939 VSS 0.012354f
C20660 VDD.n2428 VSS 0.038675f
C20661 VDD.t3951 VSS 0.012354f
C20662 VDD.t3947 VSS 0.012354f
C20663 VDD.n2429 VSS 0.040145f
C20664 VDD.n2430 VSS 0.059265f
C20665 VDD.t1626 VSS 0.017476f
C20666 VDD.t1630 VSS 0.004807f
C20667 VDD.t1628 VSS 0.004807f
C20668 VDD.n2431 VSS 0.010696f
C20669 VDD.n2432 VSS 0.099623f
C20670 VDD.n2433 VSS 0.036461f
C20671 VDD.t909 VSS 0.017476f
C20672 VDD.t3465 VSS 0.004807f
C20673 VDD.t3463 VSS 0.004807f
C20674 VDD.n2434 VSS 0.010696f
C20675 VDD.n2435 VSS 0.098224f
C20676 VDD.n2436 VSS 0.048045f
C20677 VDD.t3941 VSS 0.017462f
C20678 VDD.t300 VSS 0.017474f
C20679 VDD.t298 VSS 0.004807f
C20680 VDD.t302 VSS 0.004807f
C20681 VDD.n2437 VSS 0.010696f
C20682 VDD.n2438 VSS 0.097619f
C20683 VDD.t4096 VSS 0.052737f
C20684 VDD.t4106 VSS 0.017476f
C20685 VDD.t4110 VSS 0.004807f
C20686 VDD.t4097 VSS 0.004807f
C20687 VDD.n2439 VSS 0.010696f
C20688 VDD.n2440 VSS 0.099623f
C20689 VDD.n2441 VSS 0.194608f
C20690 VDD.t1728 VSS 0.010856f
C20691 VDD.t1740 VSS 0.012354f
C20692 VDD.n2442 VSS 0.038675f
C20693 VDD.t1732 VSS 0.012354f
C20694 VDD.t1730 VSS 0.012354f
C20695 VDD.n2443 VSS 0.040145f
C20696 VDD.n2444 VSS 0.059265f
C20697 VDD.t1551 VSS 0.012354f
C20698 VDD.t1553 VSS 0.012354f
C20699 VDD.n2445 VSS 0.040938f
C20700 VDD.t1555 VSS 0.012354f
C20701 VDD.t1557 VSS 0.010856f
C20702 VDD.n2446 VSS 0.038523f
C20703 VDD.n2447 VSS 0.058757f
C20704 VDD.t884 VSS 0.088051f
C20705 VDD.t93 VSS 0.010856f
C20706 VDD.t89 VSS 0.012354f
C20707 VDD.n2448 VSS 0.038675f
C20708 VDD.t87 VSS 0.012354f
C20709 VDD.t91 VSS 0.012354f
C20710 VDD.n2449 VSS 0.040145f
C20711 VDD.n2450 VSS 0.059265f
C20712 VDD.t266 VSS 0.017476f
C20713 VDD.t546 VSS 0.004807f
C20714 VDD.t542 VSS 0.004807f
C20715 VDD.n2451 VSS 0.010696f
C20716 VDD.n2452 VSS 0.099623f
C20717 VDD.n2453 VSS 0.036461f
C20718 VDD.t448 VSS 0.017476f
C20719 VDD.t446 VSS 0.004807f
C20720 VDD.t444 VSS 0.004807f
C20721 VDD.n2454 VSS 0.010696f
C20722 VDD.n2455 VSS 0.098224f
C20723 VDD.n2456 VSS 0.048045f
C20724 VDD.t95 VSS 0.017462f
C20725 VDD.t2467 VSS 0.017474f
C20726 VDD.t2471 VSS 0.004807f
C20727 VDD.t2469 VSS 0.004807f
C20728 VDD.n2457 VSS 0.010696f
C20729 VDD.n2458 VSS 0.097619f
C20730 VDD.t4202 VSS 0.052737f
C20731 VDD.t4207 VSS 0.017476f
C20732 VDD.t4205 VSS 0.004807f
C20733 VDD.t4203 VSS 0.004807f
C20734 VDD.n2459 VSS 0.010696f
C20735 VDD.n2460 VSS 0.099623f
C20736 VDD.n2461 VSS 0.538951f
C20737 VDD.t1328 VSS 0.017476f
C20738 VDD.t2540 VSS 0.004807f
C20739 VDD.t2538 VSS 0.004807f
C20740 VDD.n2462 VSS 0.010696f
C20741 VDD.n2463 VSS 0.098224f
C20742 VDD.n2464 VSS 0.048045f
C20743 VDD.t806 VSS 0.017462f
C20744 VDD.t749 VSS 0.017474f
C20745 VDD.t753 VSS 0.004807f
C20746 VDD.t751 VSS 0.004807f
C20747 VDD.n2465 VSS 0.010696f
C20748 VDD.n2466 VSS 0.097619f
C20749 VDD.t2219 VSS 0.052737f
C20750 VDD.t2224 VSS 0.017476f
C20751 VDD.t2222 VSS 0.004807f
C20752 VDD.t2220 VSS 0.004807f
C20753 VDD.n2467 VSS 0.010696f
C20754 VDD.n2468 VSS 0.099623f
C20755 VDD.t1825 VSS 0.017474f
C20756 VDD.t1827 VSS 0.004807f
C20757 VDD.t1823 VSS 0.004807f
C20758 VDD.n2469 VSS 0.010696f
C20759 VDD.n2470 VSS 0.097975f
C20760 VDD.n2471 VSS 0.048045f
C20761 VDD.t1776 VSS 0.017462f
C20762 VDD.t2257 VSS 0.017474f
C20763 VDD.t2255 VSS 0.004807f
C20764 VDD.t2253 VSS 0.004807f
C20765 VDD.n2472 VSS 0.010696f
C20766 VDD.n2473 VSS 0.097619f
C20767 VDD.t1824 VSS 0.19396f
C20768 VDD.t1826 VSS 0.067957f
C20769 VDD.t1822 VSS 0.052737f
C20770 VDD.t3402 VSS 0.017474f
C20771 VDD.t3404 VSS 0.004807f
C20772 VDD.t3406 VSS 0.004807f
C20773 VDD.n2474 VSS 0.010696f
C20774 VDD.n2475 VSS 0.099162f
C20775 VDD.n2476 VSS 0.02587f
C20776 VDD.n2477 VSS 0.006536f
C20777 VDD.t3403 VSS 0.049198f
C20778 VDD.t3405 VSS 0.067957f
C20779 VDD.t3401 VSS 0.176263f
C20780 VDD.t1775 VSS 0.176263f
C20781 VDD.t1769 VSS 0.067957f
C20782 VDD.t1761 VSS 0.052737f
C20783 VDD.t2221 VSS 0.067957f
C20784 VDD.t2223 VSS 0.256608f
C20785 VDD.t2256 VSS 0.256608f
C20786 VDD.t2252 VSS 0.067957f
C20787 VDD.t2254 VSS 0.049198f
C20788 VDD.n2478 VSS 0.006536f
C20789 VDD.n2479 VSS 0.024888f
C20790 VDD.t1770 VSS 0.004807f
C20791 VDD.t1762 VSS 0.004807f
C20792 VDD.n2480 VSS 0.010696f
C20793 VDD.n2481 VSS 0.036584f
C20794 VDD.n2482 VSS 0.092113f
C20795 VDD.n2483 VSS 0.194608f
C20796 VDD.t1802 VSS 0.010856f
C20797 VDD.t1752 VSS 0.012354f
C20798 VDD.n2484 VSS 0.038675f
C20799 VDD.t1768 VSS 0.012354f
C20800 VDD.t1794 VSS 0.012354f
C20801 VDD.n2485 VSS 0.040145f
C20802 VDD.n2486 VSS 0.059265f
C20803 VDD.t2261 VSS 0.012354f
C20804 VDD.t2259 VSS 0.012354f
C20805 VDD.n2487 VSS 0.040938f
C20806 VDD.t2265 VSS 0.012354f
C20807 VDD.t2263 VSS 0.010856f
C20808 VDD.n2488 VSS 0.038523f
C20809 VDD.n2489 VSS 0.058757f
C20810 VDD.t1801 VSS 0.192225f
C20811 VDD.t1751 VSS 0.116575f
C20812 VDD.t1767 VSS 0.119055f
C20813 VDD.t1793 VSS 0.119055f
C20814 VDD.t2393 VSS 0.119055f
C20815 VDD.t1441 VSS 0.119055f
C20816 VDD.t3378 VSS 0.088051f
C20817 VDD.t886 VSS 0.119055f
C20818 VDD.t885 VSS 0.119055f
C20819 VDD.t90 VSS 0.119055f
C20820 VDD.t86 VSS 0.119055f
C20821 VDD.t88 VSS 0.116575f
C20822 VDD.t92 VSS 0.362126f
C20823 VDD.t4146 VSS 0.362126f
C20824 VDD.t4144 VSS 0.116575f
C20825 VDD.t4140 VSS 0.119055f
C20826 VDD.t4142 VSS 0.119055f
C20827 VDD.t797 VSS 0.119055f
C20828 VDD.t798 VSS 0.119055f
C20829 VDD.t799 VSS 0.090532f
C20830 VDD.t4222 VSS 0.010856f
C20831 VDD.t4200 VSS 0.012354f
C20832 VDD.n2490 VSS 0.038675f
C20833 VDD.t4226 VSS 0.012354f
C20834 VDD.t4233 VSS 0.012354f
C20835 VDD.n2491 VSS 0.040145f
C20836 VDD.n2492 VSS 0.059265f
C20837 VDD.t4143 VSS 0.012354f
C20838 VDD.t4141 VSS 0.012354f
C20839 VDD.n2493 VSS 0.040938f
C20840 VDD.t4145 VSS 0.012354f
C20841 VDD.t4147 VSS 0.010856f
C20842 VDD.n2494 VSS 0.038523f
C20843 VDD.n2495 VSS 0.058757f
C20844 VDD.n2496 VSS 0.22487f
C20845 VDD.n2497 VSS 0.479072f
C20846 VDD.n2498 VSS -0.041546f
C20847 VDD.t3380 VSS 0.088051f
C20848 VDD.t1182 VSS 0.119055f
C20849 VDD.t1183 VSS 0.119055f
C20850 VDD.t4232 VSS 0.119055f
C20851 VDD.t4225 VSS 0.119055f
C20852 VDD.t4199 VSS 0.116575f
C20853 VDD.t4221 VSS 0.254852f
C20854 VDD.t758 VSS 0.254852f
C20855 VDD.t760 VSS 0.116575f
C20856 VDD.t754 VSS 0.119055f
C20857 VDD.t756 VSS 0.119055f
C20858 VDD.t1542 VSS 0.119055f
C20859 VDD.t1624 VSS 0.119055f
C20860 VDD.t1543 VSS 0.090532f
C20861 VDD.t2627 VSS 0.010856f
C20862 VDD.t2625 VSS 0.012354f
C20863 VDD.n2499 VSS 0.038675f
C20864 VDD.t2631 VSS 0.012354f
C20865 VDD.t2629 VSS 0.012354f
C20866 VDD.n2500 VSS 0.040145f
C20867 VDD.n2501 VSS 0.059265f
C20868 VDD.n2502 VSS 0.31205f
C20869 VDD.t757 VSS 0.012354f
C20870 VDD.t755 VSS 0.012354f
C20871 VDD.n2503 VSS 0.040938f
C20872 VDD.t761 VSS 0.012354f
C20873 VDD.t759 VSS 0.010856f
C20874 VDD.n2504 VSS 0.038523f
C20875 VDD.n2505 VSS 0.058757f
C20876 VDD.n2506 VSS 0.479072f
C20877 VDD.n2507 VSS -0.041546f
C20878 VDD.t2267 VSS 0.088051f
C20879 VDD.t178 VSS 0.119055f
C20880 VDD.t2266 VSS 0.119055f
C20881 VDD.t2628 VSS 0.119055f
C20882 VDD.t2630 VSS 0.119055f
C20883 VDD.t2624 VSS 0.116575f
C20884 VDD.t2626 VSS 0.362126f
C20885 VDD.t2086 VSS 0.362126f
C20886 VDD.t2094 VSS 0.116575f
C20887 VDD.t2082 VSS 0.119055f
C20888 VDD.t2088 VSS 0.119055f
C20889 VDD.t582 VSS 0.119055f
C20890 VDD.t2554 VSS 0.119055f
C20891 VDD.t581 VSS 0.090532f
C20892 VDD.t2228 VSS 0.010856f
C20893 VDD.t1678 VSS 0.012354f
C20894 VDD.n2508 VSS 0.038675f
C20895 VDD.t2245 VSS 0.012354f
C20896 VDD.t2232 VSS 0.012354f
C20897 VDD.n2509 VSS 0.040145f
C20898 VDD.n2510 VSS 0.059265f
C20899 VDD.n2511 VSS 0.22487f
C20900 VDD.t2089 VSS 0.012354f
C20901 VDD.t2083 VSS 0.012354f
C20902 VDD.n2512 VSS 0.040938f
C20903 VDD.t2095 VSS 0.012354f
C20904 VDD.t2087 VSS 0.010856f
C20905 VDD.n2513 VSS 0.038523f
C20906 VDD.n2514 VSS 0.058757f
C20907 VDD.n2515 VSS 0.479072f
C20908 VDD.n2516 VSS -0.041546f
C20909 VDD.t1254 VSS 0.088051f
C20910 VDD.t1252 VSS 0.119055f
C20911 VDD.t1253 VSS 0.119055f
C20912 VDD.t2231 VSS 0.119055f
C20913 VDD.t2244 VSS 0.119055f
C20914 VDD.t1677 VSS 0.116575f
C20915 VDD.t2227 VSS 0.254852f
C20916 VDD.t2262 VSS 0.254852f
C20917 VDD.t2264 VSS 0.116575f
C20918 VDD.t2258 VSS 0.119055f
C20919 VDD.t2260 VSS 0.119055f
C20920 VDD.t3120 VSS 0.119055f
C20921 VDD.t3119 VSS 0.119055f
C20922 VDD.t3121 VSS 0.090532f
C20923 VDD.n2517 VSS -0.041546f
C20924 VDD.n2518 VSS 0.479072f
C20925 VDD.n2519 VSS 0.31205f
C20926 VDD.n2520 VSS 0.538951f
C20927 VDD.n2521 VSS 0.392773f
C20928 VDD.n2522 VSS 0.036461f
C20929 VDD.t2085 VSS 0.017474f
C20930 VDD.t2093 VSS 0.004807f
C20931 VDD.t2091 VSS 0.004807f
C20932 VDD.n2523 VSS 0.010696f
C20933 VDD.n2524 VSS 0.099467f
C20934 VDD.n2525 VSS 0.025249f
C20935 VDD.n2526 VSS 0.006536f
C20936 VDD.t2092 VSS 0.049198f
C20937 VDD.t2090 VSS 0.067957f
C20938 VDD.t2084 VSS 0.324211f
C20939 VDD.t1327 VSS 0.324211f
C20940 VDD.t2539 VSS 0.067957f
C20941 VDD.t2537 VSS 0.052737f
C20942 VDD.t1359 VSS 0.017474f
C20943 VDD.t1363 VSS 0.004807f
C20944 VDD.t1361 VSS 0.004807f
C20945 VDD.n2527 VSS 0.010696f
C20946 VDD.n2528 VSS 0.099162f
C20947 VDD.n2529 VSS 0.02587f
C20948 VDD.n2530 VSS 0.006536f
C20949 VDD.t1362 VSS 0.049198f
C20950 VDD.t1360 VSS 0.067957f
C20951 VDD.t1358 VSS 0.176263f
C20952 VDD.t805 VSS 0.176263f
C20953 VDD.t803 VSS 0.067957f
C20954 VDD.t801 VSS 0.052737f
C20955 VDD.t4204 VSS 0.067957f
C20956 VDD.t4206 VSS 0.256608f
C20957 VDD.t748 VSS 0.256608f
C20958 VDD.t750 VSS 0.067957f
C20959 VDD.t752 VSS 0.049198f
C20960 VDD.n2531 VSS 0.006536f
C20961 VDD.n2532 VSS 0.024888f
C20962 VDD.t804 VSS 0.004807f
C20963 VDD.t802 VSS 0.004807f
C20964 VDD.n2533 VSS 0.010696f
C20965 VDD.n2534 VSS 0.036584f
C20966 VDD.n2535 VSS 0.092113f
C20967 VDD.n2536 VSS 0.194608f
C20968 VDD.n2537 VSS 0.392773f
C20969 VDD.n2538 VSS 0.036461f
C20970 VDD.t4139 VSS 0.017474f
C20971 VDD.t4137 VSS 0.004807f
C20972 VDD.t4135 VSS 0.004807f
C20973 VDD.n2539 VSS 0.010696f
C20974 VDD.n2540 VSS 0.099467f
C20975 VDD.n2541 VSS 0.025249f
C20976 VDD.n2542 VSS 0.006536f
C20977 VDD.t4136 VSS 0.049198f
C20978 VDD.t4134 VSS 0.067957f
C20979 VDD.t4138 VSS 0.324211f
C20980 VDD.t447 VSS 0.324211f
C20981 VDD.t445 VSS 0.067957f
C20982 VDD.t443 VSS 0.052737f
C20983 VDD.t3325 VSS 0.017474f
C20984 VDD.t3329 VSS 0.004807f
C20985 VDD.t3327 VSS 0.004807f
C20986 VDD.n2543 VSS 0.010696f
C20987 VDD.n2544 VSS 0.099162f
C20988 VDD.n2545 VSS 0.02587f
C20989 VDD.n2546 VSS 0.006536f
C20990 VDD.t3328 VSS 0.049198f
C20991 VDD.t3326 VSS 0.067957f
C20992 VDD.t3324 VSS 0.176263f
C20993 VDD.t94 VSS 0.176263f
C20994 VDD.t84 VSS 0.067957f
C20995 VDD.t82 VSS 0.052737f
C20996 VDD.t4109 VSS 0.067957f
C20997 VDD.t4105 VSS 0.256608f
C20998 VDD.t1562 VSS 0.256608f
C20999 VDD.t1560 VSS 0.067957f
C21000 VDD.t1558 VSS 0.049198f
C21001 VDD.t1734 VSS 0.017462f
C21002 VDD.n2547 VSS 0.092113f
C21003 VDD.t1738 VSS 0.004807f
C21004 VDD.t1736 VSS 0.004807f
C21005 VDD.n2548 VSS 0.010696f
C21006 VDD.n2549 VSS 0.036584f
C21007 VDD.t1563 VSS 0.017474f
C21008 VDD.t1559 VSS 0.004807f
C21009 VDD.t1561 VSS 0.004807f
C21010 VDD.n2550 VSS 0.010696f
C21011 VDD.n2551 VSS 0.097619f
C21012 VDD.n2552 VSS 0.024888f
C21013 VDD.n2553 VSS 0.006536f
C21014 VDD.t1735 VSS 0.052737f
C21015 VDD.t1737 VSS 0.067957f
C21016 VDD.t1733 VSS 0.176263f
C21017 VDD.t1858 VSS 0.176263f
C21018 VDD.t1854 VSS 0.067957f
C21019 VDD.t1856 VSS 0.049198f
C21020 VDD.t2190 VSS 0.017476f
C21021 VDD.t2188 VSS 0.004807f
C21022 VDD.t2186 VSS 0.004807f
C21023 VDD.n2554 VSS 0.010696f
C21024 VDD.n2555 VSS 0.098224f
C21025 VDD.n2556 VSS 0.048045f
C21026 VDD.t1859 VSS 0.017474f
C21027 VDD.t1857 VSS 0.004807f
C21028 VDD.t1855 VSS 0.004807f
C21029 VDD.n2557 VSS 0.010696f
C21030 VDD.n2558 VSS 0.099162f
C21031 VDD.n2559 VSS 0.02587f
C21032 VDD.n2560 VSS 0.006536f
C21033 VDD.t2185 VSS 0.052737f
C21034 VDD.t2187 VSS 0.067957f
C21035 VDD.t2189 VSS 0.323857f
C21036 VDD.t337 VSS 0.323857f
C21037 VDD.t341 VSS 0.067957f
C21038 VDD.t343 VSS 0.049198f
C21039 VDD.t338 VSS 0.017474f
C21040 VDD.t344 VSS 0.004807f
C21041 VDD.t342 VSS 0.004807f
C21042 VDD.n2561 VSS 0.010696f
C21043 VDD.n2562 VSS 0.099467f
C21044 VDD.n2563 VSS 0.025249f
C21045 VDD.n2564 VSS 0.006536f
C21046 VDD.t541 VSS 0.052737f
C21047 VDD.t545 VSS 0.067957f
C21048 VDD.t265 VSS 0.256608f
C21049 VDD.t2466 VSS 0.256608f
C21050 VDD.t2468 VSS 0.067957f
C21051 VDD.t2470 VSS 0.049198f
C21052 VDD.n2565 VSS 0.006536f
C21053 VDD.n2566 VSS 0.024888f
C21054 VDD.t85 VSS 0.004807f
C21055 VDD.t83 VSS 0.004807f
C21056 VDD.n2567 VSS 0.010696f
C21057 VDD.n2568 VSS 0.036584f
C21058 VDD.n2569 VSS 0.092113f
C21059 VDD.n2570 VSS 0.194608f
C21060 VDD.n2571 VSS 0.392773f
C21061 VDD.n2572 VSS 0.538951f
C21062 VDD.n2573 VSS 0.31205f
C21063 VDD.t2463 VSS 0.012354f
C21064 VDD.t2461 VSS 0.012354f
C21065 VDD.n2574 VSS 0.040938f
C21066 VDD.t2436 VSS 0.012354f
C21067 VDD.t2465 VSS 0.010856f
C21068 VDD.n2575 VSS 0.038523f
C21069 VDD.n2576 VSS 0.058757f
C21070 VDD.n2577 VSS 0.479072f
C21071 VDD.n2578 VSS -0.041546f
C21072 VDD.t1231 VSS 0.090532f
C21073 VDD.t3379 VSS 0.119055f
C21074 VDD.t1230 VSS 0.119055f
C21075 VDD.t2462 VSS 0.119055f
C21076 VDD.t2460 VSS 0.119055f
C21077 VDD.t2435 VSS 0.116575f
C21078 VDD.t2464 VSS 0.254852f
C21079 VDD.t261 VSS 0.254852f
C21080 VDD.t529 VSS 0.116575f
C21081 VDD.t267 VSS 0.119055f
C21082 VDD.t549 VSS 0.119055f
C21083 VDD.t335 VSS 0.119055f
C21084 VDD.t334 VSS 0.119055f
C21085 VDD.t336 VSS 0.088051f
C21086 VDD.t262 VSS 0.010856f
C21087 VDD.t530 VSS 0.012354f
C21088 VDD.n2579 VSS 0.038675f
C21089 VDD.t268 VSS 0.012354f
C21090 VDD.t550 VSS 0.012354f
C21091 VDD.n2580 VSS 0.040145f
C21092 VDD.n2581 VSS 0.059265f
C21093 VDD.t346 VSS 0.012354f
C21094 VDD.t340 VSS 0.012354f
C21095 VDD.n2582 VSS 0.040938f
C21096 VDD.t879 VSS 0.012354f
C21097 VDD.t877 VSS 0.010856f
C21098 VDD.n2583 VSS 0.038523f
C21099 VDD.n2584 VSS 0.058757f
C21100 VDD.n2585 VSS 0.22487f
C21101 VDD.n2586 VSS 0.479072f
C21102 VDD.n2587 VSS -0.041546f
C21103 VDD.t1518 VSS 0.090532f
C21104 VDD.t1517 VSS 0.119055f
C21105 VDD.t227 VSS 0.119055f
C21106 VDD.t345 VSS 0.119055f
C21107 VDD.t339 VSS 0.119055f
C21108 VDD.t878 VSS 0.116575f
C21109 VDD.t876 VSS 0.361506f
C21110 VDD.t1727 VSS 0.361506f
C21111 VDD.t1739 VSS 0.116575f
C21112 VDD.t1731 VSS 0.119055f
C21113 VDD.t1729 VSS 0.119055f
C21114 VDD.t2183 VSS 0.119055f
C21115 VDD.t333 VSS 0.119055f
C21116 VDD.t2184 VSS 0.088051f
C21117 VDD.t774 VSS 0.119055f
C21118 VDD.t772 VSS 0.119055f
C21119 VDD.t3946 VSS 0.119055f
C21120 VDD.t3950 VSS 0.119055f
C21121 VDD.t3938 VSS 0.116575f
C21122 VDD.t3948 VSS 0.362126f
C21123 VDD.t619 VSS 0.362126f
C21124 VDD.t621 VSS 0.116575f
C21125 VDD.t609 VSS 0.119055f
C21126 VDD.t617 VSS 0.119055f
C21127 VDD.t1576 VSS 0.119055f
C21128 VDD.t1577 VSS 0.119055f
C21129 VDD.t1575 VSS 0.090532f
C21130 VDD.t4100 VSS 0.010856f
C21131 VDD.t4122 VSS 0.012354f
C21132 VDD.n2588 VSS 0.038675f
C21133 VDD.t4102 VSS 0.012354f
C21134 VDD.t4084 VSS 0.012354f
C21135 VDD.n2589 VSS 0.040145f
C21136 VDD.n2590 VSS 0.059265f
C21137 VDD.t618 VSS 0.012354f
C21138 VDD.t610 VSS 0.012354f
C21139 VDD.n2591 VSS 0.040938f
C21140 VDD.t622 VSS 0.012354f
C21141 VDD.t620 VSS 0.010856f
C21142 VDD.n2592 VSS 0.038523f
C21143 VDD.n2593 VSS 0.058757f
C21144 VDD.n2594 VSS 0.22487f
C21145 VDD.n2595 VSS 0.479072f
C21146 VDD.n2596 VSS -0.041546f
C21147 VDD.t953 VSS 0.088051f
C21148 VDD.t954 VSS 0.119055f
C21149 VDD.t955 VSS 0.119055f
C21150 VDD.t4083 VSS 0.119055f
C21151 VDD.t4101 VSS 0.119055f
C21152 VDD.t4121 VSS 0.116575f
C21153 VDD.t4099 VSS 0.254852f
C21154 VDD.t1556 VSS 0.254852f
C21155 VDD.t1554 VSS 0.116575f
C21156 VDD.t1552 VSS 0.119055f
C21157 VDD.t1550 VSS 0.119055f
C21158 VDD.t1565 VSS 0.119055f
C21159 VDD.t1564 VSS 0.119055f
C21160 VDD.t1566 VSS 0.090532f
C21161 VDD.n2597 VSS -0.041546f
C21162 VDD.n2598 VSS 0.479072f
C21163 VDD.n2599 VSS 0.31205f
C21164 VDD.n2600 VSS 0.538951f
C21165 VDD.n2601 VSS 0.392773f
C21166 VDD.n2602 VSS 0.036461f
C21167 VDD.t612 VSS 0.017474f
C21168 VDD.t616 VSS 0.004807f
C21169 VDD.t614 VSS 0.004807f
C21170 VDD.n2603 VSS 0.010696f
C21171 VDD.n2604 VSS 0.099467f
C21172 VDD.n2605 VSS 0.025249f
C21173 VDD.n2606 VSS 0.006536f
C21174 VDD.t615 VSS 0.049198f
C21175 VDD.t613 VSS 0.067957f
C21176 VDD.t611 VSS 0.324211f
C21177 VDD.t908 VSS 0.324211f
C21178 VDD.t3464 VSS 0.067957f
C21179 VDD.t3462 VSS 0.052737f
C21180 VDD.t3995 VSS 0.017474f
C21181 VDD.t3999 VSS 0.004807f
C21182 VDD.t3997 VSS 0.004807f
C21183 VDD.n2607 VSS 0.010696f
C21184 VDD.n2608 VSS 0.099162f
C21185 VDD.n2609 VSS 0.02587f
C21186 VDD.n2610 VSS 0.006536f
C21187 VDD.t3998 VSS 0.049198f
C21188 VDD.t3996 VSS 0.067957f
C21189 VDD.t3994 VSS 0.176263f
C21190 VDD.t3940 VSS 0.176263f
C21191 VDD.t3944 VSS 0.067957f
C21192 VDD.t3942 VSS 0.052737f
C21193 VDD.t407 VSS 0.067957f
C21194 VDD.t403 VSS 0.256608f
C21195 VDD.t3908 VSS 0.256608f
C21196 VDD.t3910 VSS 0.067957f
C21197 VDD.t3906 VSS 0.049198f
C21198 VDD.t2757 VSS 0.017462f
C21199 VDD.n2611 VSS 0.092113f
C21200 VDD.t2761 VSS 0.004807f
C21201 VDD.t2759 VSS 0.004807f
C21202 VDD.n2612 VSS 0.010696f
C21203 VDD.n2613 VSS 0.036584f
C21204 VDD.t3909 VSS 0.017474f
C21205 VDD.t3907 VSS 0.004807f
C21206 VDD.t3911 VSS 0.004807f
C21207 VDD.n2614 VSS 0.010696f
C21208 VDD.n2615 VSS 0.097619f
C21209 VDD.n2616 VSS 0.024888f
C21210 VDD.n2617 VSS 0.006536f
C21211 VDD.t2758 VSS 0.052737f
C21212 VDD.t2760 VSS 0.067957f
C21213 VDD.t2756 VSS 0.176263f
C21214 VDD.t1847 VSS 0.176263f
C21215 VDD.t1849 VSS 0.067957f
C21216 VDD.t1851 VSS 0.049198f
C21217 VDD.t2701 VSS 0.017476f
C21218 VDD.t2705 VSS 0.004807f
C21219 VDD.t2703 VSS 0.004807f
C21220 VDD.n2618 VSS 0.010696f
C21221 VDD.n2619 VSS 0.098224f
C21222 VDD.n2620 VSS 0.048045f
C21223 VDD.t1848 VSS 0.017474f
C21224 VDD.t1852 VSS 0.004807f
C21225 VDD.t1850 VSS 0.004807f
C21226 VDD.n2621 VSS 0.010696f
C21227 VDD.n2622 VSS 0.099162f
C21228 VDD.n2623 VSS 0.02587f
C21229 VDD.n2624 VSS 0.006536f
C21230 VDD.t2702 VSS 0.052737f
C21231 VDD.t2704 VSS 0.067957f
C21232 VDD.t2700 VSS 0.324211f
C21233 VDD.t1435 VSS 0.324211f
C21234 VDD.t1433 VSS 0.067957f
C21235 VDD.t1431 VSS 0.049198f
C21236 VDD.t1436 VSS 0.017474f
C21237 VDD.t1432 VSS 0.004807f
C21238 VDD.t1434 VSS 0.004807f
C21239 VDD.n2625 VSS 0.010696f
C21240 VDD.n2626 VSS 0.099467f
C21241 VDD.n2627 VSS 0.025249f
C21242 VDD.n2628 VSS 0.006536f
C21243 VDD.t1627 VSS 0.052737f
C21244 VDD.t1629 VSS 0.067957f
C21245 VDD.t1625 VSS 0.256608f
C21246 VDD.t299 VSS 0.256608f
C21247 VDD.t301 VSS 0.067957f
C21248 VDD.t297 VSS 0.049198f
C21249 VDD.n2629 VSS 0.006536f
C21250 VDD.n2630 VSS 0.024888f
C21251 VDD.t3945 VSS 0.004807f
C21252 VDD.t3943 VSS 0.004807f
C21253 VDD.n2631 VSS 0.010696f
C21254 VDD.n2632 VSS 0.036584f
C21255 VDD.n2633 VSS 0.092113f
C21256 VDD.n2634 VSS 0.194608f
C21257 VDD.n2635 VSS 0.392773f
C21258 VDD.n2636 VSS 0.538951f
C21259 VDD.n2637 VSS 0.31205f
C21260 VDD.t348 VSS 0.012354f
C21261 VDD.t304 VSS 0.012354f
C21262 VDD.n2638 VSS 0.040938f
C21263 VDD.t352 VSS 0.012354f
C21264 VDD.t350 VSS 0.010856f
C21265 VDD.n2639 VSS 0.038523f
C21266 VDD.n2640 VSS 0.058757f
C21267 VDD.n2641 VSS 0.479072f
C21268 VDD.n2642 VSS -0.041546f
C21269 VDD.t1164 VSS 0.090532f
C21270 VDD.t2076 VSS 0.119055f
C21271 VDD.t2747 VSS 0.119055f
C21272 VDD.t347 VSS 0.119055f
C21273 VDD.t303 VSS 0.119055f
C21274 VDD.t351 VSS 0.116575f
C21275 VDD.t349 VSS 0.254852f
C21276 VDD.t1638 VSS 0.254852f
C21277 VDD.t2201 VSS 0.116575f
C21278 VDD.t2191 VSS 0.119055f
C21279 VDD.t1635 VSS 0.119055f
C21280 VDD.t557 VSS 0.119055f
C21281 VDD.t559 VSS 0.119055f
C21282 VDD.t558 VSS 0.088051f
C21283 VDD.t1639 VSS 0.010856f
C21284 VDD.t2202 VSS 0.012354f
C21285 VDD.n2643 VSS 0.038675f
C21286 VDD.t2192 VSS 0.012354f
C21287 VDD.t1636 VSS 0.012354f
C21288 VDD.n2644 VSS 0.040145f
C21289 VDD.n2645 VSS 0.059265f
C21290 VDD.t1428 VSS 0.012354f
C21291 VDD.t1430 VSS 0.012354f
C21292 VDD.n2646 VSS 0.040938f
C21293 VDD.t1438 VSS 0.012354f
C21294 VDD.t1426 VSS 0.010856f
C21295 VDD.n2647 VSS 0.038523f
C21296 VDD.n2648 VSS 0.058757f
C21297 VDD.n2649 VSS 0.22487f
C21298 VDD.n2650 VSS 0.479072f
C21299 VDD.n2651 VSS -0.041546f
C21300 VDD.t3375 VSS 0.090532f
C21301 VDD.t3377 VSS 0.119055f
C21302 VDD.t3376 VSS 0.119055f
C21303 VDD.t1427 VSS 0.119055f
C21304 VDD.t1429 VSS 0.119055f
C21305 VDD.t1437 VSS 0.116575f
C21306 VDD.t1425 VSS 0.362126f
C21307 VDD.t2752 VSS 0.362126f
C21308 VDD.t2748 VSS 0.116575f
C21309 VDD.t2754 VSS 0.119055f
C21310 VDD.t2750 VSS 0.119055f
C21311 VDD.t1483 VSS 0.119055f
C21312 VDD.t1485 VSS 0.119055f
C21313 VDD.t1484 VSS 0.088051f
C21314 VDD.t1448 VSS 0.119055f
C21315 VDD.t1449 VSS 0.119055f
C21316 VDD.t1146 VSS 0.119055f
C21317 VDD.t1123 VSS 0.119055f
C21318 VDD.t1144 VSS 0.116575f
C21319 VDD.t1115 VSS 0.362126f
C21320 VDD.t2884 VSS 0.362126f
C21321 VDD.t2874 VSS 0.116575f
C21322 VDD.t2872 VSS 0.119055f
C21323 VDD.t2876 VSS 0.119055f
C21324 VDD.t3897 VSS 0.119055f
C21325 VDD.t3898 VSS 0.119055f
C21326 VDD.t3899 VSS 0.090532f
C21327 VDD.t392 VSS 0.010856f
C21328 VDD.t388 VSS 0.012354f
C21329 VDD.n2652 VSS 0.038675f
C21330 VDD.t380 VSS 0.012354f
C21331 VDD.t396 VSS 0.012354f
C21332 VDD.n2653 VSS 0.040145f
C21333 VDD.n2654 VSS 0.059265f
C21334 VDD.t2877 VSS 0.012354f
C21335 VDD.t2873 VSS 0.012354f
C21336 VDD.n2655 VSS 0.040938f
C21337 VDD.t2875 VSS 0.012354f
C21338 VDD.t2885 VSS 0.010856f
C21339 VDD.n2656 VSS 0.038523f
C21340 VDD.n2657 VSS 0.058757f
C21341 VDD.n2658 VSS 0.22487f
C21342 VDD.n2659 VSS 0.479072f
C21343 VDD.n2660 VSS -0.041546f
C21344 VDD.t2047 VSS 0.088051f
C21345 VDD.t2045 VSS 0.119055f
C21346 VDD.t2046 VSS 0.119055f
C21347 VDD.t395 VSS 0.119055f
C21348 VDD.t379 VSS 0.119055f
C21349 VDD.t387 VSS 0.116575f
C21350 VDD.t391 VSS 0.254852f
C21351 VDD.t3902 VSS 0.254852f
C21352 VDD.t3912 VSS 0.116575f
C21353 VDD.t3900 VSS 0.119055f
C21354 VDD.t3904 VSS 0.119055f
C21355 VDD.t141 VSS 0.119055f
C21356 VDD.t139 VSS 0.119055f
C21357 VDD.t140 VSS 0.090532f
C21358 VDD.n2661 VSS -0.041546f
C21359 VDD.n2662 VSS 0.479072f
C21360 VDD.n2663 VSS 0.31205f
C21361 VDD.n2664 VSS 0.538951f
C21362 VDD.n2665 VSS 0.392773f
C21363 VDD.n2666 VSS 0.036461f
C21364 VDD.t2881 VSS 0.017474f
C21365 VDD.t2879 VSS 0.004807f
C21366 VDD.t2883 VSS 0.004807f
C21367 VDD.n2667 VSS 0.010696f
C21368 VDD.n2668 VSS 0.099467f
C21369 VDD.n2669 VSS 0.025249f
C21370 VDD.n2670 VSS 0.006536f
C21371 VDD.t2878 VSS 0.049198f
C21372 VDD.t2882 VSS 0.067957f
C21373 VDD.t2880 VSS 0.324211f
C21374 VDD.t2472 VSS 0.324211f
C21375 VDD.t2476 VSS 0.067957f
C21376 VDD.t2474 VSS 0.052737f
C21377 VDD.t1585 VSS 0.017474f
C21378 VDD.t1583 VSS 0.004807f
C21379 VDD.t1587 VSS 0.004807f
C21380 VDD.n2671 VSS 0.010696f
C21381 VDD.n2672 VSS 0.099162f
C21382 VDD.n2673 VSS 0.02587f
C21383 VDD.n2674 VSS 0.006536f
C21384 VDD.t1582 VSS 0.049198f
C21385 VDD.t1586 VSS 0.067957f
C21386 VDD.t1584 VSS 0.176263f
C21387 VDD.t1119 VSS 0.176263f
C21388 VDD.t1117 VSS 0.067957f
C21389 VDD.t1121 VSS 0.052737f
C21390 VDD.t2690 VSS 0.049198f
C21391 VDD.t1841 VSS 0.017476f
C21392 VDD.t1845 VSS 0.004807f
C21393 VDD.t1843 VSS 0.004807f
C21394 VDD.n2675 VSS 0.010696f
C21395 VDD.n2676 VSS 0.098224f
C21396 VDD.n2677 VSS 0.392773f
C21397 VDD.t171 VSS 0.017462f
C21398 VDD.t3476 VSS 0.017474f
C21399 VDD.t3474 VSS 0.004807f
C21400 VDD.t3480 VSS 0.004807f
C21401 VDD.n2678 VSS 0.010696f
C21402 VDD.n2679 VSS 0.097619f
C21403 VDD.t2694 VSS 0.067957f
C21404 VDD.t2692 VSS 0.176263f
C21405 VDD.t170 VSS 0.176263f
C21406 VDD.t1878 VSS 0.067957f
C21407 VDD.t1880 VSS 0.052737f
C21408 VDD.t3647 VSS 0.454462f
C21409 VDD.t3649 VSS 0.067957f
C21410 VDD.t3643 VSS 0.049198f
C21411 VDD.t3433 VSS 0.017476f
C21412 VDD.t3431 VSS 0.004807f
C21413 VDD.t3437 VSS 0.004807f
C21414 VDD.n2680 VSS 0.010696f
C21415 VDD.n2681 VSS 0.099623f
C21416 VDD.n2682 VSS 0.036461f
C21417 VDD.t3648 VSS 0.017474f
C21418 VDD.t3644 VSS 0.004807f
C21419 VDD.t3650 VSS 0.004807f
C21420 VDD.n2683 VSS 0.010696f
C21421 VDD.n2684 VSS 0.099467f
C21422 VDD.n2685 VSS 0.025249f
C21423 VDD.n2686 VSS 0.006536f
C21424 VDD.t3436 VSS 0.052737f
C21425 VDD.t3430 VSS 0.067957f
C21426 VDD.t3432 VSS 0.256608f
C21427 VDD.t3475 VSS 0.256608f
C21428 VDD.t3479 VSS 0.067957f
C21429 VDD.t3473 VSS 0.049198f
C21430 VDD.n2687 VSS 0.006536f
C21431 VDD.n2688 VSS 0.024888f
C21432 VDD.t1879 VSS 0.004807f
C21433 VDD.t1881 VSS 0.004807f
C21434 VDD.n2689 VSS 0.010696f
C21435 VDD.n2690 VSS 0.036584f
C21436 VDD.n2691 VSS 0.092113f
C21437 VDD.n2692 VSS 0.194608f
C21438 VDD.n2693 VSS 0.048045f
C21439 VDD.t2693 VSS 0.017474f
C21440 VDD.t2691 VSS 0.004807f
C21441 VDD.t2695 VSS 0.004807f
C21442 VDD.n2694 VSS 0.010696f
C21443 VDD.n2695 VSS 0.099162f
C21444 VDD.n2696 VSS 0.02587f
C21445 VDD.n2697 VSS 0.006536f
C21446 VDD.t1842 VSS 0.052737f
C21447 VDD.t1844 VSS 0.067957f
C21448 VDD.t1840 VSS 0.324211f
C21449 VDD.t3240 VSS 0.324211f
C21450 VDD.t3242 VSS 0.067957f
C21451 VDD.t3238 VSS 0.049198f
C21452 VDD.t2837 VSS 0.017476f
C21453 VDD.t2842 VSS 0.004807f
C21454 VDD.t2840 VSS 0.004807f
C21455 VDD.n2698 VSS 0.010696f
C21456 VDD.n2699 VSS 0.099623f
C21457 VDD.n2700 VSS 0.033339f
C21458 VDD.t3241 VSS 0.017474f
C21459 VDD.t3239 VSS 0.004807f
C21460 VDD.t3243 VSS 0.004807f
C21461 VDD.n2701 VSS 0.010696f
C21462 VDD.n2702 VSS 0.099467f
C21463 VDD.n2703 VSS 0.025249f
C21464 VDD.n2704 VSS 0.006536f
C21465 VDD.t2839 VSS 0.052737f
C21466 VDD.t2841 VSS 0.067957f
C21467 VDD.t2836 VSS 0.256608f
C21468 VDD.t2405 VSS 0.256608f
C21469 VDD.t2407 VSS 0.067957f
C21470 VDD.t2401 VSS 0.049198f
C21471 VDD.n2705 VSS 0.006536f
C21472 VDD.n2706 VSS 0.024888f
C21473 VDD.t1118 VSS 0.004807f
C21474 VDD.t1122 VSS 0.004807f
C21475 VDD.n2707 VSS 0.010696f
C21476 VDD.n2708 VSS 0.036584f
C21477 VDD.n2709 VSS 0.092113f
C21478 VDD.n2710 VSS 0.194608f
C21479 VDD.n2711 VSS 0.249152f
C21480 VDD.n2712 VSS 0.538951f
C21481 VDD.n2713 VSS 0.31205f
C21482 VDD.t2400 VSS 0.012354f
C21483 VDD.t823 VSS 0.012354f
C21484 VDD.n2714 VSS 0.040938f
C21485 VDD.t2410 VSS 0.012354f
C21486 VDD.t2404 VSS 0.010856f
C21487 VDD.n2715 VSS 0.038523f
C21488 VDD.n2716 VSS 0.058757f
C21489 VDD.n2717 VSS 0.479072f
C21490 VDD.n2718 VSS -0.041546f
C21491 VDD.t2648 VSS 0.090532f
C21492 VDD.t1544 VSS 0.119055f
C21493 VDD.t1494 VSS 0.119055f
C21494 VDD.t2399 VSS 0.119055f
C21495 VDD.t822 VSS 0.119055f
C21496 VDD.t2409 VSS 0.116575f
C21497 VDD.t2403 VSS 0.254852f
C21498 VDD.t2823 VSS 0.254852f
C21499 VDD.t2817 VSS 0.116575f
C21500 VDD.t2834 VSS 0.119055f
C21501 VDD.t2827 VSS 0.119055f
C21502 VDD.t1216 VSS 0.119055f
C21503 VDD.t1215 VSS 0.119055f
C21504 VDD.t1217 VSS 0.088051f
C21505 VDD.t2824 VSS 0.010856f
C21506 VDD.t2818 VSS 0.012354f
C21507 VDD.n2719 VSS 0.038675f
C21508 VDD.t2835 VSS 0.012354f
C21509 VDD.t2828 VSS 0.012354f
C21510 VDD.n2720 VSS 0.040145f
C21511 VDD.n2721 VSS 0.059265f
C21512 VDD.t3233 VSS 0.012354f
C21513 VDD.t3237 VSS 0.012354f
C21514 VDD.n2722 VSS 0.040938f
C21515 VDD.t3235 VSS 0.012354f
C21516 VDD.t3245 VSS 0.010856f
C21517 VDD.n2723 VSS 0.038523f
C21518 VDD.n2724 VSS 0.058757f
C21519 VDD.n2725 VSS 0.22487f
C21520 VDD.n2726 VSS 0.479072f
C21521 VDD.n2727 VSS -0.041546f
C21522 VDD.t1196 VSS 0.090532f
C21523 VDD.t724 VSS 0.119055f
C21524 VDD.t1195 VSS 0.119055f
C21525 VDD.t3232 VSS 0.119055f
C21526 VDD.t3236 VSS 0.119055f
C21527 VDD.t3234 VSS 0.116575f
C21528 VDD.t3244 VSS 0.362126f
C21529 VDD.t1876 VSS 0.362126f
C21530 VDD.t1874 VSS 0.116575f
C21531 VDD.t1872 VSS 0.119055f
C21532 VDD.t172 VSS 0.119055f
C21533 VDD.t1618 VSS 0.119055f
C21534 VDD.t1617 VSS 0.119055f
C21535 VDD.t1619 VSS 0.088051f
C21536 VDD.t1877 VSS 0.010856f
C21537 VDD.t1875 VSS 0.012354f
C21538 VDD.n2728 VSS 0.038675f
C21539 VDD.t1873 VSS 0.012354f
C21540 VDD.t173 VSS 0.012354f
C21541 VDD.n2729 VSS 0.040145f
C21542 VDD.n2730 VSS 0.059265f
C21543 VDD.n2731 VSS 0.31205f
C21544 VDD.t3478 VSS 0.012354f
C21545 VDD.t3470 VSS 0.012354f
C21546 VDD.n2732 VSS 0.040938f
C21547 VDD.t3472 VSS 0.012354f
C21548 VDD.t3468 VSS 0.010856f
C21549 VDD.n2733 VSS 0.038523f
C21550 VDD.n2734 VSS 0.058757f
C21551 VDD.n2735 VSS 0.479072f
C21552 VDD.n2736 VSS -0.041546f
C21553 VDD.t2488 VSS 0.090532f
C21554 VDD.t2487 VSS 0.119055f
C21555 VDD.t2489 VSS 0.119055f
C21556 VDD.t3477 VSS 0.119055f
C21557 VDD.t3469 VSS 0.119055f
C21558 VDD.t3471 VSS 0.116575f
C21559 VDD.t3467 VSS 0.254852f
C21560 VDD.t3440 VSS 0.254852f
C21561 VDD.t3427 VSS 0.116575f
C21562 VDD.t3421 VSS 0.119055f
C21563 VDD.t3444 VSS 0.119055f
C21564 VDD.t3882 VSS 0.119055f
C21565 VDD.t3881 VSS 0.119055f
C21566 VDD.t3880 VSS 0.088051f
C21567 VDD.t3651 VSS 0.532028f
C21568 VDD.t3641 VSS 0.116575f
C21569 VDD.t3645 VSS 0.119055f
C21570 VDD.t3639 VSS 0.119055f
C21571 VDD.t58 VSS 0.119055f
C21572 VDD.t3466 VSS 0.119055f
C21573 VDD.t57 VSS 0.090532f
C21574 VDD.n2737 VSS -0.041546f
C21575 VDD.t3640 VSS 0.012354f
C21576 VDD.t3646 VSS 0.012354f
C21577 VDD.n2738 VSS 0.040938f
C21578 VDD.t3642 VSS 0.012354f
C21579 VDD.t3652 VSS 0.010856f
C21580 VDD.n2739 VSS 0.038523f
C21581 VDD.n2740 VSS 0.058757f
C21582 VDD.n2741 VSS 0.479072f
C21583 VDD.n2742 VSS 0.22487f
C21584 VDD.n2743 VSS 0.282509f
C21585 VDD.t1175 VSS 0.010856f
C21586 VDD.t1409 VSS 0.012354f
C21587 VDD.n2744 VSS 0.038523f
C21588 VDD.t1405 VSS 0.012354f
C21589 VDD.t1387 VSS 0.012354f
C21590 VDD.n2745 VSS 0.040938f
C21591 VDD.n2746 VSS 0.058757f
C21592 VDD.t1174 VSS 0.189904f
C21593 VDD.t1408 VSS 0.115167f
C21594 VDD.t1404 VSS 0.117618f
C21595 VDD.t1386 VSS 0.117618f
C21596 VDD.t2413 VSS 0.117618f
C21597 VDD.t2412 VSS 0.117618f
C21598 VDD.t2411 VSS 0.089438f
C21599 VDD.t1789 VSS 0.189904f
C21600 VDD.t1771 VSS 0.115167f
C21601 VDD.t1811 VSS 0.117618f
C21602 VDD.t1745 VSS 0.117618f
C21603 VDD.t3698 VSS 0.117618f
C21604 VDD.t3699 VSS 0.117618f
C21605 VDD.t3697 VSS 0.086988f
C21606 VDD.n2747 VSS -0.042265f
C21607 VDD.t1746 VSS 0.012354f
C21608 VDD.t1812 VSS 0.012354f
C21609 VDD.n2748 VSS 0.040145f
C21610 VDD.t1772 VSS 0.012354f
C21611 VDD.t1790 VSS 0.010856f
C21612 VDD.n2749 VSS 0.038675f
C21613 VDD.n2750 VSS 0.059265f
C21614 VDD.n2751 VSS 0.479072f
C21615 VDD.n2752 VSS 0.216809f
C21616 VDD.n2753 VSS 0.684805f
C21617 VDD.n2754 VSS 0.801769f
C21618 VDD.t3530 VSS 0.010856f
C21619 VDD.t3555 VSS 0.012354f
C21620 VDD.n2755 VSS 0.038523f
C21621 VDD.t3534 VSS 0.012354f
C21622 VDD.t3565 VSS 0.012354f
C21623 VDD.n2756 VSS 0.040938f
C21624 VDD.n2757 VSS 0.058757f
C21625 VDD.t3529 VSS 0.189904f
C21626 VDD.t3554 VSS 0.115167f
C21627 VDD.t3533 VSS 0.117618f
C21628 VDD.t3564 VSS 0.117618f
C21629 VDD.t2689 VSS 0.117618f
C21630 VDD.t2688 VSS 0.117618f
C21631 VDD.t2687 VSS 0.089438f
C21632 VDD.t1753 VSS 0.189904f
C21633 VDD.t1765 VSS 0.115167f
C21634 VDD.t1807 VSS 0.117618f
C21635 VDD.t766 VSS 0.117618f
C21636 VDD.t4276 VSS 0.117618f
C21637 VDD.t4277 VSS 0.117618f
C21638 VDD.t4278 VSS 0.086988f
C21639 VDD.n2758 VSS -0.042265f
C21640 VDD.t767 VSS 0.012354f
C21641 VDD.t1808 VSS 0.012354f
C21642 VDD.n2759 VSS 0.040145f
C21643 VDD.t1766 VSS 0.012354f
C21644 VDD.t1754 VSS 0.010856f
C21645 VDD.n2760 VSS 0.038675f
C21646 VDD.n2761 VSS 0.059265f
C21647 VDD.n2762 VSS 0.479072f
C21648 VDD.n2763 VSS 0.216809f
C21649 VDD.n2764 VSS 0.684805f
C21650 VDD.n2765 VSS 0.801769f
C21651 VDD.t3973 VSS 0.010856f
C21652 VDD.t3967 VSS 0.012354f
C21653 VDD.n2766 VSS 0.038523f
C21654 VDD.t892 VSS 0.012354f
C21655 VDD.t3982 VSS 0.012354f
C21656 VDD.n2767 VSS 0.040938f
C21657 VDD.n2768 VSS 0.058757f
C21658 VDD.t3972 VSS 0.189904f
C21659 VDD.t3966 VSS 0.115167f
C21660 VDD.t891 VSS 0.117618f
C21661 VDD.t3981 VSS 0.117618f
C21662 VDD.t2855 VSS 0.117618f
C21663 VDD.t2886 VSS 0.117618f
C21664 VDD.t2856 VSS 0.089438f
C21665 VDD.t777 VSS 0.189904f
C21666 VDD.t1773 VSS 0.115167f
C21667 VDD.t1797 VSS 0.117618f
C21668 VDD.t1809 VSS 0.117618f
C21669 VDD.t2854 VSS 0.117618f
C21670 VDD.t1143 VSS 0.117618f
C21671 VDD.t1142 VSS 0.086988f
C21672 VDD.n2769 VSS -0.042265f
C21673 VDD.t1810 VSS 0.012354f
C21674 VDD.t1798 VSS 0.012354f
C21675 VDD.n2770 VSS 0.040145f
C21676 VDD.t1774 VSS 0.012354f
C21677 VDD.t778 VSS 0.010856f
C21678 VDD.n2771 VSS 0.038675f
C21679 VDD.n2772 VSS 0.059265f
C21680 VDD.n2773 VSS 0.479072f
C21681 VDD.n2774 VSS 0.216809f
C21682 VDD.n2775 VSS 0.480721f
C21683 VDD.n2776 VSS 0.460498f
C21684 VDD.t3597 VSS 0.010856f
C21685 VDD.t3603 VSS 0.012354f
C21686 VDD.n2777 VSS 0.038523f
C21687 VDD.t3583 VSS 0.012354f
C21688 VDD.t3616 VSS 0.012354f
C21689 VDD.n2778 VSS 0.040938f
C21690 VDD.n2779 VSS 0.058757f
C21691 VDD.t3596 VSS 0.189904f
C21692 VDD.t3602 VSS 0.115167f
C21693 VDD.t3582 VSS 0.117618f
C21694 VDD.t3615 VSS 0.117618f
C21695 VDD.t2730 VSS 0.117618f
C21696 VDD.t2731 VSS 0.117618f
C21697 VDD.t2729 VSS 0.089438f
C21698 VDD.t1813 VSS 0.189904f
C21699 VDD.t1747 VSS 0.115167f
C21700 VDD.t1795 VSS 0.117618f
C21701 VDD.t1785 VSS 0.117618f
C21702 VDD.t1614 VSS 0.117618f
C21703 VDD.t1531 VSS 0.117618f
C21704 VDD.t1613 VSS 0.086988f
C21705 VDD.n2780 VSS -0.042265f
C21706 VDD.t1786 VSS 0.012354f
C21707 VDD.t1796 VSS 0.012354f
C21708 VDD.n2781 VSS 0.040145f
C21709 VDD.t1748 VSS 0.012354f
C21710 VDD.t1814 VSS 0.010856f
C21711 VDD.n2782 VSS 0.038675f
C21712 VDD.n2783 VSS 0.059265f
C21713 VDD.n2784 VSS 0.479072f
C21714 VDD.n2785 VSS 0.216809f
C21715 VDD.n2786 VSS 0.684805f
C21716 VDD.n2787 VSS 0.801769f
C21717 VDD.t2156 VSS 0.010856f
C21718 VDD.t2131 VSS 0.012354f
C21719 VDD.n2788 VSS 0.038523f
C21720 VDD.t2120 VSS 0.012354f
C21721 VDD.t2169 VSS 0.012354f
C21722 VDD.n2789 VSS 0.040938f
C21723 VDD.n2790 VSS 0.058757f
C21724 VDD.t2155 VSS 0.189904f
C21725 VDD.t2130 VSS 0.115167f
C21726 VDD.t2119 VSS 0.117618f
C21727 VDD.t2168 VSS 0.117618f
C21728 VDD.t684 VSS 0.117618f
C21729 VDD.t683 VSS 0.117618f
C21730 VDD.t685 VSS 0.089438f
C21731 VDD.t1757 VSS 0.189904f
C21732 VDD.t1805 VSS 0.115167f
C21733 VDD.t779 VSS 0.117618f
C21734 VDD.t1779 VSS 0.117618f
C21735 VDD.t3381 VSS 0.117618f
C21736 VDD.t1446 VSS 0.117618f
C21737 VDD.t1447 VSS 0.086988f
C21738 VDD.n2791 VSS -0.042265f
C21739 VDD.t1780 VSS 0.012354f
C21740 VDD.t780 VSS 0.012354f
C21741 VDD.n2792 VSS 0.040145f
C21742 VDD.t1806 VSS 0.012354f
C21743 VDD.t1758 VSS 0.010856f
C21744 VDD.n2793 VSS 0.038675f
C21745 VDD.n2794 VSS 0.059265f
C21746 VDD.n2795 VSS 0.479072f
C21747 VDD.n2796 VSS 0.216809f
C21748 VDD.n2797 VSS 0.684592f
C21749 VDD.n2798 VSS 0.801557f
C21750 VDD.t2574 VSS 0.010856f
C21751 VDD.t2604 VSS 0.012354f
C21752 VDD.n2799 VSS 0.038523f
C21753 VDD.t2595 VSS 0.012354f
C21754 VDD.t2580 VSS 0.012354f
C21755 VDD.n2800 VSS 0.040938f
C21756 VDD.n2801 VSS 0.058757f
C21757 VDD.t2573 VSS 0.189904f
C21758 VDD.t2603 VSS 0.115167f
C21759 VDD.t2594 VSS 0.117618f
C21760 VDD.t2579 VSS 0.117618f
C21761 VDD.t3986 VSS 0.117618f
C21762 VDD.t3985 VSS 0.117618f
C21763 VDD.t3987 VSS 0.089438f
C21764 VDD.t762 VSS 0.189904f
C21765 VDD.t1783 VSS 0.115167f
C21766 VDD.t1803 VSS 0.117618f
C21767 VDD.t1755 VSS 0.117618f
C21768 VDD.t3959 VSS 0.117618f
C21769 VDD.t3960 VSS 0.117618f
C21770 VDD.t3958 VSS 0.086988f
C21771 VDD.n2802 VSS -0.042265f
C21772 VDD.t1756 VSS 0.012354f
C21773 VDD.t1804 VSS 0.012354f
C21774 VDD.n2803 VSS 0.040145f
C21775 VDD.t1784 VSS 0.012354f
C21776 VDD.t763 VSS 0.010856f
C21777 VDD.n2804 VSS 0.038675f
C21778 VDD.n2805 VSS 0.059265f
C21779 VDD.n2806 VSS 0.479072f
C21780 VDD.n2807 VSS 0.216809f
C21781 VDD.n2808 VSS 0.684805f
C21782 VDD.n2809 VSS 0.801769f
C21783 VDD.t1834 VSS 0.010856f
C21784 VDD.t2354 VSS 0.012354f
C21785 VDD.n2810 VSS 0.038523f
C21786 VDD.t2342 VSS 0.012354f
C21787 VDD.t2325 VSS 0.012354f
C21788 VDD.n2811 VSS 0.040938f
C21789 VDD.n2812 VSS 0.058757f
C21790 VDD.t1833 VSS 0.189904f
C21791 VDD.t2353 VSS 0.115167f
C21792 VDD.t2341 VSS 0.117618f
C21793 VDD.t2324 VSS 0.117618f
C21794 VDD.t1199 VSS 0.117618f
C21795 VDD.t1198 VSS 0.117618f
C21796 VDD.t1200 VSS 0.089438f
C21797 VDD.t781 VSS 0.189904f
C21798 VDD.t1777 VSS 0.115167f
C21799 VDD.t1799 VSS 0.117618f
C21800 VDD.t1749 VSS 0.117618f
C21801 VDD.t4185 VSS 0.117618f
C21802 VDD.t3952 VSS 0.117618f
C21803 VDD.t3953 VSS 0.086988f
C21804 VDD.n2813 VSS -0.042265f
C21805 VDD.t1750 VSS 0.012354f
C21806 VDD.t1800 VSS 0.012354f
C21807 VDD.n2814 VSS 0.040145f
C21808 VDD.t1778 VSS 0.012354f
C21809 VDD.t782 VSS 0.010856f
C21810 VDD.n2815 VSS 0.038675f
C21811 VDD.n2816 VSS 0.059265f
C21812 VDD.n2817 VSS 0.479072f
C21813 VDD.n2818 VSS 0.216809f
C21814 VDD.n2819 VSS 0.684805f
C21815 VDD.n2820 VSS 0.801769f
C21816 VDD.t586 VSS 0.010856f
C21817 VDD.t1005 VSS 0.012354f
C21818 VDD.n2821 VSS 0.038523f
C21819 VDD.t994 VSS 0.012354f
C21820 VDD.t1033 VSS 0.012354f
C21821 VDD.n2822 VSS 0.040938f
C21822 VDD.n2823 VSS 0.058757f
C21823 VDD.t585 VSS 0.189904f
C21824 VDD.t1004 VSS 0.115167f
C21825 VDD.t993 VSS 0.117618f
C21826 VDD.t1032 VSS 0.117618f
C21827 VDD.t2081 VSS 0.117618f
C21828 VDD.t1645 VSS 0.117618f
C21829 VDD.t1644 VSS 0.089438f
C21830 VDD.t775 VSS 0.189904f
C21831 VDD.t1763 VSS 0.115167f
C21832 VDD.t1791 VSS 0.117618f
C21833 VDD.t764 VSS 0.117618f
C21834 VDD.t918 VSS 0.117618f
C21835 VDD.t919 VSS 0.117618f
C21836 VDD.t920 VSS 0.086988f
C21837 VDD.n2824 VSS -0.042265f
C21838 VDD.t765 VSS 0.012354f
C21839 VDD.t1792 VSS 0.012354f
C21840 VDD.n2825 VSS 0.040145f
C21841 VDD.t1764 VSS 0.012354f
C21842 VDD.t776 VSS 0.010856f
C21843 VDD.n2826 VSS 0.038675f
C21844 VDD.n2827 VSS 0.059265f
C21845 VDD.n2828 VSS 0.479072f
C21846 VDD.n2829 VSS 0.216809f
C21847 VDD.n2830 VSS 1.22927f
C21848 VDD.n2831 VSS 1.17052f
C21849 VDD.n2832 VSS 0.22487f
C21850 VDD.t2293 VSS 0.012354f
C21851 VDD.t3418 VSS 0.012354f
C21852 VDD.n2833 VSS 0.040938f
C21853 VDD.t3426 VSS 0.012354f
C21854 VDD.t3451 VSS 0.010856f
C21855 VDD.n2834 VSS 0.038523f
C21856 VDD.n2835 VSS 0.058757f
C21857 VDD.n2836 VSS 0.479072f
C21858 VDD.n2837 VSS -0.0422f
C21859 VDD.t2771 VSS 0.087085f
C21860 VDD.t2770 VSS 0.117748f
C21861 VDD.t2769 VSS 0.117748f
C21862 VDD.t1384 VSS 0.117748f
C21863 VDD.t1410 VSS 0.117748f
C21864 VDD.t1406 VSS 0.115295f
C21865 VDD.t1391 VSS 0.280879f
C21866 VDD.t1781 VSS 0.280879f
C21867 VDD.t783 VSS 0.115295f
C21868 VDD.t1787 VSS 0.117748f
C21869 VDD.t1759 VSS 0.117748f
C21870 VDD.t1096 VSS 0.117748f
C21871 VDD.t1098 VSS 0.117748f
C21872 VDD.t1097 VSS 0.089538f
C21873 VDD.t979 VSS 0.010856f
C21874 VDD.t981 VSS 0.012354f
C21875 VDD.n2838 VSS 0.038675f
C21876 VDD.t975 VSS 0.012354f
C21877 VDD.t977 VSS 0.012354f
C21878 VDD.n2839 VSS 0.040145f
C21879 VDD.n2840 VSS 0.059265f
C21880 VDD.n2841 VSS 0.22487f
C21881 VDD.t1760 VSS 0.012354f
C21882 VDD.t1788 VSS 0.012354f
C21883 VDD.n2842 VSS 0.040938f
C21884 VDD.t784 VSS 0.012354f
C21885 VDD.t1782 VSS 0.010856f
C21886 VDD.n2843 VSS 0.038523f
C21887 VDD.n2844 VSS 0.058757f
C21888 VDD.n2845 VSS 0.479072f
C21889 VDD.n2846 VSS -0.0422f
C21890 VDD.t488 VSS 0.087085f
C21891 VDD.t487 VSS 0.117748f
C21892 VDD.t489 VSS 0.117748f
C21893 VDD.t976 VSS 0.117748f
C21894 VDD.t974 VSS 0.117748f
C21895 VDD.t980 VSS 0.115295f
C21896 VDD.t978 VSS 0.340811f
C21897 VDD.t3423 VSS 0.340811f
C21898 VDD.t3447 VSS 0.115295f
C21899 VDD.t3438 VSS 0.117748f
C21900 VDD.t2294 VSS 0.117748f
C21901 VDD.t1907 VSS 0.117748f
C21902 VDD.t1906 VSS 0.117748f
C21903 VDD.t2106 VSS 0.089538f
C21904 VDD.n2847 VSS -0.0422f
C21905 VDD.t2295 VSS 0.012354f
C21906 VDD.t3439 VSS 0.012354f
C21907 VDD.n2848 VSS 0.040938f
C21908 VDD.t3448 VSS 0.012354f
C21909 VDD.t3424 VSS 0.010856f
C21910 VDD.n2849 VSS 0.038523f
C21911 VDD.n2850 VSS 0.058757f
C21912 VDD.n2851 VSS 0.323668f
C21913 VDD.n2852 VSS 0.22487f
C21914 VDD.n2853 VSS 1.03891f
C21915 VDD.n2854 VSS 10.9661f
C21916 VDD.n2855 VSS 0.580841f
C21917 VDD.n2856 VSS 0.734784f
C21918 VDD.t1502 VSS 0.027215f
C21919 VDD.t1069 VSS 0.007233f
C21920 VDD.t1500 VSS 0.007233f
C21921 VDD.n2857 VSS 0.016652f
C21922 VDD.n2858 VSS 0.129639f
C21923 VDD.t1255 VSS -0.019301f
C21924 VDD.t1257 VSS 0.075145f
C21925 VDD.t2066 VSS 0.075145f
C21926 VDD.t2068 VSS 0.063403f
C21927 VDD.t1965 VSS 0.027215f
C21928 VDD.t1923 VSS 0.007233f
C21929 VDD.t2924 VSS 0.007233f
C21930 VDD.n2859 VSS 0.016652f
C21931 VDD.n2860 VSS 0.132756f
C21932 VDD.t3077 VSS 0.007233f
C21933 VDD.t647 VSS 0.007233f
C21934 VDD.n2861 VSS 0.016652f
C21935 VDD.n2862 VSS 0.047679f
C21936 VDD.t655 VSS 0.007233f
C21937 VDD.t3794 VSS 0.007233f
C21938 VDD.n2863 VSS 0.016652f
C21939 VDD.n2864 VSS 0.073624f
C21940 VDD.t646 VSS 0.04195f
C21941 VDD.t650 VSS 0.075275f
C21942 VDD.t3759 VSS 0.075275f
C21943 VDD.t3785 VSS 0.139181f
C21944 VDD.t1950 VSS 0.139181f
C21945 VDD.t1908 VSS 0.075275f
C21946 VDD.t848 VSS 0.075275f
C21947 VDD.t850 VSS 0.063514f
C21948 VDD.t3820 VSS 0.027188f
C21949 VDD.n2865 VSS 0.07466f
C21950 VDD.t2512 VSS 0.027188f
C21951 VDD.n2866 VSS 0.074656f
C21952 VDD.t2514 VSS 0.007233f
C21953 VDD.t3047 VSS 0.007233f
C21954 VDD.n2867 VSS 0.016652f
C21955 VDD.n2868 VSS 0.076601f
C21956 VDD.t2932 VSS 0.007233f
C21957 VDD.t4342 VSS 0.007233f
C21958 VDD.n2869 VSS 0.016652f
C21959 VDD.n2870 VSS 0.047822f
C21960 VDD.t3781 VSS 0.027215f
C21961 VDD.t4494 VSS 0.007233f
C21962 VDD.t3873 VSS 0.007233f
C21963 VDD.n2871 VSS 0.016652f
C21964 VDD.n2872 VSS 0.130541f
C21965 VDD.t4341 VSS 0.04195f
C21966 VDD.t4472 VSS 0.075275f
C21967 VDD.t3840 VSS 0.075275f
C21968 VDD.t3870 VSS 0.145846f
C21969 VDD.t1683 VSS 0.145846f
C21970 VDD.t1685 VSS 0.075275f
C21971 VDD.t860 VSS 0.075275f
C21972 VDD.t846 VSS 0.063514f
C21973 VDD.t3780 VSS 0.126243f
C21974 VDD.t3872 VSS 0.075275f
C21975 VDD.t4493 VSS 0.075275f
C21976 VDD.t4375 VSS 0.04195f
C21977 VDD.n2873 VSS 0.064751f
C21978 VDD.n2874 VSS 0.07665f
C21979 VDD.t847 VSS 0.007233f
C21980 VDD.t4376 VSS 0.007233f
C21981 VDD.n2875 VSS 0.016652f
C21982 VDD.n2876 VSS 0.047822f
C21983 VDD.t1686 VSS 0.007233f
C21984 VDD.t861 VSS 0.007233f
C21985 VDD.n2877 VSS 0.016652f
C21986 VDD.n2878 VSS 0.076601f
C21987 VDD.t1684 VSS 0.027188f
C21988 VDD.n2879 VSS 0.076624f
C21989 VDD.t3871 VSS 0.027188f
C21990 VDD.n2880 VSS 0.076629f
C21991 VDD.t4473 VSS 0.007233f
C21992 VDD.t3841 VSS 0.007233f
C21993 VDD.n2881 VSS 0.016652f
C21994 VDD.n2882 VSS 0.073624f
C21995 VDD.n2883 VSS 0.07665f
C21996 VDD.n2884 VSS 0.064751f
C21997 VDD.t2931 VSS 0.063514f
C21998 VDD.t3046 VSS 0.075275f
C21999 VDD.t2513 VSS 0.075275f
C22000 VDD.t2511 VSS 0.141141f
C22001 VDD.t3819 VSS 0.141141f
C22002 VDD.t3793 VSS 0.075275f
C22003 VDD.t654 VSS 0.075275f
C22004 VDD.t652 VSS 0.04195f
C22005 VDD.n2885 VSS 0.064751f
C22006 VDD.n2886 VSS 0.07665f
C22007 VDD.t851 VSS 0.007233f
C22008 VDD.t653 VSS 0.007233f
C22009 VDD.n2887 VSS 0.016652f
C22010 VDD.n2888 VSS 0.047822f
C22011 VDD.t1909 VSS 0.007233f
C22012 VDD.t849 VSS 0.007233f
C22013 VDD.n2889 VSS 0.016652f
C22014 VDD.n2890 VSS 0.076601f
C22015 VDD.t1951 VSS 0.027188f
C22016 VDD.n2891 VSS 0.073849f
C22017 VDD.t3786 VSS 0.027188f
C22018 VDD.n2892 VSS 0.073656f
C22019 VDD.t651 VSS 0.007233f
C22020 VDD.t3760 VSS 0.007233f
C22021 VDD.n2893 VSS 0.016652f
C22022 VDD.n2894 VSS 0.073375f
C22023 VDD.n2895 VSS 0.076519f
C22024 VDD.n2896 VSS 0.064751f
C22025 VDD.t3076 VSS 0.063514f
C22026 VDD.t2923 VSS 0.075275f
C22027 VDD.t1922 VSS 0.075275f
C22028 VDD.t1964 VSS 0.137602f
C22029 VDD.t1501 VSS 0.137365f
C22030 VDD.t1499 VSS 0.075145f
C22031 VDD.t1068 VSS 0.075145f
C22032 VDD.t1070 VSS 0.041877f
C22033 VDD.n2897 VSS 0.064693f
C22034 VDD.n2898 VSS 0.076519f
C22035 VDD.t2069 VSS 0.007233f
C22036 VDD.t1071 VSS 0.007233f
C22037 VDD.n2899 VSS 0.016652f
C22038 VDD.n2900 VSS 0.047679f
C22039 VDD.t1258 VSS 0.007233f
C22040 VDD.t2067 VSS 0.007233f
C22041 VDD.n2901 VSS 0.016652f
C22042 VDD.n2902 VSS 0.07634f
C22043 VDD.t1256 VSS 0.027188f
C22044 VDD.n2903 VSS 0.256185f
C22045 VDD.n2904 VSS 0.965405f
C22046 VDD.n2905 VSS 2.17391f
C22047 VDD.n2906 VSS 0.836811f
C22048 VDD.t3295 VSS 0.004807f
C22049 VDD.t3293 VSS 0.004807f
C22050 VDD.n2907 VSS 0.010736f
C22051 VDD.t3297 VSS 0.017466f
C22052 VDD.n2908 VSS 0.056287f
C22053 VDD.n2909 VSS 0.020342f
C22054 VDD.n2910 VSS 0.030311f
C22055 VDD.t3292 VSS 0.089594f
C22056 VDD.n2911 VSS 0.035424f
C22057 VDD.t3294 VSS 0.05332f
C22058 VDD.t3296 VSS 0.027493f
C22059 VDD.n2912 VSS 0.067089f
C22060 VDD.n2913 VSS 0.044915f
C22061 VDD.t3124 VSS 0.081296f
C22062 VDD.t3126 VSS 0.075406f
C22063 VDD.t3122 VSS 0.075406f
C22064 VDD.t3123 VSS 0.075406f
C22065 VDD.t3125 VSS 0.075406f
C22066 VDD.t3502 VSS 0.075406f
C22067 VDD.t3506 VSS 0.075406f
C22068 VDD.t3508 VSS 0.058518f
C22069 VDD.t3504 VSS 0.126462f
C22070 VDD.t3510 VSS 0.05459f
C22071 VDD.n2914 VSS 2.52e-19
C22072 VDD.t3503 VSS 0.00575f
C22073 VDD.t3507 VSS 0.00575f
C22074 VDD.n2915 VSS 0.0115f
C22075 VDD.n2916 VSS 0.012479f
C22076 VDD.t3509 VSS 0.00575f
C22077 VDD.t3511 VSS 0.00575f
C22078 VDD.n2917 VSS 0.0115f
C22079 VDD.n2918 VSS 0.007448f
C22080 VDD.n2919 VSS 0.076419f
C22081 VDD.t3505 VSS 0.01978f
C22082 VDD.n2920 VSS 0.014195f
C22083 VDD.n2921 VSS -0.011842f
C22084 VDD.n2922 VSS 0.077508f
C22085 SEL0.t131 VSS 0.046783f
C22086 SEL0.t40 VSS 0.065305f
C22087 SEL0.t87 VSS 0.065305f
C22088 SEL0.n0 VSS 0.204544f
C22089 SEL0.t110 VSS 0.071515f
C22090 SEL0.t57 VSS 0.072046f
C22091 SEL0.t94 VSS 0.222308f
C22092 SEL0.t25 VSS 0.082991f
C22093 SEL0.n1 VSS 0.278959f
C22094 SEL0.n2 VSS 0.05928f
C22095 SEL0.n3 VSS 0.551386f
C22096 SEL0.t115 VSS 0.072046f
C22097 SEL0.t64 VSS 0.222308f
C22098 SEL0.t55 VSS 0.082991f
C22099 SEL0.n4 VSS 0.278959f
C22100 SEL0.n5 VSS 0.059313f
C22101 SEL0.n6 VSS 0.518954f
C22102 SEL0.n7 VSS 2.16941f
C22103 SEL0.t23 VSS 0.072046f
C22104 SEL0.t99 VSS 0.222308f
C22105 SEL0.t143 VSS 0.082991f
C22106 SEL0.n8 VSS 0.278959f
C22107 SEL0.n9 VSS 0.059328f
C22108 SEL0.n10 VSS 0.553868f
C22109 SEL0.t138 VSS 0.072046f
C22110 SEL0.t50 VSS 0.222308f
C22111 SEL0.t49 VSS 0.082991f
C22112 SEL0.n11 VSS 0.278959f
C22113 SEL0.n12 VSS 0.059326f
C22114 SEL0.n13 VSS 0.49804f
C22115 SEL0.n14 VSS 2.4348f
C22116 SEL0.n15 VSS 2.10974f
C22117 SEL0.n16 VSS 0.664253f
C22118 SEL0.n17 VSS 0.146203f
C22119 SEL0.n18 VSS 0.158543f
C22120 SEL0.n19 VSS 0.146854f
C22121 SEL0.t84 VSS 0.046783f
C22122 SEL0.t78 VSS 0.065305f
C22123 SEL0.t128 VSS 0.065305f
C22124 SEL0.n20 VSS 0.204544f
C22125 SEL0.t7 VSS 0.071515f
C22126 SEL0.t132 VSS 0.072046f
C22127 SEL0.t102 VSS 0.222308f
C22128 SEL0.t126 VSS 0.082991f
C22129 SEL0.n21 VSS 0.278959f
C22130 SEL0.n22 VSS 0.05928f
C22131 SEL0.n23 VSS 0.551386f
C22132 SEL0.t124 VSS 0.072046f
C22133 SEL0.t109 VSS 0.222308f
C22134 SEL0.t74 VSS 0.082991f
C22135 SEL0.n24 VSS 0.278959f
C22136 SEL0.n25 VSS 0.059313f
C22137 SEL0.n26 VSS 0.518954f
C22138 SEL0.n27 VSS 2.16941f
C22139 SEL0.t90 VSS 0.072046f
C22140 SEL0.t15 VSS 0.222308f
C22141 SEL0.t85 VSS 0.082991f
C22142 SEL0.n28 VSS 0.278959f
C22143 SEL0.n29 VSS 0.059328f
C22144 SEL0.n30 VSS 0.553868f
C22145 SEL0.t32 VSS 0.072046f
C22146 SEL0.t75 VSS 0.222308f
C22147 SEL0.t107 VSS 0.082991f
C22148 SEL0.n31 VSS 0.278959f
C22149 SEL0.n32 VSS 0.059326f
C22150 SEL0.n33 VSS 0.49804f
C22151 SEL0.n34 VSS 2.4348f
C22152 SEL0.n35 VSS 2.10974f
C22153 SEL0.n36 VSS 0.664253f
C22154 SEL0.n37 VSS 0.146203f
C22155 SEL0.n38 VSS 0.158543f
C22156 SEL0.n39 VSS 0.147094f
C22157 SEL0.n40 VSS 1.13281f
C22158 SEL0.t83 VSS 0.046783f
C22159 SEL0.t37 VSS 0.065305f
C22160 SEL0.t92 VSS 0.065305f
C22161 SEL0.n41 VSS 0.204544f
C22162 SEL0.t19 VSS 0.071515f
C22163 SEL0.t125 VSS 0.072046f
C22164 SEL0.t6 VSS 0.222308f
C22165 SEL0.t111 VSS 0.082991f
C22166 SEL0.n42 VSS 0.278959f
C22167 SEL0.n43 VSS 0.05928f
C22168 SEL0.n44 VSS 0.551386f
C22169 SEL0.t108 VSS 0.072046f
C22170 SEL0.t14 VSS 0.222308f
C22171 SEL0.t67 VSS 0.082991f
C22172 SEL0.n45 VSS 0.278959f
C22173 SEL0.n46 VSS 0.059313f
C22174 SEL0.n47 VSS 0.518954f
C22175 SEL0.n48 VSS 2.16941f
C22176 SEL0.t27 VSS 0.072046f
C22177 SEL0.t52 VSS 0.222308f
C22178 SEL0.t16 VSS 0.082991f
C22179 SEL0.n49 VSS 0.278959f
C22180 SEL0.n50 VSS 0.059328f
C22181 SEL0.n51 VSS 0.553868f
C22182 SEL0.t68 VSS 0.072046f
C22183 SEL0.t98 VSS 0.222308f
C22184 SEL0.t3 VSS 0.082991f
C22185 SEL0.n52 VSS 0.278959f
C22186 SEL0.n53 VSS 0.059326f
C22187 SEL0.n54 VSS 0.49804f
C22188 SEL0.n55 VSS 2.4348f
C22189 SEL0.n56 VSS 2.10974f
C22190 SEL0.n57 VSS 0.664253f
C22191 SEL0.n58 VSS 0.146203f
C22192 SEL0.n59 VSS 0.158543f
C22193 SEL0.n60 VSS 0.147926f
C22194 SEL0.n61 VSS 4.60662f
C22195 SEL0.t120 VSS 0.046783f
C22196 SEL0.t77 VSS 0.065305f
C22197 SEL0.t127 VSS 0.065305f
C22198 SEL0.n62 VSS 0.204544f
C22199 SEL0.t88 VSS 0.071515f
C22200 SEL0.t70 VSS 0.072046f
C22201 SEL0.t140 VSS 0.222308f
C22202 SEL0.t63 VSS 0.082991f
C22203 SEL0.n63 VSS 0.278959f
C22204 SEL0.n64 VSS 0.05928f
C22205 SEL0.n65 VSS 0.551386f
C22206 SEL0.t60 VSS 0.072046f
C22207 SEL0.t2 VSS 0.222308f
C22208 SEL0.t141 VSS 0.082991f
C22209 SEL0.n66 VSS 0.278959f
C22210 SEL0.n67 VSS 0.059313f
C22211 SEL0.n68 VSS 0.518954f
C22212 SEL0.n69 VSS 2.16941f
C22213 SEL0.t129 VSS 0.072046f
C22214 SEL0.t10 VSS 0.222308f
C22215 SEL0.t122 VSS 0.082991f
C22216 SEL0.n70 VSS 0.278959f
C22217 SEL0.n71 VSS 0.059328f
C22218 SEL0.n72 VSS 0.553868f
C22219 SEL0.t29 VSS 0.072046f
C22220 SEL0.t73 VSS 0.222308f
C22221 SEL0.t105 VSS 0.082991f
C22222 SEL0.n73 VSS 0.278959f
C22223 SEL0.n74 VSS 0.059326f
C22224 SEL0.n75 VSS 0.49804f
C22225 SEL0.n76 VSS 2.4348f
C22226 SEL0.n77 VSS 2.10974f
C22227 SEL0.n78 VSS 0.664253f
C22228 SEL0.n79 VSS 0.146203f
C22229 SEL0.n80 VSS 0.158543f
C22230 SEL0.n81 VSS 0.147087f
C22231 SEL0.n82 VSS 0.182733f
C22232 SEL0.n83 VSS 3.63158f
C22233 SEL0.t80 VSS 0.046783f
C22234 SEL0.t33 VSS 0.065305f
C22235 SEL0.t134 VSS 0.065305f
C22236 SEL0.n84 VSS 0.204544f
C22237 SEL0.t53 VSS 0.071515f
C22238 SEL0.t28 VSS 0.072046f
C22239 SEL0.t34 VSS 0.222308f
C22240 SEL0.t17 VSS 0.082991f
C22241 SEL0.n85 VSS 0.278959f
C22242 SEL0.n86 VSS 0.05928f
C22243 SEL0.n87 VSS 0.551386f
C22244 SEL0.t12 VSS 0.072046f
C22245 SEL0.t43 VSS 0.222308f
C22246 SEL0.t96 VSS 0.082991f
C22247 SEL0.n88 VSS 0.278959f
C22248 SEL0.n89 VSS 0.059313f
C22249 SEL0.n90 VSS 0.518954f
C22250 SEL0.n91 VSS 2.16941f
C22251 SEL0.t24 VSS 0.072046f
C22252 SEL0.t81 VSS 0.222308f
C22253 SEL0.t11 VSS 0.082991f
C22254 SEL0.n92 VSS 0.278959f
C22255 SEL0.n93 VSS 0.059328f
C22256 SEL0.n94 VSS 0.553868f
C22257 SEL0.t66 VSS 0.072046f
C22258 SEL0.t137 VSS 0.222308f
C22259 SEL0.t1 VSS 0.082991f
C22260 SEL0.n95 VSS 0.278959f
C22261 SEL0.n96 VSS 0.059326f
C22262 SEL0.n97 VSS 0.49804f
C22263 SEL0.n98 VSS 2.4348f
C22264 SEL0.n99 VSS 2.10974f
C22265 SEL0.n100 VSS 0.664253f
C22266 SEL0.n101 VSS 0.146203f
C22267 SEL0.n102 VSS 0.158543f
C22268 SEL0.n103 VSS 0.146587f
C22269 SEL0.n104 VSS 0.181695f
C22270 SEL0.n105 VSS 3.64277f
C22271 SEL0.t8 VSS 0.046783f
C22272 SEL0.t5 VSS 0.065305f
C22273 SEL0.t65 VSS 0.065305f
C22274 SEL0.n106 VSS 0.204544f
C22275 SEL0.t86 VSS 0.071515f
C22276 SEL0.t69 VSS 0.072046f
C22277 SEL0.t41 VSS 0.222308f
C22278 SEL0.t59 VSS 0.082991f
C22279 SEL0.n107 VSS 0.278959f
C22280 SEL0.n108 VSS 0.05928f
C22281 SEL0.n109 VSS 0.551386f
C22282 SEL0.t58 VSS 0.072046f
C22283 SEL0.t48 VSS 0.222308f
C22284 SEL0.t139 VSS 0.082991f
C22285 SEL0.n110 VSS 0.278959f
C22286 SEL0.n111 VSS 0.059313f
C22287 SEL0.n112 VSS 0.518954f
C22288 SEL0.n113 VSS 2.16941f
C22289 SEL0.t21 VSS 0.072046f
C22290 SEL0.t45 VSS 0.222308f
C22291 SEL0.t9 VSS 0.082991f
C22292 SEL0.n114 VSS 0.278959f
C22293 SEL0.n115 VSS 0.059328f
C22294 SEL0.n116 VSS 0.553868f
C22295 SEL0.t62 VSS 0.072046f
C22296 SEL0.t95 VSS 0.222308f
C22297 SEL0.t142 VSS 0.082991f
C22298 SEL0.n117 VSS 0.278959f
C22299 SEL0.n118 VSS 0.059326f
C22300 SEL0.n119 VSS 0.49804f
C22301 SEL0.n120 VSS 2.4348f
C22302 SEL0.n121 VSS 2.10974f
C22303 SEL0.n122 VSS 0.664253f
C22304 SEL0.n123 VSS 0.146203f
C22305 SEL0.n124 VSS 0.158543f
C22306 SEL0.n125 VSS 0.147341f
C22307 SEL0.n126 VSS 0.188832f
C22308 SEL0.n127 VSS 3.64321f
C22309 SEL0.t35 VSS 0.046783f
C22310 SEL0.t31 VSS 0.065305f
C22311 SEL0.t82 VSS 0.065305f
C22312 SEL0.n128 VSS 0.204544f
C22313 SEL0.t13 VSS 0.071515f
C22314 SEL0.t130 VSS 0.072046f
C22315 SEL0.t101 VSS 0.222308f
C22316 SEL0.t123 VSS 0.082991f
C22317 SEL0.n129 VSS 0.278959f
C22318 SEL0.n130 VSS 0.05928f
C22319 SEL0.n131 VSS 0.551386f
C22320 SEL0.t121 VSS 0.072046f
C22321 SEL0.t106 VSS 0.222308f
C22322 SEL0.t71 VSS 0.082991f
C22323 SEL0.n132 VSS 0.278959f
C22324 SEL0.n133 VSS 0.059313f
C22325 SEL0.n134 VSS 0.518954f
C22326 SEL0.n135 VSS 2.16941f
C22327 SEL0.t56 VSS 0.072046f
C22328 SEL0.t116 VSS 0.222308f
C22329 SEL0.t47 VSS 0.082991f
C22330 SEL0.n136 VSS 0.278959f
C22331 SEL0.n137 VSS 0.059328f
C22332 SEL0.n138 VSS 0.553868f
C22333 SEL0.t135 VSS 0.072046f
C22334 SEL0.t36 VSS 0.222308f
C22335 SEL0.t79 VSS 0.082991f
C22336 SEL0.n139 VSS 0.278959f
C22337 SEL0.n140 VSS 0.059326f
C22338 SEL0.n141 VSS 0.49804f
C22339 SEL0.n142 VSS 2.4348f
C22340 SEL0.n143 VSS 2.10974f
C22341 SEL0.n144 VSS 0.664253f
C22342 SEL0.n145 VSS 0.146203f
C22343 SEL0.n146 VSS 0.158543f
C22344 SEL0.n147 VSS 0.146488f
C22345 SEL0.n148 VSS 0.180702f
C22346 SEL0.n149 VSS 3.66813f
C22347 SEL0.t20 VSS 0.046783f
C22348 SEL0.t104 VSS 0.065305f
C22349 SEL0.t26 VSS 0.065305f
C22350 SEL0.n150 VSS 0.204544f
C22351 SEL0.t117 VSS 0.071515f
C22352 SEL0.t0 VSS 0.072046f
C22353 SEL0.t118 VSS 0.222308f
C22354 SEL0.t22 VSS 0.082991f
C22355 SEL0.n151 VSS 0.278959f
C22356 SEL0.n152 VSS 0.05928f
C22357 SEL0.n153 VSS 0.551386f
C22358 SEL0.t38 VSS 0.072046f
C22359 SEL0.t100 VSS 0.222308f
C22360 SEL0.t89 VSS 0.082991f
C22361 SEL0.n154 VSS 0.278959f
C22362 SEL0.n155 VSS 0.059313f
C22363 SEL0.n156 VSS 0.518954f
C22364 SEL0.n157 VSS 2.16941f
C22365 SEL0.t97 VSS 0.072046f
C22366 SEL0.t30 VSS 0.222308f
C22367 SEL0.t113 VSS 0.082991f
C22368 SEL0.n158 VSS 0.278959f
C22369 SEL0.n159 VSS 0.059328f
C22370 SEL0.n160 VSS 0.553868f
C22371 SEL0.t44 VSS 0.072046f
C22372 SEL0.t61 VSS 0.222308f
C22373 SEL0.t91 VSS 0.082991f
C22374 SEL0.n161 VSS 0.278959f
C22375 SEL0.n162 VSS 0.059326f
C22376 SEL0.n163 VSS 0.49804f
C22377 SEL0.n164 VSS 2.4348f
C22378 SEL0.n165 VSS 2.10974f
C22379 SEL0.n166 VSS 0.664253f
C22380 SEL0.n167 VSS 0.146203f
C22381 SEL0.n168 VSS 0.158543f
C22382 SEL0.n169 VSS 0.146392f
C22383 SEL0.n170 VSS 0.179739f
C22384 SEL0.n171 VSS 3.63704f
C22385 SEL0.t42 VSS 0.046783f
C22386 SEL0.t136 VSS 0.065305f
C22387 SEL0.t46 VSS 0.065305f
C22388 SEL0.n172 VSS 0.204544f
C22389 SEL0.t114 VSS 0.071515f
C22390 SEL0.t39 VSS 0.072046f
C22391 SEL0.t103 VSS 0.222308f
C22392 SEL0.t54 VSS 0.082991f
C22393 SEL0.n173 VSS 0.278959f
C22394 SEL0.n174 VSS 0.05928f
C22395 SEL0.n175 VSS 0.551386f
C22396 SEL0.t72 VSS 0.072046f
C22397 SEL0.t93 VSS 0.222308f
C22398 SEL0.t112 VSS 0.082991f
C22399 SEL0.n176 VSS 0.278959f
C22400 SEL0.n177 VSS 0.059313f
C22401 SEL0.n178 VSS 0.518954f
C22402 SEL0.n179 VSS 2.16941f
C22403 SEL0.t133 VSS 0.072046f
C22404 SEL0.t18 VSS 0.222308f
C22405 SEL0.t4 VSS 0.082991f
C22406 SEL0.n180 VSS 0.278959f
C22407 SEL0.n181 VSS 0.059328f
C22408 SEL0.n182 VSS 0.553868f
C22409 SEL0.t76 VSS 0.072046f
C22410 SEL0.t51 VSS 0.222308f
C22411 SEL0.t119 VSS 0.082991f
C22412 SEL0.n183 VSS 0.278959f
C22413 SEL0.n184 VSS 0.059326f
C22414 SEL0.n185 VSS 0.49804f
C22415 SEL0.n186 VSS 2.4348f
C22416 SEL0.n187 VSS 2.10974f
C22417 SEL0.n188 VSS 0.664253f
C22418 SEL0.n189 VSS 0.146203f
C22419 SEL0.n190 VSS 0.158543f
C22420 SEL0.n191 VSS 0.146587f
C22421 SEL0.n192 VSS 0.181695f
C22422 SEL0.n193 VSS 4.55348f
C22423 SEL0.n194 VSS 1.10748f
C22424 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t12 VSS 0.013766f
C22425 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t18 VSS 0.027698f
C22426 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t19 VSS 0.027354f
C22427 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t21 VSS 0.027354f
C22428 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t22 VSS 0.027354f
C22429 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t23 VSS 0.005684f
C22430 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t20 VSS 0.005684f
C22431 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t13 VSS 0.005684f
C22432 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n0 VSS 0.168523f
C22433 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n1 VSS 0.124125f
C22434 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n2 VSS 0.067647f
C22435 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n3 VSS 0.066457f
C22436 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n4 VSS 0.040879f
C22437 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n5 VSS 0.05311f
C22438 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t14 VSS 0.030151f
C22439 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t16 VSS 0.009818f
C22440 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t17 VSS 0.013559f
C22441 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n6 VSS 0.014622f
C22442 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t15 VSS 0.010094f
C22443 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n7 VSS 0.025612f
C22444 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n8 VSS 0.044927f
C22445 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t1 VSS 0.004926f
C22446 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t0 VSS 0.004926f
C22447 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n9 VSS 0.011915f
C22448 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t8 VSS 0.004926f
C22449 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t7 VSS 0.004926f
C22450 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n10 VSS 0.011914f
C22451 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n11 VSS 0.085433f
C22452 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t2 VSS 0.004926f
C22453 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t10 VSS 0.004926f
C22454 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n12 VSS 0.009853f
C22455 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n13 VSS 0.00774f
C22456 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t3 VSS 0.020843f
C22457 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t6 VSS 0.020843f
C22458 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n14 VSS 0.041685f
C22459 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n15 VSS 0.016575f
C22460 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t5 VSS 0.020843f
C22461 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t4 VSS 0.020843f
C22462 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n16 VSS 0.041685f
C22463 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n17 VSS 0.018334f
C22464 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n18 VSS 0.188757f
C22465 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t11 VSS 0.020843f
C22466 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.t9 VSS 0.020843f
C22467 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n19 VSS 0.041685f
C22468 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n20 VSS 0.018362f
C22469 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n21 VSS 0.12106f
C22470 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n22 VSS 0.027282f
C22471 8bit_ADDER_0.FULL_ADDER_XORED_4.XOR2_1.A.n23 VSS 0.119748f
C22472 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t7 VSS 0.007073f
C22473 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t8 VSS 0.007073f
C22474 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n0 VSS 0.017105f
C22475 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t9 VSS 0.007073f
C22476 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t11 VSS 0.007073f
C22477 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n1 VSS 0.017107f
C22478 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n2 VSS 0.122656f
C22479 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t6 VSS 0.007073f
C22480 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t10 VSS 0.007073f
C22481 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n3 VSS 0.014146f
C22482 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n4 VSS 0.011112f
C22483 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t3 VSS 0.029924f
C22484 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t1 VSS 0.029924f
C22485 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n5 VSS 0.059848f
C22486 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n6 VSS 0.023796f
C22487 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t4 VSS 0.029924f
C22488 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t5 VSS 0.029924f
C22489 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n7 VSS 0.059848f
C22490 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n8 VSS 0.026362f
C22491 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n9 VSS 0.271f
C22492 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t0 VSS 0.029924f
C22493 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t2 VSS 0.029924f
C22494 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n10 VSS 0.059848f
C22495 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n11 VSS 0.026322f
C22496 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n12 VSS 0.173808f
C22497 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n13 VSS 0.03917f
C22498 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n14 VSS 0.172104f
C22499 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t12 VSS 0.043288f
C22500 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t15 VSS 0.014096f
C22501 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t16 VSS 0.019467f
C22502 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n15 VSS 0.020992f
C22503 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t14 VSS 0.014492f
C22504 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n16 VSS 0.036772f
C22505 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n17 VSS 0.064505f
C22506 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t17 VSS 0.019764f
C22507 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t22 VSS 0.039767f
C22508 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t13 VSS 0.039272f
C22509 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t19 VSS 0.039272f
C22510 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t21 VSS 0.039272f
C22511 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t18 VSS 0.008161f
C22512 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t23 VSS 0.008161f
C22513 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.t20 VSS 0.008161f
C22514 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n18 VSS 0.24195f
C22515 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n19 VSS 0.178207f
C22516 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n20 VSS 0.097121f
C22517 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n21 VSS 0.095413f
C22518 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n22 VSS 0.05869f
C22519 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n23 VSS 0.076991f
C22520 8bit_ADDER_0.FULL_ADDER_XORED_3.XOR2_2.Y.n24 VSS 1.26966f
.ends

