magic
tech sky130B
magscale 1 2
timestamp 1735579975
<< error_p >>
rect -365 -208 -307 -202
rect -173 -208 -115 -202
rect 19 -208 77 -202
rect 211 -208 269 -202
rect -365 -242 -353 -208
rect -173 -242 -161 -208
rect 19 -242 31 -208
rect 211 -242 223 -208
rect -365 -248 -307 -242
rect -173 -248 -115 -242
rect 19 -248 77 -242
rect 211 -248 269 -242
<< nwell >>
rect -449 -223 449 223
rect -449 -261 353 -223
<< pmos >>
rect -351 -161 -321 161
rect -255 -161 -225 161
rect -159 -161 -129 161
rect -63 -161 -33 161
rect 33 -161 63 161
rect 129 -161 159 161
rect 225 -161 255 161
rect 321 -161 351 161
<< pdiff >>
rect -413 149 -351 161
rect -413 -149 -401 149
rect -367 -149 -351 149
rect -413 -161 -351 -149
rect -321 149 -255 161
rect -321 -149 -305 149
rect -271 -149 -255 149
rect -321 -161 -255 -149
rect -225 149 -159 161
rect -225 -149 -209 149
rect -175 -149 -159 149
rect -225 -161 -159 -149
rect -129 149 -63 161
rect -129 -149 -113 149
rect -79 -149 -63 149
rect -129 -161 -63 -149
rect -33 149 33 161
rect -33 -149 -17 149
rect 17 -149 33 149
rect -33 -161 33 -149
rect 63 149 129 161
rect 63 -149 79 149
rect 113 -149 129 149
rect 63 -161 129 -149
rect 159 149 225 161
rect 159 -149 175 149
rect 209 -149 225 149
rect 159 -161 225 -149
rect 255 149 321 161
rect 255 -149 271 149
rect 305 -149 321 149
rect 255 -161 321 -149
rect 351 149 413 161
rect 351 -149 367 149
rect 401 -149 413 149
rect 351 -161 413 -149
<< pdiffc >>
rect -401 -149 -367 149
rect -305 -149 -271 149
rect -209 -149 -175 149
rect -113 -149 -79 149
rect -17 -149 17 149
rect 79 -149 113 149
rect 175 -149 209 149
rect 271 -149 305 149
rect 367 -149 401 149
<< poly >>
rect -351 161 -321 187
rect -255 161 -225 187
rect -159 161 -129 187
rect -63 161 -33 187
rect 33 161 63 187
rect 129 161 159 187
rect 225 161 255 187
rect 321 161 351 187
rect -351 -192 -321 -161
rect -255 -192 -225 -161
rect -159 -192 -129 -161
rect -63 -192 -33 -161
rect 33 -192 63 -161
rect 129 -192 159 -161
rect 225 -192 255 -161
rect 321 -192 351 -161
rect -369 -208 -225 -192
rect -369 -242 -353 -208
rect -319 -242 -225 -208
rect -369 -258 -225 -242
rect -177 -208 -33 -192
rect -177 -242 -161 -208
rect -127 -242 -33 -208
rect -177 -258 -33 -242
rect 15 -208 159 -192
rect 15 -242 31 -208
rect 65 -242 159 -208
rect 15 -258 159 -242
rect 207 -208 351 -192
rect 207 -242 223 -208
rect 257 -242 351 -208
rect 207 -258 351 -242
<< polycont >>
rect -353 -242 -319 -208
rect -161 -242 -127 -208
rect 31 -242 65 -208
rect 223 -242 257 -208
<< locali >>
rect -401 149 -367 165
rect -305 149 -271 165
rect -401 -165 -367 -149
rect -305 -165 -271 -154
rect -209 149 -175 165
rect -209 -165 -175 -149
rect -113 149 -79 165
rect -17 149 17 165
rect -113 -165 -79 -154
rect -17 -165 17 -149
rect 79 149 113 165
rect 175 149 209 165
rect 79 -165 113 -154
rect 175 -165 209 -149
rect 271 149 305 165
rect 367 149 401 165
rect 271 -165 305 -154
rect 367 -165 401 -149
rect -369 -242 -353 -208
rect -319 -242 -303 -208
rect -177 -242 -161 -208
rect -127 -242 -111 -208
rect 15 -242 31 -208
rect 65 -242 81 -208
rect 207 -242 223 -208
rect 257 -242 273 -208
<< viali >>
rect -401 36 -367 146
rect -306 -149 -305 -42
rect -305 -149 -271 -42
rect -306 -154 -271 -149
rect -209 36 -175 146
rect -17 36 17 146
rect -113 -149 -79 -42
rect -79 -149 -78 -42
rect -113 -154 -78 -149
rect 175 36 209 146
rect 79 -149 113 -42
rect 113 -149 114 -42
rect 79 -154 114 -149
rect 367 36 401 146
rect 271 -149 305 -42
rect 305 -149 306 -42
rect 271 -154 306 -149
rect -353 -242 -319 -208
rect -161 -242 -127 -208
rect 31 -242 65 -208
rect 223 -242 257 -208
<< metal1 >>
rect -413 146 413 161
rect -413 36 -401 146
rect -367 36 -209 146
rect -175 36 -17 146
rect 17 36 175 146
rect 209 36 367 146
rect 401 36 413 146
rect -413 27 413 36
rect -413 -42 413 -27
rect -413 -154 -306 -42
rect -271 -154 -113 -42
rect -78 -154 79 -42
rect 114 -154 271 -42
rect 306 -154 413 -42
rect -413 -161 413 -154
rect -365 -208 -307 -202
rect -365 -242 -353 -208
rect -319 -242 -307 -208
rect -365 -248 -307 -242
rect -173 -208 -115 -202
rect -173 -242 -161 -208
rect -127 -242 -115 -208
rect -173 -248 -115 -242
rect 19 -208 77 -202
rect 19 -242 31 -208
rect 65 -242 77 -208
rect 19 -248 77 -242
rect 211 -208 269 -202
rect 211 -242 223 -208
rect 257 -242 269 -208
rect 211 -248 269 -242
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.605 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
