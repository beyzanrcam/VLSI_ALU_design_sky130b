magic
tech sky130B
magscale 1 2
timestamp 1735226356
<< error_s >>
rect 878 683 6842 684
rect 123 266 6842 683
rect 123 265 6087 266
rect 199 139 399 197
rect 578 139 778 197
rect 1051 139 1251 197
rect 1430 139 1630 197
rect 1903 139 2103 197
rect 2282 139 2482 197
rect 2755 139 2955 197
rect 3134 139 3334 197
rect 3607 139 3807 197
rect 3986 139 4186 197
rect 4459 139 4659 197
rect 4838 139 5038 197
rect 5311 140 5511 198
rect 5690 140 5890 198
rect 6163 140 6363 198
rect 6542 140 6742 198
rect 199 51 399 109
rect 578 51 778 109
rect 1051 51 1251 109
rect 1430 51 1630 109
rect 1903 51 2103 109
rect 2282 51 2482 109
rect 2755 51 2955 109
rect 3134 51 3334 109
rect 3607 51 3807 109
rect 3986 51 4186 109
rect 4459 51 4659 109
rect 4838 51 5038 109
rect 5311 52 5511 110
rect 5690 52 5890 110
rect 6163 52 6363 110
rect 6542 52 6742 110
rect 333 18 653 42
rect 1185 18 1505 42
rect 2037 18 2357 42
rect 2889 18 3209 42
rect 3741 18 4061 42
rect 4593 18 4913 42
rect 5445 19 5765 43
rect 6297 19 6617 43
rect 333 -254 357 18
rect 1185 -254 1209 18
rect 2037 -254 2061 18
rect 2889 -254 2913 18
rect 3741 -254 3765 18
rect 4593 -254 4617 18
rect 5445 -253 5469 19
rect 6297 -253 6321 19
rect 333 -278 653 -254
rect 1185 -278 1505 -254
rect 2037 -278 2357 -254
rect 2889 -278 3209 -254
rect 3741 -278 4061 -254
rect 4593 -278 4913 -254
rect 5445 -277 5765 -253
rect 6297 -277 6617 -253
<< nwell >>
rect 878 265 6087 684
<< metal1 >>
rect 809 858 878 859
rect 809 683 975 858
rect 1661 684 1827 859
rect 2513 685 2679 860
rect 809 603 878 683
rect 1661 603 1730 684
rect 2513 603 2582 685
rect 3365 684 3531 859
rect 4217 684 4383 859
rect 5069 684 5235 859
rect 5921 684 6087 859
rect 6773 684 6939 859
rect 3365 603 3434 684
rect 4217 603 4286 684
rect 5069 603 5138 684
rect 5921 604 5990 684
rect 6773 604 6842 684
rect 54 6 123 603
rect 906 6 975 603
rect 1758 6 1827 603
rect 2610 6 2679 603
rect 3462 6 3531 603
rect 4314 6 4383 603
rect -43 -278 123 6
rect 809 -278 975 6
rect 1661 -278 1827 6
rect 2513 -278 2679 6
rect 3365 -278 3531 6
rect 4217 -278 4383 6
rect 5166 -1 5235 596
rect 6018 7 6087 604
rect 5069 -277 5235 -1
rect 5921 -277 6087 7
rect 6677 -277 6843 16
use buffer  buffer_0 ~/Documents/Dersler/VLSI/vlsi_sky130b/design/mag/inv
timestamp 1735226356
transform -1 0 8314 0 1 313
box 1472 -590 2227 547
use buffer  buffer_1
timestamp 1735226356
transform -1 0 2350 0 1 312
box 1472 -590 2227 547
use buffer  buffer_2
timestamp 1735226356
transform -1 0 3202 0 1 312
box 1472 -590 2227 547
use buffer  buffer_3
timestamp 1735226356
transform -1 0 4054 0 1 312
box 1472 -590 2227 547
use buffer  buffer_4
timestamp 1735226356
transform -1 0 4906 0 1 312
box 1472 -590 2227 547
use buffer  buffer_5
timestamp 1735226356
transform -1 0 5758 0 1 312
box 1472 -590 2227 547
use buffer  buffer_6
timestamp 1735226356
transform -1 0 6610 0 1 312
box 1472 -590 2227 547
use buffer  buffer_7
timestamp 1735226356
transform -1 0 7462 0 1 313
box 1472 -590 2227 547
<< end >>
