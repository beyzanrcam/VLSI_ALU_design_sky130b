magic
tech sky130B
magscale 1 2
timestamp 1732804393
<< nwell >>
rect 0 366 376 418
rect 101 347 104 366
rect 223 290 343 338
rect 326 288 343 290
<< poly >>
rect 3 -124 70 -108
rect 3 -158 19 -124
rect 53 -126 70 -124
rect 53 -156 75 -126
rect 53 -158 70 -156
rect 3 -174 70 -158
<< polycont >>
rect 19 -158 53 -124
<< locali >>
rect 3 -124 53 339
rect 3 -158 19 -124
rect 3 -174 53 -158
<< viali >>
rect 19 -158 53 -124
<< metal1 >>
rect 0 366 376 418
rect 101 347 104 366
rect 0 80 53 338
rect 223 82 376 338
rect 0 -124 69 80
rect 100 -114 376 82
rect 0 -158 19 -124
rect 53 -158 69 -124
rect 0 -175 69 -158
rect 100 -203 300 -161
rect 328 -175 376 -114
rect 0 -250 376 -203
use efepmos_W107-L15-F3  efepmos_W107-L15-F3_0 ~/Documents/vlsi/vlsi_sky130b/design/mag
timestamp 1732803117
transform 0 1 207 -1 0 209
box -209 -207 209 169
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0 ~/Documents/vlsi/vlsi_sky130b/design/mag
timestamp 1732515081
transform 0 1 200 -1 0 -141
box -73 -126 73 126
<< labels >>
rlabel metal1 376 -31 376 -31 3 Y
port 2 e
rlabel metal1 0 -31 0 -31 7 A
rlabel metal1 144 418 144 418 1 vss
port 1 n
rlabel metal1 201 -250 201 -250 5 VSS
port 3 s
<< end >>
