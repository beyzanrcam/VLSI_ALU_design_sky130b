magic
tech sky130B
magscale 1 2
timestamp 1734121007
<< error_p >>
rect -401 383 401 421
rect -497 -421 497 383
<< nwell >>
rect -401 383 401 421
rect -497 -421 497 383
<< pmos >>
rect -399 -321 -369 321
rect -303 -321 -273 321
rect -207 -321 -177 321
rect -111 -321 -81 321
rect -15 -321 15 321
rect 81 -321 111 321
rect 177 -321 207 321
rect 273 -321 303 321
rect 369 -321 399 321
<< pdiff >>
rect -461 309 -399 321
rect -461 -309 -449 309
rect -415 -309 -399 309
rect -461 -321 -399 -309
rect -369 309 -303 321
rect -369 -309 -353 309
rect -319 -309 -303 309
rect -369 -321 -303 -309
rect -273 309 -207 321
rect -273 -309 -257 309
rect -223 -309 -207 309
rect -273 -321 -207 -309
rect -177 309 -111 321
rect -177 -309 -161 309
rect -127 -309 -111 309
rect -177 -321 -111 -309
rect -81 309 -15 321
rect -81 -309 -65 309
rect -31 -309 -15 309
rect -81 -321 -15 -309
rect 15 309 81 321
rect 15 -309 31 309
rect 65 -309 81 309
rect 15 -321 81 -309
rect 111 309 177 321
rect 111 -309 127 309
rect 161 -309 177 309
rect 111 -321 177 -309
rect 207 309 273 321
rect 207 -309 223 309
rect 257 -309 273 309
rect 207 -321 273 -309
rect 303 309 369 321
rect 303 -309 319 309
rect 353 -309 369 309
rect 303 -321 369 -309
rect 399 309 461 321
rect 399 -309 415 309
rect 449 -309 461 309
rect 399 -321 461 -309
<< pdiffc >>
rect -449 -309 -415 309
rect -353 -309 -319 309
rect -257 -309 -223 309
rect -161 -309 -127 309
rect -65 -309 -31 309
rect 31 -309 65 309
rect 127 -309 161 309
rect 223 -309 257 309
rect 319 -309 353 309
rect 415 -309 449 309
<< poly >>
rect -399 321 -369 347
rect -303 321 -273 347
rect -207 321 -177 347
rect -111 321 -81 347
rect -15 321 15 347
rect 81 321 111 347
rect 177 321 207 347
rect 273 321 303 347
rect 369 321 399 347
rect -399 -352 -369 -321
rect -303 -352 -273 -321
rect -207 -352 -177 -321
rect -399 -382 -177 -352
rect -111 -352 -81 -321
rect -15 -352 15 -321
rect 81 -352 111 -321
rect -111 -382 111 -352
rect 177 -352 207 -321
rect 273 -352 303 -321
rect 369 -352 399 -321
rect 177 -382 399 -352
<< locali >>
rect -449 309 -415 325
rect -449 -325 -415 -309
rect -353 309 -319 325
rect -353 -325 -319 -309
rect -257 309 -223 325
rect -257 -325 -223 -309
rect -161 309 -127 325
rect -161 -325 -127 -309
rect -65 309 -31 325
rect -65 -325 -31 -309
rect 31 309 65 325
rect 31 -325 65 -309
rect 127 309 161 325
rect 127 -325 161 -309
rect 223 309 257 325
rect 223 -325 257 -309
rect 319 309 353 325
rect 319 -325 353 -309
rect 415 309 449 325
rect 415 -325 449 -309
<< viali >>
rect -449 17 -415 309
rect -353 -309 -319 -37
rect -257 17 -223 309
rect -161 -309 -127 -37
rect -65 17 -31 309
rect 31 -309 65 -37
rect 127 17 161 309
rect 223 -309 257 -37
rect 319 17 353 309
rect 415 -309 449 -37
<< metal1 >>
rect -455 309 -409 321
rect -455 17 -449 309
rect -415 17 -409 309
rect -263 309 -217 321
rect -263 17 -257 309
rect -223 17 -217 309
rect -71 309 -25 321
rect -71 17 -65 309
rect -31 17 -25 309
rect 121 309 167 321
rect 121 17 127 309
rect 161 17 167 309
rect 313 309 359 321
rect 313 17 319 309
rect 353 17 359 309
rect -359 -309 -353 -37
rect -319 -309 -313 -37
rect -359 -321 -313 -309
rect -167 -309 -161 -37
rect -127 -309 -121 -37
rect -167 -321 -121 -309
rect 25 -309 31 -37
rect 65 -309 71 -37
rect 25 -321 71 -309
rect 217 -309 223 -37
rect 257 -309 263 -37
rect 217 -321 263 -309
rect 409 -309 415 -37
rect 449 -309 455 -37
rect 409 -321 455 -309
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.21 l 0.15 m 1 nf 9 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
