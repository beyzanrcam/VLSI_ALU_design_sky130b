* NGSPICE file created from NAND4.ext - technology: sky130B

.subckt nmos4_fingered a_n63_n227# a_n33_n200# a_n265_n299# a_n413_n200# a_n159_n226#
+ a_n413_n382# a_351_n200# VSUBS
X0 a_n33_n200# a_n63_n227# a_n129_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1 a_351_n200# a_n413_n382# a_255_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2 a_255_n200# a_n265_n299# a_159_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3 a_n321_n200# a_n413_n382# a_n413_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X4 a_159_n200# a_n159_n226# a_63_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X5 a_n225_n200# a_n265_n299# a_n321_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X6 a_63_n200# a_n63_n227# a_n33_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X7 a_n129_n200# a_n159_n226# a_n225_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
.ends

.subckt pmos4_f2 a_n177_n258# a_n413_n161# a_207_n258# w_n449_n261# a_n369_n258# a_n321_n161#
+ a_15_n258#
X0 a_n321_n161# a_207_n258# a_n413_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X1 a_n321_n161# a_n369_n258# a_n413_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.4991 ps=3.84 w=1.61 l=0.15
X2 a_n413_n161# a_15_n258# a_n321_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X3 a_n413_n161# a_n369_n258# a_n321_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X4 a_n321_n161# a_15_n258# a_n413_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X5 a_n321_n161# a_n177_n258# a_n413_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X6 a_n413_n161# a_n177_n258# a_n321_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.26565 pd=1.94 as=0.26565 ps=1.94 w=1.61 l=0.15
X7 a_n413_n161# a_207_n258# a_n321_n161# w_n449_n261# sky130_fd_pr__pfet_01v8 ad=0.4991 pd=3.84 as=0.26565 ps=1.94 w=1.61 l=0.15
.ends

.subckt NAND4 A B C D VSS VDD Y
Xsky130_fd_pr__nfet_01v8_V69YKH_0 D Y B VSS C A VSS VSS nmos4_fingered
Xsky130_fd_pr__pfet_01v8_NFZE9G_0 B VDD D VDD A Y C pmos4_f2
.ends

