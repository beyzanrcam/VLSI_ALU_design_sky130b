magic
tech sky130B
magscale 1 2
timestamp 1734125383
<< nwell >>
rect -205 775 789 1745
<< nmos >>
rect 181 296 211 496
rect 277 296 307 496
rect 373 296 403 496
<< pmos >>
rect -107 875 -77 1517
rect -11 875 19 1517
rect 85 875 115 1517
rect 181 875 211 1517
rect 277 875 307 1517
rect 373 875 403 1517
rect 469 875 499 1517
rect 565 875 595 1517
rect 661 875 691 1517
<< ndiff >>
rect 119 484 181 496
rect 119 308 131 484
rect 165 308 181 484
rect 119 296 181 308
rect 211 484 277 496
rect 211 308 227 484
rect 261 308 277 484
rect 211 296 277 308
rect 307 484 373 496
rect 307 308 323 484
rect 357 308 373 484
rect 307 296 373 308
rect 403 484 465 496
rect 403 308 419 484
rect 453 308 465 484
rect 403 296 465 308
<< pdiff >>
rect -169 1505 -107 1517
rect -169 887 -157 1505
rect -123 887 -107 1505
rect -169 875 -107 887
rect -77 1505 -11 1517
rect -77 887 -61 1505
rect -27 887 -11 1505
rect -77 875 -11 887
rect 19 1505 85 1517
rect 19 887 35 1505
rect 69 887 85 1505
rect 19 875 85 887
rect 115 1505 181 1517
rect 115 887 131 1505
rect 165 887 181 1505
rect 115 875 181 887
rect 211 1505 277 1517
rect 211 887 227 1505
rect 261 887 277 1505
rect 211 875 277 887
rect 307 1505 373 1517
rect 307 887 323 1505
rect 357 887 373 1505
rect 307 875 373 887
rect 403 1505 469 1517
rect 403 887 419 1505
rect 453 887 469 1505
rect 403 875 469 887
rect 499 1505 565 1517
rect 499 887 515 1505
rect 549 887 565 1505
rect 499 875 565 887
rect 595 1505 661 1517
rect 595 887 611 1505
rect 645 887 661 1505
rect 595 875 661 887
rect 691 1505 753 1517
rect 691 887 707 1505
rect 741 887 753 1505
rect 691 875 753 887
<< ndiffc >>
rect 131 308 165 484
rect 227 308 261 484
rect 323 308 357 484
rect 419 308 453 484
<< pdiffc >>
rect -157 887 -123 1505
rect -61 887 -27 1505
rect 35 887 69 1505
rect 131 887 165 1505
rect 227 887 261 1505
rect 323 887 357 1505
rect 419 887 453 1505
rect 515 887 549 1505
rect 611 887 645 1505
rect 707 887 741 1505
<< psubdiff >>
rect 119 219 465 240
rect 119 101 144 219
rect 420 101 465 219
rect 119 79 465 101
<< nsubdiff >>
rect -162 1694 753 1709
rect -162 1600 -135 1694
rect 78 1600 753 1694
rect -162 1582 753 1600
<< psubdiffcont >>
rect 144 101 420 219
<< nsubdiffcont >>
rect -135 1600 78 1694
<< poly >>
rect -107 1517 -77 1543
rect -11 1517 19 1543
rect 85 1517 115 1543
rect 181 1517 211 1543
rect 277 1517 307 1543
rect 373 1517 403 1543
rect 469 1517 499 1543
rect 565 1517 595 1543
rect 661 1517 691 1543
rect -107 844 -77 875
rect -11 844 19 875
rect 85 844 115 875
rect -107 814 115 844
rect 181 844 211 875
rect 277 844 307 875
rect 373 844 403 875
rect 181 814 403 844
rect 469 844 499 875
rect 565 844 595 875
rect 661 844 691 875
rect 469 814 691 844
rect 49 799 115 814
rect 49 765 65 799
rect 99 765 115 799
rect 49 748 115 765
rect 85 661 115 748
rect 277 718 307 814
rect 259 702 325 718
rect 259 668 275 702
rect 309 668 325 702
rect 85 631 211 661
rect 259 652 325 668
rect 181 496 211 631
rect 277 496 307 652
rect 469 590 499 814
rect 373 574 499 590
rect 373 540 389 574
rect 423 560 499 574
rect 423 540 439 560
rect 373 524 439 540
rect 373 496 403 524
rect 181 270 211 296
rect 277 270 307 296
rect 373 270 403 296
<< polycont >>
rect 65 765 99 799
rect 275 668 309 702
rect 389 540 423 574
<< locali >>
rect -162 1694 753 1702
rect -162 1600 -135 1694
rect 78 1600 753 1694
rect -162 1590 753 1600
rect -157 1505 -123 1521
rect -157 871 -123 887
rect -61 1505 -27 1521
rect -61 871 -27 887
rect 35 1505 69 1521
rect 35 871 69 887
rect 131 1505 165 1521
rect 131 871 165 887
rect 227 1505 261 1521
rect 227 871 261 887
rect 323 1505 357 1521
rect 323 871 357 887
rect 419 1505 453 1521
rect 419 871 453 887
rect 515 1505 549 1521
rect 515 871 549 887
rect 611 1505 645 1521
rect 611 871 645 887
rect 707 1505 741 1521
rect 707 871 741 887
rect 49 765 65 799
rect 99 765 115 799
rect 259 668 275 702
rect 309 668 325 702
rect 373 540 389 574
rect 423 540 439 574
rect 131 484 165 500
rect 131 228 165 308
rect 227 484 261 500
rect 227 292 261 308
rect 323 484 357 500
rect 323 228 357 308
rect 419 484 453 500
rect 419 292 453 308
rect 119 219 465 228
rect 119 101 144 219
rect 420 101 465 219
rect 119 91 465 101
<< viali >>
rect -135 1600 78 1694
rect -157 1213 -123 1505
rect -61 887 -27 1159
rect 35 1213 69 1505
rect 131 887 165 1159
rect 227 1213 261 1505
rect 323 887 357 1159
rect 419 1213 453 1505
rect 515 887 549 1159
rect 611 1213 645 1505
rect 707 887 741 1159
rect 65 765 99 799
rect 275 668 309 702
rect 389 540 423 574
rect 227 308 261 484
rect 419 308 453 484
<< metal1 >>
rect -147 1694 90 1701
rect -147 1600 -135 1694
rect 78 1600 90 1694
rect -147 1593 90 1600
rect -147 1517 57 1593
rect -163 1505 75 1517
rect -163 1213 -157 1505
rect -123 1213 35 1505
rect 69 1213 75 1505
rect -163 1201 75 1213
rect 221 1505 651 1517
rect 221 1213 227 1505
rect 261 1213 419 1505
rect 453 1213 611 1505
rect 645 1213 651 1505
rect 221 1201 651 1213
rect -67 1159 363 1171
rect -67 887 -61 1159
rect -27 887 131 1159
rect 165 887 323 1159
rect 357 887 363 1159
rect -67 875 363 887
rect 509 1159 747 1171
rect 509 887 515 1159
rect 549 887 707 1159
rect 741 887 747 1159
rect 509 875 747 887
rect -310 799 115 814
rect -310 765 65 799
rect 99 765 115 799
rect -310 747 115 765
rect -310 702 325 718
rect -310 668 275 702
rect 309 668 325 702
rect -310 652 325 668
rect -310 574 439 590
rect -310 540 389 574
rect 423 540 439 574
rect -310 524 439 540
rect 595 496 747 875
rect 221 484 747 496
rect 221 308 227 484
rect 261 308 419 484
rect 453 308 747 484
rect 221 296 747 308
<< labels >>
rlabel metal1 -310 778 -310 778 7 A
port 1 w
rlabel metal1 -310 684 -310 684 7 B
port 2 w
rlabel metal1 -310 559 -310 559 3 C
port 3 e
rlabel psubdiffcont 246 158 246 158 1 VSS
port 4 n
rlabel viali -29 1648 -29 1648 5 VDD
port 5 s
rlabel metal1 676 638 676 638 3 Y
port 6 e
<< end >>
