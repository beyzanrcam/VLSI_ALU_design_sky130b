magic
tech sky130B
magscale 1 2
timestamp 1733174445
<< error_p >>
rect -206 114 -148 120
rect -88 114 -30 120
rect 30 114 88 120
rect 148 114 206 120
rect -206 80 -194 114
rect -88 80 -76 114
rect 30 80 42 114
rect 148 80 160 114
rect -206 74 -148 80
rect -88 74 -30 80
rect 30 74 88 80
rect 148 74 206 80
rect -206 -80 -148 -74
rect -88 -80 -30 -74
rect 30 -80 88 -74
rect 148 -80 206 -74
rect -206 -114 -194 -80
rect -88 -114 -76 -80
rect 30 -114 42 -80
rect 148 -114 160 -80
rect -206 -120 -148 -114
rect -88 -120 -30 -114
rect 30 -120 88 -114
rect 148 -120 206 -114
<< pwell >>
rect -403 -252 403 252
<< nmos >>
rect -207 -42 -147 42
rect -89 -42 -29 42
rect 29 -42 89 42
rect 147 -42 207 42
<< ndiff >>
rect -265 30 -207 42
rect -265 -30 -253 30
rect -219 -30 -207 30
rect -265 -42 -207 -30
rect -147 30 -89 42
rect -147 -30 -135 30
rect -101 -30 -89 30
rect -147 -42 -89 -30
rect -29 30 29 42
rect -29 -30 -17 30
rect 17 -30 29 30
rect -29 -42 29 -30
rect 89 30 147 42
rect 89 -30 101 30
rect 135 -30 147 30
rect 89 -42 147 -30
rect 207 30 265 42
rect 207 -30 219 30
rect 253 -30 265 30
rect 207 -42 265 -30
<< ndiffc >>
rect -253 -30 -219 30
rect -135 -30 -101 30
rect -17 -30 17 30
rect 101 -30 135 30
rect 219 -30 253 30
<< psubdiff >>
rect -367 182 -271 216
rect 271 182 367 216
rect -367 120 -333 182
rect 333 120 367 182
rect -367 -182 -333 -120
rect 333 -182 367 -120
rect -367 -216 -271 -182
rect 271 -216 367 -182
<< psubdiffcont >>
rect -271 182 271 216
rect -367 -120 -333 120
rect 333 -120 367 120
rect -271 -216 271 -182
<< poly >>
rect -210 114 -144 130
rect -210 80 -194 114
rect -160 80 -144 114
rect -210 64 -144 80
rect -92 114 -26 130
rect -92 80 -76 114
rect -42 80 -26 114
rect -92 64 -26 80
rect 26 114 92 130
rect 26 80 42 114
rect 76 80 92 114
rect 26 64 92 80
rect 144 114 210 130
rect 144 80 160 114
rect 194 80 210 114
rect 144 64 210 80
rect -207 42 -147 64
rect -89 42 -29 64
rect 29 42 89 64
rect 147 42 207 64
rect -207 -64 -147 -42
rect -89 -64 -29 -42
rect 29 -64 89 -42
rect 147 -64 207 -42
rect -210 -80 -144 -64
rect -210 -114 -194 -80
rect -160 -114 -144 -80
rect -210 -130 -144 -114
rect -92 -80 -26 -64
rect -92 -114 -76 -80
rect -42 -114 -26 -80
rect -92 -130 -26 -114
rect 26 -80 92 -64
rect 26 -114 42 -80
rect 76 -114 92 -80
rect 26 -130 92 -114
rect 144 -80 210 -64
rect 144 -114 160 -80
rect 194 -114 210 -80
rect 144 -130 210 -114
<< polycont >>
rect -194 80 -160 114
rect -76 80 -42 114
rect 42 80 76 114
rect 160 80 194 114
rect -194 -114 -160 -80
rect -76 -114 -42 -80
rect 42 -114 76 -80
rect 160 -114 194 -80
<< locali >>
rect -367 182 -271 216
rect 271 182 367 216
rect -367 120 -333 182
rect 333 120 367 182
rect -210 80 -194 114
rect -160 80 -144 114
rect -92 80 -76 114
rect -42 80 -26 114
rect 26 80 42 114
rect 76 80 92 114
rect 144 80 160 114
rect 194 80 210 114
rect -253 30 -219 46
rect -253 -46 -219 -30
rect -135 30 -101 46
rect -135 -46 -101 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 101 30 135 46
rect 101 -46 135 -30
rect 219 30 253 46
rect 219 -46 253 -30
rect -210 -114 -194 -80
rect -160 -114 -144 -80
rect -92 -114 -76 -80
rect -42 -114 -26 -80
rect 26 -114 42 -80
rect 76 -114 92 -80
rect 144 -114 160 -80
rect 194 -114 210 -80
rect -367 -182 -333 -120
rect 333 -182 367 -120
rect -367 -216 -271 -182
rect 271 -216 367 -182
<< viali >>
rect -194 80 -160 114
rect -76 80 -42 114
rect 42 80 76 114
rect 160 80 194 114
rect -253 -30 -219 30
rect -135 -30 -101 30
rect -17 -30 17 30
rect 101 -30 135 30
rect 219 -30 253 30
rect -194 -114 -160 -80
rect -76 -114 -42 -80
rect 42 -114 76 -80
rect 160 -114 194 -80
<< metal1 >>
rect -206 114 -148 120
rect -206 80 -194 114
rect -160 80 -148 114
rect -206 74 -148 80
rect -88 114 -30 120
rect -88 80 -76 114
rect -42 80 -30 114
rect -88 74 -30 80
rect 30 114 88 120
rect 30 80 42 114
rect 76 80 88 114
rect 30 74 88 80
rect 148 114 206 120
rect 148 80 160 114
rect 194 80 206 114
rect 148 74 206 80
rect -259 30 -213 42
rect -259 -30 -253 30
rect -219 -30 -213 30
rect -259 -42 -213 -30
rect -141 30 -95 42
rect -141 -30 -135 30
rect -101 -30 -95 30
rect -141 -42 -95 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 95 30 141 42
rect 95 -30 101 30
rect 135 -30 141 30
rect 95 -42 141 -30
rect 213 30 259 42
rect 213 -30 219 30
rect 253 -30 259 30
rect 213 -42 259 -30
rect -206 -80 -148 -74
rect -206 -114 -194 -80
rect -160 -114 -148 -80
rect -206 -120 -148 -114
rect -88 -80 -30 -74
rect -88 -114 -76 -80
rect -42 -114 -30 -80
rect -88 -120 -30 -114
rect 30 -80 88 -74
rect 30 -114 42 -80
rect 76 -114 88 -80
rect 30 -120 88 -114
rect 148 -80 206 -74
rect 148 -114 160 -80
rect 194 -114 206 -80
rect 148 -120 206 -114
<< properties >>
string FIXED_BBOX -350 -199 350 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.30 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
