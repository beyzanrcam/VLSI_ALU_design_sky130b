magic
tech sky130B
magscale 1 2
timestamp 1736682680
<< nwell >>
rect -3439 3542 3242 4070
rect -3388 1730 -2206 2288
rect -1652 1730 -524 2272
rect -3388 438 -2260 980
rect -1652 438 -524 980
rect -3388 -1535 -2260 -993
rect -1651 -1535 -523 -993
rect -3388 -2827 -2260 -2285
rect -1652 -2827 -524 -2285
rect -3388 -4799 -2260 -4257
rect -1651 -4799 -523 -4257
rect -3388 -6091 -2260 -5549
rect -1651 -6091 -523 -5549
<< locali >>
rect 154 1006 264 1634
rect 154 942 596 1006
<< metal1 >>
rect -2584 4006 -2370 4028
rect -3404 3904 -2770 3938
rect -2584 3927 -2561 4006
rect -2392 3927 -2370 4006
rect -564 4006 -350 4028
rect -2584 3908 -2370 3927
rect -3404 3764 -3366 3904
rect -2812 3764 -2770 3904
rect -3404 3725 -2770 3764
rect -1367 3904 -733 3938
rect -564 3927 -541 4006
rect -372 3927 -350 4006
rect 1177 4006 1391 4028
rect -564 3908 -350 3927
rect -1367 3764 -1329 3904
rect -775 3764 -733 3904
rect -1367 3725 -733 3764
rect 363 3904 997 3938
rect 1177 3927 1200 4006
rect 1369 3927 1391 4006
rect 2956 4006 3170 4028
rect 1177 3908 1391 3927
rect 363 3764 401 3904
rect 955 3764 997 3904
rect 363 3725 997 3764
rect 2123 3904 2757 3938
rect 2956 3927 2979 4006
rect 3148 3927 3170 4006
rect 2956 3908 3170 3927
rect 2123 3764 2161 3904
rect 2715 3764 2757 3904
rect 2123 3725 2757 3764
rect -3597 3440 -3591 3583
rect -3448 3440 -3357 3583
rect -2781 3422 -2683 3696
rect -1749 3574 -1335 3576
rect -1749 3557 -1330 3574
rect -2305 3484 -2010 3524
rect -3544 3291 -3388 3372
rect -2584 3353 -2384 3381
rect -3559 3244 -3350 3291
rect -3559 3066 -3506 3244
rect -3384 3066 -3350 3244
rect -3169 3248 -2769 3276
rect -3169 3174 -3140 3248
rect -2800 3174 -2769 3248
rect -2584 3257 -2557 3353
rect -2408 3257 -2384 3353
rect -2305 3365 -2209 3484
rect -2077 3365 -2010 3484
rect -1749 3464 -1687 3557
rect -1369 3470 -1330 3557
rect -1369 3464 -1335 3470
rect -1749 3440 -1335 3464
rect -712 3422 -664 3696
rect 92 3556 400 3579
rect 92 3459 155 3556
rect 362 3459 400 3556
rect -2305 3320 -2010 3365
rect -1583 3379 -1356 3412
rect -2584 3231 -2384 3257
rect -3169 3153 -2769 3174
rect -1583 3151 -1550 3379
rect -1387 3151 -1356 3379
rect -564 3353 -364 3381
rect -336 3372 -249 3456
rect -165 3452 -159 3456
rect -165 3372 -158 3452
rect 92 3439 400 3459
rect 1030 3422 1078 3696
rect 1933 3558 2137 3578
rect 1933 3451 2001 3558
rect -336 3368 -158 3372
rect -1132 3248 -732 3276
rect -1132 3174 -1103 3248
rect -763 3174 -732 3248
rect -564 3257 -537 3353
rect -388 3257 -364 3353
rect 100 3265 328 3411
rect 1177 3353 1377 3381
rect 1405 3367 1489 3451
rect 1573 3367 1579 3451
rect 1933 3439 2137 3451
rect 2792 3422 2856 3696
rect 3218 3535 3508 3553
rect -564 3231 -364 3257
rect -1132 3153 -732 3174
rect 99 3189 328 3265
rect 598 3248 998 3276
rect -1583 3118 -1356 3151
rect -3559 3037 -3350 3066
rect 99 3066 127 3189
rect 303 3066 327 3189
rect 598 3174 627 3248
rect 967 3174 998 3248
rect 1177 3257 1204 3353
rect 1353 3257 1377 3353
rect 1177 3231 1377 3257
rect 1752 3297 2088 3411
rect 598 3153 998 3174
rect 1752 3144 1803 3297
rect 2001 3144 2088 3297
rect 2956 3353 3156 3381
rect 3218 3379 3351 3535
rect 3465 3379 3508 3535
rect 3218 3366 3508 3379
rect 2358 3248 2758 3276
rect 2358 3174 2387 3248
rect 2727 3174 2758 3248
rect 2956 3257 2983 3353
rect 3132 3257 3156 3353
rect 2956 3231 3156 3257
rect 2358 3153 2758 3174
rect 1752 3116 2088 3144
rect 99 3043 327 3066
rect -2260 2840 8008 2924
rect -3817 2215 -3534 2234
rect -3818 2167 -3534 2215
rect -3818 1894 -3763 2167
rect -3574 1894 -3534 2167
rect -2540 2194 -2326 2216
rect -3353 2092 -2719 2126
rect -2540 2115 -2517 2194
rect -2348 2115 -2326 2194
rect -2540 2096 -2326 2115
rect -3353 1952 -3315 2092
rect -2761 1952 -2719 2092
rect -3353 1913 -2719 1952
rect -3818 1852 -3534 1894
rect -3818 1763 -3652 1852
rect -3818 1628 -3388 1763
rect -3818 -1502 -3652 1628
rect -2687 1610 -2639 1884
rect -2260 1615 -2166 2840
rect -2044 2693 -3 2777
rect -3571 1463 -3252 1599
rect -2540 1541 -2340 1569
rect -3571 1234 -3435 1463
rect -3118 1436 -2718 1464
rect -3118 1362 -3089 1436
rect -2749 1362 -2718 1436
rect -2540 1445 -2513 1541
rect -2364 1445 -2340 1541
rect -2540 1419 -2340 1445
rect -3118 1341 -2718 1362
rect -3571 480 -3435 1098
rect -2542 902 -2328 924
rect -3353 800 -2719 834
rect -2542 823 -2519 902
rect -2350 823 -2328 902
rect -2542 804 -2328 823
rect -3353 660 -3315 800
rect -2761 660 -2719 800
rect -2044 777 -1907 2693
rect -215 2545 -3 2629
rect -802 2194 -588 2216
rect -1617 2092 -983 2126
rect -802 2115 -779 2194
rect -610 2115 -588 2194
rect -802 2096 -588 2115
rect -1617 1952 -1579 2092
rect -1025 1952 -983 2092
rect -1617 1913 -983 1952
rect -1844 1750 -1611 1762
rect -1844 1637 -1792 1750
rect -1646 1637 -1611 1750
rect -1844 1628 -1611 1637
rect -949 1610 -901 1884
rect -215 1702 -84 2545
rect -3353 621 -2719 660
rect -3571 344 -3318 480
rect -2689 318 -2641 592
rect -3593 182 -3388 307
rect -3593 -16 -3568 182
rect -3422 -16 -3388 182
rect -2542 249 -2342 277
rect -2308 265 -1907 777
rect -1825 1463 -1516 1599
rect -802 1541 -602 1569
rect -528 1555 -84 1702
rect -1825 1240 -1689 1463
rect -1382 1436 -982 1464
rect -1382 1362 -1353 1436
rect -1013 1362 -982 1436
rect -802 1445 -775 1541
rect -626 1445 -602 1541
rect -802 1419 -602 1445
rect -1382 1341 -982 1362
rect -1825 1234 -1688 1240
rect -1825 1098 -1824 1234
rect -1825 1092 -1688 1098
rect -1825 472 -1689 1092
rect -808 902 -594 924
rect -1617 800 -983 834
rect -808 823 -785 902
rect -616 823 -594 902
rect -808 804 -594 823
rect -1617 660 -1579 800
rect -1025 660 -983 800
rect 12815 788 12906 1021
rect -1617 621 -983 660
rect -1825 336 -1570 472
rect -956 318 -908 592
rect -566 500 -260 526
rect -566 309 -516 500
rect -303 309 -260 500
rect -1868 295 -1580 307
rect -2308 263 -1968 265
rect -3118 144 -2718 172
rect -3118 70 -3089 144
rect -2749 70 -2718 144
rect -2542 153 -2515 249
rect -2366 153 -2342 249
rect -1868 185 -1840 295
rect -1608 185 -1580 295
rect -1868 172 -1580 185
rect -808 249 -608 277
rect -566 263 -260 309
rect -2542 127 -2342 153
rect -1382 144 -982 172
rect -3118 49 -2718 70
rect -1382 70 -1353 144
rect -1013 70 -982 144
rect -808 153 -781 249
rect -632 153 -608 249
rect -808 127 -608 153
rect -1382 49 -982 70
rect -3593 -31 -3388 -16
rect -2260 -341 -2166 -340
rect -2260 -425 9761 -341
rect -2541 -1071 -2327 -1049
rect -3353 -1173 -2719 -1139
rect -2541 -1150 -2518 -1071
rect -2349 -1150 -2327 -1071
rect -2541 -1169 -2327 -1150
rect -3353 -1313 -3315 -1173
rect -2761 -1313 -2719 -1173
rect -3353 -1352 -2719 -1313
rect -3818 -1637 -3388 -1502
rect -3818 -4766 -3652 -1637
rect -2688 -1655 -2640 -1381
rect -2260 -1649 -2166 -425
rect -2044 -572 -3 -488
rect -3588 -1680 -3298 -1666
rect -3588 -1784 -3567 -1680
rect -3324 -1784 -3298 -1680
rect -3588 -1802 -3298 -1784
rect -2541 -1724 -2341 -1696
rect -3118 -1829 -2718 -1801
rect -3118 -1903 -3089 -1829
rect -2749 -1903 -2718 -1829
rect -2541 -1820 -2514 -1724
rect -2365 -1820 -2341 -1724
rect -2541 -1846 -2341 -1820
rect -3118 -1924 -2718 -1903
rect -2539 -2363 -2325 -2341
rect -3353 -2465 -2719 -2431
rect -2539 -2442 -2516 -2363
rect -2347 -2442 -2325 -2363
rect -2539 -2461 -2325 -2442
rect -3353 -2605 -3315 -2465
rect -2761 -2605 -2719 -2465
rect -3353 -2644 -2719 -2605
rect -3588 -2808 -3388 -2794
rect -3588 -2915 -3557 -2808
rect -3401 -2915 -3388 -2808
rect -3588 -2929 -3388 -2915
rect -2687 -2947 -2639 -2673
rect -2044 -2674 -1907 -572
rect -215 -720 -3 -636
rect -806 -1071 -592 -1049
rect -1616 -1173 -982 -1139
rect -806 -1150 -783 -1071
rect -614 -1150 -592 -1071
rect -806 -1169 -592 -1150
rect -1616 -1313 -1578 -1173
rect -1024 -1313 -982 -1173
rect -1616 -1352 -982 -1313
rect -1798 -1518 -1623 -1502
rect -1798 -1625 -1764 -1518
rect -1644 -1625 -1623 -1518
rect -1798 -1637 -1623 -1625
rect -949 -1655 -901 -1381
rect -215 -1563 -84 -720
rect -1866 -1676 -1570 -1666
rect -1866 -1784 -1813 -1676
rect -1584 -1784 -1570 -1676
rect -1866 -1807 -1570 -1784
rect -806 -1724 -606 -1696
rect -531 -1710 -84 -1563
rect -1381 -1829 -981 -1801
rect -1381 -1903 -1352 -1829
rect -1012 -1903 -981 -1829
rect -806 -1820 -779 -1724
rect -630 -1820 -606 -1724
rect -806 -1846 -606 -1820
rect -1381 -1924 -981 -1903
rect -802 -2363 -588 -2341
rect -1617 -2465 -983 -2431
rect -802 -2442 -779 -2363
rect -610 -2442 -588 -2363
rect -802 -2461 -588 -2442
rect -1617 -2605 -1579 -2465
rect -1025 -2605 -983 -2465
rect 12859 -2477 12950 -2243
rect -1617 -2644 -983 -2605
rect -3593 -3083 -3388 -2958
rect -3593 -3281 -3568 -3083
rect -3422 -3281 -3388 -3083
rect -2539 -3016 -2339 -2988
rect -2307 -3000 -1907 -2674
rect -1866 -2795 -1644 -2794
rect -1866 -2806 -1614 -2795
rect -1866 -2917 -1841 -2806
rect -1639 -2917 -1614 -2806
rect -1866 -2929 -1614 -2917
rect -950 -2947 -902 -2673
rect -566 -2788 -260 -2739
rect -1869 -2980 -1609 -2958
rect -2307 -3002 -1968 -3000
rect -3118 -3121 -2718 -3093
rect -3118 -3195 -3089 -3121
rect -2749 -3195 -2718 -3121
rect -2539 -3112 -2512 -3016
rect -2363 -3112 -2339 -3016
rect -1869 -3072 -1847 -2980
rect -1642 -3072 -1609 -2980
rect -566 -2962 -529 -2788
rect -307 -2962 -260 -2788
rect -1869 -3094 -1609 -3072
rect -802 -3016 -602 -2988
rect -566 -3002 -260 -2962
rect -2539 -3138 -2339 -3112
rect -1382 -3121 -982 -3093
rect -3118 -3216 -2718 -3195
rect -1382 -3195 -1353 -3121
rect -1013 -3195 -982 -3121
rect -802 -3112 -775 -3016
rect -626 -3112 -602 -3016
rect -802 -3138 -602 -3112
rect -1382 -3216 -982 -3195
rect -3593 -3296 -3388 -3281
rect -2260 -3689 -3 -3605
rect -2539 -4335 -2325 -4313
rect -3353 -4437 -2719 -4403
rect -2539 -4414 -2516 -4335
rect -2347 -4414 -2325 -4335
rect -2539 -4433 -2325 -4414
rect -3353 -4577 -3315 -4437
rect -2761 -4577 -2719 -4437
rect -3353 -4616 -2719 -4577
rect -3818 -4901 -3388 -4766
rect -2687 -4919 -2639 -4645
rect -3588 -4956 -3225 -4930
rect -3588 -5047 -3519 -4956
rect -3291 -5047 -3225 -4956
rect -3588 -5066 -3225 -5047
rect -2539 -4988 -2339 -4960
rect -2260 -4974 -2167 -3689
rect -2044 -3836 -3 -3752
rect -3118 -5093 -2718 -5065
rect -3118 -5167 -3089 -5093
rect -2749 -5167 -2718 -5093
rect -2539 -5084 -2512 -4988
rect -2363 -5084 -2339 -4988
rect -2539 -5110 -2339 -5084
rect -3118 -5188 -2718 -5167
rect -2539 -5627 -2325 -5605
rect -3353 -5729 -2719 -5695
rect -2539 -5706 -2516 -5627
rect -2347 -5706 -2325 -5627
rect -2539 -5725 -2325 -5706
rect -3353 -5869 -3315 -5729
rect -2761 -5869 -2719 -5729
rect -2044 -5783 -1907 -3836
rect -215 -3984 -3 -3900
rect -806 -4335 -592 -4313
rect -1616 -4437 -982 -4403
rect -806 -4414 -783 -4335
rect -614 -4414 -592 -4335
rect -806 -4433 -592 -4414
rect -1616 -4577 -1578 -4437
rect -1024 -4577 -982 -4437
rect -1616 -4616 -982 -4577
rect -1848 -4788 -1564 -4766
rect -1848 -4882 -1788 -4788
rect -1606 -4882 -1564 -4788
rect -1848 -4900 -1564 -4882
rect -951 -4919 -903 -4645
rect -215 -4827 -84 -3984
rect -1848 -4948 -1564 -4930
rect -1848 -5044 -1804 -4948
rect -1600 -5044 -1564 -4948
rect -1848 -5066 -1564 -5044
rect -806 -4988 -606 -4960
rect -528 -4974 -84 -4827
rect -1381 -5093 -981 -5065
rect -1381 -5167 -1352 -5093
rect -1012 -5167 -981 -5093
rect -806 -5084 -779 -4988
rect -630 -5084 -606 -4988
rect -806 -5110 -606 -5084
rect -1381 -5188 -981 -5167
rect -810 -5627 -596 -5605
rect -3353 -5908 -2719 -5869
rect -3588 -6082 -3281 -6058
rect -3588 -6169 -3526 -6082
rect -3309 -6169 -3281 -6082
rect -3588 -6193 -3281 -6169
rect -2685 -6211 -2637 -5937
rect -3593 -6347 -3388 -6222
rect -3593 -6545 -3568 -6347
rect -3422 -6545 -3388 -6347
rect -2539 -6280 -2339 -6252
rect -2307 -6264 -1907 -5783
rect -1616 -5729 -982 -5695
rect -810 -5706 -787 -5627
rect -618 -5706 -596 -5627
rect -810 -5725 -596 -5706
rect -1616 -5869 -1578 -5729
rect -1024 -5869 -982 -5729
rect 12839 -5741 12930 -5505
rect -1616 -5908 -982 -5869
rect -1866 -6085 -1593 -6058
rect -1866 -6177 -1824 -6085
rect -1626 -6177 -1593 -6085
rect -1866 -6193 -1593 -6177
rect -958 -6211 -910 -5937
rect -566 -6045 -260 -6003
rect -1729 -6241 -1528 -6223
rect -2307 -6266 -1968 -6264
rect -3118 -6385 -2718 -6357
rect -3118 -6459 -3089 -6385
rect -2749 -6459 -2718 -6385
rect -2539 -6376 -2512 -6280
rect -2363 -6376 -2339 -6280
rect -1729 -6329 -1686 -6241
rect -1567 -6329 -1528 -6241
rect -566 -6231 -510 -6045
rect -311 -6231 -260 -6045
rect -1729 -6358 -1528 -6329
rect -810 -6280 -610 -6252
rect -566 -6266 -260 -6231
rect -2539 -6402 -2339 -6376
rect -1381 -6385 -981 -6357
rect -3118 -6480 -2718 -6459
rect -1381 -6459 -1352 -6385
rect -1012 -6459 -981 -6385
rect -810 -6376 -783 -6280
rect -634 -6376 -610 -6280
rect -810 -6402 -610 -6376
rect -1381 -6480 -981 -6459
rect -3593 -6560 -3388 -6545
<< via1 >>
rect -2561 3927 -2392 4006
rect -3366 3764 -2812 3904
rect -541 3927 -372 4006
rect -1329 3764 -775 3904
rect 1200 3927 1369 4006
rect 401 3764 955 3904
rect 2979 3927 3148 4006
rect 2161 3764 2715 3904
rect -3591 3440 -3448 3583
rect -3506 3066 -3384 3244
rect -3140 3174 -2800 3248
rect -2557 3257 -2408 3353
rect -2209 3365 -2077 3484
rect -1687 3464 -1369 3557
rect 155 3459 362 3556
rect -1550 3151 -1387 3379
rect -249 3372 -165 3456
rect 2001 3451 2150 3558
rect -1103 3174 -763 3248
rect -537 3257 -388 3353
rect 1489 3367 1573 3451
rect 127 3066 303 3189
rect 627 3174 967 3248
rect 1204 3257 1353 3353
rect 1803 3144 2001 3297
rect 3351 3379 3465 3535
rect 2387 3174 2727 3248
rect 2983 3257 3132 3353
rect -3763 1894 -3574 2167
rect -2517 2115 -2348 2194
rect -3315 1952 -2761 2092
rect -3089 1362 -2749 1436
rect -2513 1445 -2364 1541
rect -3571 1098 -3435 1234
rect -2519 823 -2350 902
rect -3315 660 -2761 800
rect -779 2115 -610 2194
rect -1579 1952 -1025 2092
rect -1792 1637 -1646 1750
rect -3568 -16 -3422 182
rect -1353 1362 -1013 1436
rect -775 1445 -626 1541
rect -1824 1098 -1688 1234
rect -785 823 -616 902
rect -1579 660 -1025 800
rect -516 309 -303 500
rect -3089 70 -2749 144
rect -2515 153 -2366 249
rect -1840 185 -1608 295
rect -1353 70 -1013 144
rect -781 153 -632 249
rect -2518 -1150 -2349 -1071
rect -3315 -1313 -2761 -1173
rect -3567 -1784 -3324 -1680
rect -3089 -1903 -2749 -1829
rect -2514 -1820 -2365 -1724
rect -2516 -2442 -2347 -2363
rect -3315 -2605 -2761 -2465
rect -3557 -2915 -3401 -2808
rect -783 -1150 -614 -1071
rect -1578 -1313 -1024 -1173
rect -1764 -1625 -1644 -1518
rect -1813 -1784 -1584 -1676
rect -1352 -1903 -1012 -1829
rect -779 -1820 -630 -1724
rect -779 -2442 -610 -2363
rect -1579 -2605 -1025 -2465
rect -3568 -3281 -3422 -3083
rect -1841 -2917 -1639 -2806
rect -3089 -3195 -2749 -3121
rect -2512 -3112 -2363 -3016
rect -1847 -3072 -1642 -2980
rect -529 -2962 -307 -2788
rect -1353 -3195 -1013 -3121
rect -775 -3112 -626 -3016
rect -2516 -4414 -2347 -4335
rect -3315 -4577 -2761 -4437
rect -3519 -5047 -3291 -4956
rect -3089 -5167 -2749 -5093
rect -2512 -5084 -2363 -4988
rect -2516 -5706 -2347 -5627
rect -3315 -5869 -2761 -5729
rect -783 -4414 -614 -4335
rect -1578 -4577 -1024 -4437
rect -1788 -4882 -1606 -4788
rect -1804 -5044 -1600 -4948
rect -1352 -5167 -1012 -5093
rect -779 -5084 -630 -4988
rect -3526 -6169 -3309 -6082
rect -3568 -6545 -3422 -6347
rect -787 -5706 -618 -5627
rect -1578 -5869 -1024 -5729
rect -1824 -6177 -1626 -6085
rect -3089 -6459 -2749 -6385
rect -2512 -6376 -2363 -6280
rect -1686 -6329 -1567 -6241
rect -510 -6231 -311 -6045
rect -1352 -6459 -1012 -6385
rect -783 -6376 -634 -6280
<< metal2 >>
rect -3591 4118 2084 4255
rect -3591 3583 -3448 4118
rect -2584 4006 -2370 4028
rect -3404 3904 -2770 3938
rect -2584 3927 -2561 4006
rect -2392 3927 -2370 4006
rect -2584 3908 -2370 3927
rect -3404 3764 -3366 3904
rect -2812 3764 -2770 3904
rect -3404 3725 -2770 3764
rect -1749 3576 -1606 4118
rect -564 4006 -350 4028
rect -1367 3904 -733 3938
rect -564 3927 -541 4006
rect -372 3927 -350 4006
rect -564 3908 -350 3927
rect -1367 3764 -1329 3904
rect -775 3764 -733 3904
rect -1367 3725 -733 3764
rect 92 3579 235 4118
rect 1177 4006 1391 4028
rect 363 3904 997 3938
rect 1177 3927 1200 4006
rect 1369 3927 1391 4006
rect 1177 3908 1391 3927
rect 363 3764 401 3904
rect 955 3764 997 3904
rect 363 3725 997 3764
rect -1749 3557 -1335 3576
rect -3591 3434 -3448 3440
rect -2251 3511 -2177 3515
rect -2251 3484 -2030 3511
rect -2584 3353 -2384 3381
rect -3559 3244 -3350 3291
rect -3559 3066 -3506 3244
rect -3384 3066 -3350 3244
rect -3169 3248 -2769 3276
rect -3169 3174 -3140 3248
rect -2800 3174 -2769 3248
rect -2584 3257 -2557 3353
rect -2408 3257 -2384 3353
rect -2251 3365 -2209 3484
rect -2077 3365 -2030 3484
rect -1749 3464 -1687 3557
rect -1369 3464 -1335 3557
rect 92 3556 400 3579
rect -1749 3440 -1335 3464
rect -275 3511 -244 3515
rect -275 3456 -135 3511
rect -2251 3324 -2030 3365
rect -2584 3231 -2384 3257
rect -3169 3153 -2769 3174
rect -3559 3037 -3350 3066
rect -2216 2727 -2030 3324
rect -1583 3379 -1356 3412
rect -1583 3151 -1550 3379
rect -1387 3151 -1356 3379
rect -564 3353 -364 3381
rect -1132 3248 -732 3276
rect -1132 3174 -1103 3248
rect -763 3174 -732 3248
rect -564 3257 -537 3353
rect -388 3257 -364 3353
rect -564 3231 -364 3257
rect -275 3372 -249 3456
rect -165 3372 -135 3456
rect 92 3459 155 3556
rect 362 3459 400 3556
rect 1933 3578 2076 4118
rect 2956 4006 3170 4028
rect 2123 3904 2757 3938
rect 2956 3927 2979 4006
rect 3148 3927 3170 4006
rect 2956 3908 3170 3927
rect 2123 3764 2161 3904
rect 2715 3764 2757 3904
rect 2123 3725 2757 3764
rect 1933 3558 2238 3578
rect 92 3439 400 3459
rect 1477 3510 1516 3515
rect 1477 3451 1600 3510
rect -1132 3153 -732 3174
rect -1583 3118 -1356 3151
rect -275 2833 -135 3372
rect 1177 3353 1377 3381
rect 598 3248 998 3276
rect 100 3189 318 3210
rect 100 3066 127 3189
rect 303 3066 318 3189
rect 598 3174 627 3248
rect 967 3174 998 3248
rect 1177 3257 1204 3353
rect 1353 3257 1377 3353
rect 1477 3367 1489 3451
rect 1573 3367 1600 3451
rect 1933 3451 2001 3558
rect 2150 3451 2238 3558
rect 1933 3439 2238 3451
rect 3318 3535 3608 3554
rect 1477 3327 1600 3367
rect 1177 3231 1377 3257
rect 598 3153 998 3174
rect 100 3045 318 3066
rect 1505 2985 1600 3327
rect 2956 3353 3156 3381
rect 3318 3379 3351 3535
rect 3465 3379 3608 3535
rect 3318 3367 3608 3379
rect 1752 3297 2032 3323
rect 1752 3144 1803 3297
rect 2001 3144 2032 3297
rect 2358 3248 2758 3276
rect 2358 3174 2387 3248
rect 2727 3174 2758 3248
rect 2956 3257 2983 3353
rect 3132 3257 3156 3353
rect 2956 3231 3156 3257
rect 2358 3153 2758 3174
rect 3453 3186 3608 3367
rect 1752 3116 2032 3144
rect 3453 3064 13159 3186
rect 3458 3036 13159 3064
rect 1505 2984 10159 2985
rect 1505 2876 10170 2984
rect -1285 2727 -968 2736
rect -2216 2666 -968 2727
rect -285 2722 6879 2833
rect -2216 2614 3582 2666
rect -1285 2553 3582 2614
rect -1285 2544 -968 2553
rect -1869 2517 -1700 2527
rect -1869 2489 -1407 2517
rect -1869 2383 -1556 2489
rect -1432 2383 -1407 2489
rect 3458 2408 3581 2553
rect -1869 2354 -1407 2383
rect 6750 2376 6878 2722
rect 10028 2388 10170 2876
rect -3817 2167 -3534 2234
rect -3817 1894 -3763 2167
rect -3574 1894 -3534 2167
rect -2540 2194 -2326 2216
rect -3353 2092 -2719 2126
rect -2540 2115 -2517 2194
rect -2348 2115 -2326 2194
rect -2540 2096 -2326 2115
rect -3353 1952 -3315 2092
rect -2761 1952 -2719 2092
rect -3353 1913 -2719 1952
rect -3817 1852 -3534 1894
rect -1869 1763 -1700 2354
rect -802 2194 -588 2216
rect -1617 2092 -983 2126
rect -802 2115 -779 2194
rect -610 2115 -588 2194
rect -802 2096 -588 2115
rect -1617 1952 -1579 2092
rect -1025 1952 -983 2092
rect -1617 1913 -983 1952
rect -2166 1762 -1692 1763
rect -2166 1751 -1611 1762
rect -2166 1637 -2151 1751
rect -2020 1750 -1611 1751
rect -2020 1637 -1792 1750
rect -1646 1637 -1611 1750
rect -2166 1628 -1611 1637
rect -2540 1541 -2340 1569
rect -3118 1436 -2718 1464
rect -3118 1362 -3089 1436
rect -2749 1362 -2718 1436
rect -2540 1445 -2513 1541
rect -2364 1445 -2340 1541
rect -802 1541 -602 1569
rect -2540 1419 -2340 1445
rect -1382 1436 -982 1464
rect -3118 1341 -2718 1362
rect -1382 1362 -1353 1436
rect -1013 1362 -982 1436
rect -802 1445 -775 1541
rect -626 1445 -602 1541
rect -312 1468 -3 1475
rect -802 1419 -602 1445
rect -1382 1341 -982 1362
rect -351 1335 -3 1468
rect -3578 1234 -3428 1242
rect -3578 1098 -3571 1234
rect -3435 1098 -1824 1234
rect -1688 1098 -1682 1234
rect -3578 1090 -3428 1098
rect -2542 902 -2328 924
rect -3353 800 -2719 834
rect -2542 823 -2519 902
rect -2350 823 -2328 902
rect -808 902 -594 924
rect -2542 804 -2328 823
rect -3353 660 -3315 800
rect -2761 660 -2719 800
rect -3353 621 -2719 660
rect -1617 800 -983 834
rect -808 823 -785 902
rect -616 823 -594 902
rect -808 804 -594 823
rect -1617 660 -1579 800
rect -1025 660 -983 800
rect -1617 621 -983 660
rect -518 526 -433 528
rect -351 526 -260 1335
rect -566 500 -260 526
rect -566 309 -516 500
rect -303 309 -260 500
rect -1868 295 -1580 307
rect -2542 249 -2342 277
rect -3593 182 -3395 211
rect -3593 -16 -3568 182
rect -3422 -16 -3395 182
rect -3118 144 -2718 172
rect -3118 70 -3089 144
rect -2749 70 -2718 144
rect -2542 153 -2515 249
rect -2366 153 -2342 249
rect -2542 127 -2342 153
rect -1868 185 -1840 295
rect -1608 185 -1580 295
rect -3118 49 -2718 70
rect -3593 -31 -3395 -16
rect -1868 -210 -1818 185
rect -1729 172 -1580 185
rect -808 249 -608 277
rect -566 263 -260 309
rect -1729 -108 -1692 172
rect -1382 144 -982 172
rect -1382 70 -1353 144
rect -1013 70 -982 144
rect -808 153 -781 249
rect -632 153 -608 249
rect -808 127 -608 153
rect -1382 49 -982 70
rect -1729 -210 -1693 -108
rect -1868 -254 -1693 -210
rect 10 -200 287 -196
rect 10 -401 315 -200
rect 3275 -213 3407 -128
rect 6574 -187 6881 -83
rect 3275 -343 3638 -213
rect 3342 -344 3638 -343
rect -3604 -447 -299 -427
rect -3604 -453 -471 -447
rect -3604 -593 -3575 -453
rect -3446 -587 -471 -453
rect -342 -587 -299 -447
rect -3446 -593 -299 -587
rect -3604 -614 -299 -593
rect 171 -822 315 -401
rect 3452 -848 3636 -344
rect 6755 -863 6878 -187
rect 9870 -241 9997 -101
rect 13154 -136 13282 56
rect 10040 -241 10168 -240
rect 9865 -397 10168 -241
rect 9870 -398 9997 -397
rect 10040 -839 10168 -397
rect -2541 -1071 -2327 -1049
rect -3353 -1173 -2719 -1139
rect -2541 -1150 -2518 -1071
rect -2349 -1150 -2327 -1071
rect -806 -1071 -592 -1049
rect -2541 -1169 -2327 -1150
rect -3353 -1313 -3315 -1173
rect -2761 -1313 -2719 -1173
rect -3353 -1352 -2719 -1313
rect -1616 -1173 -982 -1139
rect -806 -1150 -783 -1071
rect -614 -1150 -592 -1071
rect -806 -1169 -592 -1150
rect -1616 -1313 -1578 -1173
rect -1024 -1313 -982 -1173
rect -1616 -1352 -982 -1313
rect -2166 -1512 -1623 -1502
rect -2166 -1626 -2154 -1512
rect -2023 -1514 -1623 -1512
rect -2020 -1518 -1623 -1514
rect -2020 -1625 -1764 -1518
rect -1644 -1625 -1623 -1518
rect -2166 -1628 -2151 -1626
rect -2020 -1628 -1623 -1625
rect -2166 -1637 -1623 -1628
rect -3588 -1680 -3298 -1666
rect -3588 -1784 -3567 -1680
rect -3324 -1784 -3298 -1680
rect -1866 -1676 -1570 -1666
rect -3588 -1802 -3298 -1784
rect -2541 -1724 -2341 -1696
rect -3588 -2061 -3412 -1802
rect -3118 -1829 -2718 -1801
rect -3118 -1903 -3089 -1829
rect -2749 -1903 -2718 -1829
rect -2541 -1820 -2514 -1724
rect -2365 -1820 -2341 -1724
rect -2541 -1846 -2341 -1820
rect -1866 -1784 -1813 -1676
rect -1584 -1784 -1570 -1676
rect -1866 -1807 -1570 -1784
rect -806 -1724 -606 -1696
rect -3118 -1924 -2718 -1903
rect -1866 -2061 -1690 -1807
rect -1381 -1829 -981 -1801
rect -1381 -1903 -1352 -1829
rect -1012 -1903 -981 -1829
rect -806 -1820 -779 -1724
rect -630 -1820 -606 -1724
rect -312 -1797 -3 -1790
rect -806 -1846 -606 -1820
rect -1381 -1924 -981 -1903
rect -3590 -2196 -1690 -2061
rect -3588 -2794 -3412 -2196
rect -2539 -2363 -2325 -2341
rect -3353 -2465 -2719 -2431
rect -2539 -2442 -2516 -2363
rect -2347 -2442 -2325 -2363
rect -2539 -2461 -2325 -2442
rect -3353 -2605 -3315 -2465
rect -2761 -2605 -2719 -2465
rect -3353 -2644 -2719 -2605
rect -1866 -2794 -1690 -2196
rect -351 -1930 -3 -1797
rect -802 -2363 -588 -2341
rect -1617 -2465 -983 -2431
rect -802 -2442 -779 -2363
rect -610 -2442 -588 -2363
rect -802 -2461 -588 -2442
rect -1617 -2605 -1579 -2465
rect -1025 -2605 -983 -2465
rect -1617 -2644 -983 -2605
rect -518 -2739 -433 -2737
rect -351 -2739 -260 -1930
rect -566 -2788 -260 -2739
rect -3588 -2808 -3388 -2794
rect -3588 -2915 -3557 -2808
rect -3401 -2915 -3388 -2808
rect -3588 -2929 -3388 -2915
rect -1866 -2795 -1644 -2794
rect -1866 -2806 -1614 -2795
rect -1866 -2917 -1841 -2806
rect -1639 -2917 -1614 -2806
rect -1866 -2929 -1614 -2917
rect -1869 -2980 -1609 -2958
rect -2539 -3016 -2339 -2988
rect -3593 -3083 -3395 -3054
rect -3593 -3281 -3568 -3083
rect -3422 -3281 -3395 -3083
rect -3118 -3121 -2718 -3093
rect -3118 -3195 -3089 -3121
rect -2749 -3195 -2718 -3121
rect -2539 -3112 -2512 -3016
rect -2363 -3112 -2339 -3016
rect -1869 -3072 -1847 -2980
rect -1642 -3072 -1609 -2980
rect -566 -2962 -529 -2788
rect -307 -2962 -260 -2788
rect -1869 -3094 -1822 -3072
rect -2539 -3138 -2339 -3112
rect -3118 -3216 -2718 -3195
rect -3593 -3296 -3395 -3281
rect -1867 -3454 -1822 -3094
rect -1729 -3094 -1609 -3072
rect -802 -3016 -602 -2988
rect -566 -3002 -260 -2962
rect -1729 -3373 -1692 -3094
rect -1382 -3121 -982 -3093
rect -1382 -3195 -1353 -3121
rect -1013 -3195 -982 -3121
rect -802 -3112 -775 -3016
rect -626 -3112 -602 -3016
rect -802 -3138 -602 -3112
rect -1382 -3216 -982 -3195
rect -1867 -3475 -1818 -3454
rect -1729 -3475 -1693 -3373
rect -1867 -3519 -1693 -3475
rect -11 -3621 314 -3495
rect 3281 -3497 3615 -3375
rect 169 -4142 299 -3621
rect 3456 -4161 3592 -3497
rect 6570 -3532 6886 -3387
rect 9874 -3505 10165 -3369
rect 13156 -3414 13288 -3296
rect 6744 -4189 6874 -3532
rect 10040 -4161 10164 -3505
rect -2539 -4335 -2325 -4313
rect -3353 -4437 -2719 -4403
rect -2539 -4414 -2516 -4335
rect -2347 -4414 -2325 -4335
rect -806 -4335 -592 -4313
rect -2539 -4433 -2325 -4414
rect -3353 -4577 -3315 -4437
rect -2761 -4577 -2719 -4437
rect -3353 -4616 -2719 -4577
rect -1616 -4437 -982 -4403
rect -806 -4414 -783 -4335
rect -614 -4414 -592 -4335
rect -806 -4433 -592 -4414
rect -1616 -4577 -1578 -4437
rect -1024 -4577 -982 -4437
rect -1616 -4616 -982 -4577
rect -2166 -4776 -1533 -4766
rect -2166 -4890 -2154 -4776
rect -2017 -4788 -1533 -4776
rect -2017 -4882 -1788 -4788
rect -1606 -4882 -1533 -4788
rect -2017 -4890 -1533 -4882
rect -2166 -4892 -2151 -4890
rect -2020 -4892 -1533 -4890
rect -2166 -4901 -1533 -4892
rect -3588 -4956 -3225 -4930
rect -3588 -5047 -3519 -4956
rect -3291 -5047 -3225 -4956
rect -1866 -4948 -1547 -4930
rect -3588 -5066 -3225 -5047
rect -2539 -4988 -2339 -4960
rect -3588 -5325 -3412 -5066
rect -3118 -5093 -2718 -5065
rect -3118 -5167 -3089 -5093
rect -2749 -5167 -2718 -5093
rect -2539 -5084 -2512 -4988
rect -2363 -5084 -2339 -4988
rect -2539 -5110 -2339 -5084
rect -1866 -5044 -1804 -4948
rect -1600 -5044 -1547 -4948
rect -1866 -5066 -1547 -5044
rect -806 -4988 -606 -4960
rect -3118 -5188 -2718 -5167
rect -1866 -5325 -1690 -5066
rect -1381 -5093 -981 -5065
rect -1381 -5167 -1352 -5093
rect -1012 -5167 -981 -5093
rect -806 -5084 -779 -4988
rect -630 -5084 -606 -4988
rect -312 -5061 -3 -5054
rect -806 -5110 -606 -5084
rect -1381 -5188 -981 -5167
rect -3590 -5460 -1690 -5325
rect -3588 -6058 -3412 -5460
rect -2539 -5627 -2325 -5605
rect -3353 -5729 -2719 -5695
rect -2539 -5706 -2516 -5627
rect -2347 -5706 -2325 -5627
rect -2539 -5725 -2325 -5706
rect -3353 -5869 -3315 -5729
rect -2761 -5869 -2719 -5729
rect -3353 -5908 -2719 -5869
rect -1866 -6058 -1690 -5460
rect -351 -5194 -3 -5061
rect -810 -5627 -596 -5605
rect -1616 -5729 -982 -5695
rect -810 -5706 -787 -5627
rect -618 -5706 -596 -5627
rect -810 -5725 -596 -5706
rect -1616 -5869 -1578 -5729
rect -1024 -5869 -982 -5729
rect -1616 -5908 -982 -5869
rect -518 -6003 -433 -6001
rect -351 -6003 -260 -5194
rect -566 -6045 -260 -6003
rect -3588 -6082 -3281 -6058
rect -3588 -6169 -3526 -6082
rect -3309 -6169 -3281 -6082
rect -3588 -6193 -3281 -6169
rect -1866 -6085 -1593 -6058
rect -1866 -6177 -1824 -6085
rect -1626 -6177 -1593 -6085
rect -1866 -6193 -1593 -6177
rect -1867 -6229 -1528 -6223
rect -1868 -6241 -1528 -6229
rect -2539 -6280 -2339 -6252
rect -3593 -6347 -3395 -6318
rect -3593 -6545 -3568 -6347
rect -3422 -6545 -3395 -6347
rect -3118 -6385 -2718 -6357
rect -3118 -6459 -3089 -6385
rect -2749 -6459 -2718 -6385
rect -2539 -6376 -2512 -6280
rect -2363 -6376 -2339 -6280
rect -2539 -6402 -2339 -6376
rect -1868 -6272 -1686 -6241
rect -1868 -6287 -1822 -6272
rect -3118 -6480 -2718 -6459
rect -3593 -6560 -3395 -6545
rect -1868 -6733 -1825 -6287
rect -1733 -6293 -1686 -6272
rect -1729 -6329 -1686 -6293
rect -1567 -6329 -1528 -6241
rect -566 -6231 -510 -6045
rect -311 -6231 -260 -6045
rect -1729 -6358 -1528 -6329
rect -810 -6280 -610 -6252
rect -566 -6266 -260 -6231
rect -1729 -6637 -1692 -6358
rect -1381 -6385 -981 -6357
rect -1381 -6459 -1352 -6385
rect -1012 -6459 -981 -6385
rect -810 -6376 -783 -6280
rect -634 -6376 -610 -6280
rect -810 -6402 -610 -6376
rect -1381 -6480 -981 -6459
rect -1868 -6739 -1818 -6733
rect -1729 -6739 -1693 -6637
rect -1868 -6783 -1693 -6739
rect 5 -6819 190 -6596
rect 3288 -6679 3396 -6550
rect 6579 -6679 6688 -6554
rect 9870 -6679 9978 -6550
rect 13156 -6678 13288 -6560
<< via2 >>
rect -2561 3927 -2392 4006
rect -3366 3764 -2812 3904
rect -541 3927 -372 4006
rect -1329 3764 -775 3904
rect 1200 3927 1369 4006
rect 401 3764 955 3904
rect -3506 3066 -3384 3244
rect -3140 3174 -2800 3248
rect -2557 3257 -2408 3353
rect -1550 3151 -1387 3379
rect -1103 3174 -763 3248
rect -537 3257 -388 3353
rect 2979 3927 3148 4006
rect 2161 3764 2715 3904
rect 127 3066 303 3189
rect 627 3174 967 3248
rect 1204 3257 1353 3353
rect 1803 3144 2001 3297
rect 2387 3174 2727 3248
rect 2983 3257 3132 3353
rect -1556 2383 -1432 2489
rect -3763 1894 -3574 2167
rect -2517 2115 -2348 2194
rect -3315 1952 -2761 2092
rect -779 2115 -610 2194
rect -1579 1952 -1025 2092
rect -2151 1637 -2020 1751
rect -3089 1362 -2749 1436
rect -2513 1445 -2364 1541
rect -1353 1362 -1013 1436
rect -775 1445 -626 1541
rect -2519 823 -2350 902
rect -3315 660 -2761 800
rect -785 823 -616 902
rect -1579 660 -1025 800
rect -3568 -16 -3422 182
rect -3089 70 -2749 144
rect -2515 153 -2366 249
rect -1818 185 -1729 236
rect -1818 -210 -1729 185
rect -1353 70 -1013 144
rect -781 153 -632 249
rect -3575 -593 -3446 -453
rect -471 -587 -342 -447
rect -2518 -1150 -2349 -1071
rect -3315 -1313 -2761 -1173
rect -783 -1150 -614 -1071
rect -1578 -1313 -1024 -1173
rect -2154 -1514 -2023 -1512
rect -2154 -1626 -2020 -1514
rect -2151 -1628 -2020 -1626
rect -3089 -1903 -2749 -1829
rect -2514 -1820 -2365 -1724
rect -1352 -1903 -1012 -1829
rect -779 -1820 -630 -1724
rect -2516 -2442 -2347 -2363
rect -3315 -2605 -2761 -2465
rect -779 -2442 -610 -2363
rect -1579 -2605 -1025 -2465
rect -3568 -3281 -3422 -3083
rect -3089 -3195 -2749 -3121
rect -2512 -3112 -2363 -3016
rect -1822 -3029 -1733 -3008
rect -1822 -3072 -1729 -3029
rect -1822 -3454 -1729 -3072
rect -1353 -3195 -1013 -3121
rect -775 -3112 -626 -3016
rect -1818 -3475 -1729 -3454
rect -2516 -4414 -2347 -4335
rect -3315 -4577 -2761 -4437
rect -783 -4414 -614 -4335
rect -1578 -4577 -1024 -4437
rect -2154 -4890 -2017 -4776
rect -2151 -4892 -2020 -4890
rect -3089 -5167 -2749 -5093
rect -2512 -5084 -2363 -4988
rect -1352 -5167 -1012 -5093
rect -779 -5084 -630 -4988
rect -2516 -5706 -2347 -5627
rect -3315 -5869 -2761 -5729
rect -787 -5706 -618 -5627
rect -1578 -5869 -1024 -5729
rect -3568 -6545 -3422 -6347
rect -3089 -6459 -2749 -6385
rect -2512 -6376 -2363 -6280
rect -1822 -6287 -1733 -6272
rect -1825 -6293 -1733 -6287
rect -1825 -6733 -1729 -6293
rect -1352 -6459 -1012 -6385
rect -783 -6376 -634 -6280
rect -1818 -6739 -1729 -6733
<< metal3 >>
rect -3817 4255 -3635 4259
rect -3817 4090 1969 4255
rect -3817 2234 -3635 4090
rect -2584 4006 -2370 4028
rect -3404 3904 -2770 3938
rect -2584 3927 -2561 4006
rect -2392 3927 -2370 4006
rect -564 4006 -350 4028
rect -2584 3908 -2370 3927
rect -3404 3764 -3366 3904
rect -2812 3764 -2770 3904
rect -3404 3725 -2770 3764
rect -1367 3904 -733 3938
rect -564 3927 -541 4006
rect -372 3927 -350 4006
rect 1177 4006 1391 4028
rect -564 3908 -350 3927
rect -1367 3764 -1329 3904
rect -775 3764 -733 3904
rect -1367 3725 -733 3764
rect 363 3904 997 3938
rect 1177 3927 1200 4006
rect 1369 3927 1391 4006
rect 1177 3908 1391 3927
rect 363 3764 401 3904
rect 955 3764 997 3904
rect 363 3725 997 3764
rect -3544 3291 -3354 3372
rect -2584 3353 -2384 3381
rect -3559 3244 -3350 3291
rect -3559 3066 -3506 3244
rect -3384 3066 -3350 3244
rect -3169 3248 -2769 3276
rect -3169 3174 -3140 3248
rect -2800 3174 -2769 3248
rect -2584 3257 -2557 3353
rect -2408 3257 -2384 3353
rect -2584 3231 -2384 3257
rect -1583 3379 -1356 3412
rect -3169 3153 -2769 3174
rect -3559 3037 -3350 3066
rect -1583 3151 -1550 3379
rect -1387 3151 -1356 3379
rect -564 3353 -364 3381
rect -1132 3248 -732 3276
rect -1132 3174 -1103 3248
rect -763 3174 -732 3248
rect -564 3257 -537 3353
rect -388 3257 -364 3353
rect 1177 3353 1377 3381
rect -564 3231 -364 3257
rect 598 3248 998 3276
rect -1132 3153 -732 3174
rect 100 3189 318 3210
rect -1583 3118 -1356 3151
rect -3542 2836 -3358 3037
rect -3542 2832 -1710 2836
rect -3542 2636 -1708 2832
rect -3817 2167 -3534 2234
rect -3817 1894 -3763 2167
rect -3574 1894 -3534 2167
rect -2540 2194 -2326 2216
rect -3353 2092 -2719 2126
rect -2540 2115 -2517 2194
rect -2348 2115 -2326 2194
rect -2540 2096 -2326 2115
rect -3353 1952 -3315 2092
rect -2761 1952 -2719 2092
rect -3353 1913 -2719 1952
rect -3817 1852 -3534 1894
rect -2166 1751 -2007 1796
rect -2166 1637 -2151 1751
rect -2020 1637 -2007 1751
rect -2540 1541 -2340 1569
rect -3118 1436 -2718 1464
rect -3118 1362 -3089 1436
rect -2749 1362 -2718 1436
rect -2540 1445 -2513 1541
rect -2364 1445 -2340 1541
rect -2540 1419 -2340 1445
rect -3118 1341 -2718 1362
rect -2542 902 -2328 924
rect -3353 800 -2719 834
rect -2542 823 -2519 902
rect -2350 823 -2328 902
rect -2542 804 -2328 823
rect -3353 660 -3315 800
rect -2761 660 -2719 800
rect -3353 621 -2719 660
rect -3607 211 -3416 332
rect -2542 249 -2342 277
rect -3607 182 -3395 211
rect -3607 -16 -3568 182
rect -3422 -16 -3395 182
rect -3118 144 -2718 172
rect -3118 70 -3089 144
rect -2749 70 -2718 144
rect -2542 153 -2515 249
rect -2366 153 -2342 249
rect -2542 127 -2342 153
rect -3118 49 -2718 70
rect -3607 -31 -3395 -16
rect -3607 -453 -3416 -31
rect -3607 -593 -3575 -453
rect -3446 -593 -3416 -453
rect -3607 -3054 -3416 -593
rect -2541 -1071 -2327 -1049
rect -3353 -1173 -2719 -1139
rect -2541 -1150 -2518 -1071
rect -2349 -1150 -2327 -1071
rect -2541 -1169 -2327 -1150
rect -3353 -1313 -3315 -1173
rect -2761 -1313 -2719 -1173
rect -3353 -1352 -2719 -1313
rect -2166 -1512 -2007 1637
rect -2166 -1626 -2154 -1512
rect -2023 -1514 -2007 -1512
rect -2166 -1628 -2151 -1626
rect -2020 -1628 -2007 -1514
rect -2541 -1724 -2341 -1696
rect -3118 -1829 -2718 -1801
rect -3118 -1903 -3089 -1829
rect -2749 -1903 -2718 -1829
rect -2541 -1820 -2514 -1724
rect -2365 -1820 -2341 -1724
rect -2541 -1846 -2341 -1820
rect -3118 -1924 -2718 -1903
rect -2539 -2363 -2325 -2341
rect -3353 -2465 -2719 -2431
rect -2539 -2442 -2516 -2363
rect -2347 -2442 -2325 -2363
rect -2539 -2461 -2325 -2442
rect -3353 -2605 -3315 -2465
rect -2761 -2605 -2719 -2465
rect -3353 -2644 -2719 -2605
rect -2539 -3016 -2339 -2988
rect -3607 -3083 -3395 -3054
rect -3607 -3281 -3568 -3083
rect -3422 -3281 -3395 -3083
rect -3118 -3121 -2718 -3093
rect -3118 -3195 -3089 -3121
rect -2749 -3195 -2718 -3121
rect -2539 -3112 -2512 -3016
rect -2363 -3112 -2339 -3016
rect -2539 -3138 -2339 -3112
rect -3118 -3216 -2718 -3195
rect -3607 -3296 -3395 -3281
rect -3607 -6318 -3416 -3296
rect -2539 -4335 -2325 -4313
rect -3353 -4437 -2719 -4403
rect -2539 -4414 -2516 -4335
rect -2347 -4414 -2325 -4335
rect -2539 -4433 -2325 -4414
rect -3353 -4577 -3315 -4437
rect -2761 -4577 -2719 -4437
rect -3353 -4616 -2719 -4577
rect -2166 -4776 -2007 -1628
rect -2166 -4890 -2154 -4776
rect -2017 -4890 -2007 -4776
rect -2166 -4892 -2151 -4890
rect -2020 -4892 -2007 -4890
rect -2166 -4901 -2007 -4892
rect -1893 236 -1708 2636
rect -1583 2489 -1415 3118
rect 100 3066 127 3189
rect 303 3066 318 3189
rect 598 3174 627 3248
rect 967 3174 998 3248
rect 1177 3257 1204 3353
rect 1353 3257 1377 3353
rect 1177 3231 1377 3257
rect 1752 3323 1969 4090
rect 2956 4006 3170 4028
rect 2123 3904 2757 3938
rect 2956 3927 2979 4006
rect 3148 3927 3170 4006
rect 2956 3908 3170 3927
rect 2123 3764 2161 3904
rect 2715 3764 2757 3904
rect 2123 3725 2757 3764
rect 2956 3353 3156 3381
rect 1752 3297 2032 3323
rect 598 3153 998 3174
rect 1752 3144 1803 3297
rect 2001 3144 2032 3297
rect 2358 3248 2758 3276
rect 2358 3174 2387 3248
rect 2727 3174 2758 3248
rect 2956 3257 2983 3353
rect 3132 3257 3156 3353
rect 2956 3231 3156 3257
rect 2358 3153 2758 3174
rect 1752 3116 2032 3144
rect 100 3052 318 3066
rect -480 3045 318 3052
rect -480 3033 271 3045
rect -1583 2383 -1556 2489
rect -1432 2383 -1415 2489
rect -1583 2362 -1415 2383
rect -481 2868 271 3033
rect -481 2858 265 2868
rect -802 2194 -588 2216
rect -1617 2092 -983 2126
rect -802 2115 -779 2194
rect -610 2115 -588 2194
rect -802 2096 -588 2115
rect -1617 1952 -1579 2092
rect -1025 1952 -983 2092
rect -1617 1913 -983 1952
rect -802 1541 -602 1569
rect -1382 1436 -982 1464
rect -1382 1362 -1353 1436
rect -1013 1362 -982 1436
rect -802 1445 -775 1541
rect -626 1445 -602 1541
rect -802 1419 -602 1445
rect -1382 1341 -982 1362
rect -808 902 -594 924
rect -1617 800 -983 834
rect -808 823 -785 902
rect -616 823 -594 902
rect -808 804 -594 823
rect -1617 660 -1579 800
rect -1025 660 -983 800
rect -1617 621 -983 660
rect -1893 -210 -1818 236
rect -1729 -210 -1708 236
rect -808 249 -608 277
rect -1382 144 -982 172
rect -1382 70 -1353 144
rect -1013 70 -982 144
rect -808 153 -781 249
rect -632 153 -608 249
rect -808 127 -608 153
rect -1382 49 -982 70
rect -1893 -3008 -1708 -210
rect -481 -447 -301 2858
rect -481 -587 -471 -447
rect -342 -587 -301 -447
rect -481 -623 -301 -587
rect -806 -1071 -592 -1049
rect -1616 -1173 -982 -1139
rect -806 -1150 -783 -1071
rect -614 -1150 -592 -1071
rect -806 -1169 -592 -1150
rect -1616 -1313 -1578 -1173
rect -1024 -1313 -982 -1173
rect -1616 -1352 -982 -1313
rect -806 -1724 -606 -1696
rect -1381 -1829 -981 -1801
rect -1381 -1903 -1352 -1829
rect -1012 -1903 -981 -1829
rect -806 -1820 -779 -1724
rect -630 -1820 -606 -1724
rect -806 -1846 -606 -1820
rect -1381 -1924 -981 -1903
rect -802 -2363 -588 -2341
rect -1617 -2465 -983 -2431
rect -802 -2442 -779 -2363
rect -610 -2442 -588 -2363
rect -802 -2461 -588 -2442
rect -1617 -2605 -1579 -2465
rect -1025 -2605 -983 -2465
rect -1617 -2644 -983 -2605
rect -1893 -3454 -1822 -3008
rect -1733 -3029 -1708 -3008
rect -1893 -3475 -1818 -3454
rect -1729 -3475 -1708 -3029
rect -802 -3016 -602 -2988
rect -1382 -3121 -982 -3093
rect -1382 -3195 -1353 -3121
rect -1013 -3195 -982 -3121
rect -802 -3112 -775 -3016
rect -626 -3112 -602 -3016
rect -802 -3138 -602 -3112
rect -1382 -3216 -982 -3195
rect -1893 -4788 -1708 -3475
rect -806 -4335 -592 -4313
rect -1616 -4437 -982 -4403
rect -806 -4414 -783 -4335
rect -614 -4414 -592 -4335
rect -806 -4433 -592 -4414
rect -1616 -4577 -1578 -4437
rect -1024 -4577 -982 -4437
rect -1616 -4616 -982 -4577
rect -1893 -4882 -1606 -4788
rect -1893 -4948 -1708 -4882
rect -2539 -4988 -2339 -4960
rect -3118 -5093 -2718 -5065
rect -3118 -5167 -3089 -5093
rect -2749 -5167 -2718 -5093
rect -2539 -5084 -2512 -4988
rect -2363 -5084 -2339 -4988
rect -2539 -5110 -2339 -5084
rect -1893 -5044 -1600 -4948
rect -806 -4988 -606 -4960
rect -3118 -5188 -2718 -5167
rect -2539 -5627 -2325 -5605
rect -3353 -5729 -2719 -5695
rect -2539 -5706 -2516 -5627
rect -2347 -5706 -2325 -5627
rect -2539 -5725 -2325 -5706
rect -3353 -5869 -3315 -5729
rect -2761 -5869 -2719 -5729
rect -3353 -5908 -2719 -5869
rect -2539 -6280 -2339 -6252
rect -3607 -6347 -3395 -6318
rect -3607 -6545 -3568 -6347
rect -3422 -6545 -3395 -6347
rect -3118 -6385 -2718 -6357
rect -3118 -6459 -3089 -6385
rect -2749 -6459 -2718 -6385
rect -2539 -6376 -2512 -6280
rect -2363 -6376 -2339 -6280
rect -2539 -6402 -2339 -6376
rect -1893 -6272 -1708 -5044
rect -1381 -5093 -981 -5065
rect -1381 -5167 -1352 -5093
rect -1012 -5167 -981 -5093
rect -806 -5084 -779 -4988
rect -630 -5084 -606 -4988
rect -806 -5110 -606 -5084
rect -1381 -5188 -981 -5167
rect -810 -5627 -596 -5605
rect -1616 -5729 -982 -5695
rect -810 -5706 -787 -5627
rect -618 -5706 -596 -5627
rect -810 -5725 -596 -5706
rect -1616 -5869 -1578 -5729
rect -1024 -5869 -982 -5729
rect -1616 -5908 -982 -5869
rect -1893 -6287 -1822 -6272
rect -3118 -6480 -2718 -6459
rect -3607 -6560 -3395 -6545
rect -3607 -6772 -3416 -6560
rect -1893 -6733 -1825 -6287
rect -1733 -6293 -1708 -6272
rect -1893 -6739 -1818 -6733
rect -1729 -6739 -1708 -6293
rect -810 -6280 -610 -6252
rect -1381 -6385 -981 -6357
rect -1381 -6459 -1352 -6385
rect -1012 -6459 -981 -6385
rect -810 -6376 -783 -6280
rect -634 -6376 -610 -6280
rect -810 -6402 -610 -6376
rect -1381 -6480 -981 -6459
rect -1893 -6782 -1708 -6739
<< via3 >>
rect -2561 3927 -2392 4006
rect -3366 3764 -2812 3904
rect -541 3927 -372 4006
rect -1329 3764 -775 3904
rect 1200 3927 1369 4006
rect 401 3764 955 3904
rect -3140 3174 -2800 3248
rect -2557 3257 -2408 3353
rect -1103 3174 -763 3248
rect -537 3257 -388 3353
rect -2517 2115 -2348 2194
rect -3315 1952 -2761 2092
rect -3089 1362 -2749 1436
rect -2513 1445 -2364 1541
rect -2519 823 -2350 902
rect -3315 660 -2761 800
rect -3089 70 -2749 144
rect -2515 153 -2366 249
rect -2518 -1150 -2349 -1071
rect -3315 -1313 -2761 -1173
rect -3089 -1903 -2749 -1829
rect -2514 -1820 -2365 -1724
rect -2516 -2442 -2347 -2363
rect -3315 -2605 -2761 -2465
rect -3089 -3195 -2749 -3121
rect -2512 -3112 -2363 -3016
rect -2516 -4414 -2347 -4335
rect -3315 -4577 -2761 -4437
rect 627 3174 967 3248
rect 1204 3257 1353 3353
rect 2979 3927 3148 4006
rect 2161 3764 2715 3904
rect 2387 3174 2727 3248
rect 2983 3257 3132 3353
rect -779 2115 -610 2194
rect -1579 1952 -1025 2092
rect -1353 1362 -1013 1436
rect -775 1445 -626 1541
rect -785 823 -616 902
rect -1579 660 -1025 800
rect -1353 70 -1013 144
rect -781 153 -632 249
rect -783 -1150 -614 -1071
rect -1578 -1313 -1024 -1173
rect -1352 -1903 -1012 -1829
rect -779 -1820 -630 -1724
rect -779 -2442 -610 -2363
rect -1579 -2605 -1025 -2465
rect -1353 -3195 -1013 -3121
rect -775 -3112 -626 -3016
rect -783 -4414 -614 -4335
rect -1578 -4577 -1024 -4437
rect -3089 -5167 -2749 -5093
rect -2512 -5084 -2363 -4988
rect -2516 -5706 -2347 -5627
rect -3315 -5869 -2761 -5729
rect -3089 -6459 -2749 -6385
rect -2512 -6376 -2363 -6280
rect -1352 -5167 -1012 -5093
rect -779 -5084 -630 -4988
rect -787 -5706 -618 -5627
rect -1578 -5869 -1024 -5729
rect -1352 -6459 -1012 -6385
rect -783 -6376 -634 -6280
<< metal4 >>
rect -3405 4141 3263 4142
rect -3405 4006 3690 4141
rect -3405 3927 -2561 4006
rect -2392 3927 -541 4006
rect -372 3927 1200 4006
rect 1369 3927 2979 4006
rect 3148 3927 3690 4006
rect -3405 3904 3690 3927
rect -3405 3764 -3366 3904
rect -2812 3764 -1329 3904
rect -775 3764 401 3904
rect 955 3764 2161 3904
rect 2715 3764 3690 3904
rect -3405 3725 3690 3764
rect -3204 3353 -328 3446
rect -3204 3348 -2557 3353
rect -2408 3348 -537 3353
rect -3204 3248 -2943 3348
rect -673 3257 -537 3348
rect -388 3257 -328 3353
rect -3204 3174 -3140 3248
rect -3204 3040 -2943 3174
rect -673 3040 -328 3257
rect -3204 2982 -328 3040
rect -51 2524 282 3725
rect 3243 3724 3690 3725
rect 559 3353 3193 3412
rect 559 3317 1204 3353
rect 1353 3317 2983 3353
rect 559 3248 797 3317
rect 3132 3257 3193 3353
rect 559 3174 627 3248
rect 559 3009 797 3174
rect 3067 3009 3193 3257
rect 559 2934 3193 3009
rect 3354 2524 3687 3724
rect -584 2499 13069 2524
rect -3355 2305 13069 2499
rect -3355 2194 -550 2305
rect -3355 2115 -2517 2194
rect -2348 2115 -779 2194
rect -610 2115 -550 2194
rect -3355 2092 -550 2115
rect -3355 1952 -3315 2092
rect -2761 1952 -1579 2092
rect -1025 1952 -550 2092
rect -3355 1912 -550 1952
rect -3166 1619 -569 1704
rect -3166 1436 -2963 1619
rect -693 1541 -569 1619
rect -626 1445 -569 1541
rect -3166 1362 -3089 1436
rect -3166 1311 -2963 1362
rect -693 1311 -569 1445
rect -3166 1247 -569 1311
rect -3359 902 -592 925
rect -3359 823 -2519 902
rect -2350 823 -785 902
rect -616 823 -592 902
rect -3359 800 -592 823
rect -3359 684 -3315 800
rect -3362 660 -3315 684
rect -2761 660 -1579 800
rect -1025 684 -592 800
rect -51 684 282 2305
rect 3354 684 3687 2305
rect 6623 684 6956 2305
rect 9928 684 10261 2305
rect -1025 660 12843 684
rect -3362 535 12843 660
rect -3163 255 -566 339
rect -3163 144 -2964 255
rect -694 249 -566 255
rect -632 153 -566 249
rect -3163 70 -3089 144
rect -3163 -53 -2964 70
rect -694 -53 -566 153
rect -3163 -118 -566 -53
rect -51 -774 282 535
rect 3354 -774 3687 535
rect 6623 -774 6956 535
rect 9928 -774 10261 535
rect -3359 -1031 13051 -774
rect -3359 -1071 -588 -1031
rect -3359 -1150 -2518 -1071
rect -2349 -1150 -783 -1071
rect -614 -1150 -588 -1071
rect -3359 -1173 -588 -1150
rect -3359 -1313 -3315 -1173
rect -2761 -1313 -1578 -1173
rect -1024 -1313 -588 -1173
rect -3359 -1352 -588 -1313
rect -3163 -1639 -566 -1572
rect -3163 -1829 -3002 -1639
rect -732 -1724 -566 -1639
rect -630 -1820 -566 -1724
rect -3163 -1903 -3089 -1829
rect -3163 -1947 -3002 -1903
rect -732 -1947 -566 -1820
rect -3163 -2029 -566 -1947
rect -3354 -2363 -587 -2341
rect -3354 -2442 -2516 -2363
rect -2347 -2442 -779 -2363
rect -610 -2442 -587 -2363
rect -3354 -2465 -587 -2442
rect -3354 -2605 -3315 -2465
rect -2761 -2605 -1579 -2465
rect -1025 -2584 -587 -2465
rect -51 -2584 282 -1031
rect 3354 -2584 3687 -1031
rect 6623 -2584 6956 -1031
rect 9928 -2584 10261 -1031
rect -1025 -2605 12851 -2584
rect -3354 -2733 12851 -2605
rect -3156 -3016 -559 -2947
rect -3156 -3017 -2512 -3016
rect -2363 -3017 -775 -3016
rect -3156 -3121 -3016 -3017
rect -626 -3112 -559 -3016
rect -3156 -3195 -3089 -3121
rect -3156 -3325 -3016 -3195
rect -746 -3325 -559 -3112
rect -3156 -3404 -559 -3325
rect -3356 -4043 -585 -4040
rect -51 -4043 282 -2733
rect 3354 -4043 3687 -2733
rect 6623 -4043 6956 -2733
rect 9928 -4043 10261 -2733
rect -3356 -4300 13039 -4043
rect -3356 -4335 -585 -4300
rect -3356 -4414 -2516 -4335
rect -2347 -4414 -783 -4335
rect -614 -4414 -585 -4335
rect -3356 -4437 -585 -4414
rect -3356 -4577 -3315 -4437
rect -2761 -4577 -1578 -4437
rect -1024 -4577 -585 -4437
rect -3356 -4618 -585 -4577
rect -3163 -4971 -566 -4907
rect -3163 -5093 -2974 -4971
rect -704 -4988 -566 -4971
rect -630 -5084 -566 -4988
rect -3163 -5167 -3089 -5093
rect -3163 -5279 -2974 -5167
rect -704 -5279 -566 -5084
rect -3163 -5364 -566 -5279
rect -3353 -5627 -586 -5603
rect -3353 -5706 -2516 -5627
rect -2347 -5706 -787 -5627
rect -618 -5706 -586 -5627
rect -3353 -5729 -586 -5706
rect -3353 -5845 -3315 -5729
rect -3355 -5869 -3315 -5845
rect -2761 -5869 -1578 -5729
rect -1024 -5845 -586 -5729
rect -51 -5845 282 -4300
rect 3354 -5845 3687 -4300
rect 6623 -5845 6956 -4300
rect 9928 -5845 10261 -4300
rect -1024 -5869 12850 -5845
rect -3355 -5994 12850 -5869
rect -3130 -6280 -592 -6214
rect -3130 -6304 -2512 -6280
rect -2363 -6304 -783 -6280
rect -3130 -6385 -2985 -6304
rect -634 -6376 -592 -6280
rect -3130 -6459 -3089 -6385
rect -3130 -6612 -2985 -6459
rect -715 -6612 -592 -6376
rect -3130 -6681 -592 -6612
<< via4 >>
rect -2943 3257 -2557 3348
rect -2557 3257 -2408 3348
rect -2408 3257 -673 3348
rect -2943 3248 -673 3257
rect -2943 3174 -2800 3248
rect -2800 3174 -1103 3248
rect -1103 3174 -763 3248
rect -763 3174 -673 3248
rect -2943 3040 -673 3174
rect 797 3257 1204 3317
rect 1204 3257 1353 3317
rect 1353 3257 2983 3317
rect 2983 3257 3067 3317
rect 797 3248 3067 3257
rect 797 3174 967 3248
rect 967 3174 2387 3248
rect 2387 3174 2727 3248
rect 2727 3174 3067 3248
rect 797 3009 3067 3174
rect -2963 1541 -693 1619
rect -2963 1445 -2513 1541
rect -2513 1445 -2364 1541
rect -2364 1445 -775 1541
rect -775 1445 -693 1541
rect -2963 1436 -693 1445
rect -2963 1362 -2749 1436
rect -2749 1362 -1353 1436
rect -1353 1362 -1013 1436
rect -1013 1362 -693 1436
rect -2963 1311 -693 1362
rect -2964 249 -694 255
rect -2964 153 -2515 249
rect -2515 153 -2366 249
rect -2366 153 -781 249
rect -781 153 -694 249
rect -2964 144 -694 153
rect -2964 70 -2749 144
rect -2749 70 -1353 144
rect -1353 70 -1013 144
rect -1013 70 -694 144
rect -2964 -53 -694 70
rect -3002 -1724 -732 -1639
rect -3002 -1820 -2514 -1724
rect -2514 -1820 -2365 -1724
rect -2365 -1820 -779 -1724
rect -779 -1820 -732 -1724
rect -3002 -1829 -732 -1820
rect -3002 -1903 -2749 -1829
rect -2749 -1903 -1352 -1829
rect -1352 -1903 -1012 -1829
rect -1012 -1903 -732 -1829
rect -3002 -1947 -732 -1903
rect -3016 -3112 -2512 -3017
rect -2512 -3112 -2363 -3017
rect -2363 -3112 -775 -3017
rect -775 -3112 -746 -3017
rect -3016 -3121 -746 -3112
rect -3016 -3195 -2749 -3121
rect -2749 -3195 -1353 -3121
rect -1353 -3195 -1013 -3121
rect -1013 -3195 -746 -3121
rect -3016 -3325 -746 -3195
rect -2974 -4988 -704 -4971
rect -2974 -5084 -2512 -4988
rect -2512 -5084 -2363 -4988
rect -2363 -5084 -779 -4988
rect -779 -5084 -704 -4988
rect -2974 -5093 -704 -5084
rect -2974 -5167 -2749 -5093
rect -2749 -5167 -1352 -5093
rect -1352 -5167 -1012 -5093
rect -1012 -5167 -704 -5093
rect -2974 -5279 -704 -5167
rect -2985 -6376 -2512 -6304
rect -2512 -6376 -2363 -6304
rect -2363 -6376 -783 -6304
rect -783 -6376 -715 -6304
rect -2985 -6385 -715 -6376
rect -2985 -6459 -2749 -6385
rect -2749 -6459 -1352 -6385
rect -1352 -6459 -1012 -6385
rect -1012 -6459 -715 -6385
rect -2985 -6612 -715 -6459
<< metal5 >>
rect -3818 3348 13360 4259
rect -3818 3040 -2943 3348
rect -673 3317 13360 3348
rect -673 3040 797 3317
rect -3818 3009 797 3040
rect 3067 3009 13360 3317
rect -3818 1619 13360 3009
rect -3818 1311 -2963 1619
rect -693 1311 13360 1619
rect -3818 255 13360 1311
rect -3818 -53 -2964 255
rect -694 -53 13360 255
rect -3818 -1639 13360 -53
rect -3818 -1947 -3002 -1639
rect -732 -1947 13360 -1639
rect -3818 -3017 13360 -1947
rect -3818 -3325 -3016 -3017
rect -746 -3325 13360 -3017
rect -3818 -4971 13360 -3325
rect -3818 -5279 -2974 -4971
rect -704 -5279 13360 -4971
rect -3818 -6304 13360 -5279
rect -3818 -6612 -2985 -6304
rect -715 -6612 13360 -6304
rect -3818 -7001 13360 -6612
use 4bit_ADDER  4bit_ADDER_0
timestamp 1736680159
transform 1 0 171 0 1 -165
box -174 -307 13189 3089
use 4bit_ADDER  4bit_ADDER_1
timestamp 1736680159
transform 1 0 171 0 1 -3430
box -174 -307 13189 3089
use 4bit_ADDER  4bit_ADDER_2
timestamp 1736680159
transform 1 0 171 0 1 -6694
box -174 -307 13189 3089
use NAND2  NAND2_0 ~/Desktop/vlsi_sky130b/design/mag/NAND/NAND2
timestamp 1736620191
transform 1 0 -3795 0 1 3170
box 356 -17 1062 804
use NAND2  NAND2_1
timestamp 1736620191
transform 1 0 -1758 0 1 3170
box 356 -17 1062 804
use NAND2  NAND2_2
timestamp 1736620191
transform 1 0 -28 0 1 3170
box 356 -17 1062 804
use NAND2  NAND2_3
timestamp 1736620191
transform 1 0 1732 0 1 3170
box 356 -17 1062 804
use NAND2  NAND2_4
timestamp 1736620191
transform 1 0 -3744 0 1 1358
box 356 -17 1062 804
use NAND2  NAND2_5
timestamp 1736620191
transform 1 0 -3744 0 1 66
box 356 -17 1062 804
use NAND2  NAND2_6
timestamp 1736620191
transform 1 0 -3744 0 1 -1907
box 356 -17 1062 804
use NAND2  NAND2_7
timestamp 1736620191
transform 1 0 -3744 0 1 -3199
box 356 -17 1062 804
use NAND2  NAND2_8
timestamp 1736620191
transform 1 0 -3744 0 1 -5171
box 356 -17 1062 804
use NAND2  NAND2_9
timestamp 1736620191
transform 1 0 -3744 0 1 -6463
box 356 -17 1062 804
use NAND2  NAND2_10
timestamp 1736620191
transform 1 0 -2008 0 1 1358
box 356 -17 1062 804
use NAND2  NAND2_11
timestamp 1736620191
transform 1 0 -2008 0 1 66
box 356 -17 1062 804
use NAND2  NAND2_12
timestamp 1736620191
transform 1 0 -2007 0 1 -1907
box 356 -17 1062 804
use NAND2  NAND2_13
timestamp 1736620191
transform 1 0 -2008 0 1 -3199
box 356 -17 1062 804
use NAND2  NAND2_14
timestamp 1736620191
transform 1 0 -2007 0 1 -5171
box 356 -17 1062 804
use NAND2  NAND2_15
timestamp 1736620191
transform 1 0 -2007 0 1 -6463
box 356 -17 1062 804
use inv  inv_0 ~/Desktop/vlsi_sky130b/design/mag/inv
timestamp 1736620191
transform 1 0 -2684 0 1 3542
box 0 -311 412 486
use inv  inv_1
timestamp 1736620191
transform 1 0 -664 0 1 3542
box 0 -311 412 486
use inv  inv_2
timestamp 1736620191
transform 1 0 1077 0 1 3542
box 0 -311 412 486
use inv  inv_3
timestamp 1736620191
transform 1 0 2856 0 1 3542
box 0 -311 412 486
use inv  inv_4
timestamp 1736620191
transform 1 0 -2642 0 1 438
box 0 -311 412 486
use inv  inv_5
timestamp 1736620191
transform 1 0 -2640 0 1 1730
box 0 -311 412 486
use inv  inv_6
timestamp 1736620191
transform 1 0 -2640 0 1 -1535
box 0 -311 412 486
use inv  inv_7
timestamp 1736620191
transform 1 0 -2639 0 1 -2827
box 0 -311 412 486
use inv  inv_8
timestamp 1736620191
transform 1 0 -2639 0 1 -4799
box 0 -311 412 486
use inv  inv_9
timestamp 1736620191
transform 1 0 -2639 0 1 -6091
box 0 -311 412 486
use inv  inv_10
timestamp 1736620191
transform 1 0 -902 0 1 1730
box 0 -311 412 486
use inv  inv_11
timestamp 1736620191
transform 1 0 -908 0 1 438
box 0 -311 412 486
use inv  inv_12
timestamp 1736620191
transform 1 0 -906 0 1 -1535
box 0 -311 412 486
use inv  inv_13
timestamp 1736620191
transform 1 0 -902 0 1 -2827
box 0 -311 412 486
use inv  inv_14
timestamp 1736620191
transform 1 0 -906 0 1 -4799
box 0 -311 412 486
use inv  inv_15
timestamp 1736620191
transform 1 0 -910 0 1 -6091
box 0 -311 412 486
<< labels >>
flabel metal2 -3228 -2190 -3108 -2070 1 FreeSerif 160 0 0 0 B2
port 7 n
flabel metal2 -3220 -5452 -3100 -5332 1 FreeSerif 160 0 0 0 B3
port 9 n
flabel metal2 -2952 -576 -2832 -456 1 FreeSerif 160 0 0 0 A1
port 11 n
flabel metal2 12820 3054 12940 3174 1 FreeSerif 160 0 0 0 SO
port 13 n
flabel metal3 -2146 -202 -2026 -82 1 FreeSerif 160 0 0 0 A2
port 10 n
flabel metal1 -3794 1646 -3674 1766 1 FreeSerif 160 0 0 0 A0
port 6 n
flabel metal3 -3190 2678 -3070 2798 1 FreeSerif 160 0 0 0 A3
port 12 n
flabel metal2 -3584 3886 -3464 4006 1 FreeSerif 160 0 0 0 B0
port 8 n
flabel metal2 54 -6728 150 -6642 1 FreeSerif 160 0 0 0 S7
port 19 n
flabel metal2 13182 -6664 13278 -6578 1 FreeSerif 160 0 0 0 S3
port 18 n
flabel metal2 9878 -6670 9974 -6584 1 FreeSerif 160 0 0 0 S4
port 17 n
flabel metal2 6586 -6668 6682 -6582 1 FreeSerif 160 0 0 0 S5
port 16 n
flabel metal2 13182 -3394 13278 -3308 1 FreeSerif 160 0 0 0 S2
port 15 n
flabel metal2 13166 -32 13262 54 1 FreeSerif 160 0 0 0 S1
port 14 n
flabel metal2 3294 -6664 3390 -6578 1 FreeSerif 160 0 0 0 S6
port 20 n
flabel metal5 5976 -6948 8074 -5352 0 FreeSans 160 0 0 0 VSS
port 21 nsew
flabel metal4 6690 2324 6822 2418 0 FreeSans 160 0 0 0 VDD
port 22 nsew
flabel metal2 -3562 1108 -3448 1226 0 FreeSans 160 0 0 0 B1
port 23 nsew
<< end >>
