magic
tech sky130B
magscale 1 2
timestamp 1732960014
<< nwell >>
rect -241 746 -208 765
<< ndiff >>
rect -62 224 185 524
<< poly >>
rect -172 801 -164 812
rect -172 796 -109 801
rect -356 602 -241 746
rect -172 713 -108 796
rect -174 707 -108 713
rect -356 568 -295 602
rect -258 568 -241 602
rect -356 550 -241 568
rect -198 705 -108 707
rect -198 671 -158 705
rect -121 671 -108 705
rect 21 699 97 812
rect -198 654 -108 671
rect -198 550 -145 654
rect -56 592 97 699
rect -56 588 48 592
rect 21 552 48 588
<< polycont >>
rect -295 568 -258 602
rect -158 671 -121 705
<< locali >>
rect -174 705 -105 796
rect -174 671 -158 705
rect -121 671 -105 705
rect -174 668 -105 671
rect -311 568 -295 602
rect -258 568 -242 602
<< viali >>
rect 37 762 71 796
rect -158 671 -121 705
rect -295 568 -258 602
<< metal1 >>
rect -407 1165 228 1227
rect 125 969 176 988
rect 125 847 181 969
rect 125 843 219 847
rect 298 843 351 989
rect -443 796 -121 815
rect 24 796 97 815
rect -443 746 -108 796
rect 24 762 37 796
rect 71 762 97 796
rect 24 741 97 762
rect -443 649 -410 718
rect -172 705 -108 718
rect -172 671 -158 705
rect -121 671 -108 705
rect -172 668 -108 671
rect 125 599 351 843
rect 125 524 198 599
rect -442 220 -318 225
rect -62 224 198 524
rect 226 332 351 524
rect 226 224 350 332
rect 275 223 350 224
rect -442 16 -340 220
rect 281 16 350 223
rect -442 -53 350 16
use efefetn  sky130_fd_pr__nfet_01v8_FBA633_0
timestamp 1732914314
transform 1 0 -39 0 1 374
box -404 -329 317 441
use efemosp  sky130_fd_pr__pfet_01v8_KFRNSS_0
timestamp 1732912614
transform 1 0 -90 0 1 1004
box -353 -261 410 223
<< labels >>
rlabel metal1 -443 779 -443 779 7 A
port 1 w
rlabel metal1 -443 649 -410 718 7 B
port 2 w
rlabel metal1 -442 552 -409 568 7 C
port 3 w
rlabel metal1 -442 -53 350 16 5 VSS
port 4 s
rlabel metal1 -407 1166 228 1227 1 VDD
port 5 n
rlabel metal1 298 599 351 989 3 Y
port 6 e
<< end >>
