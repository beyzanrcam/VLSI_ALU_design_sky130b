* NGSPICE file created from nor2_fix_pex.ext - technology: sky130B

.subckt nor2 A B VSS VDD Y
X0 VSS.t3 B.t0 Y.t4 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X1 Y.t0 A.t0 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X2 a_224_100.t2 A.t1 a_128_100.t1 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3 a_320_100.t0 A.t2 a_224_100.t1 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4 VDD.t6 A.t3 a_320_100.t1 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X5 a_512_100.t1 A.t4 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X6 a_704_100.t0 B.t1 a_224_100.t5 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X7 Y.t1 B.t2 a_704_100.t1 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X8 a_224_100.t0 A.t5 a_512_100.t0 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X9 a_896_100.t1 B.t3 Y.t2 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X10 a_224_100.t3 B.t4 a_896_100.t0 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X11 a_1088_100.t0 B.t5 a_224_100.t4 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X12 Y.t3 B.t6 a_1088_100.t1 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X13 a_128_100.t0 A.t6 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
R0 B.n0 B.t6 291.829
R1 B.n5 B.t0 239.393
R2 B.n4 B.t1 221.72
R3 B.n0 B.t5 221.72
R4 B.n1 B.t4 221.72
R5 B.n2 B.t3 221.72
R6 B.n3 B.t2 221.72
R7 B B.n5 162.648
R8 B.n5 B.n4 91.5805
R9 B.n1 B.n0 70.1096
R10 B.n2 B.n1 70.1096
R11 B.n3 B.n2 70.1096
R12 B.n4 B.n3 70.1096
R13 Y.n1 Y.t3 230.113
R14 Y.n1 Y.n0 198.593
R15 Y Y.n2 66.4022
R16 Y.n0 Y.t2 30.379
R17 Y.n0 Y.t1 30.379
R18 Y.n2 Y.t4 19.8005
R19 Y.n2 Y.t0 19.8005
R20 Y Y.n1 0.46012
R21 VSS.n1 VSS.t0 439.139
R22 VSS.n1 VSS.t2 387.476
R23 VSS VSS.n2 292.5
R24 VSS.n2 VSS.n1 292.5
R25 VSS VSS.t3 157.514
R26 VSS VSS.t1 153.499
R27 VSS.n2 VSS.n0 56.2862
R28 A.n0 A.t0 388.813
R29 A.n1 A.t6 291.829
R30 A.n4 A.t4 221.72
R31 A.n0 A.t5 221.72
R32 A.n3 A.t3 221.72
R33 A.n2 A.t2 221.72
R34 A.n1 A.t1 221.72
R35 A A.n4 162.286
R36 A.n4 A.n0 70.1096
R37 A.n4 A.n3 70.1096
R38 A.n3 A.n2 70.1096
R39 A.n2 A.n1 70.1096
R40 a_128_100.t0 a_128_100.t1 60.7575
R41 a_224_100.n2 a_224_100.n1 199.529
R42 a_224_100.n2 a_224_100.n0 199.529
R43 a_224_100.n3 a_224_100.n2 198.548
R44 a_224_100.n1 a_224_100.t1 30.379
R45 a_224_100.n1 a_224_100.t2 30.379
R46 a_224_100.n0 a_224_100.t4 30.379
R47 a_224_100.n0 a_224_100.t3 30.379
R48 a_224_100.n3 a_224_100.t5 30.379
R49 a_224_100.t0 a_224_100.n3 30.379
R50 VDD.n1 VDD.t1 317.539
R51 VDD.n1 VDD.n0 311.053
R52 VDD.n2 VDD.n1 185
R53 VDD.t10 VDD.t9 158.609
R54 VDD.t11 VDD.t10 158.609
R55 VDD.t12 VDD.t11 158.609
R56 VDD.t13 VDD.t12 158.609
R57 VDD.t14 VDD.t13 158.609
R58 VDD.t2 VDD.t14 158.609
R59 VDD.t3 VDD.t2 158.609
R60 VDD.t5 VDD.t3 158.609
R61 VDD.t7 VDD.t5 158.609
R62 VDD.t8 VDD.t7 158.609
R63 VDD.n2 VDD.t8 59.4788
R64 VDD.n0 VDD.t4 30.379
R65 VDD.n0 VDD.t6 30.379
R66 VDD VDD.n2 24.7831
R67 VDD VDD.t0 11.5657
R68 a_320_100.t0 a_320_100.t1 60.7575
R69 a_512_100.t0 a_512_100.t1 60.7575
R70 a_704_100.t0 a_704_100.t1 60.7575
R71 a_896_100.t0 a_896_100.t1 60.7575
R72 a_1088_100.t0 a_1088_100.t1 60.7575
C0 Y VDD 0.050931f
C1 Y B 0.261602f
C2 A VDD 0.216912f
C3 B A 0.636145f
C4 Y A 0.017971f
C5 B VDD 0.012666f
C6 Y VSS 0.698431f
C7 B VSS 0.602316f
C8 A VSS 0.428038f
C9 VDD VSS 2.4645f
.ends

