* NGSPICE file created from nor3_pex.ext - technology: sky130B

.subckt nor3 A B C VSS VDD Y
X0 a_329_726.t3 B.t0 a_683_726.t2 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.9309 pd=6.71 as=0.9309 ps=6.71 w=6.42 l=0.3
X1 VSS.t7 B.t1 Y.t3 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 VSS.t9 C.t0 Y.t5 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X3 a_683_726.t3 B.t2 a_329_726.t2 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.9309 pd=6.71 as=0.9309 ps=6.71 w=6.42 l=0.3
X4 Y.t1 C.t1 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X5 VDD.t11 A.t0 a_329_726.t5 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.9309 pd=6.71 as=0.9309 ps=6.71 w=6.42 l=0.3
X6 Y.t4 B.t3 VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X7 a_329_726.t0 A.t1 VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.9309 pd=6.71 as=0.9309 ps=6.71 w=6.42 l=0.3
X8 VSS.t11 A.t2 Y.t8 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X9 a_329_726.t4 A.t3 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.9309 pd=6.71 as=1.8618 ps=13.42 w=6.42 l=0.3
X10 Y.t2 A.t4 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X11 a_683_726.t0 C.t2 Y.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.9309 pd=6.71 as=0.9309 ps=6.71 w=6.42 l=0.3
X12 Y.t6 C.t3 a_683_726.t4 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.9309 pd=6.71 as=0.9309 ps=6.71 w=6.42 l=0.3
X13 Y.t7 C.t4 a_683_726.t5 VDD.t7 sky130_fd_pr__pfet_01v8 ad=1.8618 pd=13.42 as=0.9309 ps=6.71 w=6.42 l=0.3
X14 a_683_726.t1 B.t4 a_329_726.t1 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.9309 pd=6.71 as=0.9309 ps=6.71 w=6.42 l=0.3
R0 B.n0 B.t2 761.168
R1 B.n0 B.t4 761.168
R2 B.n0 B.t0 716.744
R3 B.n1 B.t3 296.695
R4 B.n1 B.t1 295.942
R5 B.n2 B.n0 80.7588
R6 B.n2 B.n1 72.1
R7 B B.n2 9.91402
R8 a_683_726.n2 a_683_726.n0 161.131
R9 a_683_726.n3 a_683_726.n2 161.131
R10 a_683_726.n2 a_683_726.n1 161.082
R11 a_683_726.n0 a_683_726.t2 4.44988
R12 a_683_726.n0 a_683_726.t3 4.44988
R13 a_683_726.n1 a_683_726.t4 4.44988
R14 a_683_726.n1 a_683_726.t1 4.44988
R15 a_683_726.n3 a_683_726.t5 4.44988
R16 a_683_726.t0 a_683_726.n3 4.44988
R17 a_329_726.n2 a_329_726.n0 153.799
R18 a_329_726.n2 a_329_726.n1 153.799
R19 a_329_726.n3 a_329_726.n2 153.799
R20 a_329_726.n0 a_329_726.t5 4.44988
R21 a_329_726.n0 a_329_726.t4 4.44988
R22 a_329_726.n1 a_329_726.t2 4.44988
R23 a_329_726.n1 a_329_726.t0 4.44988
R24 a_329_726.n3 a_329_726.t1 4.44988
R25 a_329_726.t3 a_329_726.n3 4.44988
R26 VDD.n2 VDD.n1 189.907
R27 VDD.n1 VDD.t9 165.531
R28 VDD.n1 VDD.n0 161.082
R29 VDD.t0 VDD.t7 62.8368
R30 VDD.t6 VDD.t0 62.8368
R31 VDD.t3 VDD.t6 62.8368
R32 VDD.t5 VDD.t3 62.8368
R33 VDD.t4 VDD.t5 62.8368
R34 VDD.t1 VDD.t4 62.8368
R35 VDD.t10 VDD.t1 62.8368
R36 VDD.n2 VDD.t10 46.329
R37 VDD VDD.t8 15.9758
R38 VDD.t8 VDD 11.7157
R39 VDD.n0 VDD.t2 4.44988
R40 VDD.n0 VDD.t11 4.44988
R41 VDD VDD.n2 0.533011
R42 Y.n1 Y.t7 158.25
R43 Y.n1 Y.n0 153.799
R44 Y.n4 Y.n2 66.4647
R45 Y.n4 Y.n3 66.3172
R46 Y.n6 Y.n5 66.3172
R47 Y.n2 Y.t8 17.4005
R48 Y.n2 Y.t2 17.4005
R49 Y.n3 Y.t3 17.4005
R50 Y.n3 Y.t4 17.4005
R51 Y.n5 Y.t5 17.4005
R52 Y.n5 Y.t1 17.4005
R53 Y.n0 Y.t0 4.44988
R54 Y.n0 Y.t6 4.44988
R55 Y Y.n6 0.361734
R56 Y Y.n1 0.279907
R57 Y.n6 Y.n4 0.148
R58 VSS.t0 VSS.t8 621.797
R59 VSS.t6 VSS.t0 621.797
R60 VSS.t4 VSS.t10 621.797
R61 VSS.t10 VSS.t2 621.797
R62 VSS.n2 VSS.t4 326.707
R63 VSS.n2 VSS.t6 295.091
R64 VSS.n5 VSS.n2 292.5
R65 VSS.n1 VSS.t9 173.957
R66 VSS.n4 VSS.t3 173.957
R67 VSS.n1 VSS.n0 126.043
R68 VSS.n4 VSS.n3 126.043
R69 VSS.n0 VSS.t1 17.4005
R70 VSS.n0 VSS.t7 17.4005
R71 VSS.n3 VSS.t5 17.4005
R72 VSS.n3 VSS.t11 17.4005
R73 VSS.n5 VSS.n4 15.6449
R74 VSS.n5 VSS.n1 14.8692
R75 VSS.n6 VSS.n5 2.3255
R76 VSS.n6 VSS 0.0106351
R77 VSS VSS.n6 0.0102128
R78 C.n0 C.t4 761.168
R79 C.n1 C.t3 716.744
R80 C.n0 C.t2 716.744
R81 C.n2 C.t1 296.695
R82 C.n2 C.t0 295.942
R83 C.n3 C.n2 111.812
R84 C.n1 C.n0 44.424
R85 C.n3 C.n1 41.4123
R86 C C.n3 10.2163
R87 A.n0 A.t3 761.168
R88 A.n0 A.t0 716.744
R89 A.n1 A.t1 716.744
R90 A.n2 A.t4 296.695
R91 A.n2 A.t2 295.942
R92 A.n3 A.n1 134.024
R93 A.n1 A.n0 44.424
R94 A.n3 A.n2 19.2005
R95 A A.n3 9.6181
C0 B C 0.999727f
C1 B VDD 0.044503f
C2 A C 0.090416f
C3 VDD A 0.212404f
C4 VDD C 0.071587f
C5 B Y 0.162988f
C6 A Y 0.104708f
C7 Y C 0.402085f
C8 VDD Y 0.061055f
C9 B A 0.554303f
C10 Y VSS 1.74713f
C11 C VSS 0.723721f
C12 B VSS 0.637601f
C13 A VSS 0.7537f
C14 VDD VSS 7.45947f
.ends

