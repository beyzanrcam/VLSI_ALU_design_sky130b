magic
tech sky130B
magscale 1 2
timestamp 1733246765
<< error_p >>
rect -773 -920 773 954
<< nwell >>
rect -773 -920 773 954
<< pmos >>
rect -679 -820 -619 892
rect -561 -820 -501 892
rect -443 -820 -383 892
rect -325 -820 -265 892
rect -207 -820 -147 892
rect -89 -820 -29 892
rect 29 -820 89 892
rect 147 -820 207 892
rect 265 -820 325 892
rect 383 -820 443 892
rect 501 -820 561 892
rect 619 -820 679 892
<< pdiff >>
rect -737 880 -679 892
rect -737 -808 -725 880
rect -691 -808 -679 880
rect -737 -820 -679 -808
rect -619 880 -561 892
rect -619 -808 -607 880
rect -573 -808 -561 880
rect -619 -820 -561 -808
rect -501 880 -443 892
rect -501 -808 -489 880
rect -455 -808 -443 880
rect -501 -820 -443 -808
rect -383 880 -325 892
rect -383 -808 -371 880
rect -337 -808 -325 880
rect -383 -820 -325 -808
rect -265 880 -207 892
rect -265 -808 -253 880
rect -219 -808 -207 880
rect -265 -820 -207 -808
rect -147 880 -89 892
rect -147 -808 -135 880
rect -101 -808 -89 880
rect -147 -820 -89 -808
rect -29 880 29 892
rect -29 -808 -17 880
rect 17 -808 29 880
rect -29 -820 29 -808
rect 89 880 147 892
rect 89 -808 101 880
rect 135 -808 147 880
rect 89 -820 147 -808
rect 207 880 265 892
rect 207 -808 219 880
rect 253 -808 265 880
rect 207 -820 265 -808
rect 325 880 383 892
rect 325 -808 337 880
rect 371 -808 383 880
rect 325 -820 383 -808
rect 443 880 501 892
rect 443 -808 455 880
rect 489 -808 501 880
rect 443 -820 501 -808
rect 561 880 619 892
rect 561 -808 573 880
rect 607 -808 619 880
rect 561 -820 619 -808
rect 679 880 737 892
rect 679 -808 691 880
rect 725 -808 737 880
rect 679 -820 737 -808
<< pdiffc >>
rect -725 -808 -691 880
rect -607 -808 -573 880
rect -489 -808 -455 880
rect -371 -808 -337 880
rect -253 -808 -219 880
rect -135 -808 -101 880
rect -17 -808 17 880
rect 101 -808 135 880
rect 219 -808 253 880
rect 337 -808 371 880
rect 455 -808 489 880
rect 573 -808 607 880
rect 691 -808 725 880
<< poly >>
rect -679 892 -619 918
rect -561 892 -501 918
rect -443 892 -383 918
rect -325 892 -265 918
rect -207 892 -147 918
rect -89 892 -29 918
rect 29 892 89 918
rect 147 892 207 918
rect 265 892 325 918
rect 383 892 443 918
rect 501 892 561 918
rect 619 892 679 918
rect -679 -851 -619 -820
rect -561 -851 -501 -820
rect -443 -851 -383 -820
rect -325 -851 -265 -820
rect -207 -851 -147 -820
rect -89 -851 -29 -820
rect 29 -851 89 -820
rect 147 -851 207 -820
rect 265 -851 325 -820
rect 383 -851 443 -820
rect 501 -851 561 -820
rect 619 -851 679 -820
rect -682 -867 -616 -851
rect -682 -901 -666 -867
rect -632 -901 -616 -867
rect -682 -917 -616 -901
rect -564 -867 -498 -851
rect -564 -901 -548 -867
rect -514 -901 -498 -867
rect -564 -917 -498 -901
rect -446 -867 -380 -851
rect -446 -901 -430 -867
rect -396 -901 -380 -867
rect -446 -917 -380 -901
rect -328 -867 -262 -851
rect -328 -901 -312 -867
rect -278 -901 -262 -867
rect -328 -917 -262 -901
rect -210 -867 -144 -851
rect -210 -901 -194 -867
rect -160 -901 -144 -867
rect -210 -917 -144 -901
rect -92 -867 -26 -851
rect -92 -901 -76 -867
rect -42 -901 -26 -867
rect -92 -917 -26 -901
rect 26 -867 92 -851
rect 26 -901 42 -867
rect 76 -901 92 -867
rect 26 -917 92 -901
rect 144 -867 210 -851
rect 144 -901 160 -867
rect 194 -901 210 -867
rect 144 -917 210 -901
rect 262 -867 328 -851
rect 262 -901 278 -867
rect 312 -901 328 -867
rect 262 -917 328 -901
rect 380 -867 446 -851
rect 380 -901 396 -867
rect 430 -901 446 -867
rect 380 -917 446 -901
rect 498 -867 564 -851
rect 498 -901 514 -867
rect 548 -901 564 -867
rect 498 -917 564 -901
rect 616 -867 682 -851
rect 616 -901 632 -867
rect 666 -901 682 -867
rect 616 -917 682 -901
<< polycont >>
rect -666 -901 -632 -867
rect -548 -901 -514 -867
rect -430 -901 -396 -867
rect -312 -901 -278 -867
rect -194 -901 -160 -867
rect -76 -901 -42 -867
rect 42 -901 76 -867
rect 160 -901 194 -867
rect 278 -901 312 -867
rect 396 -901 430 -867
rect 514 -901 548 -867
rect 632 -901 666 -867
<< locali >>
rect -725 880 -691 896
rect -725 -824 -691 -808
rect -607 880 -573 896
rect -607 -824 -573 -808
rect -489 880 -455 896
rect -489 -824 -455 -808
rect -371 880 -337 896
rect -371 -824 -337 -808
rect -253 880 -219 896
rect -253 -824 -219 -808
rect -135 880 -101 896
rect -135 -824 -101 -808
rect -17 880 17 896
rect -17 -824 17 -808
rect 101 880 135 896
rect 101 -824 135 -808
rect 219 880 253 896
rect 219 -824 253 -808
rect 337 880 371 896
rect 337 -824 371 -808
rect 455 880 489 896
rect 455 -824 489 -808
rect 573 880 607 896
rect 573 -824 607 -808
rect 691 880 725 896
rect 691 -824 725 -808
rect -682 -901 -666 -867
rect -632 -901 -616 -867
rect -564 -901 -548 -867
rect -514 -901 -498 -867
rect -446 -901 -430 -867
rect -396 -901 -380 -867
rect -328 -901 -312 -867
rect -278 -901 -262 -867
rect -210 -901 -194 -867
rect -160 -901 -144 -867
rect -92 -901 -76 -867
rect -42 -901 -26 -867
rect 26 -901 42 -867
rect 76 -901 92 -867
rect 144 -901 160 -867
rect 194 -901 210 -867
rect 262 -901 278 -867
rect 312 -901 328 -867
rect 380 -901 396 -867
rect 430 -901 446 -867
rect 498 -901 514 -867
rect 548 -901 564 -867
rect 616 -901 632 -867
rect 666 -901 682 -867
<< viali >>
rect -725 37 -691 880
rect -607 -808 -573 -45
rect -489 37 -455 880
rect -371 -808 -337 -45
rect -253 37 -219 880
rect -135 -808 -101 -45
rect -17 37 17 880
rect 101 -808 135 -45
rect 219 37 253 880
rect 337 -808 371 -45
rect 455 37 489 880
rect 573 -808 607 -45
rect 691 37 725 880
<< metal1 >>
rect -731 880 -685 892
rect -731 37 -725 880
rect -691 37 -685 880
rect -495 880 -449 892
rect -495 37 -489 880
rect -455 37 -449 880
rect -259 880 -213 892
rect -259 37 -253 880
rect -219 37 -213 880
rect -23 880 23 892
rect -23 37 -17 880
rect 17 37 23 880
rect 213 880 259 892
rect 213 37 219 880
rect 253 37 259 880
rect 449 880 495 892
rect 449 37 455 880
rect 489 37 495 880
rect 685 880 731 892
rect 685 37 691 880
rect 725 37 731 880
rect -613 -808 -607 -45
rect -573 -808 -567 -45
rect -613 -820 -567 -808
rect -377 -808 -371 -45
rect -337 -808 -331 -45
rect -377 -820 -331 -808
rect -141 -808 -135 -45
rect -101 -808 -95 -45
rect -141 -820 -95 -808
rect 95 -808 101 -45
rect 135 -808 141 -45
rect 95 -820 141 -808
rect 331 -808 337 -45
rect 371 -808 377 -45
rect 331 -820 377 -808
rect 567 -808 573 -45
rect 607 -808 613 -45
rect 567 -820 613 -808
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.56 l 0.30 m 1 nf 12 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
