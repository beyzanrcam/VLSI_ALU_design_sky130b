magic
tech sky130B
magscale 1 2
timestamp 1736595726
<< nwell >>
rect -76 872 3696 928
rect -76 510 3660 872
rect 311 509 417 510
rect 311 506 461 509
rect 336 398 461 506
rect 815 400 908 510
rect 1275 386 1541 510
rect 1731 386 1997 510
rect 2213 386 2479 510
rect 2713 386 2979 510
rect 3193 386 3459 510
<< metal1 >>
rect -76 736 -7 1143
rect 77 1074 129 1080
rect 77 876 129 1022
rect 404 735 473 1143
rect 558 1078 610 1084
rect 558 876 610 1026
rect 864 723 933 1143
rect 1023 1080 1075 1086
rect 1023 870 1075 1028
rect 1324 722 1393 1143
rect 1480 1082 1532 1088
rect 1480 867 1532 1030
rect 1804 719 1873 1143
rect 1949 1085 2001 1091
rect 1949 868 2001 1033
rect 2304 718 2373 1143
rect 2471 1085 2523 1091
rect 2471 867 2523 1033
rect 2784 721 2853 1143
rect 2954 1085 3006 1091
rect 2954 868 3006 1033
rect 3284 718 3353 1143
rect 3463 1079 3515 1085
rect 3463 869 3515 1027
rect 122 -195 211 89
rect 122 -290 211 -284
rect 288 -501 336 223
rect 603 -201 692 89
rect 603 -296 692 -290
rect 768 -501 816 237
rect 1045 -201 1134 89
rect 1045 -296 1134 -290
rect 1228 -501 1276 220
rect 1497 -196 1586 89
rect 1497 -291 1586 -285
rect 1688 -501 1736 219
rect 1972 -195 2061 89
rect 1972 -290 2061 -284
rect 2168 -501 2216 216
rect 2479 -199 2568 89
rect 2479 -294 2568 -288
rect 2668 -501 2716 219
rect 2965 -200 3054 89
rect 2965 -295 3054 -289
rect 3148 -501 3196 219
rect 3458 -207 3547 89
rect 3458 -302 3547 -296
rect 3648 -501 3696 229
<< via1 >>
rect 77 1022 129 1074
rect 558 1026 610 1078
rect 1023 1028 1075 1080
rect 1480 1030 1532 1082
rect 1949 1033 2001 1085
rect 2471 1033 2523 1085
rect 2954 1033 3006 1085
rect 3463 1027 3515 1079
rect 122 -284 211 -195
rect 603 -290 692 -201
rect 1045 -290 1134 -201
rect 1497 -285 1586 -196
rect 1972 -284 2061 -195
rect 2479 -288 2568 -199
rect 2965 -289 3054 -200
rect 3458 -296 3547 -207
<< metal2 >>
rect 62 1078 144 1089
rect 62 1018 73 1078
rect 133 1018 144 1078
rect 62 1007 144 1018
rect 543 1082 625 1093
rect 543 1022 554 1082
rect 614 1022 625 1082
rect 543 1011 625 1022
rect 1008 1084 1090 1095
rect 1008 1024 1019 1084
rect 1079 1024 1090 1084
rect 1008 1013 1090 1024
rect 1465 1086 1547 1097
rect 1465 1026 1476 1086
rect 1536 1026 1547 1086
rect 1465 1015 1547 1026
rect 1934 1089 2016 1100
rect 1934 1029 1945 1089
rect 2005 1029 2016 1089
rect 1934 1018 2016 1029
rect 2456 1089 2538 1100
rect 2456 1029 2467 1089
rect 2527 1029 2538 1089
rect 2456 1018 2538 1029
rect 2939 1089 3021 1100
rect 2939 1029 2950 1089
rect 3010 1029 3021 1089
rect 2939 1018 3021 1029
rect 3448 1083 3530 1094
rect 3448 1023 3459 1083
rect 3519 1023 3530 1083
rect 3448 1012 3530 1023
rect 113 -284 122 -195
rect 211 -284 220 -195
rect 598 -201 697 -190
rect 1040 -201 1139 -190
rect 1492 -196 1591 -185
rect 1967 -195 2066 -184
rect 597 -290 603 -201
rect 692 -290 698 -201
rect 1039 -290 1045 -201
rect 1134 -290 1140 -201
rect 1491 -285 1497 -196
rect 1586 -285 1592 -196
rect 1966 -284 1972 -195
rect 2061 -284 2067 -195
rect 2474 -199 2573 -188
rect 598 -301 697 -290
rect 1040 -301 1139 -290
rect 1492 -296 1591 -285
rect 1967 -295 2066 -284
rect 2473 -288 2479 -199
rect 2568 -288 2574 -199
rect 2960 -200 3059 -189
rect 2474 -299 2573 -288
rect 2959 -289 2965 -200
rect 3054 -289 3060 -200
rect 3453 -207 3552 -196
rect 2960 -300 3059 -289
rect 3452 -296 3458 -207
rect 3547 -296 3553 -207
rect 3453 -307 3552 -296
<< via2 >>
rect 73 1074 133 1078
rect 73 1022 77 1074
rect 77 1022 129 1074
rect 129 1022 133 1074
rect 73 1018 133 1022
rect 554 1078 614 1082
rect 554 1026 558 1078
rect 558 1026 610 1078
rect 610 1026 614 1078
rect 554 1022 614 1026
rect 1019 1080 1079 1084
rect 1019 1028 1023 1080
rect 1023 1028 1075 1080
rect 1075 1028 1079 1080
rect 1019 1024 1079 1028
rect 1476 1082 1536 1086
rect 1476 1030 1480 1082
rect 1480 1030 1532 1082
rect 1532 1030 1536 1082
rect 1476 1026 1536 1030
rect 1945 1085 2005 1089
rect 1945 1033 1949 1085
rect 1949 1033 2001 1085
rect 2001 1033 2005 1085
rect 1945 1029 2005 1033
rect 2467 1085 2527 1089
rect 2467 1033 2471 1085
rect 2471 1033 2523 1085
rect 2523 1033 2527 1085
rect 2467 1029 2527 1033
rect 2950 1085 3010 1089
rect 2950 1033 2954 1085
rect 2954 1033 3006 1085
rect 3006 1033 3010 1085
rect 2950 1029 3010 1033
rect 3459 1079 3519 1083
rect 3459 1027 3463 1079
rect 3463 1027 3515 1079
rect 3515 1027 3519 1079
rect 3459 1023 3519 1027
rect 122 -284 211 -195
rect 603 -290 692 -201
rect 1045 -290 1134 -201
rect 1497 -285 1586 -196
rect 1972 -284 2061 -195
rect 2479 -288 2568 -199
rect 2965 -289 3054 -200
rect 3458 -296 3547 -207
<< metal3 >>
rect 27 1083 191 1119
rect 27 1013 68 1083
rect 138 1013 191 1083
rect 27 980 191 1013
rect 527 1087 638 1102
rect 527 1017 549 1087
rect 619 1017 638 1087
rect 527 1002 638 1017
rect 991 1089 1106 1109
rect 991 1019 1014 1089
rect 1084 1019 1106 1089
rect 991 998 1106 1019
rect 1433 1091 1588 1114
rect 1433 1021 1471 1091
rect 1541 1021 1588 1091
rect 1433 997 1588 1021
rect 1903 1094 2054 1124
rect 1903 1024 1940 1094
rect 2010 1024 2054 1094
rect 1903 997 2054 1024
rect 2419 1094 2588 1124
rect 2419 1024 2462 1094
rect 2532 1024 2588 1094
rect 2419 997 2588 1024
rect 2907 1094 3062 1124
rect 2907 1024 2945 1094
rect 3015 1024 3062 1094
rect 2907 997 3062 1024
rect 3404 1088 3570 1122
rect 3404 1018 3454 1088
rect 3524 1018 3570 1088
rect 3404 997 3570 1018
rect 92 -190 242 -168
rect 92 -289 117 -190
rect 216 -289 242 -190
rect 92 -315 242 -289
rect 592 -295 598 -196
rect 697 -295 703 -196
rect 1034 -295 1040 -196
rect 1139 -295 1145 -196
rect 1486 -290 1492 -191
rect 1591 -290 1597 -191
rect 1961 -289 1967 -190
rect 2066 -289 2072 -190
rect 2468 -293 2474 -194
rect 2573 -293 2579 -194
rect 2954 -294 2960 -195
rect 3059 -294 3065 -195
rect 3447 -301 3453 -202
rect 3552 -301 3558 -202
<< via3 >>
rect 68 1078 138 1083
rect 68 1018 73 1078
rect 73 1018 133 1078
rect 133 1018 138 1078
rect 68 1013 138 1018
rect 549 1082 619 1087
rect 549 1022 554 1082
rect 554 1022 614 1082
rect 614 1022 619 1082
rect 549 1017 619 1022
rect 1014 1084 1084 1089
rect 1014 1024 1019 1084
rect 1019 1024 1079 1084
rect 1079 1024 1084 1084
rect 1014 1019 1084 1024
rect 1471 1086 1541 1091
rect 1471 1026 1476 1086
rect 1476 1026 1536 1086
rect 1536 1026 1541 1086
rect 1471 1021 1541 1026
rect 1940 1089 2010 1094
rect 1940 1029 1945 1089
rect 1945 1029 2005 1089
rect 2005 1029 2010 1089
rect 1940 1024 2010 1029
rect 2462 1089 2532 1094
rect 2462 1029 2467 1089
rect 2467 1029 2527 1089
rect 2527 1029 2532 1089
rect 2462 1024 2532 1029
rect 2945 1089 3015 1094
rect 2945 1029 2950 1089
rect 2950 1029 3010 1089
rect 3010 1029 3015 1089
rect 2945 1024 3015 1029
rect 3454 1083 3524 1088
rect 3454 1023 3459 1083
rect 3459 1023 3519 1083
rect 3519 1023 3524 1083
rect 3454 1018 3524 1023
rect 117 -195 216 -190
rect 117 -284 122 -195
rect 122 -284 211 -195
rect 211 -284 216 -195
rect 117 -289 216 -284
rect 598 -201 697 -196
rect 598 -290 603 -201
rect 603 -290 692 -201
rect 692 -290 697 -201
rect 598 -295 697 -290
rect 1040 -201 1139 -196
rect 1040 -290 1045 -201
rect 1045 -290 1134 -201
rect 1134 -290 1139 -201
rect 1040 -295 1139 -290
rect 1492 -196 1591 -191
rect 1492 -285 1497 -196
rect 1497 -285 1586 -196
rect 1586 -285 1591 -196
rect 1492 -290 1591 -285
rect 1967 -195 2066 -190
rect 1967 -284 1972 -195
rect 1972 -284 2061 -195
rect 2061 -284 2066 -195
rect 1967 -289 2066 -284
rect 2474 -199 2573 -194
rect 2474 -288 2479 -199
rect 2479 -288 2568 -199
rect 2568 -288 2573 -199
rect 2474 -293 2573 -288
rect 2960 -200 3059 -195
rect 2960 -289 2965 -200
rect 2965 -289 3054 -200
rect 3054 -289 3059 -200
rect 2960 -294 3059 -289
rect 3453 -207 3552 -202
rect 3453 -296 3458 -207
rect 3458 -296 3547 -207
rect 3547 -296 3552 -207
rect 3453 -301 3552 -296
<< metal4 >>
rect 27 1094 3570 1143
rect 27 1091 1940 1094
rect 27 1089 1471 1091
rect 27 1087 1014 1089
rect 27 1083 549 1087
rect 27 1013 68 1083
rect 138 1017 549 1083
rect 619 1019 1014 1087
rect 1084 1021 1471 1089
rect 1541 1024 1940 1091
rect 2010 1024 2462 1094
rect 2532 1024 2945 1094
rect 3015 1088 3570 1094
rect 3015 1024 3454 1088
rect 1541 1021 3454 1024
rect 1084 1019 3454 1021
rect 619 1018 3454 1019
rect 3524 1018 3570 1088
rect 619 1017 3570 1018
rect 138 1013 3570 1017
rect 27 997 3570 1013
rect 27 980 3568 997
<< via4 >>
rect 7 -190 327 -79
rect 7 -289 117 -190
rect 117 -289 216 -190
rect 216 -289 327 -190
rect 7 -399 327 -289
rect 488 -196 808 -85
rect 488 -295 598 -196
rect 598 -295 697 -196
rect 697 -295 808 -196
rect 488 -405 808 -295
rect 930 -196 1250 -85
rect 930 -295 1040 -196
rect 1040 -295 1139 -196
rect 1139 -295 1250 -196
rect 930 -405 1250 -295
rect 1382 -191 1702 -80
rect 1382 -290 1492 -191
rect 1492 -290 1591 -191
rect 1591 -290 1702 -191
rect 1382 -400 1702 -290
rect 1857 -190 2177 -79
rect 1857 -289 1967 -190
rect 1967 -289 2066 -190
rect 2066 -289 2177 -190
rect 1857 -399 2177 -289
rect 2364 -194 2684 -83
rect 2364 -293 2474 -194
rect 2474 -293 2573 -194
rect 2573 -293 2684 -194
rect 2364 -403 2684 -293
rect 2850 -195 3170 -84
rect 2850 -294 2960 -195
rect 2960 -294 3059 -195
rect 3059 -294 3170 -195
rect 2850 -404 3170 -294
rect 3343 -202 3663 -91
rect 3343 -301 3453 -202
rect 3453 -301 3552 -202
rect 3552 -301 3663 -202
rect 3343 -411 3663 -301
<< metal5 >>
rect -110 -24 435 -22
rect -110 -79 3853 -24
rect -110 -399 7 -79
rect 327 -80 1857 -79
rect 327 -85 1382 -80
rect 327 -399 488 -85
rect -110 -405 488 -399
rect 808 -405 930 -85
rect 1250 -400 1382 -85
rect 1702 -399 1857 -80
rect 2177 -83 3853 -79
rect 2177 -399 2364 -83
rect 1702 -400 2364 -399
rect 1250 -403 2364 -400
rect 2684 -84 3853 -83
rect 2684 -403 2850 -84
rect 1250 -404 2850 -403
rect 3170 -91 3853 -84
rect 3170 -404 3343 -91
rect 1250 -405 3343 -404
rect -110 -411 3343 -405
rect 3663 -411 3853 -91
rect -110 -501 3853 -411
use inv  inv_0 ~/Documents/vlsi/vlsi_sky130b/design/mag/inv
timestamp 1735843251
transform 1 0 1804 0 1 386
box 0 -311 412 486
use inv  inv_1
timestamp 1735843251
transform 1 0 -76 0 1 398
box 0 -311 412 486
use inv  inv_2
timestamp 1735843251
transform 1 0 404 0 1 400
box 0 -311 412 486
use inv  inv_3
timestamp 1735843251
transform 1 0 864 0 1 386
box 0 -311 412 486
use inv  inv_4
timestamp 1735843251
transform 1 0 1324 0 1 386
box 0 -311 412 486
use inv  inv_5
timestamp 1735843251
transform 1 0 2304 0 1 386
box 0 -311 412 486
use inv  inv_6
timestamp 1735843251
transform 1 0 2784 0 1 385
box 0 -311 412 486
use inv  inv_7
timestamp 1735843251
transform 1 0 3284 0 1 386
box 0 -311 412 486
<< labels >>
rlabel metal1 3652 -495 3687 -462 1 S0
port 9 n
rlabel metal1 3153 -488 3188 -455 1 S1
port 10 n
rlabel metal1 2674 -495 2709 -462 1 S2
port 11 n
rlabel metal1 2174 -496 2209 -463 1 S3
port 12 n
rlabel metal1 1694 -496 1729 -463 1 S4
port 13 n
rlabel metal1 1235 -496 1270 -463 1 S5
port 14 n
rlabel metal1 774 -496 809 -463 1 S6
port 15 n
rlabel metal1 294 -495 329 -462 1 S7
port 16 n
rlabel metal1 3293 1088 3344 1135 5 A0
port 8 s
rlabel metal1 2793 1090 2844 1137 5 A1
port 7 s
rlabel metal1 2312 1091 2363 1138 5 A2
port 6 s
rlabel metal1 1813 1090 1864 1137 5 A3
port 5 s
rlabel metal1 1332 1089 1383 1136 5 A4
port 4 s
rlabel metal1 872 1088 923 1135 5 A5
port 3 s
rlabel metal1 413 1091 464 1138 5 A6
port 2 s
rlabel metal1 -68 1091 -17 1138 5 A7
port 1 s
<< end >>
