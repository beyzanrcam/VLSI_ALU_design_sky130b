magic
tech sky130B
magscale 1 2
timestamp 1735598892
<< nwell >>
rect 2355 900 7564 1048
rect 8019 900 8528 1048
rect 2355 562 7528 900
rect 8088 562 8528 900
<< locali >>
rect 3121 900 3171 901
rect 3940 900 3990 901
rect 4759 900 4809 901
rect 5578 900 5628 901
rect 6397 900 6447 901
rect 7216 900 7266 901
rect 8035 900 8085 901
<< metal1 >>
rect 2286 980 2452 1164
rect 3105 980 3271 1164
rect 3924 980 4090 1164
rect 4743 980 4909 1164
rect 5562 980 5728 1164
rect 6381 980 6547 1164
rect 7200 980 7366 1164
rect 8019 980 8185 1164
rect 8255 1026 8261 1142
rect 8377 1048 8383 1142
rect 8377 1026 8528 1048
rect 8365 985 8528 1026
rect 2286 900 2355 980
rect 3105 900 3174 980
rect 3924 900 3993 980
rect 4743 900 4812 980
rect 5562 900 5631 980
rect 6381 900 6450 980
rect 7200 900 7269 980
rect 8019 900 8088 980
rect 8459 899 8528 985
rect 8466 891 8528 899
rect 3271 387 3286 448
rect 1564 74 1648 387
rect 2383 74 2467 387
rect 3202 74 3286 387
rect 4021 74 4105 387
rect 4840 74 4924 387
rect 5659 74 5743 387
rect 6478 74 6562 387
rect 7297 74 7381 387
rect 8116 348 8200 471
rect 8019 251 8200 348
rect 8019 74 8103 251
rect 1467 -110 1648 74
rect 2286 -110 2467 74
rect 3105 -110 3286 74
rect 3924 -110 4105 74
rect 4743 -110 4924 74
rect 5562 -110 5743 74
rect 6381 -110 6562 74
rect 7200 -110 7381 74
rect 7922 -110 8103 74
rect 8284 120 8381 251
rect 8284 17 8381 23
<< via1 >>
rect 8261 1026 8377 1142
rect 8284 23 8381 120
<< metal2 >>
rect 8255 1026 8261 1142
rect 8377 1026 8383 1142
rect 8275 23 8284 120
rect 8381 23 8390 120
<< via2 >>
rect 8266 1031 8372 1137
rect 8284 23 8381 120
<< metal3 >>
rect 8262 1142 8376 1147
rect 8261 1141 8377 1142
rect 8261 1027 8262 1141
rect 8376 1027 8377 1141
rect 8261 1026 8377 1027
rect 8262 1021 8376 1026
rect 8279 125 8386 131
rect 8279 12 8386 18
<< via3 >>
rect 8262 1137 8376 1141
rect 8262 1031 8266 1137
rect 8266 1031 8372 1137
rect 8372 1031 8376 1137
rect 8262 1027 8376 1031
rect 8279 120 8386 125
rect 8279 23 8284 120
rect 8284 23 8381 120
rect 8381 23 8386 120
rect 8279 18 8386 23
<< metal4 >>
rect 1901 1141 8377 1142
rect 1901 1027 8262 1141
rect 8376 1027 8377 1141
rect 1901 1026 8377 1027
<< via4 >>
rect 8196 125 8468 208
rect 8196 18 8279 125
rect 8279 18 8386 125
rect 8386 18 8468 125
rect 8196 -64 8468 18
<< metal5 >>
rect 1731 208 8511 251
rect 1731 -64 8196 208
rect 8468 -64 8511 208
rect 1731 -110 8511 -64
use buffer  buffer_0 ~/Documents/Dersler/VLSI/vlsi_sky130b/design/mag/inv
timestamp 1735596573
transform -1 0 6445 0 1 312
box -5 -422 786 852
use buffer  buffer_1
timestamp 1735596573
transform -1 0 2350 0 1 312
box -5 -422 786 852
use buffer  buffer_2
timestamp 1735596573
transform -1 0 3169 0 1 312
box -5 -422 786 852
use buffer  buffer_3
timestamp 1735596573
transform -1 0 3988 0 1 312
box -5 -422 786 852
use buffer  buffer_4
timestamp 1735596573
transform -1 0 4807 0 1 312
box -5 -422 786 852
use buffer  buffer_5
timestamp 1735596573
transform -1 0 5626 0 1 312
box -5 -422 786 852
use buffer  buffer_6
timestamp 1735596573
transform -1 0 8083 0 1 312
box -5 -422 786 852
use buffer  buffer_7
timestamp 1735596573
transform -1 0 7264 0 1 312
box -5 -422 786 852
use inv  inv_0 ~/Documents/Dersler/VLSI/vlsi_sky130b/design/mag/inv
timestamp 1735590487
transform -1 0 8528 0 1 562
box 0 -311 412 486
<< labels >>
rlabel metal1 8104 1164 8104 1164 5 A0
port 1 s
rlabel metal1 7282 1164 7282 1164 5 A1
port 2 s
rlabel metal1 6468 1164 6468 1164 5 A2
port 3 s
rlabel metal1 5646 1164 5646 1164 5 A3
port 4 s
rlabel metal1 4822 1164 4822 1164 5 A4
port 5 s
rlabel metal1 4003 1164 4003 1164 5 A5
port 6 s
rlabel metal1 3187 1164 3187 1164 5 A6
port 7 s
rlabel metal1 2373 1164 2373 1164 5 A7
port 8 s
rlabel metal1 8003 -110 8003 -110 5 S0
port 9 s
rlabel metal1 7289 -110 7289 -110 5 S1
port 10 s
rlabel metal1 6472 -110 6472 -110 5 S2
port 11 s
rlabel metal1 5653 -110 5653 -110 5 S3
port 12 s
rlabel metal1 4836 -110 4836 -110 5 S4
port 13 s
rlabel metal1 4017 -110 4017 -110 5 S5
port 14 s
rlabel metal1 3180 -110 3180 -110 5 S6
port 15 s
rlabel metal1 2385 -110 2385 -110 5 S7
port 16 s
rlabel metal1 1566 -110 1566 -110 5 C
port 17 s
rlabel metal4 4822 1142 4822 1142 5 VDD
port 18 s
rlabel metal5 4819 -110 4819 -110 5 VSS
port 19 s
<< end >>
