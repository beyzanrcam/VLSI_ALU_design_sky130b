magic
tech sky130B
magscale 1 2
timestamp 1733166153
<< error_p >>
rect -383 -131 -325 69
rect -265 -131 -207 69
rect -147 -131 -89 69
rect -29 -131 29 69
rect 89 -131 147 69
rect 207 -131 265 69
rect 325 -131 383 69
<< nmos >>
rect -325 -131 -265 69
rect -207 -131 -147 69
rect -89 -131 -29 69
rect 29 -131 89 69
rect 147 -131 207 69
rect 265 -131 325 69
<< ndiff >>
rect -383 57 -325 69
rect -383 -119 -371 57
rect -337 -119 -325 57
rect -383 -131 -325 -119
rect -265 57 -207 69
rect -265 -119 -253 57
rect -219 -119 -207 57
rect -265 -131 -207 -119
rect -147 57 -89 69
rect -147 -119 -135 57
rect -101 -119 -89 57
rect -147 -131 -89 -119
rect -29 57 29 69
rect -29 -119 -17 57
rect 17 -119 29 57
rect -29 -131 29 -119
rect 89 57 147 69
rect 89 -119 101 57
rect 135 -119 147 57
rect 89 -131 147 -119
rect 207 57 265 69
rect 207 -119 219 57
rect 253 -119 265 57
rect 207 -131 265 -119
rect 325 57 383 69
rect 325 -119 337 57
rect 371 -119 383 57
rect 325 -131 383 -119
<< ndiffc >>
rect -371 -119 -337 57
rect -253 -119 -219 57
rect -135 -119 -101 57
rect -17 -119 17 57
rect 101 -119 135 57
rect 219 -119 253 57
rect 337 -119 371 57
<< poly >>
rect -328 141 -262 157
rect -328 107 -312 141
rect -278 107 -262 141
rect -328 91 -262 107
rect -210 141 -144 157
rect -210 107 -194 141
rect -160 107 -144 141
rect -210 91 -144 107
rect -92 141 -26 157
rect -92 107 -76 141
rect -42 107 -26 141
rect -92 91 -26 107
rect 26 141 92 157
rect 26 107 42 141
rect 76 107 92 141
rect 26 91 92 107
rect 144 141 210 157
rect 144 107 160 141
rect 194 107 210 141
rect 144 91 210 107
rect 262 141 328 157
rect 262 107 278 141
rect 312 107 328 141
rect 262 91 328 107
rect -325 69 -265 91
rect -207 69 -147 91
rect -89 69 -29 91
rect 29 69 89 91
rect 147 69 207 91
rect 265 69 325 91
rect -325 -157 -265 -131
rect -207 -157 -147 -131
rect -89 -157 -29 -131
rect 29 -157 89 -131
rect 147 -157 207 -131
rect 265 -157 325 -131
<< polycont >>
rect -312 107 -278 141
rect -194 107 -160 141
rect -76 107 -42 141
rect 42 107 76 141
rect 160 107 194 141
rect 278 107 312 141
<< locali >>
rect -328 107 -312 141
rect -278 107 -262 141
rect -210 107 -194 141
rect -160 107 -144 141
rect -92 107 -76 141
rect -42 107 -26 141
rect 26 107 42 141
rect 76 107 92 141
rect 144 107 160 141
rect 194 107 210 141
rect 262 107 278 141
rect 312 107 328 141
rect -371 57 -337 73
rect -371 -135 -337 -119
rect -253 57 -219 73
rect -253 -135 -219 -119
rect -135 57 -101 73
rect -135 -135 -101 -119
rect -17 57 17 73
rect -17 -135 17 -119
rect 101 57 135 73
rect 101 -135 135 -119
rect 219 57 253 73
rect 219 -135 253 -119
rect 337 57 371 73
rect 337 -135 371 -119
<< viali >>
rect -371 -119 -337 57
rect -253 -119 -219 57
rect -135 -119 -101 57
rect -17 -119 17 57
rect 101 -119 135 57
rect 219 -119 253 57
rect 337 -119 371 57
<< metal1 >>
rect -377 57 -331 69
rect -377 -119 -371 57
rect -337 -119 -331 57
rect -377 -131 -331 -119
rect -259 57 -213 69
rect -259 -119 -253 57
rect -219 -119 -213 57
rect -259 -131 -213 -119
rect -141 57 -95 69
rect -141 -119 -135 57
rect -101 -119 -95 57
rect -141 -131 -95 -119
rect -23 57 23 69
rect -23 -119 -17 57
rect 17 -119 23 57
rect -23 -131 23 -119
rect 95 57 141 69
rect 95 -119 101 57
rect 135 -119 141 57
rect 95 -131 141 -119
rect 213 57 259 69
rect 213 -119 219 57
rect 253 -119 259 57
rect 213 -131 259 -119
rect 331 57 377 69
rect 331 -119 337 57
rect 371 -119 377 57
rect 331 -131 377 -119
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.30 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
