magic
tech sky130B
magscale 1 2
timestamp 1733249719
<< nwell >>
rect -530 1895 1099 3113
rect -530 1788 1013 1895
rect 1038 1788 1099 1895
rect -530 907 1099 1788
<< psubdiff >>
rect 17 -69 547 -1
rect 17 -182 81 -69
rect 467 -182 547 -69
rect 17 -258 547 -182
<< nsubdiff >>
rect -457 2941 -128 2989
rect -457 2868 -412 2941
rect -199 2868 -128 2941
rect -457 2813 -128 2868
<< psubdiffcont >>
rect 81 -182 467 -69
<< nsubdiffcont >>
rect -412 2868 -199 2941
<< locali >>
rect -457 2941 -128 2953
rect -457 2868 -412 2941
rect -199 2868 -128 2941
rect -457 2851 -128 2868
rect -400 966 -98 1000
rect -46 966 256 1000
rect 308 966 610 1000
rect 662 966 964 1000
rect -282 556 -216 966
rect 72 849 138 966
rect 426 849 492 966
rect 72 792 256 849
rect 190 671 256 792
rect 190 617 195 671
rect 247 617 256 671
rect -282 551 138 556
rect -282 497 -273 551
rect -221 497 138 551
rect -282 491 138 497
rect 190 491 256 617
rect 308 792 492 849
rect 780 911 846 966
rect 780 863 788 911
rect 839 863 846 911
rect 308 789 374 792
rect 308 735 316 789
rect 368 735 374 789
rect 308 491 374 735
rect 780 556 846 863
rect 426 491 846 556
rect 29 -1 63 49
rect 265 -1 299 49
rect 501 -1 535 49
rect 29 -69 535 -1
rect 29 -182 81 -69
rect 467 -182 535 -69
rect 29 -230 535 -182
<< viali >>
rect -412 2868 -199 2941
rect 195 617 247 671
rect -273 497 -221 551
rect 788 863 839 911
rect 316 735 368 789
<< metal1 >>
rect -450 2941 -167 2947
rect -450 2868 -412 2941
rect -199 2868 -167 2941
rect -450 2750 -167 2868
rect -449 1892 -167 2750
rect 23 1892 541 2759
rect 730 1892 1013 2759
rect -331 1047 187 1834
rect 377 1047 895 1834
rect -600 911 851 928
rect -600 863 788 911
rect 839 863 851 911
rect -600 846 851 863
rect -600 789 374 803
rect -600 735 316 789
rect 368 735 374 789
rect -600 715 374 735
rect -600 714 -485 715
rect -601 671 258 685
rect -601 617 195 671
rect 247 617 258 671
rect -601 597 258 617
rect -602 551 -198 568
rect -602 497 -273 551
rect -221 497 -198 551
rect -602 479 -198 497
rect 924 454 1013 1892
rect 369 453 1013 454
rect 141 231 1013 453
use sky130_fd_pr__nfet_01v8_VPSDAV  sky130_fd_pr__nfet_01v8_VPSDAV_0
timestamp 1733174963
transform 1 0 282 0 1 284
box -265 -257 265 257
use sky130_fd_pr__pfet_01v8_L8XZE7  sky130_fd_pr__pfet_01v8_L8XZE7_0
timestamp 1733246765
transform 1 0 282 0 1 1867
box -773 -920 773 954
<< labels >>
flabel metal1 -590 488 -523 557 1 FreeSerif 320 0 0 0 A
port 1 n
flabel metal1 -590 608 -523 677 1 FreeSerif 320 0 0 0 B
port 2 n
flabel metal1 -589 723 -522 792 1 FreeSerif 320 0 0 0 C
port 3 n
flabel metal1 -589 853 -522 922 1 FreeSerif 320 0 0 0 D
port 4 n
flabel metal1 869 297 997 427 1 FreeSerif 320 0 0 0 Y
port 5 n
flabel nwell -369 2833 -242 2945 1 FreeSerif 320 0 0 0 VDD
port 6 n
flabel psubdiffcont 218 -182 345 -70 1 FreeSerif 320 0 0 0 VSS
port 7 n
<< end >>
