magic
tech sky130B
magscale 1 2
timestamp 1734985533
<< nwell >>
rect -87 864 1371 1645
<< nmos >>
rect 7 367 37 497
rect 99 367 129 497
rect 195 367 225 497
rect 291 367 321 497
rect 387 367 417 497
rect 483 367 513 497
rect 579 367 609 497
rect 675 367 705 497
rect 771 367 801 497
rect 867 367 897 497
rect 963 367 993 497
rect 1059 367 1089 497
rect 1155 367 1185 497
rect 1247 367 1277 497
<< pmos >>
rect 7 987 37 1537
rect 99 987 129 1537
rect 195 987 225 1537
rect 291 987 321 1537
rect 387 987 417 1537
rect 483 987 513 1537
rect 579 987 609 1537
rect 675 987 705 1537
rect 771 987 801 1537
rect 867 987 897 1537
rect 963 987 993 1537
rect 1059 987 1089 1537
rect 1155 987 1185 1537
rect 1247 987 1277 1537
<< ndiff >>
rect -51 485 7 497
rect -51 379 -39 485
rect -5 379 7 485
rect -51 367 7 379
rect 37 485 99 497
rect 37 379 49 485
rect 83 379 99 485
rect 37 367 99 379
rect 129 485 195 497
rect 129 379 145 485
rect 179 379 195 485
rect 129 367 195 379
rect 225 485 291 497
rect 225 379 241 485
rect 275 379 291 485
rect 225 367 291 379
rect 321 485 387 497
rect 321 379 337 485
rect 371 379 387 485
rect 321 367 387 379
rect 417 485 483 497
rect 417 379 433 485
rect 467 379 483 485
rect 417 367 483 379
rect 513 485 579 497
rect 513 379 529 485
rect 563 379 579 485
rect 513 367 579 379
rect 609 485 675 497
rect 609 379 625 485
rect 659 379 675 485
rect 609 367 675 379
rect 705 485 771 497
rect 705 379 721 485
rect 755 379 771 485
rect 705 367 771 379
rect 801 485 867 497
rect 801 379 817 485
rect 851 379 867 485
rect 801 367 867 379
rect 897 485 963 497
rect 897 379 913 485
rect 947 379 963 485
rect 897 367 963 379
rect 993 485 1059 497
rect 993 379 1009 485
rect 1043 379 1059 485
rect 993 367 1059 379
rect 1089 485 1155 497
rect 1089 379 1105 485
rect 1139 379 1155 485
rect 1089 367 1155 379
rect 1185 485 1247 497
rect 1185 379 1201 485
rect 1235 379 1247 485
rect 1185 367 1247 379
rect 1277 485 1335 497
rect 1277 379 1289 485
rect 1323 379 1335 485
rect 1277 367 1335 379
<< pdiff >>
rect -51 1525 7 1537
rect -51 999 -39 1525
rect -5 999 7 1525
rect -51 987 7 999
rect 37 1525 99 1537
rect 37 999 49 1525
rect 83 999 99 1525
rect 37 987 99 999
rect 129 1525 195 1537
rect 129 999 145 1525
rect 179 999 195 1525
rect 129 987 195 999
rect 225 1525 291 1537
rect 225 999 241 1525
rect 275 999 291 1525
rect 225 987 291 999
rect 321 1525 387 1537
rect 321 999 337 1525
rect 371 999 387 1525
rect 321 987 387 999
rect 417 1525 483 1537
rect 417 999 433 1525
rect 467 999 483 1525
rect 417 987 483 999
rect 513 1525 579 1537
rect 513 999 529 1525
rect 563 999 579 1525
rect 513 987 579 999
rect 609 1525 675 1537
rect 609 999 625 1525
rect 659 999 675 1525
rect 609 987 675 999
rect 705 1525 771 1537
rect 705 999 721 1525
rect 755 999 771 1525
rect 705 987 771 999
rect 801 1525 867 1537
rect 801 999 817 1525
rect 851 999 867 1525
rect 801 987 867 999
rect 897 1525 963 1537
rect 897 999 913 1525
rect 947 999 963 1525
rect 897 987 963 999
rect 993 1525 1059 1537
rect 993 999 1009 1525
rect 1043 999 1059 1525
rect 993 987 1059 999
rect 1089 1525 1155 1537
rect 1089 999 1105 1525
rect 1139 999 1155 1525
rect 1089 987 1155 999
rect 1185 1525 1247 1537
rect 1185 999 1201 1525
rect 1235 999 1247 1525
rect 1185 987 1247 999
rect 1277 1525 1335 1537
rect 1277 999 1289 1525
rect 1323 999 1335 1525
rect 1277 987 1335 999
<< ndiffc >>
rect -39 379 -5 485
rect 49 379 83 485
rect 145 379 179 485
rect 241 379 275 485
rect 337 379 371 485
rect 433 379 467 485
rect 529 379 563 485
rect 625 379 659 485
rect 721 379 755 485
rect 817 379 851 485
rect 913 379 947 485
rect 1009 379 1043 485
rect 1105 379 1139 485
rect 1201 379 1235 485
rect 1289 379 1323 485
<< pdiffc >>
rect -39 999 -5 1525
rect 49 999 83 1525
rect 145 999 179 1525
rect 241 999 275 1525
rect 337 999 371 1525
rect 433 999 467 1525
rect 529 999 563 1525
rect 625 999 659 1525
rect 721 999 755 1525
rect 817 999 851 1525
rect 913 999 947 1525
rect 1009 999 1043 1525
rect 1105 999 1139 1525
rect 1201 999 1235 1525
rect 1289 999 1323 1525
<< poly >>
rect 7 1537 37 1563
rect 99 1537 129 1568
rect 195 1537 225 1568
rect 291 1537 321 1568
rect 387 1537 417 1568
rect 483 1537 513 1568
rect 579 1537 609 1568
rect 675 1537 705 1568
rect 771 1537 801 1568
rect 867 1537 897 1568
rect 963 1537 993 1568
rect 1059 1537 1089 1568
rect 1155 1537 1185 1568
rect 1247 1537 1277 1563
rect 7 956 37 987
rect 99 956 129 987
rect 195 956 225 987
rect 291 956 321 987
rect 387 957 417 987
rect 483 957 513 987
rect 579 957 609 987
rect -26 806 323 956
rect 387 928 609 957
rect 387 883 417 928
rect 547 883 609 928
rect 387 864 609 883
rect 675 956 705 987
rect 771 956 801 987
rect 867 956 897 987
rect 675 926 897 956
rect 675 888 739 926
rect 866 888 897 926
rect 675 863 897 888
rect 963 956 993 987
rect 1059 956 1089 987
rect 1155 956 1185 987
rect 963 890 1185 956
rect -87 697 897 806
rect -26 522 50 697
rect 99 607 321 632
rect 99 572 128 607
rect 300 572 321 607
rect 7 497 37 522
rect 99 519 321 572
rect 99 497 129 519
rect 195 497 225 519
rect 291 497 321 519
rect 387 599 609 627
rect 387 554 425 599
rect 555 554 609 599
rect 387 519 609 554
rect 387 497 417 519
rect 483 497 513 519
rect 579 497 609 519
rect 675 519 897 697
rect 675 497 705 519
rect 771 497 801 519
rect 867 497 897 519
rect 963 667 1107 890
rect 1247 841 1277 987
rect 1162 822 1277 841
rect 1162 750 1186 822
rect 1232 750 1277 822
rect 1162 732 1277 750
rect 963 592 1000 667
rect 1082 592 1107 667
rect 963 586 1107 592
rect 963 519 1185 586
rect 963 497 993 519
rect 1059 497 1089 519
rect 1155 497 1185 519
rect 1247 497 1277 732
rect 7 341 37 367
rect 99 341 129 367
rect 195 341 225 367
rect 291 341 321 367
rect 387 341 417 367
rect 483 341 513 367
rect 579 341 609 367
rect 675 341 705 367
rect 771 341 801 367
rect 867 341 897 367
rect 963 341 993 367
rect 1059 341 1089 367
rect 1155 341 1185 367
rect 1247 341 1277 367
<< polycont >>
rect 417 883 547 928
rect 739 888 866 926
rect 128 572 300 607
rect 425 554 555 599
rect 1186 750 1232 822
rect 1000 592 1082 667
<< locali >>
rect -39 1525 -5 1541
rect -39 938 -5 999
rect 49 1525 83 1541
rect 49 983 83 999
rect 145 1525 179 1541
rect 145 983 179 999
rect 241 1525 275 1541
rect 241 983 275 999
rect 337 1525 371 1541
rect 337 983 371 999
rect 433 1525 467 1541
rect 433 983 467 999
rect 529 1525 563 1541
rect 529 983 563 999
rect 625 1525 659 1541
rect 625 956 659 999
rect 721 1525 755 1541
rect 721 983 755 999
rect 817 1525 851 1541
rect 817 983 851 999
rect 913 1525 947 1541
rect 913 983 947 999
rect 1009 1525 1043 1541
rect 1009 983 1043 999
rect 1105 1525 1139 1541
rect 1105 983 1139 999
rect 1201 1525 1235 1541
rect 1201 983 1235 999
rect 1289 1525 1323 1541
rect -39 928 563 938
rect -39 883 417 928
rect 547 883 563 928
rect -39 869 563 883
rect -39 485 -5 869
rect 99 621 321 632
rect 99 562 118 621
rect 309 562 321 621
rect 99 547 321 562
rect 398 599 563 869
rect 398 554 425 599
rect 555 554 563 599
rect 398 537 563 554
rect 609 730 675 956
rect 721 933 1106 946
rect 721 876 733 933
rect 874 876 1106 933
rect 721 868 1106 876
rect 816 849 1106 868
rect 816 839 1249 849
rect 953 822 1249 839
rect 953 750 1186 822
rect 1232 750 1249 822
rect 609 696 777 730
rect 953 724 1249 750
rect 609 619 661 696
rect 747 619 777 696
rect 1289 683 1323 999
rect 609 591 777 619
rect 974 667 1323 683
rect 974 592 1000 667
rect 1082 592 1323 667
rect 609 526 675 591
rect 974 564 1323 592
rect -39 363 -5 379
rect 49 485 83 501
rect 49 363 83 379
rect 145 500 179 501
rect 145 363 179 379
rect 241 485 275 501
rect 241 363 275 365
rect 337 500 371 501
rect 337 363 371 379
rect 433 485 467 501
rect 433 363 467 365
rect 529 499 563 501
rect 529 363 563 379
rect 625 485 659 526
rect 625 363 659 365
rect 721 500 755 501
rect 721 363 755 379
rect 817 485 851 501
rect 817 363 851 365
rect 913 500 947 501
rect 913 363 947 379
rect 1009 485 1043 501
rect 1009 363 1043 365
rect 1105 500 1139 501
rect 1105 363 1139 379
rect 1201 485 1235 501
rect 1201 363 1235 379
rect 1289 485 1323 564
rect 1289 363 1323 379
<< viali >>
rect 49 1417 83 1519
rect 49 1022 83 1124
rect 145 1209 179 1333
rect 241 1417 275 1519
rect 241 1058 275 1124
rect 337 1209 371 1333
rect 433 1415 467 1517
rect 433 1058 467 1118
rect 529 1209 563 1333
rect 625 1414 659 1516
rect 625 1058 659 1101
rect 721 1209 755 1333
rect 817 1414 851 1516
rect 817 1058 851 1118
rect 913 1209 947 1333
rect 1009 1414 1043 1516
rect 1009 1058 1043 1125
rect 1105 1208 1139 1332
rect 1201 1414 1235 1516
rect 1201 1058 1235 1125
rect 118 607 309 621
rect 118 572 128 607
rect 128 572 300 607
rect 300 572 309 607
rect 118 562 309 572
rect 733 926 874 933
rect 733 888 739 926
rect 739 888 866 926
rect 866 888 874 926
rect 733 876 874 888
rect 661 619 747 696
rect 145 485 179 500
rect 145 466 179 485
rect 241 379 275 399
rect 241 365 275 379
rect 337 485 371 500
rect 337 466 371 485
rect 433 379 467 399
rect 433 365 467 379
rect 529 485 563 499
rect 529 465 563 485
rect 625 379 659 399
rect 625 365 659 379
rect 721 485 755 500
rect 721 466 755 485
rect 817 379 851 399
rect 817 365 851 379
rect 913 485 947 500
rect 913 466 947 485
rect 1009 379 1043 399
rect 1009 365 1043 379
rect 1105 485 1139 500
rect 1105 466 1139 485
<< metal1 >>
rect 37 1588 1247 1645
rect 37 1519 291 1588
rect 37 1417 49 1519
rect 83 1417 241 1519
rect 275 1417 291 1519
rect 37 1396 291 1417
rect 417 1517 867 1543
rect 417 1415 433 1517
rect 467 1516 867 1517
rect 467 1415 625 1516
rect 417 1414 625 1415
rect 659 1414 817 1516
rect 851 1414 867 1516
rect 417 1396 867 1414
rect 993 1516 1247 1588
rect 993 1414 1009 1516
rect 1043 1414 1201 1516
rect 1235 1414 1247 1516
rect 993 1396 1247 1414
rect 129 1333 1155 1358
rect 129 1209 145 1333
rect 179 1209 337 1333
rect 371 1209 529 1333
rect 563 1209 721 1333
rect 755 1209 913 1333
rect 947 1332 1155 1333
rect 947 1209 1105 1332
rect 129 1208 1105 1209
rect 1139 1208 1155 1332
rect 129 1179 1155 1208
rect 37 1124 291 1146
rect 37 1022 49 1124
rect 83 1058 241 1124
rect 275 1058 291 1124
rect 83 1022 291 1058
rect 417 1118 867 1135
rect 417 1058 433 1118
rect 467 1101 817 1118
rect 467 1058 625 1101
rect 659 1058 817 1101
rect 851 1058 867 1118
rect 417 1043 867 1058
rect 993 1125 1247 1146
rect 993 1058 1009 1125
rect 1043 1058 1201 1125
rect 1235 1058 1247 1125
rect 37 999 291 1022
rect 993 999 1247 1058
rect 712 933 898 949
rect 712 876 733 933
rect 874 876 898 933
rect 712 857 898 876
rect 112 769 898 857
rect 112 685 335 769
rect 648 696 1371 734
rect -87 621 336 685
rect -87 562 118 621
rect 309 562 336 621
rect 648 619 661 696
rect 747 619 1371 696
rect 648 602 1371 619
rect -87 542 336 562
rect 42 313 97 501
rect 129 500 579 512
rect 129 466 145 500
rect 179 466 337 500
rect 371 499 579 500
rect 371 466 529 499
rect 129 465 529 466
rect 563 465 579 499
rect 129 444 579 465
rect 705 500 1155 512
rect 705 466 721 500
rect 755 466 913 500
rect 947 466 1105 500
rect 1139 466 1155 500
rect 705 444 1155 466
rect 227 399 292 416
rect 227 365 241 399
rect 275 365 292 399
rect 227 313 292 365
rect 420 399 867 411
rect 420 365 433 399
rect 467 365 625 399
rect 659 365 817 399
rect 851 365 867 399
rect 420 347 867 365
rect 993 399 1058 415
rect 993 365 1009 399
rect 1043 365 1058 399
rect 993 313 1058 365
rect 1189 313 1244 501
rect 42 243 1244 313
<< end >>
