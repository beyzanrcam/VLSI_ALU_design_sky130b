* NGSPICE file created from ZFLAG.ext - technology: sky130B

.subckt sky130_fd_pr__pfet_01v8_64A2S3 a_n33_n428# a_447_n428# a_n605_n428# a_321_n484#
+ a_n543_n484# a_543_n428# a_159_n428# a_33_n484# a_n255_n484# a_255_n428# w_n641_n484#
+ a_351_n428# a_n417_n428# a_n513_n428# a_n129_n428# a_63_n428# a_n225_n428# a_n321_n428#
X0 a_447_n428# a_321_n484# a_351_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X1 a_n513_n428# a_n543_n484# a_n605_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=1.3268 ps=9.18 w=4.28 l=0.15
X2 a_63_n428# a_33_n484# a_n33_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X3 a_n129_n428# a_n255_n484# a_n225_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X4 a_n417_n428# a_n543_n484# a_n513_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X5 a_n33_n428# a_n255_n484# a_n129_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X6 a_351_n428# a_321_n484# a_255_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X7 a_255_n428# a_33_n484# a_159_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X8 a_n321_n428# a_n543_n484# a_n417_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X9 a_543_n428# a_321_n484# a_447_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=1.3268 pd=9.18 as=0.7062 ps=4.61 w=4.28 l=0.15
X10 a_159_n428# a_33_n484# a_63_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
X11 a_n225_n428# a_n255_n484# a_n321_n428# w_n641_n484# sky130_fd_pr__pfet_01v8 ad=0.7062 pd=4.61 as=0.7062 ps=4.61 w=4.28 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_S9NJ5Q a_159_n100# a_n159_n126# a_33_n126# a_n129_n100#
+ a_n221_n100# a_63_n100# a_n63_n126# a_n33_n100# a_129_n126# VSUBS
X0 a_n129_n100# a_n159_n126# a_n221_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1 a_63_n100# a_33_n126# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2 a_n33_n100# a_n63_n126# a_n129_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_159_n100# a_129_n126# a_63_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt nor4 A B C D VSS Y VDD
Xsky130_fd_pr__pfet_01v8_64A2S3_0 m1_n20_1047# m1_268_1523# VDD D A Y m1_n20_1047#
+ C B m1_268_1523# VDD Y VDD m1_n308_1523# m1_n308_1523# m1_268_1523# m1_n20_1047#
+ m1_n308_1523# sky130_fd_pr__pfet_01v8_64A2S3
Xsky130_fd_pr__nfet_01v8_S9NJ5Q_0 VSS A C Y VSS Y B VSS D VSS sky130_fd_pr__nfet_01v8_S9NJ5Q
.ends

.subckt sky130_fd_pr__nfet_01v8_6H9P4D a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt efepmos_W107-L15-F3 a_n129_n204# a_n173_n107# w_n209_n207# a_n81_n107#
X0 a_n81_n107# a_n129_n204# a_n173_n107# w_n209_n207# sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
X1 a_n81_n107# a_n129_n204# a_n173_n107# w_n209_n207# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2 a_n173_n107# a_n129_n204# a_n81_n107# w_n209_n207# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
.ends

.subckt inv A VSS VDD Y
Xsky130_fd_pr__nfet_01v8_6H9P4D_0 Y VSS A VSS sky130_fd_pr__nfet_01v8_6H9P4D
Xefepmos_W107-L15-F3_0 A VDD VDD Y efepmos_W107-L15-F3
.ends

.subckt nmos_2shared_W200-L015-F1 a_63_n200# a_n63_n226# a_n33_n200# a_33_n226# a_n125_n200#
+ VSUBS
X0 a_n33_n200# a_n63_n226# a_n125_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1 a_63_n200# a_33_n226# a_n33_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
.ends

.subckt pmos_p2-w321-L015-f3 a_n317_n107# w_n353_n143# a_n225_n107# a_33_n138# a_n255_n138#
X0 a_n225_n107# a_33_n138# a_n317_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X1 a_n225_n107# a_n255_n138# a_n317_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.3317 ps=2.76 w=1.07 l=0.15
X2 a_n317_n107# a_33_n138# a_n225_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X3 a_n317_n107# a_n255_n138# a_n225_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X4 a_n225_n107# a_n255_n138# a_n317_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.17655 ps=1.4 w=1.07 l=0.15
X5 a_n317_n107# a_33_n138# a_n225_n107# w_n353_n143# sky130_fd_pr__pfet_01v8 ad=0.3317 pd=2.76 as=0.17655 ps=1.4 w=1.07 l=0.15
.ends

.subckt NAND2 A B VSS VDD Y
Xnmos_2shared_W200-L015-F1_0 VSS B a_994_146# A Y VSS nmos_2shared_W200-L015-F1
Xpmos_p2-w321-L015-f3_0 VDD VDD Y B A pmos_p2-w321-L015-f3
.ends

.subckt ZFLAG A0 A1 A2 A3 A4 A5 A6 A7 Z VSS VDD
Xnor4_0 A3 A2 A1 A0 VSS nor4_0/Y VDD nor4
Xnor4_1 A4 A5 A6 A7 VSS nor4_1/Y VDD nor4
Xinv_0 inv_0/A VSS VDD Z inv
XNAND2_0 nor4_0/Y nor4_1/Y VSS VDD inv_0/A NAND2
.ends

